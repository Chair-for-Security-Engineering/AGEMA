/* modified netlist. Source: module AES in file /mnt/c/Users/Amir/Desktop/Papers_in_progress/AGEMA/Designs/AES_serial/AGEMA/sbox_opt3/AES.v */
/* 8 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 9 register stage(s) in total */

module AES_HPC2_AIG_Pipeline_d1 (plaintext_s0, key_s0, clk, start, plaintext_s1, key_s1, Fresh, ciphertext_s0, done, ciphertext_s1);
    input [127:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input start ;
    input [127:0] plaintext_s1 ;
    input [127:0] key_s1 ;
    input [33:0] Fresh ;
    output [127:0] ciphertext_s0 ;
    output done ;
    output [127:0] ciphertext_s1 ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_415 ;
    wire signal_416 ;
    wire signal_417 ;
    wire signal_418 ;
    wire signal_419 ;
    wire signal_420 ;
    wire signal_421 ;
    wire signal_422 ;
    wire signal_423 ;
    wire signal_424 ;
    wire signal_425 ;
    wire signal_426 ;
    wire signal_427 ;
    wire signal_428 ;
    wire signal_429 ;
    wire signal_431 ;
    wire signal_433 ;
    wire signal_435 ;
    wire signal_437 ;
    wire signal_439 ;
    wire signal_441 ;
    wire signal_444 ;
    wire signal_445 ;
    wire signal_446 ;
    wire signal_447 ;
    wire signal_448 ;
    wire signal_449 ;
    wire signal_450 ;
    wire signal_451 ;
    wire signal_452 ;
    wire signal_453 ;
    wire signal_454 ;
    wire signal_455 ;
    wire signal_456 ;
    wire signal_457 ;
    wire signal_458 ;
    wire signal_459 ;
    wire signal_460 ;
    wire signal_461 ;
    wire signal_462 ;
    wire signal_463 ;
    wire signal_464 ;
    wire signal_465 ;
    wire signal_467 ;
    wire signal_469 ;
    wire signal_471 ;
    wire signal_473 ;
    wire signal_475 ;
    wire signal_477 ;
    wire signal_479 ;
    wire signal_481 ;
    wire signal_483 ;
    wire signal_485 ;
    wire signal_487 ;
    wire signal_489 ;
    wire signal_491 ;
    wire signal_493 ;
    wire signal_495 ;
    wire signal_497 ;
    wire signal_499 ;
    wire signal_501 ;
    wire signal_503 ;
    wire signal_505 ;
    wire signal_507 ;
    wire signal_509 ;
    wire signal_511 ;
    wire signal_513 ;
    wire signal_515 ;
    wire signal_517 ;
    wire signal_519 ;
    wire signal_521 ;
    wire signal_523 ;
    wire signal_525 ;
    wire signal_527 ;
    wire signal_529 ;
    wire signal_531 ;
    wire signal_533 ;
    wire signal_535 ;
    wire signal_537 ;
    wire signal_539 ;
    wire signal_541 ;
    wire signal_543 ;
    wire signal_545 ;
    wire signal_547 ;
    wire signal_549 ;
    wire signal_551 ;
    wire signal_553 ;
    wire signal_555 ;
    wire signal_557 ;
    wire signal_559 ;
    wire signal_561 ;
    wire signal_563 ;
    wire signal_565 ;
    wire signal_567 ;
    wire signal_569 ;
    wire signal_571 ;
    wire signal_573 ;
    wire signal_575 ;
    wire signal_577 ;
    wire signal_579 ;
    wire signal_581 ;
    wire signal_583 ;
    wire signal_585 ;
    wire signal_587 ;
    wire signal_589 ;
    wire signal_591 ;
    wire signal_593 ;
    wire signal_595 ;
    wire signal_597 ;
    wire signal_599 ;
    wire signal_601 ;
    wire signal_603 ;
    wire signal_605 ;
    wire signal_607 ;
    wire signal_609 ;
    wire signal_611 ;
    wire signal_613 ;
    wire signal_615 ;
    wire signal_617 ;
    wire signal_619 ;
    wire signal_621 ;
    wire signal_623 ;
    wire signal_625 ;
    wire signal_627 ;
    wire signal_629 ;
    wire signal_631 ;
    wire signal_633 ;
    wire signal_635 ;
    wire signal_637 ;
    wire signal_639 ;
    wire signal_641 ;
    wire signal_643 ;
    wire signal_645 ;
    wire signal_647 ;
    wire signal_649 ;
    wire signal_651 ;
    wire signal_653 ;
    wire signal_655 ;
    wire signal_657 ;
    wire signal_659 ;
    wire signal_661 ;
    wire signal_663 ;
    wire signal_665 ;
    wire signal_667 ;
    wire signal_669 ;
    wire signal_671 ;
    wire signal_673 ;
    wire signal_675 ;
    wire signal_677 ;
    wire signal_679 ;
    wire signal_681 ;
    wire signal_683 ;
    wire signal_685 ;
    wire signal_687 ;
    wire signal_689 ;
    wire signal_691 ;
    wire signal_693 ;
    wire signal_695 ;
    wire signal_697 ;
    wire signal_699 ;
    wire signal_701 ;
    wire signal_703 ;
    wire signal_705 ;
    wire signal_707 ;
    wire signal_709 ;
    wire signal_711 ;
    wire signal_713 ;
    wire signal_715 ;
    wire signal_717 ;
    wire signal_719 ;
    wire signal_721 ;
    wire signal_722 ;
    wire signal_723 ;
    wire signal_724 ;
    wire signal_725 ;
    wire signal_726 ;
    wire signal_727 ;
    wire signal_728 ;
    wire signal_729 ;
    wire signal_730 ;
    wire signal_731 ;
    wire signal_732 ;
    wire signal_733 ;
    wire signal_734 ;
    wire signal_735 ;
    wire signal_736 ;
    wire signal_737 ;
    wire signal_738 ;
    wire signal_739 ;
    wire signal_740 ;
    wire signal_741 ;
    wire signal_742 ;
    wire signal_743 ;
    wire signal_744 ;
    wire signal_745 ;
    wire signal_746 ;
    wire signal_747 ;
    wire signal_748 ;
    wire signal_749 ;
    wire signal_750 ;
    wire signal_751 ;
    wire signal_752 ;
    wire signal_753 ;
    wire signal_754 ;
    wire signal_755 ;
    wire signal_756 ;
    wire signal_757 ;
    wire signal_758 ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_808 ;
    wire signal_809 ;
    wire signal_811 ;
    wire signal_812 ;
    wire signal_814 ;
    wire signal_815 ;
    wire signal_817 ;
    wire signal_818 ;
    wire signal_820 ;
    wire signal_821 ;
    wire signal_823 ;
    wire signal_824 ;
    wire signal_826 ;
    wire signal_827 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_841 ;
    wire signal_842 ;
    wire signal_844 ;
    wire signal_845 ;
    wire signal_847 ;
    wire signal_848 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_856 ;
    wire signal_857 ;
    wire signal_859 ;
    wire signal_860 ;
    wire signal_862 ;
    wire signal_863 ;
    wire signal_865 ;
    wire signal_866 ;
    wire signal_868 ;
    wire signal_869 ;
    wire signal_871 ;
    wire signal_872 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_904 ;
    wire signal_905 ;
    wire signal_907 ;
    wire signal_908 ;
    wire signal_910 ;
    wire signal_911 ;
    wire signal_913 ;
    wire signal_914 ;
    wire signal_916 ;
    wire signal_917 ;
    wire signal_919 ;
    wire signal_920 ;
    wire signal_922 ;
    wire signal_923 ;
    wire signal_925 ;
    wire signal_926 ;
    wire signal_928 ;
    wire signal_929 ;
    wire signal_931 ;
    wire signal_932 ;
    wire signal_934 ;
    wire signal_935 ;
    wire signal_937 ;
    wire signal_938 ;
    wire signal_940 ;
    wire signal_941 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1494 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1499 ;
    wire signal_1500 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1503 ;
    wire signal_1504 ;
    wire signal_1505 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1509 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1512 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1518 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1521 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1527 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1530 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1536 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1539 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1564 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1623 ;
    wire signal_1624 ;
    wire signal_1625 ;
    wire signal_1626 ;
    wire signal_1627 ;
    wire signal_1628 ;
    wire signal_1629 ;
    wire signal_1630 ;
    wire signal_1631 ;
    wire signal_1632 ;
    wire signal_1633 ;
    wire signal_1634 ;
    wire signal_1635 ;
    wire signal_1636 ;
    wire signal_1637 ;
    wire signal_1638 ;
    wire signal_1639 ;
    wire signal_1640 ;
    wire signal_1641 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1657 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1660 ;
    wire signal_1661 ;
    wire signal_1662 ;
    wire signal_1663 ;
    wire signal_1664 ;
    wire signal_1665 ;
    wire signal_1666 ;
    wire signal_1667 ;
    wire signal_1668 ;
    wire signal_1669 ;
    wire signal_1670 ;
    wire signal_1671 ;
    wire signal_1672 ;
    wire signal_1673 ;
    wire signal_1674 ;
    wire signal_1675 ;
    wire signal_1676 ;
    wire signal_1677 ;
    wire signal_1678 ;
    wire signal_1679 ;
    wire signal_1680 ;
    wire signal_1681 ;
    wire signal_1682 ;
    wire signal_1683 ;
    wire signal_1684 ;
    wire signal_1685 ;
    wire signal_1686 ;
    wire signal_1687 ;
    wire signal_1688 ;
    wire signal_1689 ;
    wire signal_1690 ;
    wire signal_1691 ;
    wire signal_1692 ;
    wire signal_1693 ;
    wire signal_1694 ;
    wire signal_1695 ;
    wire signal_1696 ;
    wire signal_1697 ;
    wire signal_1698 ;
    wire signal_1699 ;
    wire signal_1700 ;
    wire signal_1701 ;
    wire signal_1702 ;
    wire signal_1703 ;
    wire signal_1704 ;
    wire signal_1705 ;
    wire signal_1706 ;
    wire signal_1707 ;
    wire signal_1708 ;
    wire signal_1709 ;
    wire signal_1710 ;
    wire signal_1711 ;
    wire signal_1712 ;
    wire signal_1713 ;
    wire signal_1714 ;
    wire signal_1715 ;
    wire signal_1716 ;
    wire signal_1717 ;
    wire signal_1718 ;
    wire signal_1719 ;
    wire signal_1720 ;
    wire signal_1721 ;
    wire signal_1722 ;
    wire signal_1723 ;
    wire signal_1724 ;
    wire signal_1725 ;
    wire signal_1726 ;
    wire signal_1727 ;
    wire signal_1728 ;
    wire signal_1729 ;
    wire signal_1730 ;
    wire signal_1731 ;
    wire signal_1732 ;
    wire signal_1733 ;
    wire signal_1734 ;
    wire signal_1735 ;
    wire signal_1736 ;
    wire signal_1737 ;
    wire signal_1738 ;
    wire signal_1739 ;
    wire signal_1740 ;
    wire signal_1741 ;
    wire signal_1742 ;
    wire signal_1743 ;
    wire signal_1744 ;
    wire signal_1745 ;
    wire signal_1746 ;
    wire signal_1747 ;
    wire signal_1748 ;
    wire signal_1749 ;
    wire signal_1750 ;
    wire signal_1751 ;
    wire signal_1752 ;
    wire signal_1753 ;
    wire signal_1754 ;
    wire signal_1755 ;
    wire signal_1756 ;
    wire signal_1757 ;
    wire signal_1758 ;
    wire signal_1759 ;
    wire signal_1760 ;
    wire signal_1761 ;
    wire signal_1762 ;
    wire signal_1763 ;
    wire signal_1764 ;
    wire signal_1765 ;
    wire signal_1766 ;
    wire signal_1767 ;
    wire signal_1768 ;
    wire signal_1769 ;
    wire signal_1770 ;
    wire signal_1771 ;
    wire signal_1772 ;
    wire signal_1773 ;
    wire signal_1774 ;
    wire signal_1775 ;
    wire signal_1776 ;
    wire signal_1777 ;
    wire signal_1778 ;
    wire signal_1779 ;
    wire signal_1780 ;
    wire signal_1781 ;
    wire signal_1782 ;
    wire signal_1783 ;
    wire signal_1784 ;
    wire signal_1785 ;
    wire signal_1786 ;
    wire signal_1787 ;
    wire signal_1788 ;
    wire signal_1789 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1792 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1795 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1813 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1844 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1854 ;
    wire signal_1855 ;
    wire signal_1856 ;
    wire signal_1857 ;
    wire signal_1858 ;
    wire signal_1859 ;
    wire signal_1860 ;
    wire signal_1861 ;
    wire signal_1862 ;
    wire signal_1863 ;
    wire signal_1864 ;
    wire signal_1865 ;
    wire signal_1866 ;
    wire signal_1867 ;
    wire signal_1868 ;
    wire signal_1869 ;
    wire signal_1870 ;
    wire signal_1871 ;
    wire signal_1872 ;
    wire signal_1873 ;
    wire signal_1874 ;
    wire signal_1875 ;
    wire signal_1876 ;
    wire signal_1877 ;
    wire signal_1878 ;
    wire signal_1879 ;
    wire signal_1880 ;
    wire signal_1881 ;
    wire signal_1882 ;
    wire signal_1883 ;
    wire signal_1884 ;
    wire signal_1885 ;
    wire signal_1886 ;
    wire signal_1887 ;
    wire signal_1888 ;
    wire signal_1889 ;
    wire signal_1890 ;
    wire signal_1891 ;
    wire signal_1892 ;
    wire signal_1893 ;
    wire signal_1894 ;
    wire signal_1895 ;
    wire signal_1896 ;
    wire signal_1897 ;
    wire signal_1898 ;
    wire signal_1899 ;
    wire signal_1900 ;
    wire signal_1901 ;
    wire signal_1902 ;
    wire signal_1903 ;
    wire signal_1904 ;
    wire signal_1905 ;
    wire signal_1906 ;
    wire signal_1907 ;
    wire signal_1908 ;
    wire signal_1909 ;
    wire signal_1910 ;
    wire signal_1911 ;
    wire signal_1912 ;
    wire signal_1913 ;
    wire signal_1914 ;
    wire signal_1915 ;
    wire signal_1916 ;
    wire signal_1917 ;
    wire signal_1918 ;
    wire signal_1919 ;
    wire signal_1920 ;
    wire signal_1921 ;
    wire signal_1922 ;
    wire signal_1923 ;
    wire signal_1924 ;
    wire signal_1925 ;
    wire signal_1926 ;
    wire signal_1927 ;
    wire signal_1928 ;
    wire signal_1929 ;
    wire signal_1930 ;
    wire signal_1931 ;
    wire signal_1932 ;
    wire signal_1933 ;
    wire signal_1934 ;
    wire signal_1935 ;
    wire signal_1936 ;
    wire signal_1937 ;
    wire signal_1938 ;
    wire signal_1939 ;
    wire signal_1940 ;
    wire signal_1941 ;
    wire signal_1942 ;
    wire signal_1943 ;
    wire signal_1945 ;
    wire signal_1946 ;
    wire signal_1947 ;
    wire signal_1949 ;
    wire signal_1950 ;
    wire signal_1951 ;
    wire signal_1952 ;
    wire signal_1953 ;
    wire signal_1954 ;
    wire signal_1955 ;
    wire signal_1956 ;
    wire signal_1957 ;
    wire signal_1958 ;
    wire signal_1959 ;
    wire signal_1961 ;
    wire signal_1962 ;
    wire signal_1963 ;
    wire signal_1964 ;
    wire signal_1965 ;
    wire signal_1966 ;
    wire signal_1967 ;
    wire signal_1968 ;
    wire signal_1969 ;
    wire signal_1970 ;
    wire signal_1971 ;
    wire signal_1973 ;
    wire signal_1974 ;
    wire signal_1975 ;
    wire signal_1976 ;
    wire signal_1977 ;
    wire signal_1978 ;
    wire signal_1979 ;
    wire signal_1980 ;
    wire signal_1981 ;
    wire signal_1982 ;
    wire signal_1983 ;
    wire signal_1984 ;
    wire signal_1985 ;
    wire signal_1986 ;
    wire signal_1987 ;
    wire signal_1988 ;
    wire signal_1989 ;
    wire signal_1990 ;
    wire signal_1991 ;
    wire signal_1992 ;
    wire signal_1993 ;
    wire signal_1994 ;
    wire signal_1995 ;
    wire signal_1996 ;
    wire signal_1997 ;
    wire signal_1998 ;
    wire signal_1999 ;
    wire signal_2000 ;
    wire signal_2001 ;
    wire signal_2002 ;
    wire signal_2003 ;
    wire signal_2004 ;
    wire signal_2005 ;
    wire signal_2006 ;
    wire signal_2007 ;
    wire signal_2008 ;
    wire signal_2009 ;
    wire signal_2010 ;
    wire signal_2011 ;
    wire signal_2012 ;
    wire signal_2013 ;
    wire signal_2014 ;
    wire signal_2015 ;
    wire signal_2016 ;
    wire signal_2017 ;
    wire signal_2018 ;
    wire signal_2019 ;
    wire signal_2020 ;
    wire signal_2021 ;
    wire signal_2022 ;
    wire signal_2023 ;
    wire signal_2024 ;
    wire signal_2025 ;
    wire signal_2026 ;
    wire signal_2027 ;
    wire signal_2028 ;
    wire signal_2029 ;
    wire signal_2030 ;
    wire signal_2031 ;
    wire signal_2032 ;
    wire signal_2033 ;
    wire signal_2034 ;
    wire signal_2035 ;
    wire signal_2036 ;
    wire signal_2037 ;
    wire signal_2038 ;
    wire signal_2039 ;
    wire signal_2040 ;
    wire signal_2041 ;
    wire signal_2042 ;
    wire signal_2043 ;
    wire signal_2044 ;
    wire signal_2045 ;
    wire signal_2046 ;
    wire signal_2047 ;
    wire signal_2048 ;
    wire signal_2049 ;
    wire signal_2050 ;
    wire signal_2051 ;
    wire signal_2052 ;
    wire signal_2053 ;
    wire signal_2054 ;
    wire signal_2055 ;
    wire signal_2056 ;
    wire signal_2057 ;
    wire signal_2058 ;
    wire signal_2059 ;
    wire signal_2060 ;
    wire signal_2061 ;
    wire signal_2062 ;
    wire signal_2063 ;
    wire signal_2064 ;
    wire signal_2065 ;
    wire signal_2066 ;
    wire signal_2067 ;
    wire signal_2068 ;
    wire signal_2069 ;
    wire signal_2070 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2079 ;
    wire signal_2080 ;
    wire signal_2081 ;
    wire signal_2082 ;
    wire signal_2083 ;
    wire signal_2084 ;
    wire signal_2085 ;
    wire signal_2086 ;
    wire signal_2087 ;
    wire signal_2088 ;
    wire signal_2089 ;
    wire signal_2090 ;
    wire signal_2091 ;
    wire signal_2092 ;
    wire signal_2093 ;
    wire signal_2094 ;
    wire signal_2095 ;
    wire signal_2096 ;
    wire signal_2097 ;
    wire signal_2098 ;
    wire signal_2099 ;
    wire signal_2100 ;
    wire signal_2101 ;
    wire signal_2102 ;
    wire signal_2103 ;
    wire signal_2104 ;
    wire signal_2105 ;
    wire signal_2107 ;
    wire signal_2108 ;
    wire signal_2110 ;
    wire signal_2111 ;
    wire signal_2113 ;
    wire signal_2114 ;
    wire signal_2116 ;
    wire signal_2117 ;
    wire signal_2119 ;
    wire signal_2120 ;
    wire signal_2122 ;
    wire signal_2123 ;
    wire signal_2125 ;
    wire signal_2126 ;
    wire signal_2128 ;
    wire signal_2129 ;
    wire signal_2130 ;
    wire signal_2131 ;
    wire signal_2132 ;
    wire signal_2133 ;
    wire signal_2134 ;
    wire signal_2135 ;
    wire signal_2136 ;
    wire signal_2137 ;
    wire signal_2138 ;
    wire signal_2139 ;
    wire signal_2140 ;
    wire signal_2141 ;
    wire signal_2142 ;
    wire signal_2143 ;
    wire signal_2144 ;
    wire signal_2145 ;
    wire signal_2148 ;
    wire signal_2151 ;
    wire signal_2154 ;
    wire signal_2157 ;
    wire signal_2160 ;
    wire signal_2163 ;
    wire signal_2166 ;
    wire signal_2169 ;
    wire signal_2170 ;
    wire signal_2171 ;
    wire signal_2172 ;
    wire signal_2175 ;
    wire signal_2177 ;
    wire signal_2179 ;
    wire signal_2182 ;
    wire signal_2184 ;
    wire signal_2186 ;
    wire signal_2187 ;
    wire signal_2188 ;
    wire signal_2189 ;
    wire signal_2190 ;
    wire signal_2191 ;
    wire signal_2192 ;
    wire signal_2193 ;
    wire signal_2194 ;
    wire signal_2195 ;
    wire signal_2196 ;
    wire signal_2197 ;
    wire signal_2198 ;
    wire signal_2199 ;
    wire signal_2200 ;
    wire signal_2201 ;
    wire signal_2202 ;
    wire signal_2203 ;
    wire signal_2204 ;
    wire signal_2205 ;
    wire signal_2206 ;
    wire signal_2207 ;
    wire signal_2208 ;
    wire signal_2209 ;
    wire signal_2210 ;
    wire signal_2211 ;
    wire signal_2212 ;
    wire signal_2213 ;
    wire signal_2214 ;
    wire signal_2215 ;
    wire signal_2216 ;
    wire signal_2217 ;
    wire signal_2218 ;
    wire signal_2219 ;
    wire signal_2220 ;
    wire signal_2221 ;
    wire signal_2222 ;
    wire signal_2223 ;
    wire signal_2224 ;
    wire signal_2225 ;
    wire signal_2226 ;
    wire signal_2227 ;
    wire signal_2228 ;
    wire signal_2229 ;
    wire signal_2230 ;
    wire signal_2231 ;
    wire signal_2232 ;
    wire signal_2233 ;
    wire signal_2234 ;
    wire signal_2235 ;
    wire signal_2236 ;
    wire signal_2237 ;
    wire signal_2238 ;
    wire signal_2239 ;
    wire signal_2240 ;
    wire signal_2241 ;
    wire signal_2242 ;
    wire signal_2243 ;
    wire signal_2244 ;
    wire signal_2245 ;
    wire signal_2246 ;
    wire signal_2247 ;
    wire signal_2248 ;
    wire signal_2249 ;
    wire signal_2250 ;
    wire signal_2251 ;
    wire signal_2252 ;
    wire signal_2253 ;
    wire signal_2254 ;
    wire signal_2255 ;
    wire signal_2256 ;
    wire signal_2257 ;
    wire signal_2258 ;
    wire signal_2259 ;
    wire signal_2260 ;
    wire signal_2261 ;
    wire signal_2262 ;
    wire signal_2263 ;
    wire signal_2264 ;
    wire signal_2265 ;
    wire signal_2266 ;
    wire signal_2267 ;
    wire signal_2268 ;
    wire signal_2269 ;
    wire signal_2270 ;
    wire signal_2271 ;
    wire signal_2272 ;
    wire signal_2273 ;
    wire signal_2274 ;
    wire signal_2275 ;
    wire signal_2276 ;
    wire signal_2277 ;
    wire signal_2280 ;
    wire signal_2283 ;
    wire signal_2286 ;
    wire signal_2289 ;
    wire signal_2292 ;
    wire signal_2295 ;
    wire signal_2298 ;
    wire signal_2301 ;
    wire signal_2304 ;
    wire signal_2307 ;
    wire signal_2310 ;
    wire signal_2313 ;
    wire signal_2316 ;
    wire signal_2319 ;
    wire signal_2322 ;
    wire signal_2325 ;
    wire signal_2328 ;
    wire signal_2331 ;
    wire signal_2334 ;
    wire signal_2337 ;
    wire signal_2340 ;
    wire signal_2343 ;
    wire signal_2346 ;
    wire signal_2349 ;
    wire signal_2352 ;
    wire signal_2355 ;
    wire signal_2358 ;
    wire signal_2361 ;
    wire signal_2364 ;
    wire signal_2367 ;
    wire signal_2370 ;
    wire signal_2373 ;
    wire signal_2376 ;
    wire signal_2379 ;
    wire signal_2382 ;
    wire signal_2385 ;
    wire signal_2388 ;
    wire signal_2391 ;
    wire signal_2394 ;
    wire signal_2397 ;
    wire signal_2400 ;
    wire signal_2403 ;
    wire signal_2406 ;
    wire signal_2409 ;
    wire signal_2412 ;
    wire signal_2415 ;
    wire signal_2418 ;
    wire signal_2421 ;
    wire signal_2424 ;
    wire signal_2427 ;
    wire signal_2430 ;
    wire signal_2433 ;
    wire signal_2436 ;
    wire signal_2439 ;
    wire signal_2442 ;
    wire signal_2445 ;
    wire signal_2448 ;
    wire signal_2451 ;
    wire signal_2454 ;
    wire signal_2457 ;
    wire signal_2460 ;
    wire signal_2463 ;
    wire signal_2466 ;
    wire signal_2469 ;
    wire signal_2472 ;
    wire signal_2475 ;
    wire signal_2478 ;
    wire signal_2481 ;
    wire signal_2484 ;
    wire signal_2487 ;
    wire signal_2490 ;
    wire signal_2493 ;
    wire signal_2496 ;
    wire signal_2499 ;
    wire signal_2502 ;
    wire signal_2505 ;
    wire signal_2508 ;
    wire signal_2511 ;
    wire signal_2514 ;
    wire signal_2517 ;
    wire signal_2520 ;
    wire signal_2523 ;
    wire signal_2526 ;
    wire signal_2529 ;
    wire signal_2532 ;
    wire signal_2535 ;
    wire signal_2538 ;
    wire signal_2541 ;
    wire signal_2544 ;
    wire signal_2547 ;
    wire signal_2550 ;
    wire signal_2553 ;
    wire signal_2556 ;
    wire signal_2559 ;
    wire signal_2562 ;
    wire signal_2565 ;
    wire signal_2567 ;
    wire signal_2568 ;
    wire signal_2570 ;
    wire signal_2571 ;
    wire signal_2573 ;
    wire signal_2574 ;
    wire signal_2576 ;
    wire signal_2577 ;
    wire signal_2579 ;
    wire signal_2580 ;
    wire signal_2582 ;
    wire signal_2583 ;
    wire signal_2585 ;
    wire signal_2586 ;
    wire signal_2588 ;
    wire signal_2589 ;
    wire signal_2591 ;
    wire signal_2592 ;
    wire signal_2594 ;
    wire signal_2595 ;
    wire signal_2597 ;
    wire signal_2598 ;
    wire signal_2600 ;
    wire signal_2601 ;
    wire signal_2603 ;
    wire signal_2604 ;
    wire signal_2606 ;
    wire signal_2607 ;
    wire signal_2609 ;
    wire signal_2610 ;
    wire signal_2612 ;
    wire signal_2613 ;
    wire signal_2615 ;
    wire signal_2616 ;
    wire signal_2618 ;
    wire signal_2619 ;
    wire signal_2621 ;
    wire signal_2622 ;
    wire signal_2624 ;
    wire signal_2625 ;
    wire signal_2627 ;
    wire signal_2628 ;
    wire signal_2630 ;
    wire signal_2631 ;
    wire signal_2633 ;
    wire signal_2634 ;
    wire signal_2636 ;
    wire signal_2637 ;
    wire signal_2639 ;
    wire signal_2640 ;
    wire signal_2642 ;
    wire signal_2643 ;
    wire signal_2645 ;
    wire signal_2646 ;
    wire signal_2648 ;
    wire signal_2649 ;
    wire signal_2651 ;
    wire signal_2652 ;
    wire signal_2654 ;
    wire signal_2655 ;
    wire signal_2657 ;
    wire signal_2658 ;
    wire signal_2660 ;
    wire signal_2661 ;
    wire signal_2663 ;
    wire signal_2664 ;
    wire signal_2666 ;
    wire signal_2667 ;
    wire signal_2669 ;
    wire signal_2670 ;
    wire signal_2672 ;
    wire signal_2673 ;
    wire signal_2675 ;
    wire signal_2676 ;
    wire signal_2678 ;
    wire signal_2679 ;
    wire signal_2681 ;
    wire signal_2682 ;
    wire signal_2684 ;
    wire signal_2685 ;
    wire signal_2687 ;
    wire signal_2688 ;
    wire signal_2690 ;
    wire signal_2691 ;
    wire signal_2693 ;
    wire signal_2694 ;
    wire signal_2696 ;
    wire signal_2697 ;
    wire signal_2699 ;
    wire signal_2700 ;
    wire signal_2702 ;
    wire signal_2703 ;
    wire signal_2705 ;
    wire signal_2706 ;
    wire signal_2708 ;
    wire signal_2709 ;
    wire signal_2711 ;
    wire signal_2712 ;
    wire signal_2714 ;
    wire signal_2715 ;
    wire signal_2717 ;
    wire signal_2718 ;
    wire signal_2720 ;
    wire signal_2721 ;
    wire signal_2723 ;
    wire signal_2724 ;
    wire signal_2726 ;
    wire signal_2727 ;
    wire signal_2729 ;
    wire signal_2730 ;
    wire signal_2732 ;
    wire signal_2733 ;
    wire signal_2735 ;
    wire signal_2736 ;
    wire signal_2738 ;
    wire signal_2739 ;
    wire signal_2741 ;
    wire signal_2742 ;
    wire signal_2744 ;
    wire signal_2745 ;
    wire signal_2747 ;
    wire signal_2748 ;
    wire signal_2750 ;
    wire signal_2751 ;
    wire signal_2753 ;
    wire signal_2754 ;
    wire signal_2756 ;
    wire signal_2757 ;
    wire signal_2759 ;
    wire signal_2760 ;
    wire signal_2762 ;
    wire signal_2763 ;
    wire signal_2765 ;
    wire signal_2766 ;
    wire signal_2768 ;
    wire signal_2769 ;
    wire signal_2771 ;
    wire signal_2772 ;
    wire signal_2774 ;
    wire signal_2775 ;
    wire signal_2777 ;
    wire signal_2778 ;
    wire signal_2780 ;
    wire signal_2781 ;
    wire signal_2783 ;
    wire signal_2784 ;
    wire signal_2786 ;
    wire signal_2787 ;
    wire signal_2789 ;
    wire signal_2790 ;
    wire signal_2792 ;
    wire signal_2793 ;
    wire signal_2795 ;
    wire signal_2796 ;
    wire signal_2798 ;
    wire signal_2799 ;
    wire signal_2801 ;
    wire signal_2802 ;
    wire signal_2804 ;
    wire signal_2805 ;
    wire signal_2807 ;
    wire signal_2808 ;
    wire signal_2810 ;
    wire signal_2811 ;
    wire signal_2813 ;
    wire signal_2814 ;
    wire signal_2816 ;
    wire signal_2817 ;
    wire signal_2819 ;
    wire signal_2820 ;
    wire signal_2822 ;
    wire signal_2823 ;
    wire signal_2825 ;
    wire signal_2826 ;
    wire signal_2828 ;
    wire signal_2829 ;
    wire signal_2831 ;
    wire signal_2832 ;
    wire signal_2834 ;
    wire signal_2835 ;
    wire signal_2837 ;
    wire signal_2838 ;
    wire signal_2840 ;
    wire signal_2841 ;
    wire signal_2843 ;
    wire signal_2844 ;
    wire signal_2846 ;
    wire signal_2847 ;
    wire signal_2849 ;
    wire signal_2850 ;
    wire signal_2852 ;
    wire signal_2853 ;
    wire signal_2855 ;
    wire signal_2856 ;
    wire signal_2858 ;
    wire signal_2859 ;
    wire signal_2861 ;
    wire signal_2862 ;
    wire signal_2864 ;
    wire signal_2865 ;
    wire signal_2867 ;
    wire signal_2868 ;
    wire signal_2870 ;
    wire signal_2871 ;
    wire signal_2873 ;
    wire signal_2874 ;
    wire signal_2876 ;
    wire signal_2877 ;
    wire signal_2879 ;
    wire signal_2880 ;
    wire signal_2882 ;
    wire signal_2883 ;
    wire signal_2885 ;
    wire signal_2886 ;
    wire signal_2888 ;
    wire signal_2889 ;
    wire signal_2891 ;
    wire signal_2892 ;
    wire signal_2894 ;
    wire signal_2895 ;
    wire signal_2897 ;
    wire signal_2898 ;
    wire signal_2900 ;
    wire signal_2901 ;
    wire signal_2903 ;
    wire signal_2905 ;
    wire signal_2907 ;
    wire signal_2909 ;
    wire signal_2911 ;
    wire signal_2913 ;
    wire signal_2915 ;
    wire signal_2917 ;
    wire signal_2918 ;
    wire signal_2919 ;
    wire signal_2920 ;
    wire signal_2921 ;
    wire signal_2922 ;
    wire signal_2923 ;
    wire signal_2924 ;
    wire signal_2925 ;
    wire signal_2926 ;
    wire signal_2927 ;
    wire signal_2928 ;
    wire signal_2929 ;
    wire signal_2930 ;
    wire signal_2931 ;
    wire signal_2932 ;
    wire signal_2933 ;
    wire signal_2934 ;
    wire signal_2935 ;
    wire signal_2936 ;
    wire signal_2937 ;
    wire signal_2938 ;
    wire signal_2939 ;
    wire signal_2940 ;
    wire signal_2941 ;
    wire signal_2942 ;
    wire signal_2943 ;
    wire signal_2944 ;
    wire signal_2945 ;
    wire signal_2946 ;
    wire signal_2947 ;
    wire signal_2948 ;
    wire signal_2949 ;
    wire signal_2950 ;
    wire signal_2951 ;
    wire signal_2952 ;
    wire signal_2953 ;
    wire signal_2954 ;
    wire signal_2955 ;
    wire signal_2956 ;
    wire signal_2957 ;
    wire signal_2958 ;
    wire signal_2959 ;
    wire signal_2960 ;
    wire signal_2961 ;
    wire signal_2962 ;
    wire signal_2963 ;
    wire signal_2964 ;
    wire signal_2965 ;
    wire signal_2966 ;
    wire signal_2967 ;
    wire signal_2968 ;
    wire signal_2969 ;
    wire signal_2970 ;
    wire signal_2971 ;
    wire signal_2972 ;
    wire signal_2973 ;
    wire signal_2974 ;
    wire signal_2975 ;
    wire signal_2976 ;
    wire signal_2977 ;
    wire signal_2978 ;
    wire signal_2979 ;
    wire signal_2980 ;
    wire signal_2981 ;
    wire signal_2982 ;
    wire signal_2983 ;
    wire signal_2984 ;
    wire signal_2985 ;
    wire signal_2986 ;
    wire signal_2987 ;
    wire signal_2988 ;
    wire signal_2989 ;
    wire signal_2990 ;
    wire signal_2991 ;
    wire signal_2992 ;
    wire signal_2993 ;
    wire signal_2994 ;
    wire signal_2995 ;
    wire signal_2996 ;
    wire signal_2997 ;
    wire signal_2998 ;
    wire signal_2999 ;
    wire signal_3000 ;
    wire signal_3001 ;
    wire signal_3002 ;
    wire signal_3003 ;
    wire signal_3004 ;
    wire signal_3005 ;
    wire signal_3006 ;
    wire signal_3007 ;
    wire signal_3008 ;
    wire signal_3009 ;
    wire signal_3010 ;
    wire signal_3011 ;
    wire signal_3012 ;
    wire signal_3013 ;
    wire signal_3014 ;
    wire signal_3015 ;
    wire signal_3016 ;
    wire signal_3017 ;
    wire signal_3018 ;
    wire signal_3019 ;
    wire signal_3020 ;
    wire signal_3021 ;
    wire signal_3022 ;
    wire signal_3023 ;
    wire signal_3024 ;
    wire signal_3025 ;
    wire signal_3026 ;
    wire signal_3027 ;
    wire signal_3028 ;
    wire signal_3029 ;
    wire signal_3030 ;
    wire signal_3031 ;
    wire signal_3032 ;
    wire signal_3033 ;
    wire signal_3034 ;
    wire signal_3035 ;
    wire signal_3036 ;
    wire signal_3037 ;
    wire signal_3038 ;
    wire signal_3039 ;
    wire signal_3040 ;
    wire signal_3041 ;
    wire signal_3042 ;
    wire signal_3043 ;
    wire signal_3044 ;
    wire signal_3045 ;
    wire signal_3046 ;
    wire signal_3047 ;
    wire signal_3048 ;
    wire signal_3049 ;
    wire signal_3050 ;
    wire signal_3051 ;
    wire signal_3052 ;
    wire signal_3053 ;
    wire signal_3054 ;
    wire signal_3055 ;
    wire signal_3056 ;
    wire signal_3057 ;
    wire signal_3058 ;
    wire signal_3059 ;
    wire signal_3060 ;
    wire signal_3061 ;
    wire signal_3062 ;
    wire signal_3063 ;
    wire signal_3064 ;
    wire signal_3065 ;
    wire signal_3066 ;
    wire signal_3067 ;
    wire signal_3068 ;
    wire signal_3069 ;
    wire signal_3070 ;
    wire signal_3071 ;
    wire signal_3072 ;
    wire signal_3073 ;
    wire signal_3074 ;
    wire signal_3075 ;
    wire signal_3076 ;
    wire signal_3077 ;
    wire signal_3078 ;
    wire signal_3079 ;
    wire signal_3080 ;
    wire signal_3081 ;
    wire signal_3082 ;
    wire signal_3083 ;
    wire signal_3084 ;
    wire signal_3085 ;
    wire signal_3086 ;
    wire signal_3087 ;
    wire signal_3088 ;
    wire signal_3089 ;
    wire signal_3090 ;
    wire signal_3091 ;
    wire signal_3092 ;
    wire signal_3093 ;
    wire signal_3094 ;
    wire signal_3095 ;
    wire signal_3096 ;
    wire signal_3097 ;
    wire signal_3098 ;
    wire signal_3099 ;
    wire signal_3100 ;
    wire signal_3101 ;
    wire signal_3102 ;
    wire signal_3103 ;
    wire signal_3104 ;
    wire signal_3105 ;
    wire signal_3106 ;
    wire signal_3107 ;
    wire signal_3108 ;
    wire signal_3109 ;
    wire signal_3110 ;
    wire signal_3111 ;
    wire signal_3112 ;
    wire signal_3113 ;
    wire signal_3114 ;
    wire signal_3115 ;
    wire signal_3116 ;
    wire signal_3117 ;
    wire signal_3118 ;
    wire signal_3119 ;
    wire signal_3120 ;
    wire signal_3121 ;
    wire signal_3122 ;
    wire signal_3123 ;
    wire signal_3124 ;
    wire signal_3125 ;
    wire signal_3126 ;
    wire signal_3127 ;
    wire signal_3128 ;
    wire signal_3129 ;
    wire signal_3130 ;
    wire signal_3131 ;
    wire signal_3132 ;
    wire signal_3133 ;
    wire signal_3134 ;
    wire signal_3135 ;
    wire signal_3136 ;
    wire signal_3137 ;
    wire signal_3138 ;
    wire signal_3139 ;
    wire signal_3140 ;
    wire signal_3141 ;
    wire signal_3142 ;
    wire signal_3143 ;
    wire signal_3144 ;
    wire signal_3145 ;
    wire signal_3146 ;
    wire signal_3147 ;
    wire signal_3148 ;
    wire signal_3149 ;
    wire signal_3150 ;
    wire signal_3151 ;
    wire signal_3152 ;
    wire signal_3153 ;
    wire signal_3154 ;
    wire signal_3155 ;
    wire signal_3156 ;
    wire signal_3157 ;
    wire signal_3158 ;
    wire signal_3159 ;
    wire signal_3160 ;
    wire signal_3161 ;
    wire signal_3162 ;
    wire signal_3163 ;
    wire signal_3164 ;
    wire signal_3165 ;
    wire signal_3166 ;
    wire signal_3167 ;
    wire signal_3168 ;
    wire signal_3170 ;
    wire signal_3172 ;
    wire signal_3174 ;
    wire signal_3176 ;
    wire signal_3178 ;
    wire signal_3180 ;
    wire signal_3182 ;
    wire signal_3184 ;
    wire signal_3186 ;
    wire signal_3188 ;
    wire signal_3190 ;
    wire signal_3192 ;
    wire signal_3194 ;
    wire signal_3196 ;
    wire signal_3198 ;
    wire signal_3200 ;
    wire signal_3202 ;
    wire signal_3204 ;
    wire signal_3206 ;
    wire signal_3208 ;
    wire signal_3210 ;
    wire signal_3212 ;
    wire signal_3214 ;
    wire signal_3216 ;
    wire signal_3217 ;
    wire signal_3218 ;
    wire signal_3219 ;
    wire signal_3220 ;
    wire signal_3221 ;
    wire signal_3222 ;
    wire signal_3223 ;
    wire signal_3224 ;
    wire signal_3225 ;
    wire signal_3226 ;
    wire signal_3227 ;
    wire signal_3228 ;
    wire signal_3229 ;
    wire signal_3230 ;
    wire signal_3231 ;
    wire signal_3232 ;
    wire signal_3233 ;
    wire signal_3234 ;
    wire signal_3235 ;
    wire signal_3236 ;
    wire signal_3237 ;
    wire signal_3238 ;
    wire signal_3239 ;
    wire signal_3240 ;
    wire signal_3241 ;
    wire signal_3242 ;
    wire signal_3243 ;
    wire signal_3244 ;
    wire signal_3245 ;
    wire signal_3246 ;
    wire signal_3247 ;
    wire signal_3248 ;
    wire signal_3249 ;
    wire signal_3250 ;
    wire signal_3251 ;
    wire signal_3252 ;
    wire signal_3253 ;
    wire signal_3254 ;
    wire signal_3255 ;
    wire signal_3256 ;
    wire signal_3257 ;
    wire signal_3258 ;
    wire signal_3259 ;
    wire signal_3260 ;
    wire signal_3261 ;
    wire signal_3262 ;
    wire signal_3263 ;
    wire signal_3264 ;
    wire signal_3265 ;
    wire signal_3266 ;
    wire signal_3267 ;
    wire signal_3268 ;
    wire signal_3269 ;
    wire signal_3270 ;
    wire signal_3271 ;
    wire signal_3272 ;
    wire signal_3273 ;
    wire signal_3274 ;
    wire signal_3275 ;
    wire signal_3276 ;
    wire signal_3277 ;
    wire signal_3278 ;
    wire signal_3279 ;
    wire signal_3280 ;
    wire signal_3281 ;
    wire signal_3282 ;
    wire signal_3283 ;
    wire signal_3284 ;
    wire signal_3285 ;
    wire signal_3286 ;
    wire signal_3287 ;
    wire signal_3288 ;
    wire signal_3289 ;
    wire signal_3290 ;
    wire signal_3291 ;
    wire signal_3292 ;
    wire signal_3293 ;
    wire signal_3294 ;
    wire signal_3295 ;
    wire signal_3296 ;
    wire signal_3297 ;
    wire signal_3298 ;
    wire signal_3299 ;
    wire signal_3300 ;
    wire signal_3301 ;
    wire signal_3302 ;
    wire signal_3303 ;
    wire signal_3304 ;
    wire signal_3305 ;
    wire signal_3306 ;
    wire signal_3307 ;
    wire signal_3308 ;
    wire signal_3309 ;
    wire signal_3310 ;
    wire signal_3311 ;
    wire signal_3312 ;
    wire signal_3313 ;
    wire signal_3314 ;
    wire signal_3315 ;
    wire signal_3316 ;
    wire signal_3317 ;
    wire signal_3318 ;
    wire signal_3319 ;
    wire signal_3320 ;
    wire signal_3321 ;
    wire signal_3322 ;
    wire signal_3323 ;
    wire signal_3324 ;
    wire signal_3325 ;
    wire signal_3326 ;
    wire signal_3327 ;
    wire signal_3328 ;
    wire signal_3329 ;
    wire signal_3330 ;
    wire signal_3331 ;
    wire signal_3332 ;
    wire signal_3333 ;
    wire signal_3334 ;
    wire signal_3335 ;
    wire signal_3336 ;
    wire signal_3337 ;
    wire signal_3338 ;
    wire signal_3339 ;
    wire signal_3340 ;
    wire signal_3341 ;
    wire signal_3342 ;
    wire signal_3343 ;
    wire signal_3344 ;
    wire signal_3345 ;
    wire signal_3346 ;
    wire signal_3347 ;
    wire signal_3348 ;
    wire signal_3349 ;
    wire signal_3350 ;
    wire signal_3351 ;
    wire signal_3352 ;
    wire signal_3353 ;
    wire signal_3354 ;
    wire signal_3355 ;
    wire signal_3356 ;
    wire signal_3357 ;
    wire signal_3358 ;
    wire signal_3359 ;
    wire signal_3360 ;
    wire signal_3361 ;
    wire signal_3362 ;
    wire signal_3363 ;
    wire signal_3364 ;
    wire signal_3365 ;
    wire signal_3366 ;
    wire signal_3367 ;
    wire signal_3368 ;
    wire signal_3369 ;
    wire signal_3371 ;
    wire signal_3373 ;
    wire signal_3375 ;
    wire signal_3377 ;
    wire signal_3379 ;
    wire signal_3381 ;
    wire signal_3383 ;
    wire signal_3385 ;
    wire signal_3386 ;
    wire signal_3387 ;
    wire signal_3388 ;
    wire signal_3389 ;
    wire signal_3390 ;
    wire signal_3391 ;
    wire signal_3392 ;
    wire signal_3393 ;
    wire signal_3394 ;
    wire signal_3395 ;
    wire signal_3396 ;
    wire signal_3397 ;
    wire signal_3398 ;
    wire signal_3399 ;
    wire signal_3400 ;
    wire signal_3401 ;
    wire signal_3402 ;
    wire signal_3403 ;
    wire signal_3404 ;
    wire signal_3405 ;
    wire signal_3406 ;
    wire signal_3407 ;
    wire signal_3408 ;
    wire signal_3409 ;
    wire signal_3410 ;
    wire signal_3411 ;
    wire signal_3412 ;
    wire signal_3413 ;
    wire signal_3414 ;
    wire signal_3415 ;
    wire signal_3416 ;
    wire signal_3417 ;
    wire signal_3418 ;
    wire signal_3419 ;
    wire signal_3420 ;
    wire signal_3421 ;
    wire signal_3422 ;
    wire signal_3423 ;
    wire signal_3424 ;
    wire signal_3425 ;
    wire signal_3426 ;
    wire signal_3427 ;
    wire signal_3428 ;
    wire signal_3429 ;
    wire signal_3430 ;
    wire signal_3431 ;
    wire signal_3432 ;
    wire signal_3433 ;
    wire signal_3434 ;
    wire signal_3435 ;
    wire signal_3436 ;
    wire signal_3437 ;
    wire signal_3438 ;
    wire signal_3439 ;
    wire signal_3440 ;
    wire signal_3441 ;
    wire signal_3442 ;
    wire signal_3443 ;
    wire signal_3444 ;
    wire signal_3445 ;
    wire signal_3446 ;
    wire signal_3447 ;
    wire signal_3448 ;
    wire signal_3449 ;
    wire signal_3450 ;
    wire signal_3451 ;
    wire signal_3452 ;
    wire signal_3453 ;
    wire signal_3454 ;
    wire signal_3455 ;
    wire signal_3456 ;
    wire signal_3457 ;
    wire signal_3458 ;
    wire signal_3459 ;
    wire signal_3460 ;
    wire signal_3461 ;
    wire signal_3462 ;
    wire signal_3463 ;
    wire signal_3464 ;
    wire signal_3465 ;
    wire signal_3466 ;
    wire signal_3467 ;
    wire signal_3468 ;
    wire signal_3469 ;
    wire signal_3470 ;
    wire signal_3471 ;
    wire signal_3472 ;
    wire signal_3473 ;
    wire signal_3474 ;
    wire signal_3475 ;
    wire signal_3476 ;
    wire signal_3477 ;
    wire signal_3478 ;
    wire signal_3479 ;
    wire signal_3480 ;
    wire signal_3481 ;
    wire signal_3482 ;
    wire signal_3483 ;
    wire signal_3484 ;
    wire signal_3485 ;
    wire signal_3486 ;
    wire signal_3487 ;
    wire signal_3488 ;
    wire signal_3489 ;
    wire signal_3490 ;
    wire signal_3491 ;
    wire signal_3492 ;
    wire signal_3493 ;
    wire signal_3494 ;
    wire signal_3495 ;
    wire signal_3496 ;
    wire signal_3497 ;
    wire signal_3498 ;
    wire signal_3499 ;
    wire signal_3500 ;
    wire signal_3501 ;
    wire signal_3502 ;
    wire signal_3503 ;
    wire signal_3504 ;
    wire signal_3505 ;
    wire signal_3506 ;
    wire signal_3507 ;
    wire signal_3508 ;
    wire signal_3509 ;
    wire signal_3510 ;
    wire signal_3511 ;
    wire signal_3512 ;
    wire signal_3513 ;
    wire signal_3514 ;
    wire signal_3515 ;
    wire signal_3516 ;
    wire signal_3517 ;
    wire signal_3518 ;
    wire signal_3519 ;
    wire signal_3520 ;
    wire signal_3521 ;
    wire signal_3522 ;
    wire signal_3523 ;
    wire signal_3524 ;
    wire signal_3525 ;
    wire signal_3526 ;
    wire signal_3527 ;
    wire signal_3528 ;
    wire signal_3529 ;
    wire signal_3530 ;
    wire signal_3531 ;
    wire signal_3532 ;
    wire signal_3533 ;
    wire signal_3534 ;
    wire signal_3535 ;
    wire signal_3536 ;
    wire signal_3537 ;
    wire signal_3538 ;
    wire signal_3539 ;
    wire signal_3540 ;
    wire signal_3541 ;
    wire signal_3542 ;
    wire signal_3543 ;
    wire signal_3544 ;
    wire signal_3545 ;
    wire signal_3546 ;
    wire signal_3547 ;
    wire signal_3548 ;
    wire signal_3549 ;
    wire signal_3550 ;
    wire signal_3551 ;
    wire signal_3552 ;
    wire signal_3553 ;
    wire signal_3554 ;
    wire signal_3555 ;
    wire signal_3556 ;
    wire signal_3557 ;
    wire signal_3558 ;
    wire signal_3559 ;
    wire signal_3560 ;
    wire signal_3561 ;
    wire signal_3562 ;
    wire signal_3563 ;
    wire signal_3564 ;
    wire signal_3565 ;
    wire signal_3566 ;
    wire signal_3567 ;
    wire signal_3568 ;
    wire signal_3569 ;
    wire signal_3570 ;
    wire signal_3571 ;
    wire signal_3572 ;
    wire signal_3573 ;
    wire signal_3574 ;
    wire signal_3575 ;
    wire signal_3576 ;
    wire signal_3577 ;
    wire signal_3578 ;
    wire signal_3579 ;
    wire signal_3580 ;
    wire signal_3581 ;
    wire signal_3582 ;
    wire signal_3583 ;
    wire signal_3584 ;
    wire signal_3585 ;
    wire signal_3586 ;
    wire signal_3587 ;
    wire signal_3588 ;
    wire signal_3589 ;
    wire signal_3590 ;
    wire signal_3591 ;
    wire signal_3592 ;
    wire signal_3593 ;
    wire signal_3594 ;
    wire signal_3595 ;
    wire signal_3596 ;
    wire signal_3597 ;
    wire signal_3598 ;
    wire signal_3599 ;
    wire signal_3600 ;
    wire signal_3601 ;
    wire signal_3602 ;
    wire signal_3603 ;
    wire signal_3604 ;
    wire signal_3605 ;
    wire signal_3606 ;
    wire signal_3607 ;
    wire signal_3608 ;
    wire signal_3609 ;
    wire signal_3610 ;
    wire signal_3611 ;
    wire signal_3612 ;
    wire signal_3613 ;
    wire signal_3614 ;
    wire signal_3615 ;
    wire signal_3616 ;
    wire signal_3617 ;
    wire signal_3618 ;
    wire signal_3620 ;
    wire signal_3622 ;
    wire signal_3624 ;
    wire signal_3626 ;
    wire signal_3628 ;
    wire signal_3629 ;
    wire signal_3630 ;
    wire signal_3631 ;
    wire signal_3632 ;
    wire signal_3633 ;
    wire signal_3634 ;
    wire signal_3635 ;
    wire signal_3636 ;
    wire signal_3637 ;
    wire signal_3638 ;
    wire signal_3639 ;
    wire signal_3640 ;
    wire signal_3641 ;
    wire signal_3643 ;
    wire signal_3645 ;
    wire signal_3647 ;
    wire signal_3648 ;
    wire signal_3649 ;
    wire signal_3650 ;
    wire signal_3651 ;
    wire signal_3652 ;
    wire signal_3653 ;
    wire signal_3654 ;
    wire signal_3655 ;
    wire signal_3656 ;
    wire signal_3657 ;
    wire signal_3658 ;
    wire signal_3659 ;
    wire signal_3660 ;
    wire signal_3661 ;
    wire signal_3696 ;
    wire signal_3697 ;
    wire signal_3698 ;
    wire signal_3699 ;
    wire signal_3700 ;
    wire signal_3701 ;
    wire signal_3702 ;
    wire signal_3703 ;
    wire signal_3704 ;
    wire signal_3705 ;
    wire signal_3706 ;
    wire signal_3707 ;
    wire signal_3708 ;
    wire signal_3709 ;
    wire signal_3710 ;
    wire signal_3711 ;
    wire signal_3712 ;
    wire signal_3713 ;
    wire signal_3714 ;
    wire signal_3715 ;
    wire signal_3716 ;
    wire signal_3717 ;
    wire signal_3718 ;
    wire signal_3719 ;
    wire signal_3720 ;
    wire signal_3721 ;
    wire signal_3722 ;
    wire signal_3723 ;
    wire signal_3724 ;
    wire signal_3725 ;
    wire signal_3726 ;
    wire signal_3727 ;
    wire signal_3728 ;
    wire signal_3729 ;
    wire signal_3730 ;
    wire signal_3731 ;
    wire signal_3732 ;
    wire signal_3733 ;
    wire signal_3734 ;
    wire signal_3735 ;
    wire signal_3736 ;
    wire signal_3737 ;
    wire signal_3738 ;
    wire signal_3739 ;
    wire signal_3740 ;
    wire signal_3741 ;
    wire signal_3742 ;
    wire signal_3743 ;
    wire signal_3744 ;
    wire signal_3745 ;
    wire signal_3746 ;
    wire signal_3747 ;
    wire signal_3748 ;
    wire signal_3749 ;
    wire signal_3750 ;
    wire signal_3751 ;
    wire signal_3752 ;
    wire signal_3753 ;
    wire signal_3754 ;
    wire signal_3755 ;
    wire signal_3756 ;
    wire signal_3757 ;
    wire signal_3758 ;
    wire signal_3759 ;
    wire signal_3760 ;
    wire signal_3761 ;
    wire signal_3762 ;
    wire signal_3763 ;
    wire signal_3764 ;
    wire signal_3765 ;
    wire signal_3766 ;
    wire signal_3767 ;
    wire signal_3768 ;
    wire signal_3769 ;
    wire signal_3770 ;
    wire signal_3771 ;
    wire signal_3772 ;
    wire signal_3773 ;
    wire signal_3774 ;
    wire signal_3775 ;
    wire signal_3776 ;
    wire signal_3777 ;
    wire signal_3778 ;
    wire signal_3779 ;
    wire signal_3780 ;
    wire signal_3781 ;
    wire signal_3782 ;
    wire signal_3783 ;
    wire signal_3784 ;
    wire signal_3785 ;
    wire signal_3786 ;
    wire signal_3787 ;
    wire signal_3788 ;
    wire signal_3789 ;
    wire signal_3790 ;
    wire signal_3791 ;
    wire signal_3792 ;
    wire signal_3793 ;
    wire signal_3794 ;
    wire signal_3795 ;
    wire signal_3796 ;
    wire signal_3797 ;
    wire signal_3798 ;
    wire signal_3799 ;
    wire signal_3800 ;
    wire signal_3801 ;
    wire signal_3802 ;
    wire signal_3803 ;
    wire signal_3804 ;
    wire signal_3805 ;
    wire signal_3806 ;
    wire signal_3807 ;
    wire signal_3808 ;
    wire signal_3809 ;
    wire signal_3810 ;
    wire signal_3811 ;
    wire signal_3812 ;
    wire signal_3813 ;
    wire signal_3814 ;
    wire signal_3815 ;
    wire signal_3816 ;
    wire signal_3817 ;
    wire signal_3818 ;
    wire signal_3819 ;
    wire signal_3820 ;
    wire signal_3821 ;
    wire signal_3822 ;
    wire signal_3823 ;
    wire signal_3824 ;
    wire signal_3825 ;
    wire signal_3826 ;
    wire signal_3827 ;
    wire signal_3828 ;
    wire signal_3829 ;
    wire signal_3830 ;
    wire signal_3831 ;
    wire signal_3832 ;
    wire signal_3833 ;
    wire signal_3834 ;
    wire signal_3835 ;
    wire signal_3836 ;
    wire signal_3837 ;
    wire signal_3838 ;
    wire signal_3839 ;
    wire signal_3840 ;
    wire signal_3841 ;
    wire signal_3842 ;
    wire signal_3843 ;
    wire signal_3844 ;
    wire signal_3845 ;
    wire signal_3846 ;
    wire signal_3847 ;
    wire signal_3848 ;
    wire signal_3849 ;
    wire signal_3850 ;
    wire signal_3851 ;
    wire signal_3852 ;
    wire signal_3853 ;
    wire signal_3854 ;
    wire signal_3855 ;
    wire signal_3856 ;
    wire signal_3857 ;
    wire signal_3858 ;
    wire signal_3859 ;
    wire signal_3860 ;
    wire signal_3861 ;
    wire signal_3862 ;
    wire signal_3863 ;
    wire signal_3864 ;
    wire signal_3865 ;
    wire signal_3866 ;
    wire signal_3867 ;
    wire signal_3868 ;
    wire signal_3869 ;
    wire signal_3870 ;
    wire signal_3871 ;
    wire signal_3872 ;
    wire signal_3873 ;
    wire signal_3874 ;
    wire signal_3875 ;
    wire signal_3876 ;
    wire signal_3877 ;
    wire signal_3878 ;
    wire signal_3879 ;
    wire signal_3880 ;
    wire signal_3881 ;
    wire signal_3882 ;
    wire signal_3883 ;
    wire signal_3884 ;
    wire signal_3885 ;
    wire signal_3886 ;
    wire signal_3887 ;
    wire signal_3888 ;
    wire signal_3889 ;
    wire signal_3890 ;
    wire signal_3891 ;
    wire signal_3892 ;
    wire signal_3893 ;
    wire signal_3894 ;
    wire signal_3895 ;
    wire signal_3896 ;
    wire signal_3897 ;
    wire signal_3898 ;
    wire signal_3899 ;
    wire signal_3900 ;
    wire signal_3901 ;
    wire signal_3902 ;
    wire signal_3903 ;
    wire signal_3904 ;
    wire signal_3905 ;
    wire signal_3906 ;
    wire signal_3907 ;
    wire signal_3908 ;
    wire signal_3909 ;
    wire signal_3910 ;
    wire signal_3911 ;
    wire signal_3912 ;
    wire signal_3913 ;
    wire signal_3914 ;
    wire signal_3915 ;
    wire signal_3916 ;
    wire signal_3917 ;
    wire signal_3918 ;
    wire signal_3919 ;
    wire signal_3920 ;
    wire signal_3921 ;
    wire signal_3922 ;
    wire signal_3923 ;
    wire signal_3924 ;
    wire signal_3925 ;
    wire signal_3926 ;
    wire signal_3927 ;
    wire signal_3928 ;
    wire signal_3929 ;
    wire signal_3930 ;
    wire signal_3931 ;
    wire signal_3932 ;
    wire signal_3933 ;
    wire signal_3934 ;
    wire signal_3935 ;
    wire signal_3936 ;
    wire signal_3937 ;
    wire signal_3938 ;
    wire signal_3939 ;
    wire signal_3940 ;
    wire signal_3941 ;
    wire signal_3942 ;
    wire signal_3943 ;
    wire signal_3944 ;
    wire signal_3945 ;
    wire signal_3946 ;
    wire signal_3947 ;
    wire signal_3948 ;
    wire signal_3949 ;
    wire signal_3950 ;
    wire signal_3951 ;
    wire signal_3952 ;
    wire signal_3953 ;
    wire signal_3954 ;
    wire signal_3955 ;
    wire signal_3956 ;
    wire signal_3957 ;
    wire signal_3958 ;
    wire signal_3959 ;
    wire signal_3960 ;
    wire signal_3961 ;
    wire signal_3962 ;
    wire signal_3963 ;
    wire signal_3964 ;
    wire signal_3965 ;
    wire signal_3966 ;
    wire signal_3967 ;
    wire signal_3968 ;
    wire signal_3969 ;
    wire signal_3970 ;
    wire signal_3971 ;
    wire signal_3972 ;
    wire signal_3973 ;
    wire signal_3974 ;
    wire signal_3975 ;
    wire signal_3976 ;
    wire signal_3977 ;
    wire signal_3978 ;
    wire signal_3979 ;
    wire signal_3980 ;
    wire signal_3981 ;
    wire signal_3982 ;
    wire signal_3983 ;
    wire signal_3984 ;
    wire signal_3985 ;
    wire signal_3986 ;
    wire signal_3987 ;
    wire signal_3988 ;
    wire signal_3989 ;
    wire signal_3990 ;
    wire signal_3991 ;
    wire signal_3992 ;
    wire signal_3993 ;
    wire signal_3994 ;
    wire signal_3995 ;
    wire signal_3996 ;
    wire signal_3997 ;
    wire signal_3998 ;
    wire signal_3999 ;
    wire signal_4000 ;
    wire signal_4001 ;
    wire signal_4002 ;
    wire signal_4003 ;
    wire signal_4004 ;
    wire signal_4005 ;
    wire signal_4006 ;
    wire signal_4007 ;
    wire signal_4008 ;
    wire signal_4009 ;
    wire signal_4010 ;
    wire signal_4011 ;
    wire signal_4012 ;
    wire signal_4013 ;
    wire signal_4014 ;
    wire signal_4015 ;
    wire signal_4016 ;
    wire signal_4017 ;
    wire signal_4018 ;
    wire signal_4019 ;
    wire signal_4020 ;
    wire signal_4021 ;
    wire signal_4022 ;
    wire signal_4023 ;
    wire signal_4024 ;
    wire signal_4025 ;
    wire signal_4026 ;
    wire signal_4027 ;
    wire signal_4028 ;
    wire signal_4029 ;
    wire signal_4030 ;
    wire signal_4031 ;
    wire signal_4032 ;
    wire signal_4033 ;
    wire signal_4034 ;
    wire signal_4035 ;
    wire signal_4036 ;
    wire signal_4037 ;
    wire signal_4038 ;
    wire signal_4039 ;
    wire signal_4040 ;
    wire signal_4041 ;
    wire signal_4042 ;
    wire signal_4043 ;
    wire signal_4044 ;
    wire signal_4045 ;
    wire signal_4046 ;
    wire signal_4047 ;
    wire signal_4048 ;
    wire signal_4049 ;
    wire signal_4050 ;
    wire signal_4051 ;
    wire signal_4052 ;
    wire signal_4053 ;
    wire signal_4054 ;
    wire signal_4055 ;
    wire signal_4056 ;
    wire signal_4057 ;
    wire signal_4058 ;
    wire signal_4059 ;
    wire signal_4060 ;
    wire signal_4061 ;
    wire signal_4062 ;
    wire signal_4063 ;
    wire signal_4064 ;
    wire signal_4065 ;
    wire signal_4066 ;
    wire signal_4067 ;
    wire signal_4068 ;
    wire signal_4069 ;
    wire signal_4070 ;
    wire signal_4071 ;
    wire signal_4072 ;
    wire signal_4073 ;
    wire signal_4074 ;
    wire signal_4075 ;
    wire signal_4076 ;
    wire signal_4077 ;
    wire signal_4078 ;
    wire signal_4079 ;
    wire signal_4080 ;
    wire signal_4081 ;
    wire signal_4082 ;
    wire signal_4083 ;
    wire signal_4084 ;
    wire signal_4085 ;
    wire signal_4086 ;
    wire signal_4087 ;
    wire signal_4088 ;
    wire signal_4089 ;
    wire signal_4090 ;
    wire signal_4091 ;
    wire signal_4092 ;
    wire signal_4093 ;
    wire signal_4094 ;
    wire signal_4095 ;
    wire signal_4096 ;
    wire signal_4097 ;
    wire signal_4098 ;
    wire signal_4099 ;
    wire signal_4100 ;
    wire signal_4101 ;
    wire signal_4102 ;
    wire signal_4103 ;
    wire signal_4104 ;
    wire signal_4105 ;
    wire signal_4106 ;
    wire signal_4107 ;
    wire signal_4108 ;
    wire signal_4109 ;
    wire signal_4110 ;
    wire signal_4111 ;
    wire signal_4112 ;
    wire signal_4113 ;
    wire signal_4114 ;
    wire signal_4115 ;
    wire signal_4116 ;
    wire signal_4117 ;
    wire signal_4118 ;
    wire signal_4119 ;
    wire signal_4120 ;
    wire signal_4121 ;
    wire signal_4122 ;
    wire signal_4123 ;
    wire signal_4124 ;
    wire signal_4125 ;
    wire signal_4126 ;
    wire signal_4127 ;
    wire signal_4128 ;
    wire signal_4129 ;
    wire signal_4130 ;
    wire signal_4131 ;
    wire signal_4132 ;
    wire signal_4133 ;
    wire signal_4134 ;
    wire signal_4135 ;
    wire signal_4136 ;
    wire signal_4137 ;
    wire signal_4138 ;
    wire signal_4139 ;
    wire signal_4140 ;
    wire signal_4141 ;
    wire signal_4142 ;
    wire signal_4143 ;
    wire signal_4144 ;
    wire signal_4145 ;
    wire signal_4146 ;
    wire signal_4147 ;
    wire signal_4148 ;
    wire signal_4149 ;
    wire signal_4150 ;
    wire signal_4151 ;
    wire signal_4152 ;
    wire signal_4153 ;
    wire signal_4154 ;
    wire signal_4155 ;
    wire signal_4156 ;
    wire signal_4157 ;
    wire signal_4158 ;
    wire signal_4159 ;
    wire signal_4160 ;
    wire signal_4161 ;
    wire signal_4162 ;
    wire signal_4163 ;
    wire signal_4164 ;
    wire signal_4165 ;
    wire signal_4166 ;
    wire signal_4167 ;
    wire signal_4168 ;
    wire signal_4169 ;
    wire signal_4170 ;
    wire signal_4171 ;
    wire signal_4172 ;
    wire signal_4173 ;
    wire signal_4174 ;
    wire signal_4175 ;
    wire signal_4176 ;
    wire signal_4177 ;
    wire signal_4178 ;
    wire signal_4179 ;
    wire signal_4180 ;
    wire signal_4181 ;
    wire signal_4182 ;
    wire signal_4183 ;
    wire signal_4184 ;
    wire signal_4185 ;
    wire signal_4186 ;
    wire signal_4187 ;
    wire signal_4188 ;
    wire signal_4189 ;
    wire signal_4190 ;
    wire signal_4191 ;
    wire signal_4192 ;
    wire signal_4193 ;
    wire signal_4194 ;
    wire signal_4195 ;
    wire signal_4196 ;
    wire signal_4197 ;
    wire signal_4198 ;
    wire signal_4199 ;
    wire signal_4200 ;
    wire signal_4201 ;
    wire signal_4202 ;
    wire signal_4203 ;
    wire signal_4204 ;
    wire signal_4205 ;
    wire signal_4206 ;
    wire signal_4207 ;
    wire signal_4208 ;
    wire signal_4209 ;
    wire signal_4210 ;
    wire signal_4211 ;
    wire signal_4212 ;
    wire signal_4213 ;
    wire signal_4214 ;
    wire signal_4215 ;
    wire signal_4216 ;
    wire signal_4217 ;
    wire signal_4218 ;
    wire signal_4219 ;
    wire signal_4220 ;
    wire signal_4221 ;
    wire signal_4222 ;
    wire signal_4223 ;
    wire signal_4224 ;
    wire signal_4225 ;
    wire signal_4226 ;
    wire signal_4227 ;
    wire signal_4228 ;
    wire signal_4229 ;
    wire signal_4230 ;
    wire signal_4231 ;
    wire signal_4232 ;
    wire signal_4233 ;
    wire signal_4234 ;
    wire signal_4235 ;
    wire signal_4236 ;
    wire signal_4237 ;
    wire signal_4238 ;
    wire signal_4239 ;
    wire signal_4240 ;
    wire signal_4241 ;
    wire signal_4242 ;
    wire signal_4243 ;
    wire signal_4244 ;
    wire signal_4245 ;
    wire signal_4246 ;
    wire signal_4247 ;
    wire signal_4248 ;
    wire signal_4249 ;
    wire signal_4250 ;
    wire signal_4251 ;
    wire signal_4252 ;
    wire signal_4253 ;
    wire signal_4254 ;
    wire signal_4255 ;
    wire signal_4256 ;
    wire signal_4257 ;
    wire signal_4258 ;
    wire signal_4259 ;
    wire signal_4260 ;
    wire signal_4261 ;
    wire signal_4262 ;
    wire signal_4263 ;
    wire signal_4264 ;
    wire signal_4265 ;
    wire signal_4266 ;
    wire signal_4267 ;
    wire signal_4268 ;
    wire signal_4269 ;
    wire signal_4270 ;
    wire signal_4271 ;
    wire signal_4272 ;
    wire signal_4273 ;
    wire signal_4274 ;
    wire signal_4275 ;
    wire signal_4276 ;
    wire signal_4277 ;
    wire signal_4278 ;
    wire signal_4279 ;
    wire signal_4280 ;
    wire signal_4281 ;
    wire signal_4282 ;
    wire signal_4283 ;
    wire signal_4284 ;
    wire signal_4285 ;
    wire signal_4286 ;
    wire signal_4287 ;
    wire signal_4288 ;
    wire signal_4289 ;
    wire signal_4290 ;
    wire signal_4291 ;
    wire signal_4292 ;
    wire signal_4293 ;
    wire signal_4294 ;
    wire signal_4295 ;
    wire signal_4296 ;
    wire signal_4297 ;
    wire signal_4298 ;
    wire signal_4299 ;
    wire signal_4300 ;
    wire signal_4301 ;
    wire signal_4302 ;
    wire signal_4303 ;
    wire signal_4304 ;
    wire signal_4305 ;
    wire signal_4306 ;
    wire signal_4307 ;
    wire signal_4308 ;
    wire signal_4309 ;
    wire signal_4310 ;
    wire signal_4311 ;
    wire signal_4312 ;
    wire signal_4313 ;
    wire signal_4314 ;
    wire signal_4315 ;
    wire signal_4316 ;
    wire signal_4317 ;
    wire signal_4318 ;
    wire signal_4319 ;
    wire signal_4320 ;
    wire signal_4321 ;
    wire signal_4322 ;
    wire signal_4323 ;
    wire signal_4324 ;
    wire signal_4325 ;
    wire signal_4326 ;
    wire signal_4327 ;
    wire signal_4328 ;
    wire signal_4329 ;
    wire signal_4330 ;
    wire signal_4331 ;
    wire signal_4332 ;
    wire signal_4333 ;
    wire signal_4334 ;
    wire signal_4335 ;
    wire signal_4336 ;
    wire signal_4337 ;
    wire signal_4338 ;
    wire signal_4339 ;
    wire signal_4340 ;
    wire signal_4341 ;
    wire signal_4342 ;
    wire signal_4343 ;
    wire signal_4344 ;
    wire signal_4345 ;
    wire signal_4346 ;
    wire signal_4347 ;
    wire signal_4348 ;
    wire signal_4349 ;
    wire signal_4350 ;
    wire signal_4351 ;
    wire signal_4352 ;
    wire signal_4353 ;
    wire signal_4354 ;
    wire signal_4355 ;
    wire signal_4356 ;
    wire signal_4357 ;
    wire signal_4358 ;
    wire signal_4359 ;
    wire signal_4360 ;
    wire signal_4361 ;
    wire signal_4362 ;
    wire signal_4363 ;
    wire signal_4364 ;
    wire signal_4365 ;
    wire signal_4366 ;
    wire signal_4367 ;
    wire signal_4368 ;
    wire signal_4369 ;
    wire signal_4370 ;
    wire signal_4371 ;
    wire signal_4372 ;
    wire signal_4373 ;
    wire signal_4374 ;
    wire signal_4375 ;
    wire signal_4376 ;
    wire signal_4377 ;
    wire signal_4378 ;
    wire signal_4379 ;
    wire signal_4380 ;
    wire signal_4381 ;
    wire signal_4382 ;
    wire signal_4383 ;
    wire signal_4384 ;
    wire signal_4385 ;
    wire signal_4386 ;
    wire signal_4387 ;
    wire signal_4388 ;
    wire signal_4389 ;
    wire signal_4390 ;
    wire signal_4391 ;
    wire signal_4392 ;
    wire signal_4393 ;
    wire signal_4394 ;
    wire signal_4395 ;
    wire signal_4396 ;
    wire signal_4397 ;
    wire signal_4398 ;
    wire signal_4399 ;
    wire signal_4400 ;
    wire signal_4401 ;
    wire signal_4402 ;
    wire signal_4403 ;
    wire signal_4404 ;
    wire signal_4405 ;
    wire signal_4406 ;
    wire signal_4407 ;
    wire signal_4408 ;
    wire signal_4409 ;
    wire signal_4410 ;
    wire signal_4411 ;
    wire signal_4412 ;
    wire signal_4413 ;
    wire signal_4414 ;
    wire signal_4415 ;
    wire signal_4416 ;
    wire signal_4417 ;
    wire signal_4418 ;
    wire signal_4419 ;
    wire signal_4420 ;
    wire signal_4421 ;
    wire signal_4422 ;
    wire signal_4423 ;
    wire signal_4424 ;
    wire signal_4425 ;
    wire signal_4426 ;
    wire signal_4427 ;
    wire signal_4428 ;
    wire signal_4429 ;
    wire signal_4430 ;
    wire signal_4431 ;
    wire signal_4432 ;
    wire signal_4433 ;
    wire signal_4434 ;
    wire signal_4435 ;
    wire signal_4436 ;
    wire signal_4437 ;
    wire signal_4438 ;
    wire signal_4439 ;
    wire signal_4440 ;
    wire signal_4441 ;
    wire signal_4442 ;
    wire signal_4443 ;
    wire signal_4444 ;
    wire signal_4445 ;
    wire signal_4446 ;
    wire signal_4447 ;
    wire signal_4448 ;
    wire signal_4449 ;
    wire signal_4450 ;
    wire signal_4451 ;
    wire signal_4452 ;
    wire signal_4453 ;
    wire signal_4454 ;
    wire signal_4455 ;
    wire signal_4456 ;
    wire signal_4457 ;
    wire signal_4458 ;
    wire signal_4459 ;
    wire signal_4460 ;
    wire signal_4461 ;
    wire signal_4462 ;
    wire signal_4463 ;
    wire signal_4464 ;
    wire signal_4465 ;
    wire signal_4466 ;
    wire signal_4467 ;
    wire signal_4468 ;
    wire signal_4469 ;
    wire signal_4470 ;
    wire signal_4471 ;
    wire signal_4472 ;
    wire signal_4473 ;
    wire signal_4474 ;
    wire signal_4475 ;
    wire signal_4476 ;
    wire signal_4477 ;
    wire signal_4478 ;
    wire signal_4479 ;
    wire signal_4480 ;
    wire signal_4481 ;
    wire signal_4482 ;
    wire signal_4483 ;
    wire signal_4484 ;
    wire signal_4485 ;
    wire signal_4486 ;
    wire signal_4487 ;
    wire signal_4488 ;
    wire signal_4489 ;
    wire signal_4490 ;
    wire signal_4491 ;
    wire signal_4492 ;
    wire signal_4493 ;
    wire signal_4494 ;
    wire signal_4495 ;
    wire signal_4496 ;
    wire signal_4497 ;
    wire signal_4498 ;
    wire signal_4499 ;
    wire signal_4500 ;
    wire signal_4501 ;
    wire signal_4502 ;
    wire signal_4503 ;
    wire signal_4504 ;
    wire signal_4505 ;
    wire signal_4506 ;
    wire signal_4507 ;
    wire signal_4508 ;
    wire signal_4509 ;
    wire signal_4510 ;
    wire signal_4511 ;
    wire signal_4512 ;
    wire signal_4513 ;
    wire signal_4514 ;
    wire signal_4515 ;
    wire signal_4516 ;
    wire signal_4517 ;
    wire signal_4518 ;
    wire signal_4519 ;
    wire signal_4520 ;
    wire signal_4521 ;
    wire signal_4522 ;
    wire signal_4523 ;
    wire signal_4524 ;
    wire signal_4525 ;
    wire signal_4526 ;
    wire signal_4527 ;
    wire signal_4528 ;
    wire signal_4529 ;
    wire signal_4530 ;
    wire signal_4531 ;
    wire signal_4532 ;
    wire signal_4533 ;
    wire signal_4534 ;
    wire signal_4535 ;
    wire signal_4536 ;
    wire signal_4537 ;
    wire signal_4538 ;
    wire signal_4539 ;
    wire signal_4540 ;
    wire signal_4541 ;
    wire signal_4542 ;
    wire signal_4543 ;
    wire signal_4544 ;
    wire signal_4545 ;
    wire signal_4546 ;
    wire signal_4547 ;
    wire signal_4548 ;
    wire signal_4549 ;
    wire signal_4550 ;
    wire signal_4551 ;
    wire signal_4552 ;
    wire signal_4553 ;
    wire signal_4554 ;
    wire signal_4555 ;
    wire signal_4556 ;
    wire signal_4557 ;
    wire signal_4558 ;
    wire signal_4559 ;
    wire signal_4560 ;
    wire signal_4561 ;
    wire signal_4562 ;
    wire signal_4563 ;
    wire signal_4564 ;
    wire signal_4565 ;
    wire signal_4566 ;
    wire signal_4567 ;
    wire signal_4568 ;
    wire signal_4569 ;
    wire signal_4570 ;
    wire signal_4571 ;
    wire signal_4572 ;
    wire signal_4573 ;
    wire signal_4574 ;
    wire signal_4575 ;
    wire signal_4576 ;
    wire signal_4577 ;
    wire signal_4578 ;
    wire signal_4579 ;
    wire signal_4580 ;
    wire signal_4581 ;
    wire signal_4582 ;
    wire signal_4583 ;
    wire signal_4584 ;
    wire signal_4585 ;
    wire signal_4586 ;
    wire signal_4587 ;
    wire signal_4588 ;
    wire signal_4589 ;
    wire signal_4590 ;
    wire signal_4591 ;
    wire signal_4592 ;
    wire signal_4593 ;
    wire signal_4594 ;
    wire signal_4595 ;
    wire signal_4596 ;
    wire signal_4597 ;
    wire signal_4598 ;
    wire signal_4599 ;
    wire signal_4600 ;
    wire signal_4601 ;
    wire signal_4602 ;
    wire signal_4603 ;
    wire signal_4604 ;
    wire signal_4605 ;
    wire signal_4606 ;
    wire signal_4607 ;
    wire signal_4608 ;
    wire signal_4609 ;
    wire signal_4610 ;
    wire signal_4611 ;
    wire signal_4612 ;
    wire signal_4613 ;
    wire signal_4614 ;
    wire signal_4615 ;
    wire signal_4616 ;
    wire signal_4617 ;
    wire signal_4618 ;
    wire signal_4619 ;
    wire signal_4620 ;
    wire signal_4621 ;
    wire signal_4622 ;
    wire signal_4623 ;
    wire signal_4624 ;
    wire signal_4625 ;
    wire signal_4626 ;
    wire signal_4627 ;
    wire signal_4628 ;
    wire signal_4629 ;
    wire signal_4630 ;
    wire signal_4631 ;
    wire signal_4632 ;
    wire signal_4633 ;
    wire signal_4634 ;
    wire signal_4635 ;
    wire signal_4636 ;
    wire signal_4637 ;
    wire signal_4638 ;
    wire signal_4639 ;
    wire signal_4640 ;
    wire signal_4641 ;
    wire signal_4642 ;
    wire signal_4643 ;
    wire signal_4644 ;
    wire signal_4645 ;
    wire signal_4646 ;
    wire signal_4647 ;
    wire signal_4648 ;
    wire signal_4649 ;
    wire signal_4650 ;
    wire signal_4651 ;
    wire signal_4652 ;
    wire signal_4653 ;
    wire signal_4654 ;
    wire signal_4655 ;
    wire signal_4656 ;
    wire signal_4657 ;
    wire signal_4658 ;
    wire signal_4659 ;
    wire signal_4660 ;
    wire signal_4661 ;
    wire signal_4662 ;
    wire signal_4663 ;
    wire signal_4664 ;
    wire signal_4665 ;
    wire signal_4666 ;
    wire signal_4667 ;
    wire signal_4668 ;
    wire signal_4669 ;
    wire signal_4670 ;
    wire signal_4671 ;
    wire signal_4672 ;
    wire signal_4673 ;
    wire signal_4674 ;
    wire signal_4675 ;
    wire signal_4676 ;
    wire signal_4677 ;
    wire signal_4678 ;
    wire signal_4679 ;
    wire signal_4680 ;
    wire signal_4681 ;
    wire signal_4682 ;
    wire signal_4683 ;
    wire signal_4684 ;
    wire signal_4685 ;
    wire signal_4686 ;
    wire signal_4687 ;
    wire signal_4688 ;
    wire signal_4689 ;
    wire signal_4690 ;
    wire signal_4691 ;
    wire signal_4692 ;
    wire signal_4693 ;
    wire signal_4694 ;
    wire signal_4695 ;
    wire signal_4696 ;
    wire signal_4697 ;
    wire signal_4698 ;
    wire signal_4699 ;
    wire signal_4700 ;
    wire signal_4701 ;
    wire signal_4702 ;
    wire signal_4703 ;
    wire signal_4704 ;
    wire signal_4705 ;
    wire signal_4706 ;
    wire signal_4707 ;
    wire signal_4708 ;
    wire signal_4709 ;
    wire signal_4710 ;
    wire signal_4711 ;
    wire signal_4712 ;
    wire signal_4713 ;
    wire signal_4714 ;
    wire signal_4715 ;
    wire signal_4716 ;
    wire signal_4717 ;
    wire signal_4718 ;
    wire signal_4719 ;
    wire signal_4720 ;
    wire signal_4721 ;
    wire signal_4722 ;
    wire signal_4723 ;
    wire signal_4724 ;
    wire signal_4725 ;
    wire signal_4726 ;
    wire signal_4727 ;
    wire signal_4728 ;
    wire signal_4729 ;
    wire signal_4730 ;
    wire signal_4731 ;
    wire signal_4732 ;
    wire signal_4733 ;
    wire signal_4734 ;
    wire signal_4735 ;
    wire signal_4736 ;
    wire signal_4737 ;
    wire signal_4738 ;
    wire signal_4739 ;
    wire signal_4740 ;
    wire signal_4741 ;
    wire signal_4742 ;
    wire signal_4743 ;
    wire signal_4744 ;
    wire signal_4745 ;
    wire signal_4746 ;
    wire signal_4747 ;
    wire signal_4748 ;
    wire signal_4749 ;
    wire signal_4750 ;
    wire signal_4751 ;
    wire signal_4752 ;
    wire signal_4753 ;
    wire signal_4754 ;
    wire signal_4755 ;
    wire signal_4756 ;
    wire signal_4757 ;
    wire signal_4758 ;
    wire signal_4759 ;
    wire signal_4760 ;
    wire signal_4761 ;
    wire signal_4762 ;
    wire signal_4763 ;
    wire signal_4764 ;
    wire signal_4765 ;
    wire signal_4766 ;
    wire signal_4767 ;
    wire signal_4768 ;
    wire signal_4769 ;
    wire signal_4770 ;
    wire signal_4771 ;
    wire signal_4772 ;
    wire signal_4773 ;
    wire signal_4774 ;
    wire signal_4775 ;
    wire signal_4776 ;
    wire signal_4777 ;
    wire signal_4778 ;
    wire signal_4779 ;
    wire signal_4780 ;
    wire signal_4781 ;
    wire signal_4782 ;
    wire signal_4783 ;
    wire signal_4784 ;
    wire signal_4785 ;
    wire signal_4786 ;
    wire signal_4787 ;
    wire signal_4788 ;
    wire signal_4789 ;
    wire signal_4790 ;
    wire signal_4791 ;
    wire signal_4792 ;
    wire signal_4793 ;
    wire signal_4794 ;
    wire signal_4795 ;
    wire signal_4796 ;
    wire signal_4797 ;
    wire signal_4798 ;
    wire signal_4799 ;
    wire signal_4800 ;
    wire signal_4801 ;
    wire signal_4802 ;
    wire signal_4803 ;
    wire signal_4804 ;
    wire signal_4805 ;
    wire signal_4806 ;
    wire signal_4807 ;
    wire signal_4808 ;
    wire signal_4809 ;
    wire signal_4810 ;
    wire signal_4811 ;
    wire signal_4812 ;
    wire signal_4813 ;
    wire signal_4814 ;
    wire signal_4815 ;
    wire signal_4816 ;
    wire signal_4817 ;
    wire signal_4818 ;
    wire signal_4819 ;
    wire signal_4820 ;
    wire signal_4821 ;
    wire signal_4822 ;
    wire signal_4823 ;
    wire signal_4824 ;
    wire signal_4825 ;
    wire signal_4826 ;
    wire signal_4827 ;
    wire signal_4828 ;
    wire signal_4829 ;
    wire signal_4830 ;
    wire signal_4831 ;
    wire signal_4832 ;
    wire signal_4833 ;
    wire signal_4834 ;
    wire signal_4835 ;
    wire signal_4836 ;
    wire signal_4837 ;
    wire signal_4838 ;
    wire signal_4839 ;
    wire signal_4840 ;
    wire signal_4841 ;
    wire signal_4842 ;
    wire signal_4843 ;
    wire signal_4844 ;
    wire signal_4845 ;
    wire signal_4846 ;
    wire signal_4847 ;
    wire signal_4848 ;
    wire signal_4849 ;
    wire signal_4850 ;
    wire signal_4851 ;
    wire signal_4852 ;
    wire signal_4853 ;
    wire signal_4854 ;
    wire signal_4855 ;
    wire signal_4856 ;
    wire signal_4857 ;
    wire signal_4858 ;
    wire signal_4859 ;
    wire signal_4860 ;
    wire signal_4861 ;
    wire signal_4862 ;
    wire signal_4863 ;
    wire signal_4864 ;
    wire signal_4865 ;
    wire signal_4866 ;
    wire signal_4867 ;
    wire signal_4868 ;
    wire signal_4869 ;
    wire signal_4870 ;
    wire signal_4871 ;
    wire signal_4872 ;
    wire signal_4873 ;
    wire signal_4874 ;
    wire signal_4875 ;
    wire signal_4876 ;
    wire signal_4877 ;
    wire signal_4878 ;
    wire signal_4879 ;
    wire signal_4880 ;
    wire signal_4881 ;
    wire signal_4882 ;
    wire signal_4883 ;
    wire signal_4884 ;
    wire signal_4885 ;
    wire signal_4886 ;
    wire signal_4887 ;
    wire signal_4888 ;
    wire signal_4889 ;
    wire signal_4890 ;
    wire signal_4891 ;
    wire signal_4892 ;
    wire signal_4893 ;
    wire signal_4894 ;
    wire signal_4895 ;
    wire signal_4896 ;
    wire signal_4897 ;
    wire signal_4898 ;
    wire signal_4899 ;
    wire signal_4900 ;
    wire signal_4901 ;
    wire signal_4902 ;
    wire signal_4903 ;
    wire signal_4904 ;
    wire signal_4905 ;
    wire signal_4906 ;
    wire signal_4907 ;
    wire signal_4908 ;
    wire signal_4909 ;
    wire signal_4910 ;
    wire signal_4911 ;
    wire signal_4912 ;
    wire signal_4913 ;
    wire signal_4914 ;
    wire signal_4915 ;
    wire signal_4916 ;
    wire signal_4917 ;
    wire signal_4918 ;
    wire signal_4919 ;
    wire signal_4920 ;
    wire signal_4921 ;
    wire signal_4922 ;
    wire signal_4923 ;
    wire signal_4924 ;
    wire signal_4925 ;
    wire signal_4926 ;
    wire signal_4927 ;
    wire signal_4928 ;
    wire signal_4929 ;
    wire signal_4930 ;
    wire signal_4931 ;
    wire signal_4932 ;
    wire signal_4933 ;
    wire signal_4934 ;
    wire signal_4935 ;
    wire signal_4936 ;
    wire signal_4937 ;
    wire signal_4938 ;
    wire signal_4939 ;
    wire signal_4940 ;
    wire signal_4941 ;
    wire signal_4942 ;
    wire signal_4943 ;
    wire signal_4944 ;
    wire signal_4945 ;
    wire signal_4946 ;
    wire signal_4947 ;
    wire signal_4948 ;
    wire signal_4949 ;
    wire signal_4950 ;
    wire signal_4951 ;
    wire signal_4952 ;
    wire signal_4953 ;
    wire signal_4954 ;
    wire signal_4955 ;
    wire signal_4956 ;
    wire signal_4957 ;
    wire signal_4958 ;
    wire signal_4959 ;
    wire signal_4960 ;
    wire signal_4961 ;
    wire signal_4962 ;
    wire signal_4963 ;
    wire signal_4964 ;
    wire signal_4965 ;
    wire signal_4966 ;
    wire signal_4967 ;
    wire signal_4968 ;
    wire signal_4969 ;
    wire signal_4970 ;
    wire signal_4971 ;
    wire signal_4972 ;
    wire signal_4973 ;
    wire signal_4974 ;
    wire signal_4975 ;
    wire signal_4976 ;
    wire signal_4977 ;
    wire signal_4978 ;
    wire signal_4979 ;
    wire signal_4980 ;
    wire signal_4981 ;
    wire signal_4982 ;
    wire signal_4983 ;
    wire signal_4984 ;
    wire signal_4985 ;
    wire signal_4986 ;
    wire signal_4987 ;
    wire signal_4988 ;
    wire signal_4989 ;
    wire signal_4990 ;
    wire signal_4991 ;
    wire signal_4992 ;
    wire signal_4993 ;
    wire signal_4994 ;
    wire signal_4995 ;
    wire signal_4996 ;
    wire signal_4997 ;
    wire signal_4998 ;
    wire signal_4999 ;
    wire signal_5000 ;
    wire signal_5001 ;
    wire signal_5002 ;
    wire signal_5003 ;
    wire signal_5004 ;
    wire signal_5005 ;
    wire signal_5006 ;
    wire signal_5007 ;
    wire signal_5008 ;
    wire signal_5009 ;
    wire signal_5010 ;
    wire signal_5011 ;
    wire signal_5012 ;
    wire signal_5013 ;
    wire signal_5014 ;
    wire signal_5015 ;
    wire signal_5016 ;
    wire signal_5017 ;
    wire signal_5018 ;
    wire signal_5019 ;
    wire signal_5020 ;
    wire signal_5021 ;
    wire signal_5022 ;
    wire signal_5023 ;
    wire signal_5024 ;
    wire signal_5025 ;
    wire signal_5026 ;
    wire signal_5027 ;
    wire signal_5028 ;
    wire signal_5029 ;
    wire signal_5030 ;
    wire signal_5031 ;
    wire signal_5032 ;
    wire signal_5033 ;
    wire signal_5034 ;
    wire signal_5035 ;
    wire signal_5036 ;
    wire signal_5037 ;
    wire signal_5038 ;
    wire signal_5039 ;
    wire signal_5040 ;
    wire signal_5041 ;
    wire signal_5042 ;
    wire signal_5043 ;
    wire signal_5044 ;
    wire signal_5045 ;
    wire signal_5046 ;
    wire signal_5047 ;
    wire signal_5048 ;
    wire signal_5049 ;
    wire signal_5050 ;
    wire signal_5051 ;
    wire signal_5052 ;
    wire signal_5053 ;
    wire signal_5054 ;
    wire signal_5055 ;
    wire signal_5056 ;
    wire signal_5057 ;
    wire signal_5058 ;
    wire signal_5059 ;
    wire signal_5060 ;
    wire signal_5061 ;
    wire signal_5062 ;
    wire signal_5063 ;
    wire signal_5064 ;
    wire signal_5065 ;
    wire signal_5066 ;
    wire signal_5067 ;
    wire signal_5068 ;
    wire signal_5069 ;
    wire signal_5070 ;
    wire signal_5071 ;
    wire signal_5072 ;
    wire signal_5073 ;
    wire signal_5074 ;
    wire signal_5075 ;
    wire signal_5076 ;
    wire signal_5077 ;
    wire signal_5078 ;
    wire signal_5079 ;
    wire signal_5080 ;
    wire signal_5081 ;
    wire signal_5082 ;
    wire signal_5083 ;
    wire signal_5084 ;
    wire signal_5085 ;
    wire signal_5086 ;
    wire signal_5087 ;
    wire signal_5088 ;
    wire signal_5089 ;
    wire signal_5090 ;
    wire signal_5091 ;
    wire signal_5092 ;
    wire signal_5093 ;
    wire signal_5094 ;
    wire signal_5095 ;
    wire signal_5096 ;
    wire signal_5097 ;
    wire signal_5098 ;
    wire signal_5099 ;
    wire signal_5100 ;
    wire signal_5101 ;
    wire signal_5102 ;
    wire signal_5103 ;
    wire signal_5104 ;
    wire signal_5105 ;
    wire signal_5106 ;
    wire signal_5107 ;
    wire signal_5108 ;
    wire signal_5109 ;
    wire signal_5110 ;
    wire signal_5111 ;
    wire signal_5112 ;
    wire signal_5113 ;
    wire signal_5114 ;
    wire signal_5115 ;
    wire signal_5116 ;
    wire signal_5117 ;
    wire signal_5118 ;
    wire signal_5119 ;
    wire signal_5120 ;
    wire signal_5121 ;
    wire signal_5122 ;
    wire signal_5123 ;
    wire signal_5124 ;
    wire signal_5125 ;
    wire signal_5126 ;
    wire signal_5127 ;
    wire signal_5128 ;
    wire signal_5129 ;
    wire signal_5130 ;
    wire signal_5131 ;
    wire signal_5132 ;
    wire signal_5133 ;
    wire signal_5134 ;
    wire signal_5135 ;
    wire signal_5136 ;
    wire signal_5137 ;
    wire signal_5138 ;
    wire signal_5139 ;
    wire signal_5140 ;
    wire signal_5141 ;
    wire signal_5142 ;
    wire signal_5143 ;
    wire signal_5144 ;
    wire signal_5145 ;
    wire signal_5146 ;
    wire signal_5147 ;
    wire signal_5148 ;
    wire signal_5149 ;
    wire signal_5150 ;
    wire signal_5151 ;
    wire signal_5152 ;
    wire signal_5153 ;
    wire signal_5154 ;
    wire signal_5155 ;
    wire signal_5156 ;
    wire signal_5157 ;
    wire signal_5158 ;
    wire signal_5159 ;
    wire signal_5160 ;
    wire signal_5161 ;
    wire signal_5162 ;
    wire signal_5163 ;
    wire signal_5164 ;
    wire signal_5165 ;
    wire signal_5166 ;
    wire signal_5167 ;
    wire signal_5168 ;
    wire signal_5169 ;
    wire signal_5170 ;
    wire signal_5171 ;
    wire signal_5172 ;
    wire signal_5173 ;
    wire signal_5174 ;
    wire signal_5175 ;
    wire signal_5176 ;
    wire signal_5177 ;
    wire signal_5178 ;
    wire signal_5179 ;
    wire signal_5180 ;
    wire signal_5181 ;
    wire signal_5182 ;
    wire signal_5183 ;
    wire signal_5184 ;
    wire signal_5185 ;
    wire signal_5186 ;
    wire signal_5187 ;
    wire signal_5188 ;
    wire signal_5189 ;
    wire signal_5190 ;
    wire signal_5191 ;
    wire signal_5192 ;
    wire signal_5193 ;
    wire signal_5194 ;
    wire signal_5195 ;
    wire signal_5196 ;
    wire signal_5197 ;
    wire signal_5198 ;
    wire signal_5199 ;
    wire signal_5200 ;
    wire signal_5201 ;
    wire signal_5202 ;
    wire signal_5203 ;
    wire signal_5204 ;
    wire signal_5205 ;
    wire signal_5206 ;
    wire signal_5207 ;
    wire signal_5208 ;
    wire signal_5209 ;
    wire signal_5210 ;
    wire signal_5211 ;
    wire signal_5212 ;
    wire signal_5213 ;
    wire signal_5214 ;
    wire signal_5215 ;
    wire signal_5216 ;
    wire signal_5217 ;
    wire signal_5218 ;
    wire signal_5219 ;
    wire signal_5220 ;
    wire signal_5221 ;
    wire signal_5222 ;
    wire signal_5223 ;
    wire signal_5224 ;
    wire signal_5225 ;
    wire signal_5226 ;
    wire signal_5227 ;
    wire signal_5228 ;
    wire signal_5229 ;
    wire signal_5230 ;
    wire signal_5231 ;
    wire signal_5232 ;
    wire signal_5233 ;
    wire signal_5234 ;
    wire signal_5235 ;
    wire signal_5236 ;
    wire signal_5237 ;
    wire signal_5238 ;
    wire signal_5239 ;
    wire signal_5240 ;
    wire signal_5241 ;
    wire signal_5242 ;
    wire signal_5243 ;
    wire signal_5244 ;
    wire signal_5245 ;
    wire signal_5246 ;
    wire signal_5247 ;
    wire signal_5248 ;
    wire signal_5249 ;
    wire signal_5250 ;
    wire signal_5251 ;
    wire signal_5252 ;
    wire signal_5253 ;
    wire signal_5254 ;
    wire signal_5255 ;
    wire signal_5256 ;
    wire signal_5257 ;
    wire signal_5258 ;
    wire signal_5259 ;
    wire signal_5260 ;
    wire signal_5261 ;
    wire signal_5262 ;
    wire signal_5263 ;
    wire signal_5264 ;
    wire signal_5265 ;
    wire signal_5266 ;
    wire signal_5267 ;
    wire signal_5268 ;
    wire signal_5269 ;
    wire signal_5270 ;
    wire signal_5271 ;
    wire signal_5272 ;
    wire signal_5273 ;
    wire signal_5274 ;
    wire signal_5275 ;
    wire signal_5276 ;
    wire signal_5277 ;
    wire signal_5278 ;
    wire signal_5279 ;
    wire signal_5280 ;
    wire signal_5281 ;
    wire signal_5282 ;
    wire signal_5283 ;
    wire signal_5284 ;
    wire signal_5285 ;
    wire signal_5286 ;
    wire signal_5287 ;
    wire signal_5288 ;
    wire signal_5289 ;
    wire signal_5290 ;
    wire signal_5291 ;
    wire signal_5292 ;
    wire signal_5293 ;
    wire signal_5294 ;
    wire signal_5295 ;
    wire signal_5296 ;
    wire signal_5297 ;
    wire signal_5298 ;
    wire signal_5299 ;
    wire signal_5300 ;
    wire signal_5301 ;
    wire signal_5302 ;
    wire signal_5303 ;
    wire signal_5304 ;
    wire signal_5305 ;
    wire signal_5306 ;
    wire signal_5307 ;
    wire signal_5308 ;
    wire signal_5309 ;
    wire signal_5310 ;
    wire signal_5311 ;
    wire signal_5312 ;
    wire signal_5313 ;
    wire signal_5314 ;
    wire signal_5315 ;
    wire signal_5316 ;
    wire signal_5317 ;
    wire signal_5318 ;
    wire signal_5319 ;
    wire signal_5320 ;
    wire signal_5321 ;
    wire signal_5322 ;
    wire signal_5323 ;
    wire signal_5324 ;
    wire signal_5325 ;
    wire signal_5326 ;
    wire signal_5327 ;
    wire signal_5328 ;
    wire signal_5329 ;
    wire signal_5330 ;
    wire signal_5331 ;
    wire signal_5332 ;
    wire signal_5333 ;
    wire signal_5334 ;
    wire signal_5335 ;
    wire signal_5336 ;
    wire signal_5337 ;
    wire signal_5338 ;
    wire signal_5339 ;
    wire signal_5340 ;
    wire signal_5341 ;
    wire signal_5342 ;
    wire signal_5343 ;
    wire signal_5344 ;
    wire signal_5345 ;
    wire signal_5346 ;
    wire signal_5347 ;
    wire signal_5348 ;
    wire signal_5349 ;
    wire signal_5350 ;
    wire signal_5351 ;
    wire signal_5352 ;
    wire signal_5353 ;
    wire signal_5354 ;
    wire signal_5355 ;
    wire signal_5356 ;
    wire signal_5357 ;
    wire signal_5358 ;
    wire signal_5359 ;
    wire signal_5360 ;
    wire signal_5361 ;
    wire signal_5362 ;
    wire signal_5363 ;
    wire signal_5364 ;
    wire signal_5365 ;
    wire signal_5366 ;
    wire signal_5367 ;
    wire signal_5368 ;
    wire signal_5369 ;
    wire signal_5370 ;
    wire signal_5371 ;
    wire signal_5372 ;
    wire signal_5373 ;
    wire signal_5374 ;
    wire signal_5375 ;
    wire signal_5376 ;
    wire signal_5377 ;
    wire signal_5378 ;
    wire signal_5379 ;
    wire signal_5380 ;
    wire signal_5381 ;
    wire signal_5382 ;
    wire signal_5383 ;
    wire signal_5384 ;
    wire signal_5385 ;
    wire signal_5386 ;
    wire signal_5387 ;
    wire signal_5388 ;
    wire signal_5389 ;
    wire signal_5390 ;
    wire signal_5391 ;
    wire signal_5392 ;
    wire signal_5393 ;
    wire signal_5394 ;
    wire signal_5395 ;
    wire signal_5396 ;
    wire signal_5397 ;
    wire signal_5398 ;
    wire signal_5399 ;
    wire signal_5400 ;
    wire signal_5401 ;
    wire signal_5402 ;
    wire signal_5403 ;
    wire signal_5404 ;
    wire signal_5405 ;
    wire signal_5406 ;
    wire signal_5407 ;
    wire signal_5408 ;
    wire signal_5409 ;
    wire signal_5410 ;
    wire signal_5411 ;
    wire signal_5412 ;
    wire signal_5413 ;
    wire signal_5414 ;
    wire signal_5415 ;
    wire signal_5416 ;
    wire signal_5417 ;
    wire signal_5418 ;
    wire signal_5419 ;
    wire signal_5420 ;
    wire signal_5421 ;
    wire signal_5422 ;
    wire signal_5423 ;
    wire signal_5424 ;
    wire signal_5425 ;
    wire signal_5426 ;
    wire signal_5427 ;
    wire signal_5428 ;
    wire signal_5429 ;
    wire signal_5430 ;
    wire signal_5431 ;
    wire signal_5432 ;
    wire signal_5433 ;
    wire signal_5434 ;
    wire signal_5435 ;
    wire signal_5436 ;
    wire signal_5437 ;
    wire signal_5438 ;
    wire signal_5439 ;
    wire signal_5440 ;
    wire signal_5441 ;
    wire signal_5442 ;
    wire signal_5443 ;
    wire signal_5444 ;
    wire signal_5445 ;
    wire signal_5446 ;
    wire signal_5447 ;
    wire signal_5448 ;
    wire signal_5449 ;
    wire signal_5450 ;
    wire signal_5451 ;
    wire signal_5452 ;
    wire signal_5453 ;
    wire signal_5454 ;
    wire signal_5455 ;
    wire signal_5456 ;
    wire signal_5457 ;
    wire signal_5458 ;
    wire signal_5459 ;
    wire signal_5460 ;
    wire signal_5461 ;
    wire signal_5462 ;
    wire signal_5463 ;
    wire signal_5464 ;
    wire signal_5465 ;
    wire signal_5466 ;
    wire signal_5467 ;
    wire signal_5468 ;
    wire signal_5469 ;
    wire signal_5470 ;
    wire signal_5471 ;
    wire signal_5472 ;
    wire signal_5473 ;
    wire signal_5474 ;
    wire signal_5475 ;
    wire signal_5476 ;
    wire signal_5477 ;
    wire signal_5478 ;
    wire signal_5479 ;
    wire signal_5480 ;
    wire signal_5481 ;
    wire signal_5482 ;
    wire signal_5483 ;
    wire signal_5484 ;
    wire signal_5485 ;
    wire signal_5486 ;
    wire signal_5487 ;
    wire signal_5488 ;
    wire signal_5489 ;
    wire signal_5490 ;
    wire signal_5491 ;
    wire signal_5492 ;
    wire signal_5493 ;
    wire signal_5494 ;
    wire signal_5495 ;
    wire signal_5496 ;
    wire signal_5497 ;
    wire signal_5498 ;
    wire signal_5499 ;
    wire signal_5500 ;
    wire signal_5501 ;
    wire signal_5502 ;
    wire signal_5503 ;
    wire signal_5504 ;
    wire signal_5505 ;
    wire signal_5506 ;
    wire signal_5507 ;
    wire signal_5508 ;
    wire signal_5509 ;
    wire signal_5510 ;
    wire signal_5511 ;
    wire signal_5512 ;
    wire signal_5513 ;
    wire signal_5514 ;
    wire signal_5515 ;
    wire signal_5516 ;
    wire signal_5517 ;
    wire signal_5518 ;
    wire signal_5519 ;
    wire signal_5520 ;
    wire signal_5521 ;
    wire signal_5522 ;
    wire signal_5523 ;
    wire signal_5524 ;
    wire signal_5525 ;
    wire signal_5526 ;
    wire signal_5527 ;
    wire signal_5528 ;
    wire signal_5529 ;
    wire signal_5530 ;
    wire signal_5531 ;
    wire signal_5532 ;
    wire signal_5533 ;
    wire signal_5534 ;
    wire signal_5535 ;
    wire signal_5536 ;
    wire signal_5537 ;
    wire signal_5538 ;
    wire signal_5539 ;
    wire signal_5540 ;
    wire signal_5541 ;
    wire signal_5542 ;
    wire signal_5543 ;
    wire signal_5544 ;
    wire signal_5545 ;
    wire signal_5546 ;
    wire signal_5547 ;
    wire signal_5548 ;
    wire signal_5549 ;
    wire signal_5550 ;
    wire signal_5551 ;
    wire signal_5552 ;
    wire signal_5553 ;
    wire signal_5554 ;
    wire signal_5555 ;
    wire signal_5556 ;
    wire signal_5557 ;
    wire signal_5558 ;
    wire signal_5559 ;
    wire signal_5560 ;
    wire signal_5561 ;
    wire signal_5562 ;
    wire signal_5563 ;
    wire signal_5564 ;
    wire signal_5565 ;
    wire signal_5566 ;
    wire signal_5567 ;
    wire signal_5568 ;
    wire signal_5569 ;
    wire signal_5570 ;
    wire signal_5571 ;
    wire signal_5572 ;
    wire signal_5573 ;
    wire signal_5574 ;
    wire signal_5575 ;
    wire signal_5576 ;
    wire signal_5577 ;
    wire signal_5578 ;
    wire signal_5579 ;
    wire signal_5580 ;
    wire signal_5581 ;
    wire signal_5582 ;
    wire signal_5583 ;
    wire signal_5584 ;
    wire signal_5585 ;
    wire signal_5586 ;
    wire signal_5587 ;
    wire signal_5588 ;
    wire signal_5589 ;
    wire signal_5590 ;
    wire signal_5591 ;
    wire signal_5592 ;
    wire signal_5593 ;
    wire signal_5594 ;
    wire signal_5595 ;
    wire signal_5596 ;
    wire signal_5597 ;
    wire signal_5598 ;
    wire signal_5599 ;
    wire signal_5600 ;
    wire signal_5601 ;
    wire signal_5602 ;
    wire signal_5603 ;
    wire signal_5604 ;
    wire signal_5605 ;
    wire signal_5606 ;
    wire signal_5607 ;
    wire signal_5608 ;
    wire signal_5609 ;
    wire signal_5610 ;
    wire signal_5611 ;
    wire signal_5612 ;
    wire signal_5613 ;
    wire signal_5614 ;
    wire signal_5615 ;
    wire signal_5616 ;
    wire signal_5617 ;
    wire signal_5618 ;
    wire signal_5619 ;
    wire signal_5620 ;
    wire signal_5621 ;
    wire signal_5622 ;
    wire signal_5623 ;
    wire signal_5624 ;
    wire signal_5625 ;
    wire signal_5626 ;
    wire signal_5627 ;
    wire signal_5628 ;
    wire signal_5629 ;
    wire signal_5630 ;
    wire signal_5631 ;
    wire signal_5632 ;
    wire signal_5633 ;
    wire signal_5634 ;
    wire signal_5635 ;
    wire signal_5636 ;
    wire signal_5637 ;
    wire signal_5638 ;
    wire signal_5639 ;
    wire signal_5640 ;
    wire signal_5641 ;
    wire signal_5642 ;
    wire signal_5643 ;
    wire signal_5644 ;
    wire signal_5645 ;
    wire signal_5646 ;
    wire signal_5647 ;
    wire signal_5648 ;
    wire signal_5649 ;
    wire signal_5650 ;
    wire signal_5651 ;
    wire signal_5652 ;
    wire signal_5653 ;
    wire signal_5654 ;
    wire signal_5655 ;
    wire signal_5656 ;
    wire signal_5657 ;
    wire signal_5658 ;
    wire signal_5659 ;
    wire signal_5660 ;
    wire signal_5661 ;
    wire signal_5662 ;
    wire signal_5663 ;
    wire signal_5664 ;
    wire signal_5665 ;
    wire signal_5666 ;
    wire signal_5667 ;
    wire signal_5668 ;
    wire signal_5669 ;
    wire signal_5670 ;
    wire signal_5671 ;
    wire signal_5672 ;
    wire signal_5673 ;
    wire signal_5674 ;
    wire signal_5675 ;
    wire signal_5676 ;
    wire signal_5677 ;
    wire signal_5678 ;
    wire signal_5679 ;
    wire signal_5680 ;
    wire signal_5681 ;
    wire signal_5682 ;
    wire signal_5683 ;
    wire signal_5684 ;
    wire signal_5685 ;
    wire signal_5686 ;
    wire signal_5687 ;
    wire signal_5688 ;
    wire signal_5689 ;
    wire signal_5690 ;
    wire signal_5691 ;
    wire signal_5692 ;
    wire signal_5693 ;
    wire signal_5694 ;
    wire signal_5695 ;
    wire signal_5696 ;
    wire signal_5697 ;
    wire signal_5698 ;
    wire signal_5699 ;
    wire signal_5700 ;
    wire signal_5701 ;
    wire signal_5702 ;
    wire signal_5703 ;
    wire signal_5704 ;
    wire signal_5705 ;
    wire signal_5706 ;
    wire signal_5707 ;
    wire signal_5708 ;
    wire signal_5709 ;
    wire signal_5710 ;
    wire signal_5711 ;
    wire signal_5712 ;
    wire signal_5713 ;
    wire signal_5714 ;
    wire signal_5715 ;
    wire signal_5716 ;
    wire signal_5717 ;
    wire signal_5718 ;
    wire signal_5719 ;
    wire signal_5720 ;
    wire signal_5721 ;
    wire signal_5722 ;
    wire signal_5723 ;
    wire signal_5724 ;
    wire signal_5725 ;
    wire signal_5726 ;
    wire signal_5727 ;
    wire signal_5728 ;
    wire signal_5729 ;
    wire signal_5730 ;
    wire signal_5731 ;
    wire signal_5732 ;
    wire signal_5733 ;
    wire signal_5734 ;
    wire signal_5735 ;
    wire signal_5736 ;
    wire signal_5737 ;
    wire signal_5738 ;
    wire signal_5739 ;
    wire signal_5740 ;
    wire signal_5741 ;
    wire signal_5742 ;
    wire signal_5743 ;
    wire signal_5744 ;
    wire signal_5745 ;
    wire signal_5746 ;
    wire signal_5747 ;
    wire signal_5748 ;
    wire signal_5749 ;
    wire signal_5750 ;
    wire signal_5751 ;
    wire signal_5752 ;
    wire signal_5753 ;
    wire signal_5754 ;
    wire signal_5755 ;
    wire signal_5756 ;
    wire signal_5757 ;
    wire signal_5758 ;
    wire signal_5759 ;
    wire signal_5760 ;
    wire signal_5761 ;
    wire signal_5762 ;
    wire signal_5763 ;
    wire signal_5764 ;
    wire signal_5765 ;
    wire signal_5766 ;
    wire signal_5767 ;
    wire signal_5768 ;
    wire signal_5769 ;
    wire signal_5770 ;
    wire signal_5771 ;
    wire signal_5772 ;
    wire signal_5773 ;
    wire signal_5774 ;
    wire signal_5775 ;
    wire signal_5776 ;
    wire signal_5777 ;
    wire signal_5778 ;
    wire signal_5779 ;
    wire signal_5780 ;
    wire signal_5781 ;
    wire signal_5782 ;
    wire signal_5783 ;
    wire signal_5784 ;
    wire signal_5785 ;
    wire signal_5786 ;
    wire signal_5787 ;
    wire signal_5788 ;
    wire signal_5789 ;
    wire signal_5790 ;
    wire signal_5791 ;
    wire signal_5792 ;
    wire signal_5793 ;
    wire signal_5794 ;
    wire signal_5795 ;
    wire signal_5796 ;
    wire signal_5797 ;
    wire signal_5798 ;
    wire signal_5799 ;
    wire signal_5800 ;
    wire signal_5801 ;
    wire signal_5802 ;
    wire signal_5803 ;
    wire signal_5804 ;
    wire signal_5805 ;
    wire signal_5806 ;
    wire signal_5807 ;
    wire signal_5808 ;
    wire signal_5809 ;
    wire signal_5810 ;
    wire signal_5811 ;
    wire signal_5812 ;
    wire signal_5813 ;
    wire signal_5814 ;
    wire signal_5815 ;
    wire signal_5816 ;
    wire signal_5817 ;
    wire signal_5818 ;
    wire signal_5819 ;
    wire signal_5820 ;
    wire signal_5821 ;
    wire signal_5822 ;
    wire signal_5823 ;
    wire signal_5824 ;
    wire signal_5825 ;
    wire signal_5826 ;
    wire signal_5827 ;
    wire signal_5828 ;
    wire signal_5829 ;
    wire signal_5830 ;
    wire signal_5831 ;
    wire signal_5832 ;
    wire signal_5833 ;
    wire signal_5834 ;
    wire signal_5835 ;
    wire signal_5836 ;
    wire signal_5837 ;
    wire signal_5838 ;
    wire signal_5839 ;
    wire signal_5840 ;
    wire signal_5841 ;
    wire signal_5842 ;
    wire signal_5843 ;
    wire signal_5844 ;
    wire signal_5845 ;
    wire signal_5846 ;
    wire signal_5847 ;
    wire signal_5848 ;
    wire signal_5849 ;
    wire signal_5850 ;
    wire signal_5851 ;
    wire signal_5852 ;
    wire signal_5853 ;
    wire signal_5854 ;
    wire signal_5855 ;
    wire signal_5856 ;
    wire signal_5857 ;
    wire signal_5858 ;
    wire signal_5859 ;
    wire signal_5860 ;
    wire signal_5861 ;
    wire signal_5862 ;
    wire signal_5863 ;
    wire signal_5864 ;
    wire signal_5865 ;
    wire signal_5866 ;
    wire signal_5867 ;
    wire signal_5868 ;
    wire signal_5869 ;
    wire signal_5870 ;
    wire signal_5871 ;
    wire signal_5872 ;
    wire signal_5873 ;
    wire signal_5874 ;
    wire signal_5875 ;
    wire signal_5876 ;
    wire signal_5877 ;
    wire signal_5878 ;
    wire signal_5879 ;
    wire signal_5880 ;
    wire signal_5881 ;
    wire signal_5882 ;
    wire signal_5883 ;
    wire signal_5884 ;
    wire signal_5885 ;
    wire signal_5886 ;
    wire signal_5887 ;
    wire signal_5888 ;
    wire signal_5889 ;
    wire signal_5890 ;
    wire signal_5891 ;
    wire signal_5892 ;
    wire signal_5893 ;
    wire signal_5894 ;
    wire signal_5895 ;
    wire signal_5896 ;
    wire signal_5897 ;
    wire signal_5898 ;
    wire signal_5899 ;
    wire signal_5900 ;
    wire signal_5901 ;
    wire signal_5902 ;
    wire signal_5903 ;
    wire signal_5904 ;
    wire signal_5905 ;
    wire signal_5906 ;
    wire signal_5907 ;
    wire signal_5908 ;
    wire signal_5909 ;
    wire signal_5910 ;
    wire signal_5911 ;
    wire signal_5912 ;
    wire signal_5913 ;
    wire signal_5914 ;
    wire signal_5915 ;
    wire signal_5916 ;
    wire signal_5917 ;
    wire signal_5918 ;
    wire signal_5919 ;
    wire signal_5920 ;
    wire signal_5921 ;
    wire signal_5922 ;
    wire signal_5923 ;
    wire signal_5924 ;
    wire signal_5925 ;
    wire signal_5926 ;
    wire signal_5927 ;
    wire signal_5928 ;
    wire signal_5929 ;
    wire signal_5930 ;
    wire signal_5931 ;
    wire signal_5932 ;
    wire signal_5933 ;
    wire signal_5934 ;
    wire signal_5935 ;
    wire signal_5936 ;
    wire signal_5937 ;
    wire signal_5938 ;
    wire signal_5939 ;
    wire signal_5940 ;
    wire signal_5941 ;
    wire signal_5942 ;
    wire signal_5943 ;
    wire signal_5944 ;
    wire signal_5945 ;
    wire signal_5946 ;
    wire signal_5947 ;
    wire signal_5948 ;
    wire signal_5949 ;
    wire signal_5950 ;
    wire signal_5951 ;
    wire signal_5952 ;
    wire signal_5953 ;
    wire signal_5954 ;
    wire signal_5955 ;
    wire signal_5956 ;
    wire signal_5957 ;
    wire signal_5958 ;
    wire signal_5959 ;
    wire signal_5960 ;
    wire signal_5961 ;
    wire signal_5962 ;
    wire signal_5963 ;
    wire signal_5964 ;
    wire signal_5965 ;
    wire signal_5966 ;
    wire signal_5967 ;
    wire signal_5968 ;
    wire signal_5969 ;
    wire signal_5970 ;
    wire signal_5971 ;
    wire signal_5972 ;
    wire signal_5973 ;
    wire signal_5974 ;
    wire signal_5975 ;
    wire signal_5976 ;
    wire signal_5977 ;
    wire signal_5978 ;
    wire signal_5979 ;
    wire signal_5980 ;
    wire signal_5981 ;
    wire signal_5982 ;
    wire signal_5983 ;
    wire signal_5984 ;
    wire signal_5985 ;
    wire signal_5986 ;
    wire signal_5987 ;
    wire signal_5988 ;
    wire signal_5989 ;
    wire signal_5990 ;
    wire signal_5991 ;
    wire signal_5992 ;
    wire signal_5993 ;
    wire signal_5994 ;
    wire signal_5995 ;
    wire signal_5996 ;
    wire signal_5997 ;
    wire signal_5998 ;
    wire signal_5999 ;
    wire signal_6000 ;
    wire signal_6001 ;
    wire signal_6002 ;
    wire signal_6003 ;
    wire signal_6004 ;
    wire signal_6005 ;
    wire signal_6006 ;
    wire signal_6007 ;
    wire signal_6008 ;
    wire signal_6009 ;
    wire signal_6010 ;
    wire signal_6011 ;
    wire signal_6012 ;
    wire signal_6013 ;
    wire signal_6014 ;
    wire signal_6015 ;
    wire signal_6016 ;
    wire signal_6017 ;
    wire signal_6018 ;
    wire signal_6019 ;
    wire signal_6020 ;
    wire signal_6021 ;
    wire signal_6022 ;
    wire signal_6023 ;
    wire signal_6024 ;
    wire signal_6025 ;
    wire signal_6026 ;
    wire signal_6027 ;
    wire signal_6028 ;
    wire signal_6029 ;
    wire signal_6030 ;
    wire signal_6031 ;
    wire signal_6032 ;
    wire signal_6033 ;
    wire signal_6034 ;
    wire signal_6035 ;
    wire signal_6036 ;
    wire signal_6037 ;
    wire signal_6038 ;
    wire signal_6039 ;
    wire signal_6040 ;
    wire signal_6041 ;
    wire signal_6042 ;
    wire signal_6043 ;
    wire signal_6044 ;
    wire signal_6045 ;
    wire signal_6046 ;
    wire signal_6047 ;
    wire signal_6048 ;
    wire signal_6049 ;
    wire signal_6050 ;
    wire signal_6051 ;
    wire signal_6052 ;
    wire signal_6053 ;
    wire signal_6054 ;
    wire signal_6055 ;
    wire signal_6056 ;
    wire signal_6057 ;
    wire signal_6058 ;
    wire signal_6059 ;
    wire signal_6060 ;
    wire signal_6061 ;
    wire signal_6062 ;
    wire signal_6063 ;
    wire signal_6064 ;
    wire signal_6065 ;
    wire signal_6066 ;
    wire signal_6067 ;
    wire signal_6068 ;
    wire signal_6069 ;
    wire signal_6070 ;
    wire signal_6071 ;
    wire signal_6072 ;
    wire signal_6073 ;
    wire signal_6074 ;
    wire signal_6075 ;
    wire signal_6076 ;
    wire signal_6077 ;
    wire signal_6078 ;
    wire signal_6079 ;
    wire signal_6080 ;
    wire signal_6081 ;
    wire signal_6082 ;
    wire signal_6083 ;
    wire signal_6084 ;
    wire signal_6085 ;
    wire signal_6086 ;
    wire signal_6087 ;
    wire signal_6088 ;
    wire signal_6089 ;
    wire signal_6090 ;
    wire signal_6091 ;
    wire signal_6092 ;
    wire signal_6093 ;
    wire signal_6094 ;
    wire signal_6095 ;
    wire signal_6096 ;
    wire signal_6097 ;
    wire signal_6098 ;
    wire signal_6099 ;
    wire signal_6100 ;
    wire signal_6101 ;
    wire signal_6102 ;
    wire signal_6103 ;
    wire signal_6104 ;
    wire signal_6105 ;
    wire signal_6106 ;
    wire signal_6107 ;
    wire signal_6108 ;
    wire signal_6109 ;
    wire signal_6110 ;
    wire signal_6111 ;
    wire signal_6112 ;
    wire signal_6113 ;
    wire signal_6114 ;
    wire signal_6115 ;
    wire signal_6116 ;
    wire signal_6117 ;
    wire signal_6118 ;
    wire signal_6119 ;
    wire signal_6120 ;
    wire signal_6121 ;
    wire signal_6122 ;
    wire signal_6123 ;
    wire signal_6124 ;
    wire signal_6125 ;
    wire signal_6126 ;
    wire signal_6127 ;
    wire signal_6128 ;
    wire signal_6129 ;
    wire signal_6130 ;
    wire signal_6131 ;
    wire signal_6132 ;
    wire signal_6133 ;
    wire signal_6134 ;
    wire signal_6135 ;
    wire signal_6136 ;
    wire signal_6137 ;
    wire signal_6138 ;
    wire signal_6139 ;
    wire signal_6140 ;
    wire signal_6141 ;
    wire signal_6142 ;
    wire signal_6143 ;
    wire signal_6144 ;
    wire signal_6145 ;
    wire signal_6146 ;
    wire signal_6147 ;
    wire signal_6148 ;
    wire signal_6149 ;
    wire signal_6150 ;
    wire signal_6151 ;
    wire signal_6152 ;
    wire signal_6153 ;
    wire signal_6154 ;
    wire signal_6155 ;
    wire signal_6156 ;
    wire signal_6157 ;
    wire signal_6158 ;
    wire signal_6159 ;
    wire signal_6160 ;
    wire signal_6161 ;
    wire signal_6162 ;
    wire signal_6163 ;
    wire signal_6164 ;
    wire signal_6165 ;
    wire signal_6166 ;
    wire signal_6167 ;
    wire signal_6168 ;
    wire signal_6169 ;
    wire signal_6170 ;
    wire signal_6171 ;
    wire signal_6172 ;
    wire signal_6173 ;
    wire signal_6174 ;
    wire signal_6175 ;
    wire signal_6176 ;
    wire signal_6177 ;
    wire signal_6178 ;
    wire signal_6179 ;
    wire signal_6180 ;
    wire signal_6181 ;
    wire signal_6182 ;
    wire signal_6183 ;
    wire signal_6184 ;
    wire signal_6185 ;
    wire signal_6186 ;
    wire signal_6187 ;
    wire signal_6188 ;
    wire signal_6189 ;
    wire signal_6190 ;
    wire signal_6191 ;
    wire signal_6192 ;
    wire signal_6193 ;
    wire signal_6194 ;
    wire signal_6195 ;
    wire signal_6196 ;
    wire signal_6197 ;
    wire signal_6198 ;
    wire signal_6199 ;
    wire signal_6200 ;
    wire signal_6201 ;
    wire signal_6202 ;
    wire signal_6203 ;
    wire signal_6204 ;
    wire signal_6205 ;
    wire signal_6206 ;
    wire signal_6207 ;
    wire signal_6208 ;
    wire signal_6209 ;
    wire signal_6210 ;
    wire signal_6211 ;
    wire signal_6212 ;
    wire signal_6213 ;
    wire signal_6214 ;
    wire signal_6215 ;
    wire signal_6216 ;
    wire signal_6217 ;
    wire signal_6218 ;
    wire signal_6219 ;
    wire signal_6220 ;
    wire signal_6221 ;
    wire signal_6222 ;
    wire signal_6223 ;
    wire signal_6224 ;
    wire signal_6225 ;
    wire signal_6226 ;
    wire signal_6227 ;
    wire signal_6228 ;
    wire signal_6229 ;
    wire signal_6230 ;
    wire signal_6231 ;
    wire signal_6232 ;
    wire signal_6233 ;
    wire signal_6234 ;
    wire signal_6235 ;
    wire signal_6236 ;
    wire signal_6237 ;
    wire signal_6238 ;
    wire signal_6239 ;
    wire signal_6240 ;
    wire signal_6241 ;
    wire signal_6242 ;
    wire signal_6243 ;
    wire signal_6244 ;
    wire signal_6245 ;
    wire signal_6246 ;
    wire signal_6247 ;
    wire signal_6248 ;
    wire signal_6249 ;
    wire signal_6250 ;
    wire signal_6251 ;
    wire signal_6252 ;
    wire signal_6253 ;
    wire signal_6254 ;
    wire signal_6255 ;
    wire signal_6256 ;
    wire signal_6257 ;
    wire signal_6258 ;
    wire signal_6259 ;
    wire signal_6260 ;
    wire signal_6261 ;
    wire signal_6262 ;
    wire signal_6263 ;
    wire signal_6264 ;
    wire signal_6265 ;
    wire signal_6266 ;
    wire signal_6267 ;
    wire signal_6268 ;
    wire signal_6269 ;
    wire signal_6270 ;
    wire signal_6271 ;
    wire signal_6272 ;
    wire signal_6273 ;
    wire signal_6274 ;
    wire signal_6275 ;
    wire signal_6276 ;
    wire signal_6277 ;
    wire signal_6278 ;
    wire signal_6279 ;
    wire signal_6280 ;
    wire signal_6281 ;
    wire signal_6282 ;
    wire signal_6283 ;
    wire signal_6284 ;
    wire signal_6285 ;
    wire signal_6286 ;
    wire signal_6287 ;
    wire signal_6288 ;
    wire signal_6289 ;
    wire signal_6290 ;
    wire signal_6291 ;
    wire signal_6292 ;
    wire signal_6293 ;
    wire signal_6294 ;
    wire signal_6295 ;
    wire signal_6296 ;
    wire signal_6297 ;
    wire signal_6298 ;
    wire signal_6299 ;
    wire signal_6300 ;
    wire signal_6301 ;
    wire signal_6302 ;
    wire signal_6303 ;
    wire signal_6304 ;
    wire signal_6305 ;
    wire signal_6306 ;
    wire signal_6307 ;
    wire signal_6308 ;
    wire signal_6309 ;
    wire signal_6310 ;
    wire signal_6311 ;
    wire signal_6312 ;
    wire signal_6313 ;
    wire signal_6314 ;
    wire signal_6315 ;
    wire signal_6316 ;
    wire signal_6317 ;
    wire signal_6318 ;
    wire signal_6319 ;
    wire signal_6320 ;
    wire signal_6321 ;
    wire signal_6322 ;
    wire signal_6323 ;
    wire signal_6324 ;
    wire signal_6325 ;
    wire signal_6326 ;
    wire signal_6327 ;
    wire signal_6328 ;
    wire signal_6329 ;
    wire signal_6330 ;
    wire signal_6331 ;
    wire signal_6332 ;
    wire signal_6333 ;
    wire signal_6334 ;
    wire signal_6335 ;
    wire signal_6336 ;
    wire signal_6337 ;
    wire signal_6338 ;
    wire signal_6339 ;
    wire signal_6340 ;
    wire signal_6341 ;
    wire signal_6342 ;
    wire signal_6343 ;
    wire signal_6344 ;
    wire signal_6345 ;
    wire signal_6346 ;
    wire signal_6347 ;
    wire signal_6348 ;
    wire signal_6349 ;
    wire signal_6350 ;
    wire signal_6351 ;
    wire signal_6352 ;
    wire signal_6353 ;
    wire signal_6354 ;
    wire signal_6355 ;
    wire signal_6356 ;
    wire signal_6357 ;
    wire signal_6358 ;
    wire signal_6359 ;
    wire signal_6360 ;
    wire signal_6361 ;
    wire signal_6362 ;
    wire signal_6363 ;
    wire signal_6364 ;
    wire signal_6365 ;
    wire signal_6366 ;
    wire signal_6367 ;
    wire signal_6368 ;
    wire signal_6369 ;
    wire signal_6370 ;
    wire signal_6371 ;
    wire signal_6372 ;
    wire signal_6373 ;
    wire signal_6374 ;
    wire signal_6375 ;
    wire signal_6376 ;
    wire signal_6377 ;
    wire signal_6378 ;
    wire signal_6379 ;
    wire signal_6380 ;
    wire signal_6381 ;
    wire signal_6382 ;
    wire signal_6383 ;
    wire signal_6384 ;
    wire signal_6385 ;
    wire signal_6386 ;
    wire signal_6387 ;
    wire signal_6388 ;
    wire signal_6389 ;
    wire signal_6390 ;
    wire signal_6391 ;
    wire signal_6392 ;
    wire signal_6393 ;
    wire signal_6394 ;
    wire signal_6395 ;
    wire signal_6396 ;
    wire signal_6397 ;
    wire signal_6398 ;
    wire signal_6399 ;
    wire signal_6400 ;
    wire signal_6401 ;
    wire signal_6402 ;
    wire signal_6403 ;
    wire signal_6404 ;
    wire signal_6405 ;
    wire signal_6406 ;
    wire signal_6407 ;
    wire signal_6408 ;
    wire signal_6409 ;
    wire signal_6410 ;
    wire signal_6411 ;
    wire signal_6412 ;
    wire signal_6413 ;
    wire signal_6414 ;
    wire signal_6415 ;
    wire signal_6416 ;
    wire signal_6417 ;
    wire signal_6418 ;
    wire signal_6419 ;
    wire signal_6420 ;
    wire signal_6421 ;
    wire signal_6422 ;
    wire signal_6423 ;
    wire signal_6424 ;
    wire signal_6425 ;
    wire signal_6426 ;
    wire signal_6427 ;
    wire signal_6428 ;
    wire signal_6429 ;
    wire signal_6430 ;
    wire signal_6431 ;
    wire signal_6432 ;
    wire signal_6433 ;
    wire signal_6434 ;
    wire signal_6435 ;
    wire signal_6436 ;
    wire signal_6437 ;
    wire signal_6438 ;
    wire signal_6439 ;
    wire signal_6440 ;
    wire signal_6441 ;
    wire signal_6442 ;
    wire signal_6443 ;
    wire signal_6444 ;
    wire signal_6445 ;
    wire signal_6446 ;
    wire signal_6447 ;
    wire signal_6448 ;
    wire signal_6449 ;
    wire signal_6450 ;
    wire signal_6451 ;
    wire signal_6452 ;
    wire signal_6453 ;
    wire signal_6454 ;
    wire signal_6455 ;
    wire signal_6456 ;
    wire signal_6457 ;
    wire signal_6458 ;
    wire signal_6459 ;
    wire signal_6460 ;
    wire signal_6461 ;
    wire signal_6462 ;
    wire signal_6463 ;
    wire signal_6464 ;
    wire signal_6465 ;
    wire signal_6466 ;
    wire signal_6467 ;
    wire signal_6468 ;
    wire signal_6469 ;
    wire signal_6470 ;
    wire signal_6471 ;
    wire signal_6472 ;
    wire signal_6473 ;
    wire signal_6474 ;
    wire signal_6475 ;
    wire signal_6476 ;
    wire signal_6477 ;
    wire signal_6478 ;
    wire signal_6479 ;
    wire signal_6480 ;
    wire signal_6481 ;
    wire signal_6482 ;
    wire signal_6483 ;
    wire signal_6484 ;
    wire signal_6485 ;
    wire signal_6486 ;
    wire signal_6487 ;
    wire signal_6488 ;
    wire signal_6489 ;
    wire signal_6490 ;
    wire signal_6491 ;
    wire signal_6492 ;
    wire signal_6493 ;
    wire signal_6494 ;
    wire signal_6495 ;
    wire signal_6496 ;
    wire signal_6497 ;
    wire signal_6498 ;
    wire signal_6499 ;
    wire signal_6500 ;
    wire signal_6501 ;
    wire signal_6502 ;
    wire signal_6503 ;
    wire signal_6504 ;
    wire signal_6505 ;
    wire signal_6506 ;
    wire signal_6507 ;
    wire signal_6508 ;
    wire signal_6509 ;
    wire signal_6510 ;
    wire signal_6511 ;
    wire signal_6512 ;
    wire signal_6513 ;
    wire signal_6514 ;
    wire signal_6515 ;
    wire signal_6516 ;
    wire signal_6517 ;
    wire signal_6518 ;
    wire signal_6519 ;
    wire signal_6520 ;
    wire signal_6521 ;
    wire signal_6522 ;
    wire signal_6523 ;
    wire signal_6524 ;
    wire signal_6525 ;
    wire signal_6526 ;
    wire signal_6527 ;
    wire signal_6528 ;
    wire signal_6529 ;
    wire signal_6530 ;
    wire signal_6531 ;
    wire signal_6532 ;
    wire signal_6533 ;
    wire signal_6534 ;
    wire signal_6535 ;
    wire signal_6536 ;
    wire signal_6537 ;
    wire signal_6538 ;
    wire signal_6539 ;
    wire signal_6540 ;
    wire signal_6541 ;
    wire signal_6542 ;
    wire signal_6543 ;
    wire signal_6544 ;
    wire signal_6545 ;
    wire signal_6546 ;
    wire signal_6547 ;
    wire signal_6548 ;
    wire signal_6549 ;
    wire signal_6550 ;
    wire signal_6551 ;
    wire signal_6552 ;
    wire signal_6553 ;
    wire signal_6554 ;
    wire signal_6555 ;
    wire signal_6556 ;
    wire signal_6557 ;
    wire signal_6558 ;
    wire signal_6559 ;
    wire signal_6560 ;
    wire signal_6561 ;
    wire signal_6562 ;
    wire signal_6563 ;
    wire signal_6564 ;
    wire signal_6565 ;
    wire signal_6566 ;
    wire signal_6567 ;
    wire signal_6568 ;
    wire signal_6569 ;
    wire signal_6570 ;
    wire signal_6571 ;
    wire signal_6572 ;
    wire signal_6573 ;
    wire signal_6574 ;
    wire signal_6575 ;
    wire signal_6576 ;
    wire signal_6577 ;
    wire signal_6578 ;
    wire signal_6579 ;
    wire signal_6580 ;
    wire signal_6581 ;
    wire signal_6582 ;
    wire signal_6583 ;
    wire signal_6584 ;
    wire signal_6585 ;
    wire signal_6586 ;
    wire signal_6587 ;
    wire signal_6588 ;
    wire signal_6589 ;
    wire signal_6590 ;
    wire signal_6591 ;
    wire signal_6592 ;
    wire signal_6593 ;
    wire signal_6594 ;
    wire signal_6595 ;
    wire signal_6596 ;
    wire signal_6597 ;
    wire signal_6598 ;
    wire signal_6599 ;
    wire signal_6600 ;
    wire signal_6601 ;
    wire signal_6602 ;
    wire signal_6603 ;
    wire signal_6604 ;
    wire signal_6605 ;
    wire signal_6606 ;
    wire signal_6607 ;
    wire signal_6608 ;
    wire signal_6609 ;
    wire signal_6610 ;
    wire signal_6611 ;
    wire signal_6612 ;
    wire signal_6613 ;
    wire signal_6614 ;
    wire signal_6615 ;
    wire signal_6616 ;
    wire signal_6617 ;
    wire signal_6618 ;
    wire signal_6619 ;
    wire signal_6620 ;
    wire signal_6621 ;
    wire signal_6622 ;
    wire signal_6623 ;
    wire signal_6624 ;
    wire signal_6625 ;
    wire signal_6626 ;
    wire signal_6627 ;
    wire signal_6628 ;
    wire signal_6629 ;
    wire signal_6630 ;
    wire signal_6631 ;
    wire signal_6632 ;
    wire signal_6633 ;
    wire signal_6634 ;
    wire signal_6635 ;
    wire signal_6636 ;
    wire signal_6637 ;
    wire signal_6638 ;
    wire signal_6639 ;
    wire signal_6640 ;
    wire signal_6641 ;
    wire signal_6642 ;
    wire signal_6643 ;
    wire signal_6644 ;
    wire signal_6645 ;
    wire signal_6646 ;
    wire signal_6647 ;
    wire signal_6648 ;
    wire signal_6649 ;
    wire signal_6650 ;
    wire signal_6651 ;
    wire signal_6652 ;
    wire signal_6653 ;
    wire signal_6654 ;
    wire signal_6655 ;
    wire signal_6656 ;
    wire signal_6657 ;
    wire signal_6658 ;
    wire signal_6659 ;
    wire signal_6660 ;
    wire signal_6661 ;
    wire signal_6662 ;
    wire signal_6663 ;
    wire signal_6664 ;
    wire signal_6665 ;
    wire signal_6666 ;
    wire signal_6667 ;
    wire signal_6668 ;
    wire signal_6669 ;
    wire signal_6670 ;
    wire signal_6671 ;
    wire signal_6672 ;
    wire signal_6673 ;
    wire signal_6674 ;
    wire signal_6675 ;
    wire signal_6676 ;
    wire signal_6677 ;
    wire signal_6678 ;
    wire signal_6679 ;
    wire signal_6680 ;
    wire signal_6681 ;
    wire signal_6682 ;
    wire signal_6683 ;
    wire signal_6684 ;
    wire signal_6685 ;
    wire signal_6686 ;
    wire signal_6687 ;
    wire signal_6688 ;
    wire signal_6689 ;
    wire signal_6690 ;
    wire signal_6691 ;
    wire signal_6692 ;
    wire signal_6693 ;
    wire signal_6694 ;
    wire signal_6695 ;
    wire signal_6696 ;
    wire signal_6697 ;
    wire signal_6698 ;
    wire signal_6699 ;
    wire signal_6700 ;
    wire signal_6701 ;
    wire signal_6702 ;
    wire signal_6703 ;
    wire signal_6704 ;
    wire signal_6705 ;
    wire signal_6706 ;
    wire signal_6707 ;
    wire signal_6708 ;
    wire signal_6709 ;
    wire signal_6710 ;
    wire signal_6711 ;
    wire signal_6712 ;
    wire signal_6713 ;
    wire signal_6714 ;
    wire signal_6715 ;
    wire signal_6716 ;
    wire signal_6717 ;
    wire signal_6718 ;
    wire signal_6719 ;
    wire signal_6720 ;
    wire signal_6721 ;
    wire signal_6722 ;
    wire signal_6723 ;
    wire signal_6724 ;
    wire signal_6725 ;
    wire signal_6726 ;
    wire signal_6727 ;
    wire signal_6728 ;
    wire signal_6729 ;
    wire signal_6730 ;
    wire signal_6731 ;
    wire signal_6732 ;
    wire signal_6733 ;
    wire signal_6734 ;
    wire signal_6735 ;
    wire signal_6736 ;
    wire signal_6737 ;
    wire signal_6738 ;
    wire signal_6739 ;
    wire signal_6740 ;
    wire signal_6741 ;
    wire signal_6742 ;
    wire signal_6743 ;
    wire signal_6744 ;
    wire signal_6745 ;
    wire signal_6746 ;
    wire signal_6747 ;
    wire signal_6748 ;
    wire signal_6749 ;
    wire signal_6750 ;
    wire signal_6751 ;
    wire signal_6752 ;
    wire signal_6753 ;
    wire signal_6754 ;
    wire signal_6755 ;
    wire signal_6756 ;
    wire signal_6757 ;
    wire signal_6758 ;
    wire signal_6759 ;
    wire signal_6760 ;
    wire signal_6761 ;
    wire signal_6762 ;
    wire signal_6763 ;
    wire signal_6764 ;
    wire signal_6765 ;
    wire signal_6766 ;
    wire signal_6767 ;
    wire signal_6768 ;
    wire signal_6769 ;
    wire signal_6770 ;
    wire signal_6771 ;
    wire signal_6772 ;
    wire signal_6773 ;
    wire signal_6774 ;
    wire signal_6775 ;
    wire signal_6776 ;
    wire signal_6777 ;
    wire signal_6778 ;
    wire signal_6779 ;
    wire signal_6780 ;
    wire signal_6781 ;
    wire signal_6782 ;
    wire signal_6783 ;
    wire signal_6784 ;
    wire signal_6785 ;
    wire signal_6786 ;
    wire signal_6787 ;
    wire signal_6788 ;
    wire signal_6789 ;
    wire signal_6790 ;
    wire signal_6791 ;
    wire signal_6792 ;
    wire signal_6793 ;
    wire signal_6794 ;
    wire signal_6795 ;
    wire signal_6796 ;
    wire signal_6797 ;
    wire signal_6798 ;
    wire signal_6799 ;
    wire signal_6800 ;
    wire signal_6801 ;
    wire signal_6802 ;
    wire signal_6803 ;
    wire signal_6804 ;
    wire signal_6805 ;
    wire signal_6806 ;
    wire signal_6807 ;
    wire signal_6808 ;
    wire signal_6809 ;
    wire signal_6810 ;
    wire signal_6811 ;
    wire signal_6812 ;
    wire signal_6813 ;
    wire signal_6814 ;
    wire signal_6815 ;
    wire signal_6816 ;
    wire signal_6817 ;
    wire signal_6818 ;
    wire signal_6819 ;
    wire signal_6820 ;
    wire signal_6821 ;
    wire signal_6822 ;
    wire signal_6823 ;
    wire signal_6824 ;
    wire signal_6825 ;
    wire signal_6826 ;
    wire signal_6827 ;
    wire signal_6828 ;
    wire signal_6829 ;
    wire signal_6830 ;
    wire signal_6831 ;
    wire signal_6832 ;
    wire signal_6833 ;
    wire signal_6834 ;
    wire signal_6835 ;
    wire signal_6836 ;
    wire signal_6837 ;
    wire signal_6838 ;
    wire signal_6839 ;
    wire signal_6840 ;
    wire signal_6841 ;
    wire signal_6842 ;
    wire signal_6843 ;
    wire signal_6844 ;
    wire signal_6845 ;
    wire signal_6846 ;
    wire signal_6847 ;
    wire signal_6848 ;
    wire signal_6849 ;
    wire signal_6850 ;
    wire signal_6851 ;
    wire signal_6852 ;
    wire signal_6853 ;
    wire signal_6854 ;
    wire signal_6855 ;
    wire signal_6856 ;
    wire signal_6857 ;
    wire signal_6858 ;
    wire signal_6859 ;
    wire signal_6860 ;
    wire signal_6861 ;
    wire signal_6862 ;
    wire signal_6863 ;
    wire signal_6864 ;
    wire signal_6865 ;
    wire signal_6866 ;
    wire signal_6867 ;
    wire signal_6868 ;
    wire signal_6869 ;
    wire signal_6870 ;
    wire signal_6871 ;
    wire signal_6872 ;
    wire signal_6873 ;
    wire signal_6874 ;
    wire signal_6875 ;
    wire signal_6876 ;
    wire signal_6877 ;
    wire signal_6878 ;
    wire signal_6879 ;
    wire signal_6880 ;
    wire signal_6881 ;
    wire signal_6882 ;
    wire signal_6883 ;
    wire signal_6884 ;
    wire signal_6885 ;
    wire signal_6886 ;
    wire signal_6887 ;
    wire signal_6888 ;
    wire signal_6889 ;
    wire signal_6890 ;
    wire signal_6891 ;
    wire signal_6892 ;
    wire signal_6893 ;
    wire signal_6894 ;
    wire signal_6895 ;
    wire signal_6896 ;
    wire signal_6897 ;
    wire signal_6898 ;
    wire signal_6899 ;
    wire signal_6900 ;
    wire signal_6901 ;
    wire signal_6902 ;
    wire signal_6903 ;
    wire signal_6904 ;
    wire signal_6905 ;
    wire signal_6906 ;
    wire signal_6907 ;
    wire signal_6908 ;
    wire signal_6909 ;
    wire signal_6910 ;
    wire signal_6911 ;
    wire signal_6912 ;
    wire signal_6913 ;
    wire signal_6914 ;
    wire signal_6915 ;
    wire signal_6916 ;
    wire signal_6917 ;
    wire signal_6918 ;
    wire signal_6919 ;
    wire signal_6920 ;
    wire signal_6921 ;
    wire signal_6922 ;
    wire signal_6923 ;
    wire signal_6924 ;
    wire signal_6925 ;
    wire signal_6926 ;
    wire signal_6927 ;
    wire signal_6928 ;
    wire signal_6929 ;
    wire signal_6930 ;
    wire signal_6931 ;
    wire signal_6932 ;
    wire signal_6933 ;
    wire signal_6934 ;
    wire signal_6935 ;
    wire signal_6936 ;
    wire signal_6937 ;
    wire signal_6938 ;
    wire signal_6939 ;
    wire signal_6940 ;
    wire signal_6941 ;
    wire signal_6942 ;
    wire signal_6943 ;
    wire signal_6944 ;
    wire signal_6945 ;
    wire signal_6946 ;
    wire signal_6947 ;
    wire signal_6948 ;
    wire signal_6949 ;
    wire signal_6950 ;
    wire signal_6951 ;
    wire signal_6952 ;
    wire signal_6953 ;
    wire signal_6954 ;
    wire signal_6955 ;
    wire signal_6956 ;
    wire signal_6957 ;
    wire signal_6958 ;
    wire signal_6959 ;
    wire signal_6960 ;
    wire signal_6961 ;
    wire signal_6962 ;
    wire signal_6963 ;
    wire signal_6964 ;
    wire signal_6965 ;
    wire signal_6966 ;
    wire signal_6967 ;
    wire signal_6968 ;
    wire signal_6969 ;
    wire signal_6970 ;
    wire signal_6971 ;
    wire signal_6972 ;
    wire signal_6973 ;
    wire signal_6974 ;
    wire signal_6975 ;
    wire signal_6976 ;
    wire signal_6977 ;
    wire signal_6978 ;
    wire signal_6979 ;
    wire signal_6980 ;
    wire signal_6981 ;
    wire signal_6982 ;
    wire signal_6983 ;
    wire signal_6984 ;
    wire signal_6985 ;
    wire signal_6986 ;
    wire signal_6987 ;
    wire signal_6988 ;
    wire signal_6989 ;
    wire signal_6990 ;
    wire signal_6991 ;
    wire signal_6992 ;
    wire signal_6993 ;
    wire signal_6994 ;
    wire signal_6995 ;
    wire signal_6996 ;
    wire signal_6997 ;
    wire signal_6998 ;
    wire signal_6999 ;
    wire signal_7000 ;
    wire signal_7001 ;
    wire signal_7002 ;
    wire signal_7003 ;
    wire signal_7004 ;
    wire signal_7005 ;
    wire signal_7006 ;
    wire signal_7007 ;
    wire signal_7008 ;
    wire signal_7009 ;
    wire signal_7010 ;
    wire signal_7011 ;
    wire signal_7012 ;
    wire signal_7013 ;
    wire signal_7014 ;
    wire signal_7015 ;
    wire signal_7016 ;
    wire signal_7017 ;
    wire signal_7018 ;
    wire signal_7019 ;
    wire signal_7020 ;
    wire signal_7021 ;
    wire signal_7022 ;
    wire signal_7023 ;
    wire signal_7024 ;
    wire signal_7025 ;
    wire signal_7026 ;
    wire signal_7027 ;
    wire signal_7028 ;
    wire signal_7029 ;
    wire signal_7030 ;
    wire signal_7031 ;
    wire signal_7032 ;
    wire signal_7033 ;
    wire signal_7034 ;
    wire signal_7035 ;
    wire signal_7036 ;
    wire signal_7037 ;
    wire signal_7038 ;
    wire signal_7039 ;
    wire signal_7040 ;
    wire signal_7041 ;
    wire signal_7042 ;
    wire signal_7043 ;
    wire signal_7044 ;
    wire signal_7045 ;
    wire signal_7046 ;
    wire signal_7047 ;
    wire signal_7048 ;
    wire signal_7049 ;
    wire signal_7050 ;
    wire signal_7051 ;
    wire signal_7052 ;
    wire signal_7053 ;
    wire signal_7054 ;
    wire signal_7055 ;
    wire signal_7056 ;
    wire signal_7057 ;
    wire signal_7058 ;
    wire signal_7059 ;
    wire signal_7060 ;
    wire signal_7061 ;
    wire signal_7062 ;
    wire signal_7063 ;
    wire signal_7064 ;
    wire signal_7065 ;
    wire signal_7066 ;
    wire signal_7067 ;
    wire signal_7068 ;
    wire signal_7069 ;
    wire signal_7070 ;
    wire signal_7071 ;
    wire signal_7072 ;
    wire signal_7073 ;
    wire signal_7074 ;
    wire signal_7075 ;
    wire signal_7076 ;
    wire signal_7077 ;
    wire signal_7078 ;
    wire signal_7079 ;
    wire signal_7080 ;
    wire signal_7081 ;
    wire signal_7082 ;
    wire signal_7083 ;
    wire signal_7084 ;
    wire signal_7085 ;
    wire signal_7086 ;
    wire signal_7087 ;
    wire signal_7088 ;
    wire signal_7089 ;
    wire signal_7090 ;
    wire signal_7091 ;
    wire signal_7092 ;
    wire signal_7093 ;
    wire signal_7094 ;
    wire signal_7095 ;
    wire signal_7096 ;
    wire signal_7097 ;
    wire signal_7098 ;
    wire signal_7099 ;
    wire signal_7100 ;
    wire signal_7101 ;
    wire signal_7102 ;
    wire signal_7103 ;
    wire signal_7104 ;
    wire signal_7105 ;
    wire signal_7106 ;
    wire signal_7107 ;
    wire signal_7108 ;
    wire signal_7109 ;
    wire signal_7110 ;
    wire signal_7111 ;
    wire signal_7112 ;
    wire signal_7113 ;
    wire signal_7114 ;
    wire signal_7115 ;
    wire signal_7116 ;
    wire signal_7117 ;
    wire signal_7118 ;
    wire signal_7119 ;
    wire signal_7120 ;
    wire signal_7121 ;
    wire signal_7122 ;
    wire signal_7123 ;
    wire signal_7124 ;
    wire signal_7125 ;
    wire signal_7126 ;
    wire signal_7127 ;
    wire signal_7128 ;
    wire signal_7129 ;
    wire signal_7130 ;
    wire signal_7131 ;
    wire signal_7132 ;
    wire signal_7133 ;
    wire signal_7134 ;
    wire signal_7135 ;
    wire signal_7136 ;
    wire signal_7137 ;
    wire signal_7138 ;
    wire signal_7139 ;
    wire signal_7140 ;
    wire signal_7141 ;
    wire signal_7142 ;
    wire signal_7143 ;
    wire signal_7144 ;
    wire signal_7145 ;
    wire signal_7146 ;
    wire signal_7147 ;
    wire signal_7148 ;
    wire signal_7149 ;
    wire signal_7150 ;
    wire signal_7151 ;
    wire signal_7152 ;
    wire signal_7153 ;
    wire signal_7154 ;
    wire signal_7155 ;
    wire signal_7156 ;
    wire signal_7157 ;
    wire signal_7158 ;
    wire signal_7159 ;
    wire signal_7160 ;
    wire signal_7161 ;
    wire signal_7162 ;
    wire signal_7163 ;
    wire signal_7164 ;
    wire signal_7165 ;
    wire signal_7166 ;
    wire signal_7167 ;
    wire signal_7168 ;
    wire signal_7169 ;
    wire signal_7170 ;
    wire signal_7171 ;
    wire signal_7172 ;
    wire signal_7173 ;
    wire signal_7174 ;
    wire signal_7175 ;
    wire signal_7176 ;
    wire signal_7177 ;
    wire signal_7178 ;
    wire signal_7179 ;
    wire signal_7180 ;
    wire signal_7181 ;
    wire signal_7182 ;
    wire signal_7183 ;
    wire signal_7184 ;
    wire signal_7185 ;
    wire signal_7186 ;
    wire signal_7187 ;
    wire signal_7188 ;
    wire signal_7189 ;
    wire signal_7190 ;
    wire signal_7191 ;
    wire signal_7192 ;
    wire signal_7193 ;
    wire signal_7194 ;
    wire signal_7195 ;
    wire signal_7196 ;
    wire signal_7197 ;
    wire signal_7198 ;
    wire signal_7199 ;
    wire signal_7200 ;
    wire signal_7201 ;
    wire signal_7202 ;
    wire signal_7203 ;
    wire signal_7204 ;
    wire signal_7205 ;
    wire signal_7206 ;
    wire signal_7207 ;
    wire signal_7208 ;
    wire signal_7209 ;
    wire signal_7210 ;
    wire signal_7211 ;
    wire signal_7212 ;
    wire signal_7213 ;
    wire signal_7214 ;
    wire signal_7215 ;
    wire signal_7216 ;
    wire signal_7217 ;
    wire signal_7218 ;
    wire signal_7219 ;
    wire signal_7220 ;
    wire signal_7221 ;
    wire signal_7222 ;
    wire signal_7223 ;
    wire signal_7224 ;
    wire signal_7225 ;
    wire signal_7226 ;
    wire signal_7227 ;
    wire signal_7228 ;
    wire signal_7229 ;
    wire signal_7230 ;
    wire signal_7231 ;
    wire signal_7232 ;
    wire signal_7233 ;
    wire signal_7234 ;
    wire signal_7235 ;
    wire signal_7236 ;
    wire signal_7237 ;
    wire signal_7238 ;
    wire signal_7239 ;
    wire signal_7240 ;
    wire signal_7241 ;
    wire signal_7242 ;
    wire signal_7243 ;
    wire signal_7244 ;
    wire signal_7245 ;
    wire signal_7246 ;
    wire signal_7247 ;
    wire signal_7248 ;
    wire signal_7249 ;
    wire signal_7250 ;
    wire signal_7251 ;
    wire signal_7252 ;
    wire signal_7253 ;
    wire signal_7254 ;
    wire signal_7255 ;
    wire signal_7256 ;
    wire signal_7257 ;
    wire signal_7258 ;
    wire signal_7259 ;
    wire signal_7260 ;
    wire signal_7261 ;
    wire signal_7262 ;
    wire signal_7263 ;
    wire signal_7264 ;
    wire signal_7265 ;
    wire signal_7266 ;
    wire signal_7267 ;
    wire signal_7268 ;
    wire signal_7269 ;
    wire signal_7270 ;
    wire signal_7271 ;
    wire signal_7272 ;
    wire signal_7273 ;
    wire signal_7274 ;
    wire signal_7275 ;
    wire signal_7276 ;
    wire signal_7277 ;
    wire signal_7278 ;
    wire signal_7279 ;
    wire signal_7280 ;
    wire signal_7281 ;
    wire signal_7282 ;
    wire signal_7283 ;
    wire signal_7284 ;
    wire signal_7285 ;
    wire signal_7286 ;
    wire signal_7287 ;
    wire signal_7288 ;
    wire signal_7289 ;
    wire signal_7290 ;
    wire signal_7291 ;
    wire signal_7292 ;
    wire signal_7293 ;
    wire signal_7294 ;
    wire signal_7295 ;
    wire signal_7296 ;
    wire signal_7297 ;
    wire signal_7298 ;
    wire signal_7299 ;
    wire signal_7300 ;
    wire signal_7301 ;
    wire signal_7302 ;
    wire signal_7303 ;
    wire signal_7304 ;
    wire signal_7305 ;
    wire signal_7306 ;
    wire signal_7307 ;
    wire signal_7308 ;
    wire signal_7309 ;
    wire signal_7310 ;
    wire signal_7311 ;
    wire signal_7312 ;
    wire signal_7313 ;
    wire signal_7314 ;
    wire signal_7315 ;
    wire signal_7316 ;
    wire signal_7317 ;
    wire signal_7318 ;
    wire signal_7319 ;
    wire signal_7320 ;
    wire signal_7321 ;
    wire signal_7322 ;
    wire signal_7323 ;
    wire signal_7324 ;
    wire signal_7325 ;
    wire signal_7326 ;
    wire signal_7327 ;
    wire signal_7328 ;
    wire signal_7329 ;
    wire signal_7330 ;
    wire signal_7331 ;
    wire signal_7332 ;
    wire signal_7333 ;
    wire signal_7334 ;
    wire signal_7335 ;
    wire signal_7336 ;
    wire signal_7337 ;
    wire signal_7338 ;
    wire signal_7339 ;
    wire signal_7340 ;
    wire signal_7341 ;
    wire signal_7342 ;
    wire signal_7343 ;
    wire signal_7344 ;
    wire signal_7345 ;
    wire signal_7346 ;
    wire signal_7347 ;
    wire signal_7348 ;
    wire signal_7349 ;
    wire signal_7350 ;
    wire signal_7351 ;
    wire signal_7352 ;
    wire signal_7353 ;
    wire signal_7354 ;
    wire signal_7355 ;
    wire signal_7356 ;
    wire signal_7357 ;
    wire signal_7358 ;
    wire signal_7359 ;
    wire signal_7360 ;
    wire signal_7361 ;
    wire signal_7362 ;
    wire signal_7363 ;
    wire signal_7364 ;
    wire signal_7365 ;
    wire signal_7366 ;
    wire signal_7367 ;
    wire signal_7368 ;
    wire signal_7369 ;
    wire signal_7370 ;
    wire signal_7371 ;
    wire signal_7372 ;
    wire signal_7373 ;
    wire signal_7374 ;
    wire signal_7375 ;
    wire signal_7376 ;
    wire signal_7377 ;
    wire signal_7378 ;
    wire signal_7379 ;
    wire signal_7380 ;
    wire signal_7381 ;
    wire signal_7382 ;
    wire signal_7383 ;
    wire signal_7384 ;
    wire signal_7385 ;
    wire signal_7386 ;
    wire signal_7387 ;
    wire signal_7388 ;
    wire signal_7389 ;
    wire signal_7390 ;
    wire signal_7391 ;
    wire signal_7392 ;
    wire signal_7393 ;
    wire signal_7394 ;
    wire signal_7395 ;
    wire signal_7396 ;
    wire signal_7397 ;
    wire signal_7398 ;
    wire signal_7399 ;
    wire signal_7400 ;
    wire signal_7401 ;
    wire signal_7402 ;
    wire signal_7403 ;
    wire signal_7404 ;
    wire signal_7405 ;
    wire signal_7406 ;
    wire signal_7407 ;
    wire signal_7408 ;
    wire signal_7409 ;
    wire signal_7410 ;
    wire signal_7411 ;
    wire signal_7412 ;
    wire signal_7413 ;
    wire signal_7414 ;
    wire signal_7415 ;
    wire signal_7416 ;
    wire signal_7417 ;
    wire signal_7418 ;
    wire signal_7419 ;
    wire signal_7420 ;
    wire signal_7421 ;
    wire signal_7422 ;
    wire signal_7423 ;
    wire signal_7424 ;
    wire signal_7425 ;
    wire signal_7426 ;
    wire signal_7427 ;
    wire signal_7428 ;
    wire signal_7429 ;
    wire signal_7430 ;
    wire signal_7431 ;
    wire signal_7432 ;
    wire signal_7433 ;
    wire signal_7434 ;
    wire signal_7435 ;
    wire signal_7436 ;
    wire signal_7437 ;
    wire signal_7438 ;
    wire signal_7439 ;
    wire signal_7440 ;
    wire signal_7441 ;
    wire signal_7442 ;
    wire signal_7443 ;
    wire signal_7444 ;
    wire signal_7445 ;
    wire signal_7446 ;
    wire signal_7447 ;
    wire signal_7448 ;
    wire signal_7449 ;
    wire signal_7450 ;
    wire signal_7451 ;
    wire signal_7452 ;
    wire signal_7453 ;
    wire signal_7454 ;
    wire signal_7455 ;
    wire signal_7456 ;
    wire signal_7457 ;
    wire signal_7458 ;
    wire signal_7459 ;
    wire signal_7460 ;
    wire signal_7461 ;
    wire signal_7462 ;
    wire signal_7463 ;
    wire signal_7464 ;
    wire signal_7465 ;
    wire signal_7466 ;
    wire signal_7467 ;
    wire signal_7468 ;
    wire signal_7469 ;
    wire signal_7470 ;
    wire signal_7471 ;
    wire signal_7472 ;
    wire signal_7473 ;
    wire signal_7474 ;
    wire signal_7475 ;
    wire signal_7476 ;
    wire signal_7477 ;
    wire signal_7478 ;
    wire signal_7479 ;
    wire signal_7480 ;
    wire signal_7481 ;
    wire signal_7482 ;
    wire signal_7483 ;
    wire signal_7484 ;
    wire signal_7485 ;
    wire signal_7486 ;
    wire signal_7487 ;
    wire signal_7488 ;
    wire signal_7489 ;
    wire signal_7490 ;
    wire signal_7491 ;
    wire signal_7492 ;
    wire signal_7493 ;
    wire signal_7494 ;
    wire signal_7495 ;
    wire signal_7496 ;
    wire signal_7497 ;
    wire signal_7498 ;
    wire signal_7499 ;
    wire signal_7500 ;
    wire signal_7501 ;
    wire signal_7502 ;
    wire signal_7503 ;
    wire signal_7504 ;
    wire signal_7505 ;
    wire signal_7506 ;
    wire signal_7507 ;
    wire signal_7508 ;
    wire signal_7509 ;
    wire signal_7510 ;
    wire signal_7511 ;
    wire signal_7512 ;
    wire signal_7513 ;
    wire signal_7514 ;
    wire signal_7515 ;
    wire signal_7516 ;
    wire signal_7517 ;
    wire signal_7518 ;
    wire signal_7519 ;
    wire signal_7520 ;
    wire signal_7521 ;
    wire signal_7522 ;
    wire signal_7523 ;
    wire signal_7524 ;
    wire signal_7525 ;
    wire signal_7526 ;
    wire signal_7527 ;
    wire signal_7528 ;
    wire signal_7529 ;
    wire signal_7530 ;
    wire signal_7531 ;
    wire signal_7532 ;
    wire signal_7533 ;
    wire signal_7534 ;
    wire signal_7535 ;
    wire signal_7536 ;
    wire signal_7537 ;
    wire signal_7538 ;
    wire signal_7539 ;
    wire signal_7540 ;
    wire signal_7541 ;
    wire signal_7542 ;
    wire signal_7543 ;
    wire signal_7544 ;
    wire signal_7545 ;
    wire signal_7546 ;
    wire signal_7547 ;
    wire signal_7548 ;
    wire signal_7549 ;
    wire signal_7550 ;
    wire signal_7551 ;
    wire signal_7552 ;
    wire signal_7553 ;
    wire signal_7554 ;
    wire signal_7555 ;
    wire signal_7556 ;
    wire signal_7557 ;
    wire signal_7558 ;
    wire signal_7559 ;
    wire signal_7560 ;
    wire signal_7561 ;
    wire signal_7562 ;
    wire signal_7563 ;
    wire signal_7564 ;
    wire signal_7565 ;
    wire signal_7566 ;
    wire signal_7567 ;
    wire signal_7568 ;
    wire signal_7569 ;
    wire signal_7570 ;
    wire signal_7571 ;
    wire signal_7572 ;
    wire signal_7573 ;
    wire signal_7574 ;
    wire signal_7575 ;
    wire signal_7576 ;
    wire signal_7577 ;
    wire signal_7578 ;
    wire signal_7579 ;
    wire signal_7580 ;
    wire signal_7581 ;
    wire signal_7582 ;
    wire signal_7583 ;
    wire signal_7584 ;
    wire signal_7585 ;
    wire signal_7586 ;
    wire signal_7587 ;
    wire signal_7588 ;
    wire signal_7589 ;
    wire signal_7590 ;
    wire signal_7591 ;
    wire signal_7592 ;
    wire signal_7593 ;
    wire signal_7594 ;
    wire signal_7595 ;
    wire signal_7596 ;
    wire signal_7597 ;
    wire signal_7598 ;
    wire signal_7599 ;
    wire signal_7600 ;
    wire signal_7601 ;
    wire signal_7602 ;
    wire signal_7603 ;
    wire signal_7604 ;
    wire signal_7605 ;
    wire signal_7606 ;
    wire signal_7607 ;
    wire signal_7608 ;
    wire signal_7609 ;
    wire signal_7610 ;
    wire signal_7611 ;
    wire signal_7612 ;
    wire signal_7613 ;
    wire signal_7614 ;
    wire signal_7615 ;
    wire signal_7616 ;
    wire signal_7617 ;
    wire signal_7618 ;
    wire signal_7619 ;
    wire signal_7620 ;
    wire signal_7621 ;
    wire signal_7622 ;
    wire signal_7623 ;
    wire signal_7624 ;
    wire signal_7625 ;
    wire signal_7626 ;
    wire signal_7627 ;
    wire signal_7628 ;
    wire signal_7629 ;
    wire signal_7630 ;
    wire signal_7631 ;
    wire signal_7632 ;
    wire signal_7633 ;
    wire signal_7634 ;
    wire signal_7635 ;
    wire signal_7636 ;
    wire signal_7637 ;
    wire signal_7638 ;
    wire signal_7639 ;
    wire signal_7640 ;
    wire signal_7641 ;
    wire signal_7642 ;
    wire signal_7643 ;
    wire signal_7644 ;
    wire signal_7645 ;
    wire signal_7646 ;
    wire signal_7647 ;
    wire signal_7648 ;
    wire signal_7649 ;
    wire signal_7650 ;
    wire signal_7651 ;
    wire signal_7652 ;
    wire signal_7653 ;
    wire signal_7654 ;
    wire signal_7655 ;
    wire signal_7656 ;
    wire signal_7657 ;
    wire signal_7658 ;
    wire signal_7659 ;
    wire signal_7660 ;
    wire signal_7661 ;
    wire signal_7662 ;
    wire signal_7663 ;
    wire signal_7664 ;
    wire signal_7665 ;
    wire signal_7666 ;
    wire signal_7667 ;
    wire signal_7668 ;
    wire signal_7669 ;
    wire signal_7670 ;
    wire signal_7671 ;
    wire signal_7672 ;
    wire signal_7673 ;
    wire signal_7674 ;
    wire signal_7675 ;
    wire signal_7676 ;
    wire signal_7677 ;
    wire signal_7678 ;
    wire signal_7679 ;
    wire signal_7680 ;
    wire signal_7681 ;
    wire signal_7682 ;
    wire signal_7683 ;
    wire signal_7684 ;
    wire signal_7685 ;
    wire signal_7686 ;
    wire signal_7687 ;
    wire signal_7688 ;
    wire signal_7689 ;
    wire signal_7690 ;
    wire signal_7691 ;
    wire signal_7692 ;
    wire signal_7693 ;
    wire signal_7694 ;
    wire signal_7695 ;
    wire signal_7696 ;
    wire signal_7697 ;
    wire signal_7698 ;
    wire signal_7699 ;
    wire signal_7700 ;
    wire signal_7701 ;
    wire signal_7702 ;
    wire signal_7703 ;
    wire signal_7704 ;
    wire signal_7705 ;
    wire signal_7706 ;
    wire signal_7707 ;
    wire signal_7708 ;
    wire signal_7709 ;
    wire signal_7710 ;
    wire signal_7711 ;
    wire signal_7712 ;
    wire signal_7713 ;
    wire signal_7714 ;
    wire signal_7715 ;
    wire signal_7716 ;
    wire signal_7717 ;
    wire signal_7718 ;
    wire signal_7719 ;
    wire signal_7720 ;
    wire signal_7721 ;
    wire signal_7722 ;
    wire signal_7723 ;
    wire signal_7724 ;
    wire signal_7725 ;
    wire signal_7726 ;
    wire signal_7727 ;
    wire signal_7728 ;
    wire signal_7729 ;
    wire signal_7730 ;
    wire signal_7731 ;
    wire signal_7732 ;
    wire signal_7733 ;
    wire signal_7734 ;
    wire signal_7735 ;
    wire signal_7736 ;
    wire signal_7737 ;
    wire signal_7738 ;
    wire signal_7739 ;
    wire signal_7740 ;
    wire signal_7741 ;
    wire signal_7742 ;
    wire signal_7743 ;
    wire signal_7744 ;
    wire signal_7745 ;
    wire signal_7746 ;
    wire signal_7747 ;
    wire signal_7748 ;
    wire signal_7749 ;
    wire signal_7750 ;
    wire signal_7751 ;
    wire signal_7752 ;
    wire signal_7753 ;
    wire signal_7754 ;
    wire signal_7755 ;
    wire signal_7756 ;
    wire signal_7757 ;
    wire signal_7758 ;
    wire signal_7759 ;
    wire signal_7760 ;
    wire signal_7761 ;
    wire signal_7762 ;
    wire signal_7763 ;
    wire signal_7764 ;
    wire signal_7765 ;
    wire signal_7766 ;
    wire signal_7767 ;
    wire signal_7768 ;
    wire signal_7769 ;
    wire signal_7770 ;
    wire signal_7771 ;
    wire signal_7772 ;
    wire signal_7773 ;
    wire signal_7774 ;
    wire signal_7775 ;
    wire signal_7776 ;
    wire signal_7777 ;
    wire signal_7778 ;
    wire signal_7779 ;
    wire signal_7780 ;
    wire signal_7781 ;
    wire signal_7782 ;
    wire signal_7783 ;
    wire signal_7784 ;
    wire signal_7785 ;
    wire signal_7786 ;
    wire signal_7787 ;
    wire signal_7788 ;
    wire signal_7789 ;
    wire signal_7790 ;
    wire signal_7791 ;
    wire signal_7792 ;
    wire signal_7793 ;
    wire signal_7794 ;
    wire signal_7795 ;
    wire signal_7796 ;
    wire signal_7797 ;
    wire signal_7798 ;
    wire signal_7799 ;
    wire signal_7800 ;
    wire signal_7801 ;
    wire signal_7802 ;
    wire signal_7803 ;
    wire signal_7804 ;
    wire signal_7805 ;
    wire signal_7806 ;
    wire signal_7807 ;
    wire signal_7808 ;
    wire signal_7809 ;
    wire signal_7810 ;
    wire signal_7811 ;
    wire signal_7812 ;
    wire signal_7813 ;
    wire signal_7814 ;
    wire signal_7815 ;
    wire signal_7816 ;
    wire signal_7817 ;
    wire signal_7818 ;
    wire signal_7819 ;
    wire signal_7820 ;
    wire signal_7821 ;
    wire signal_7822 ;
    wire signal_7823 ;
    wire signal_7824 ;
    wire signal_7825 ;
    wire signal_7826 ;
    wire signal_7827 ;
    wire signal_7828 ;
    wire signal_7829 ;
    wire signal_7830 ;
    wire signal_7831 ;
    wire signal_7832 ;
    wire signal_7833 ;
    wire signal_7834 ;
    wire signal_7835 ;
    wire signal_7836 ;
    wire signal_7837 ;
    wire signal_7838 ;
    wire signal_7839 ;
    wire signal_7840 ;
    wire signal_7841 ;
    wire signal_7842 ;
    wire signal_7843 ;
    wire signal_7844 ;
    wire signal_7845 ;
    wire signal_7846 ;
    wire signal_7847 ;
    wire signal_7848 ;
    wire signal_7849 ;
    wire signal_7850 ;
    wire signal_7851 ;
    wire signal_7852 ;
    wire signal_7853 ;
    wire signal_7854 ;
    wire signal_7855 ;
    wire signal_7856 ;
    wire signal_7857 ;
    wire signal_7858 ;
    wire signal_7859 ;
    wire signal_7860 ;
    wire signal_7861 ;
    wire signal_7862 ;
    wire signal_7863 ;
    wire signal_7864 ;
    wire signal_7865 ;
    wire signal_7866 ;
    wire signal_7867 ;
    wire signal_7868 ;
    wire signal_7869 ;
    wire signal_7870 ;
    wire signal_7871 ;
    wire signal_7872 ;
    wire signal_7873 ;
    wire signal_7874 ;
    wire signal_7875 ;
    wire signal_7876 ;
    wire signal_7877 ;
    wire signal_7878 ;
    wire signal_7879 ;
    wire signal_7880 ;
    wire signal_7881 ;
    wire signal_7882 ;
    wire signal_7883 ;
    wire signal_7884 ;
    wire signal_7885 ;
    wire signal_7886 ;
    wire signal_7887 ;
    wire signal_7888 ;
    wire signal_7889 ;
    wire signal_7890 ;
    wire signal_7891 ;
    wire signal_7892 ;
    wire signal_7893 ;
    wire signal_7894 ;
    wire signal_7895 ;
    wire signal_7896 ;
    wire signal_7897 ;
    wire signal_7898 ;
    wire signal_7899 ;
    wire signal_7900 ;
    wire signal_7901 ;
    wire signal_7902 ;
    wire signal_7903 ;
    wire signal_7904 ;
    wire signal_7905 ;
    wire signal_7906 ;
    wire signal_7907 ;
    wire signal_7908 ;
    wire signal_7909 ;
    wire signal_7910 ;
    wire signal_7911 ;
    wire signal_7912 ;
    wire signal_7913 ;
    wire signal_7914 ;
    wire signal_7915 ;
    wire signal_7916 ;
    wire signal_7917 ;
    wire signal_7918 ;
    wire signal_7919 ;
    wire signal_7920 ;
    wire signal_7921 ;
    wire signal_7922 ;
    wire signal_7923 ;
    wire signal_7924 ;
    wire signal_7925 ;
    wire signal_7926 ;
    wire signal_7927 ;
    wire signal_7928 ;
    wire signal_7929 ;
    wire signal_7930 ;
    wire signal_7931 ;
    wire signal_7932 ;
    wire signal_7933 ;
    wire signal_7934 ;
    wire signal_7935 ;
    wire signal_7936 ;
    wire signal_7937 ;
    wire signal_7938 ;
    wire signal_7939 ;
    wire signal_7940 ;
    wire signal_7941 ;
    wire signal_7942 ;
    wire signal_7943 ;
    wire signal_7944 ;
    wire signal_7945 ;
    wire signal_7946 ;
    wire signal_7947 ;
    wire signal_7948 ;
    wire signal_7949 ;
    wire signal_7950 ;
    wire signal_7951 ;
    wire signal_7952 ;
    wire signal_7953 ;
    wire signal_7954 ;
    wire signal_7955 ;
    wire signal_7956 ;
    wire signal_7957 ;
    wire signal_7958 ;
    wire signal_7959 ;
    wire signal_7960 ;
    wire signal_7961 ;
    wire signal_7962 ;
    wire signal_7963 ;
    wire signal_7964 ;
    wire signal_7965 ;
    wire signal_7966 ;
    wire signal_7967 ;
    wire signal_7968 ;
    wire signal_7969 ;
    wire signal_7970 ;
    wire signal_7971 ;
    wire signal_7972 ;
    wire signal_7973 ;
    wire signal_7974 ;
    wire signal_7975 ;
    wire signal_7976 ;
    wire signal_7977 ;
    wire signal_7978 ;
    wire signal_7979 ;
    wire signal_7980 ;
    wire signal_7981 ;
    wire signal_7982 ;
    wire signal_7983 ;
    wire signal_7984 ;
    wire signal_7985 ;
    wire signal_7986 ;
    wire signal_7987 ;
    wire signal_7988 ;
    wire signal_7989 ;
    wire signal_7990 ;
    wire signal_7991 ;
    wire signal_7992 ;
    wire signal_7993 ;
    wire signal_7994 ;
    wire signal_7995 ;
    wire signal_7996 ;
    wire signal_7997 ;
    wire signal_7998 ;
    wire signal_7999 ;
    wire signal_8000 ;
    wire signal_8001 ;
    wire signal_8002 ;
    wire signal_8003 ;
    wire signal_8004 ;
    wire signal_8005 ;
    wire signal_8006 ;
    wire signal_8007 ;
    wire signal_8008 ;
    wire signal_8009 ;
    wire signal_8010 ;
    wire signal_8011 ;
    wire signal_8012 ;
    wire signal_8013 ;
    wire signal_8014 ;
    wire signal_8015 ;
    wire signal_8016 ;
    wire signal_8017 ;
    wire signal_8018 ;
    wire signal_8019 ;
    wire signal_8020 ;
    wire signal_8021 ;
    wire signal_8022 ;
    wire signal_8023 ;
    wire signal_8024 ;
    wire signal_8025 ;
    wire signal_8026 ;
    wire signal_8027 ;
    wire signal_8028 ;
    wire signal_8029 ;
    wire signal_8030 ;
    wire signal_8031 ;
    wire signal_8032 ;
    wire signal_8033 ;
    wire signal_8034 ;
    wire signal_8035 ;
    wire signal_8036 ;
    wire signal_8037 ;
    wire signal_8038 ;
    wire signal_8039 ;
    wire signal_8040 ;
    wire signal_8041 ;
    wire signal_8042 ;
    wire signal_8043 ;
    wire signal_8044 ;
    wire signal_8045 ;
    wire signal_8046 ;
    wire signal_8047 ;
    wire signal_8048 ;
    wire signal_8049 ;
    wire signal_8050 ;
    wire signal_8051 ;
    wire signal_8052 ;
    wire signal_8053 ;
    wire signal_8054 ;
    wire signal_8055 ;
    wire signal_8056 ;
    wire signal_8057 ;
    wire signal_8058 ;
    wire signal_8059 ;
    wire signal_8060 ;
    wire signal_8061 ;
    wire signal_8062 ;
    wire signal_8063 ;
    wire signal_8064 ;
    wire signal_8065 ;
    wire signal_8066 ;
    wire signal_8067 ;
    wire signal_8068 ;
    wire signal_8069 ;
    wire signal_8070 ;
    wire signal_8071 ;
    wire signal_8072 ;
    wire signal_8073 ;
    wire signal_8074 ;
    wire signal_8075 ;
    wire signal_8076 ;
    wire signal_8077 ;
    wire signal_8078 ;
    wire signal_8079 ;
    wire signal_8080 ;
    wire signal_8081 ;
    wire signal_8082 ;
    wire signal_8083 ;
    wire signal_8084 ;
    wire signal_8085 ;
    wire signal_8086 ;
    wire signal_8087 ;
    wire signal_8088 ;
    wire signal_8089 ;
    wire signal_8090 ;
    wire signal_8091 ;
    wire signal_8092 ;
    wire signal_8093 ;
    wire signal_8094 ;
    wire signal_8095 ;
    wire signal_8096 ;
    wire signal_8097 ;
    wire signal_8098 ;
    wire signal_8099 ;
    wire signal_8100 ;
    wire signal_8101 ;
    wire signal_8102 ;
    wire signal_8103 ;
    wire signal_8104 ;
    wire signal_8105 ;
    wire signal_8106 ;
    wire signal_8107 ;
    wire signal_8108 ;
    wire signal_8109 ;
    wire signal_8110 ;
    wire signal_8111 ;
    wire signal_8112 ;
    wire signal_8113 ;
    wire signal_8114 ;
    wire signal_8115 ;
    wire signal_8116 ;
    wire signal_8117 ;
    wire signal_8118 ;
    wire signal_8119 ;
    wire signal_8120 ;
    wire signal_8121 ;
    wire signal_8122 ;
    wire signal_8123 ;
    wire signal_8124 ;
    wire signal_8125 ;
    wire signal_8126 ;
    wire signal_8127 ;
    wire signal_8128 ;
    wire signal_8129 ;
    wire signal_8130 ;
    wire signal_8131 ;
    wire signal_8132 ;
    wire signal_8133 ;
    wire signal_8134 ;
    wire signal_8135 ;
    wire signal_8136 ;
    wire signal_8137 ;
    wire signal_8138 ;
    wire signal_8139 ;
    wire signal_8140 ;
    wire signal_8141 ;
    wire signal_8142 ;
    wire signal_8143 ;
    wire signal_8144 ;
    wire signal_8145 ;
    wire signal_8146 ;
    wire signal_8147 ;
    wire signal_8148 ;
    wire signal_8149 ;
    wire signal_8150 ;
    wire signal_8151 ;
    wire signal_8152 ;
    wire signal_8153 ;
    wire signal_8154 ;
    wire signal_8155 ;
    wire signal_8156 ;
    wire signal_8157 ;
    wire signal_8158 ;
    wire signal_8159 ;
    wire signal_8160 ;
    wire signal_8161 ;
    wire signal_8162 ;
    wire signal_8163 ;
    wire signal_8164 ;
    wire signal_8165 ;
    wire signal_8166 ;
    wire signal_8167 ;
    wire signal_8168 ;
    wire signal_8169 ;
    wire signal_8170 ;
    wire signal_8171 ;
    wire signal_8172 ;
    wire signal_8173 ;
    wire signal_8174 ;
    wire signal_8175 ;
    wire signal_8176 ;
    wire signal_8177 ;
    wire signal_8178 ;
    wire signal_8179 ;
    wire signal_8180 ;
    wire signal_8181 ;
    wire signal_8182 ;
    wire signal_8183 ;
    wire signal_8184 ;
    wire signal_8185 ;
    wire signal_8186 ;
    wire signal_8187 ;
    wire signal_8188 ;
    wire signal_8189 ;
    wire signal_8190 ;
    wire signal_8191 ;
    wire signal_8192 ;
    wire signal_8193 ;
    wire signal_8194 ;
    wire signal_8195 ;
    wire signal_8196 ;
    wire signal_8197 ;
    wire signal_8198 ;
    wire signal_8199 ;
    wire signal_8200 ;
    wire signal_8201 ;
    wire signal_8202 ;
    wire signal_8203 ;
    wire signal_8204 ;
    wire signal_8205 ;
    wire signal_8206 ;
    wire signal_8207 ;
    wire signal_8208 ;
    wire signal_8209 ;
    wire signal_8210 ;
    wire signal_8211 ;
    wire signal_8212 ;
    wire signal_8213 ;
    wire signal_8214 ;
    wire signal_8215 ;
    wire signal_8216 ;
    wire signal_8217 ;
    wire signal_8218 ;
    wire signal_8219 ;
    wire signal_8220 ;
    wire signal_8221 ;
    wire signal_8222 ;
    wire signal_8223 ;
    wire signal_8224 ;
    wire signal_8225 ;
    wire signal_8226 ;
    wire signal_8227 ;
    wire signal_8228 ;
    wire signal_8229 ;
    wire signal_8230 ;
    wire signal_8231 ;
    wire signal_8232 ;
    wire signal_8233 ;
    wire signal_8234 ;
    wire signal_8235 ;
    wire signal_8236 ;
    wire signal_8237 ;
    wire signal_8238 ;
    wire signal_8239 ;
    wire signal_8240 ;
    wire signal_8241 ;
    wire signal_8242 ;
    wire signal_8243 ;
    wire signal_8244 ;
    wire signal_8245 ;
    wire signal_8246 ;
    wire signal_8247 ;
    wire signal_8248 ;
    wire signal_8249 ;
    wire signal_8250 ;
    wire signal_8251 ;
    wire signal_8252 ;
    wire signal_8253 ;
    wire signal_8254 ;
    wire signal_8255 ;
    wire signal_8256 ;
    wire signal_8257 ;
    wire signal_8258 ;
    wire signal_8259 ;
    wire signal_8260 ;
    wire signal_8261 ;
    wire signal_8262 ;
    wire signal_8263 ;
    wire signal_8264 ;
    wire signal_8265 ;
    wire signal_8266 ;
    wire signal_8267 ;
    wire signal_8268 ;
    wire signal_8269 ;
    wire signal_8270 ;
    wire signal_8271 ;
    wire signal_8272 ;
    wire signal_8273 ;
    wire signal_8274 ;
    wire signal_8275 ;
    wire signal_8276 ;
    wire signal_8277 ;
    wire signal_8278 ;
    wire signal_8279 ;
    wire signal_8280 ;
    wire signal_8281 ;
    wire signal_8282 ;
    wire signal_8283 ;
    wire signal_8284 ;
    wire signal_8285 ;
    wire signal_8286 ;
    wire signal_8287 ;
    wire signal_8288 ;
    wire signal_8289 ;
    wire signal_8290 ;
    wire signal_8291 ;
    wire signal_8292 ;
    wire signal_8293 ;
    wire signal_8294 ;
    wire signal_8295 ;
    wire signal_8296 ;
    wire signal_8297 ;
    wire signal_8298 ;
    wire signal_8299 ;
    wire signal_8300 ;
    wire signal_8301 ;
    wire signal_8302 ;
    wire signal_8303 ;
    wire signal_8304 ;
    wire signal_8305 ;
    wire signal_8306 ;
    wire signal_8307 ;
    wire signal_8308 ;
    wire signal_8309 ;
    wire signal_8310 ;
    wire signal_8311 ;
    wire signal_8312 ;
    wire signal_8313 ;
    wire signal_8314 ;
    wire signal_8315 ;
    wire signal_8316 ;
    wire signal_8317 ;
    wire signal_8318 ;
    wire signal_8319 ;
    wire signal_8320 ;
    wire signal_8321 ;
    wire signal_8322 ;
    wire signal_8323 ;
    wire signal_8324 ;
    wire signal_8325 ;
    wire signal_8326 ;
    wire signal_8327 ;
    wire signal_8328 ;
    wire signal_8329 ;
    wire signal_8330 ;
    wire signal_8331 ;
    wire signal_8332 ;
    wire signal_8333 ;
    wire signal_8334 ;
    wire signal_8335 ;
    wire signal_8336 ;
    wire signal_8337 ;
    wire signal_8338 ;
    wire signal_8339 ;
    wire signal_8340 ;
    wire signal_8341 ;
    wire signal_8342 ;
    wire signal_8343 ;
    wire signal_8344 ;
    wire signal_8345 ;
    wire signal_8346 ;
    wire signal_8347 ;
    wire signal_8348 ;
    wire signal_8349 ;
    wire signal_8350 ;
    wire signal_8351 ;
    wire signal_8352 ;
    wire signal_8353 ;
    wire signal_8354 ;
    wire signal_8355 ;
    wire signal_8356 ;
    wire signal_8357 ;
    wire signal_8358 ;
    wire signal_8359 ;
    wire signal_8360 ;
    wire signal_8361 ;
    wire signal_8362 ;
    wire signal_8363 ;
    wire signal_8364 ;
    wire signal_8365 ;
    wire signal_8366 ;
    wire signal_8367 ;
    wire signal_8368 ;
    wire signal_8369 ;
    wire signal_8370 ;
    wire signal_8371 ;
    wire signal_8372 ;
    wire signal_8373 ;
    wire signal_8374 ;
    wire signal_8375 ;
    wire signal_8376 ;
    wire signal_8377 ;
    wire signal_8378 ;
    wire signal_8379 ;
    wire signal_8380 ;
    wire signal_8381 ;
    wire signal_8382 ;
    wire signal_8383 ;
    wire signal_8384 ;
    wire signal_8385 ;
    wire signal_8386 ;
    wire signal_8387 ;
    wire signal_8388 ;
    wire signal_8389 ;
    wire signal_8390 ;
    wire signal_8391 ;
    wire signal_8392 ;
    wire signal_8393 ;
    wire signal_8394 ;
    wire signal_8395 ;
    wire signal_8396 ;
    wire signal_8397 ;
    wire signal_8398 ;
    wire signal_8399 ;
    wire signal_8400 ;
    wire signal_8401 ;
    wire signal_8402 ;
    wire signal_8403 ;
    wire signal_8404 ;
    wire signal_8405 ;
    wire signal_8406 ;
    wire signal_8407 ;
    wire signal_8408 ;
    wire signal_8409 ;
    wire signal_8410 ;
    wire signal_8411 ;
    wire signal_8412 ;
    wire signal_8413 ;
    wire signal_8414 ;
    wire signal_8415 ;
    wire signal_8416 ;
    wire signal_8417 ;
    wire signal_8418 ;
    wire signal_8419 ;
    wire signal_8420 ;
    wire signal_8421 ;
    wire signal_8422 ;
    wire signal_8423 ;
    wire signal_8424 ;
    wire signal_8425 ;
    wire signal_8426 ;
    wire signal_8427 ;
    wire signal_8428 ;
    wire signal_8429 ;
    wire signal_8430 ;
    wire signal_8431 ;
    wire signal_8432 ;
    wire signal_8433 ;
    wire signal_8434 ;
    wire signal_8435 ;
    wire signal_8436 ;
    wire signal_8437 ;
    wire signal_8438 ;
    wire signal_8439 ;
    wire signal_8440 ;
    wire signal_8441 ;
    wire signal_8442 ;
    wire signal_8443 ;
    wire signal_8444 ;
    wire signal_8445 ;
    wire signal_8446 ;
    wire signal_8447 ;
    wire signal_8448 ;
    wire signal_8449 ;
    wire signal_8450 ;
    wire signal_8451 ;
    wire signal_8452 ;
    wire signal_8453 ;
    wire signal_8454 ;
    wire signal_8455 ;
    wire signal_8456 ;
    wire signal_8457 ;
    wire signal_8458 ;
    wire signal_8459 ;
    wire signal_8460 ;
    wire signal_8461 ;
    wire signal_8462 ;
    wire signal_8463 ;
    wire signal_8464 ;
    wire signal_8465 ;
    wire signal_8466 ;
    wire signal_8467 ;
    wire signal_8468 ;
    wire signal_8469 ;
    wire signal_8470 ;
    wire signal_8471 ;
    wire signal_8472 ;
    wire signal_8473 ;
    wire signal_8474 ;
    wire signal_8475 ;
    wire signal_8476 ;
    wire signal_8477 ;
    wire signal_8478 ;
    wire signal_8479 ;
    wire signal_8480 ;
    wire signal_8481 ;
    wire signal_8482 ;
    wire signal_8483 ;
    wire signal_8484 ;
    wire signal_8485 ;
    wire signal_8486 ;
    wire signal_8487 ;
    wire signal_8488 ;
    wire signal_8489 ;
    wire signal_8490 ;
    wire signal_8491 ;
    wire signal_8492 ;
    wire signal_8493 ;
    wire signal_8494 ;
    wire signal_8495 ;
    wire signal_8496 ;
    wire signal_8497 ;
    wire signal_8498 ;
    wire signal_8499 ;
    wire signal_8500 ;
    wire signal_8501 ;
    wire signal_8502 ;
    wire signal_8503 ;
    wire signal_8504 ;
    wire signal_8505 ;
    wire signal_8506 ;
    wire signal_8507 ;
    wire signal_8508 ;
    wire signal_8509 ;
    wire signal_8510 ;
    wire signal_8511 ;
    wire signal_8512 ;
    wire signal_8513 ;
    wire signal_8514 ;
    wire signal_8515 ;
    wire signal_8516 ;
    wire signal_8517 ;
    wire signal_8518 ;
    wire signal_8519 ;
    wire signal_8520 ;
    wire signal_8521 ;
    wire signal_8522 ;
    wire signal_8523 ;
    wire signal_8524 ;
    wire signal_8525 ;
    wire signal_8526 ;
    wire signal_8527 ;
    wire signal_8528 ;
    wire signal_8529 ;
    wire signal_8530 ;
    wire signal_8531 ;
    wire signal_8532 ;
    wire signal_8533 ;
    wire signal_8534 ;
    wire signal_8535 ;
    wire signal_8536 ;
    wire signal_8537 ;
    wire signal_8538 ;
    wire signal_8539 ;
    wire signal_8540 ;
    wire signal_8541 ;
    wire signal_8542 ;
    wire signal_8543 ;
    wire signal_8544 ;
    wire signal_8545 ;
    wire signal_8546 ;
    wire signal_8547 ;
    wire signal_8548 ;
    wire signal_8549 ;
    wire signal_8550 ;
    wire signal_8551 ;
    wire signal_8552 ;
    wire signal_8553 ;
    wire signal_8554 ;
    wire signal_8555 ;
    wire signal_8556 ;
    wire signal_8557 ;
    wire signal_8558 ;
    wire signal_8559 ;
    wire signal_8560 ;
    wire signal_8561 ;
    wire signal_8562 ;
    wire signal_8563 ;
    wire signal_8564 ;
    wire signal_8565 ;
    wire signal_8566 ;
    wire signal_8567 ;
    wire signal_8568 ;
    wire signal_8569 ;
    wire signal_8570 ;
    wire signal_8571 ;
    wire signal_8572 ;
    wire signal_8573 ;
    wire signal_8574 ;
    wire signal_8575 ;
    wire signal_8576 ;
    wire signal_8577 ;
    wire signal_8578 ;
    wire signal_8579 ;
    wire signal_8580 ;
    wire signal_8581 ;
    wire signal_8582 ;
    wire signal_8583 ;
    wire signal_8584 ;
    wire signal_8585 ;
    wire signal_8586 ;
    wire signal_8587 ;
    wire signal_8588 ;
    wire signal_8589 ;
    wire signal_8590 ;
    wire signal_8591 ;
    wire signal_8592 ;
    wire signal_8593 ;
    wire signal_8594 ;
    wire signal_8595 ;
    wire signal_8596 ;
    wire signal_8597 ;
    wire signal_8598 ;
    wire signal_8599 ;
    wire signal_8600 ;
    wire signal_8601 ;
    wire signal_8602 ;
    wire signal_8603 ;
    wire signal_8604 ;
    wire signal_8605 ;
    wire signal_8606 ;
    wire signal_8607 ;
    wire signal_8608 ;
    wire signal_8609 ;
    wire signal_8610 ;
    wire signal_8611 ;
    wire signal_8612 ;
    wire signal_8613 ;
    wire signal_8614 ;
    wire signal_8615 ;
    wire signal_8616 ;
    wire signal_8617 ;
    wire signal_8618 ;
    wire signal_8619 ;
    wire signal_8620 ;
    wire signal_8621 ;
    wire signal_8622 ;
    wire signal_8623 ;
    wire signal_8624 ;
    wire signal_8625 ;
    wire signal_8626 ;
    wire signal_8627 ;
    wire signal_8628 ;
    wire signal_8629 ;
    wire signal_8630 ;
    wire signal_8631 ;
    wire signal_8632 ;
    wire signal_8633 ;
    wire signal_8634 ;
    wire signal_8635 ;
    wire signal_8636 ;
    wire signal_8637 ;
    wire signal_8638 ;
    wire signal_8639 ;
    wire signal_8640 ;
    wire signal_8641 ;
    wire signal_8642 ;
    wire signal_8643 ;
    wire signal_8644 ;
    wire signal_8645 ;
    wire signal_8646 ;
    wire signal_8647 ;
    wire signal_8648 ;
    wire signal_8649 ;
    wire signal_8650 ;
    wire signal_8651 ;
    wire signal_8652 ;
    wire signal_8653 ;
    wire signal_8654 ;
    wire signal_8655 ;
    wire signal_8656 ;
    wire signal_8657 ;
    wire signal_8658 ;
    wire signal_8659 ;
    wire signal_8660 ;
    wire signal_8661 ;
    wire signal_8662 ;
    wire signal_8663 ;
    wire signal_8664 ;
    wire signal_8665 ;
    wire signal_8666 ;
    wire signal_8667 ;
    wire signal_8668 ;
    wire signal_8669 ;
    wire signal_8670 ;
    wire signal_8671 ;
    wire signal_8672 ;
    wire signal_8673 ;
    wire signal_8674 ;
    wire signal_8675 ;
    wire signal_8676 ;
    wire signal_8677 ;
    wire signal_8678 ;
    wire signal_8679 ;
    wire signal_8680 ;
    wire signal_8681 ;
    wire signal_8682 ;
    wire signal_8683 ;
    wire signal_8684 ;
    wire signal_8685 ;
    wire signal_8686 ;
    wire signal_8687 ;
    wire signal_8688 ;
    wire signal_8689 ;
    wire signal_8690 ;
    wire signal_8691 ;
    wire signal_8692 ;
    wire signal_8693 ;
    wire signal_8694 ;
    wire signal_8695 ;
    wire signal_8696 ;
    wire signal_8697 ;
    wire signal_8698 ;
    wire signal_8699 ;
    wire signal_8700 ;
    wire signal_8701 ;
    wire signal_8702 ;
    wire signal_8703 ;
    wire signal_8704 ;
    wire signal_8705 ;
    wire signal_8706 ;
    wire signal_8707 ;
    wire signal_8708 ;
    wire signal_8709 ;
    wire signal_8710 ;
    wire signal_8711 ;
    wire signal_8712 ;
    wire signal_8713 ;
    wire signal_8714 ;
    wire signal_8715 ;
    wire signal_8716 ;
    wire signal_8717 ;
    wire signal_8718 ;
    wire signal_8719 ;
    wire signal_8720 ;
    wire signal_8721 ;
    wire signal_8722 ;
    wire signal_8723 ;
    wire signal_8724 ;
    wire signal_8725 ;
    wire signal_8726 ;
    wire signal_8727 ;
    wire signal_8728 ;
    wire signal_8729 ;
    wire signal_8730 ;
    wire signal_8731 ;
    wire signal_8732 ;
    wire signal_8733 ;
    wire signal_8734 ;
    wire signal_8735 ;
    wire signal_8736 ;
    wire signal_8737 ;
    wire signal_8738 ;
    wire signal_8739 ;
    wire signal_8740 ;
    wire signal_8741 ;
    wire signal_8742 ;
    wire signal_8743 ;
    wire signal_8744 ;
    wire signal_8745 ;
    wire signal_8746 ;
    wire signal_8747 ;
    wire signal_8748 ;
    wire signal_8749 ;
    wire signal_8750 ;
    wire signal_8751 ;
    wire signal_8752 ;
    wire signal_8753 ;
    wire signal_8754 ;
    wire signal_8755 ;
    wire signal_8756 ;
    wire signal_8757 ;
    wire signal_8758 ;
    wire signal_8759 ;
    wire signal_8760 ;
    wire signal_8761 ;
    wire signal_8762 ;
    wire signal_8763 ;
    wire signal_8764 ;
    wire signal_8765 ;
    wire signal_8766 ;
    wire signal_8767 ;
    wire signal_8768 ;
    wire signal_8769 ;
    wire signal_8770 ;
    wire signal_8771 ;
    wire signal_8772 ;
    wire signal_8773 ;
    wire signal_8774 ;
    wire signal_8775 ;
    wire signal_8776 ;
    wire signal_8777 ;
    wire signal_8778 ;
    wire signal_8779 ;
    wire signal_8780 ;
    wire signal_8781 ;
    wire signal_8782 ;
    wire signal_8783 ;
    wire signal_8784 ;
    wire signal_8785 ;
    wire signal_8786 ;
    wire signal_8787 ;
    wire signal_8788 ;
    wire signal_8789 ;
    wire signal_8790 ;
    wire signal_8791 ;
    wire signal_8792 ;
    wire signal_8793 ;
    wire signal_8794 ;
    wire signal_8795 ;
    wire signal_8796 ;
    wire signal_8797 ;
    wire signal_8798 ;
    wire signal_8799 ;
    wire signal_8800 ;
    wire signal_8801 ;
    wire signal_8802 ;
    wire signal_8803 ;
    wire signal_8804 ;
    wire signal_8805 ;
    wire signal_8806 ;
    wire signal_8807 ;
    wire signal_8808 ;
    wire signal_8809 ;
    wire signal_8810 ;
    wire signal_8811 ;
    wire signal_8812 ;
    wire signal_8813 ;
    wire signal_8814 ;
    wire signal_8815 ;
    wire signal_8816 ;
    wire signal_8817 ;
    wire signal_8818 ;
    wire signal_8819 ;
    wire signal_8820 ;
    wire signal_8821 ;
    wire signal_8822 ;
    wire signal_8823 ;
    wire signal_8824 ;
    wire signal_8825 ;
    wire signal_8826 ;
    wire signal_8827 ;
    wire signal_8828 ;
    wire signal_8829 ;
    wire signal_8830 ;
    wire signal_8831 ;
    wire signal_8832 ;
    wire signal_8833 ;
    wire signal_8834 ;
    wire signal_8835 ;
    wire signal_8836 ;
    wire signal_8837 ;
    wire signal_8838 ;
    wire signal_8839 ;
    wire signal_8840 ;
    wire signal_8841 ;
    wire signal_8842 ;
    wire signal_8843 ;
    wire signal_8844 ;
    wire signal_8845 ;
    wire signal_8846 ;
    wire signal_8847 ;
    wire signal_8848 ;
    wire signal_8849 ;
    wire signal_8850 ;
    wire signal_8851 ;
    wire signal_8852 ;
    wire signal_8853 ;
    wire signal_8854 ;
    wire signal_8855 ;
    wire signal_8856 ;
    wire signal_8857 ;
    wire signal_8858 ;
    wire signal_8859 ;
    wire signal_8860 ;
    wire signal_8861 ;
    wire signal_8862 ;
    wire signal_8863 ;
    wire signal_8864 ;
    wire signal_8865 ;
    wire signal_8866 ;
    wire signal_8867 ;
    wire signal_8868 ;
    wire signal_8869 ;
    wire signal_8870 ;
    wire signal_8871 ;
    wire signal_8872 ;
    wire signal_8873 ;
    wire signal_8874 ;
    wire signal_8875 ;
    wire signal_8876 ;
    wire signal_8877 ;
    wire signal_8878 ;
    wire signal_8879 ;
    wire signal_8880 ;
    wire signal_8881 ;
    wire signal_8882 ;
    wire signal_8883 ;
    wire signal_8884 ;
    wire signal_8885 ;
    wire signal_8886 ;
    wire signal_8887 ;
    wire signal_8888 ;
    wire signal_8889 ;
    wire signal_8890 ;
    wire signal_8891 ;
    wire signal_8892 ;
    wire signal_8893 ;
    wire signal_8894 ;
    wire signal_8895 ;
    wire signal_8896 ;
    wire signal_8897 ;
    wire signal_8898 ;
    wire signal_8899 ;
    wire signal_8900 ;
    wire signal_8901 ;
    wire signal_8902 ;
    wire signal_8903 ;
    wire signal_8904 ;
    wire signal_8905 ;
    wire signal_8906 ;
    wire signal_8907 ;
    wire signal_8908 ;
    wire signal_8909 ;
    wire signal_8910 ;
    wire signal_8911 ;
    wire signal_8912 ;
    wire signal_8913 ;
    wire signal_8914 ;
    wire signal_8915 ;
    wire signal_8916 ;
    wire signal_8917 ;
    wire signal_8918 ;
    wire signal_8919 ;
    wire signal_8920 ;
    wire signal_8921 ;
    wire signal_8922 ;
    wire signal_8923 ;
    wire signal_8924 ;
    wire signal_8925 ;
    wire signal_8926 ;
    wire signal_8927 ;
    wire signal_8928 ;
    wire signal_8929 ;
    wire signal_8930 ;
    wire signal_8931 ;
    wire signal_8932 ;
    wire signal_8933 ;
    wire signal_8934 ;
    wire signal_8935 ;
    wire signal_8936 ;
    wire signal_8937 ;
    wire signal_8938 ;
    wire signal_8939 ;
    wire signal_8940 ;
    wire signal_8941 ;
    wire signal_8942 ;
    wire signal_8943 ;
    wire signal_8944 ;
    wire signal_8945 ;
    wire signal_8946 ;
    wire signal_8947 ;
    wire signal_8948 ;
    wire signal_8949 ;
    wire signal_8950 ;
    wire signal_8951 ;

    /* cells in depth 0 */
    INV_X1 cell_0 ( .A (signal_395), .ZN (signal_404) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({signal_2107, signal_1493}), .c ({signal_2108, signal_1413}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_2 ( .a ({ciphertext_s1[121], ciphertext_s0[121]}), .b ({signal_2110, signal_1492}), .c ({signal_2111, signal_1412}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3 ( .a ({ciphertext_s1[122], ciphertext_s0[122]}), .b ({signal_2113, signal_1491}), .c ({signal_2114, signal_1411}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4 ( .a ({ciphertext_s1[123], ciphertext_s0[123]}), .b ({signal_2116, signal_1490}), .c ({signal_2117, signal_1410}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5 ( .a ({ciphertext_s1[124], ciphertext_s0[124]}), .b ({signal_2119, signal_1489}), .c ({signal_2120, signal_1409}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6 ( .a ({ciphertext_s1[125], ciphertext_s0[125]}), .b ({signal_2122, signal_1488}), .c ({signal_2123, signal_1408}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7 ( .a ({ciphertext_s1[126], ciphertext_s0[126]}), .b ({signal_2125, signal_1487}), .c ({signal_2126, signal_1407}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_8 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({signal_2128, signal_1486}), .c ({signal_2129, signal_1406}) ) ;
    NAND2_X1 cell_9 ( .A1 (signal_399), .A2 (signal_398), .ZN (signal_405) ) ;
    NOR2_X1 cell_10 ( .A1 (signal_402), .A2 (signal_405), .ZN (done) ) ;
    AND2_X1 cell_11 ( .A1 (signal_401), .A2 (signal_396), .ZN (signal_400) ) ;
    INV_X1 cell_12 ( .A (start), .ZN (signal_403) ) ;
    NOR2_X1 cell_13 ( .A1 (signal_406), .A2 (signal_415), .ZN (signal_422) ) ;
    XNOR2_X1 cell_14 ( .A (signal_424), .B (signal_425), .ZN (signal_423) ) ;
    NOR2_X1 cell_15 ( .A1 (signal_407), .A2 (signal_408), .ZN (signal_398) ) ;
    NAND2_X1 cell_16 ( .A1 (signal_421), .A2 (signal_416), .ZN (signal_408) ) ;
    INV_X1 cell_17 ( .A (signal_406), .ZN (signal_407) ) ;
    INV_X1 cell_18 ( .A (signal_420), .ZN (signal_416) ) ;
    NAND2_X1 cell_19 ( .A1 (signal_409), .A2 (signal_410), .ZN (signal_419) ) ;
    NAND2_X1 cell_20 ( .A1 (signal_396), .A2 (signal_418), .ZN (signal_409) ) ;
    NOR2_X1 cell_21 ( .A1 (signal_427), .A2 (signal_424), .ZN (signal_413) ) ;
    NOR2_X1 cell_22 ( .A1 (signal_425), .A2 (signal_428), .ZN (signal_412) ) ;
    NOR2_X1 cell_23 ( .A1 (signal_415), .A2 (signal_414), .ZN (signal_396) ) ;
    NOR2_X1 cell_24 ( .A1 (signal_420), .A2 (signal_421), .ZN (signal_414) ) ;
    INV_X1 cell_25 ( .A (signal_393), .ZN (signal_415) ) ;
    NAND2_X1 cell_26 ( .A1 (signal_412), .A2 (signal_413), .ZN (signal_411) ) ;
    NOR2_X1 cell_27 ( .A1 (signal_426), .A2 (signal_411), .ZN (signal_406) ) ;
    NAND2_X1 cell_28 ( .A1 (signal_393), .A2 (signal_406), .ZN (signal_410) ) ;
    INV_X1 cell_29 ( .A (signal_410), .ZN (signal_395) ) ;
    NOR2_X1 cell_30 ( .A1 (signal_417), .A2 (signal_415), .ZN (signal_394) ) ;
    MUX2_X1 cell_31 ( .S (signal_393), .A (1'b1), .B (signal_423), .Z (signal_429) ) ;
    MUX2_X1 cell_34 ( .S (signal_393), .A (1'b0), .B (signal_425), .Z (signal_431) ) ;
    MUX2_X1 cell_37 ( .S (signal_393), .A (1'b1), .B (signal_426), .Z (signal_433) ) ;
    MUX2_X1 cell_40 ( .S (signal_393), .A (1'b0), .B (signal_427), .Z (signal_435) ) ;
    MUX2_X1 cell_43 ( .S (signal_393), .A (1'b1), .B (signal_428), .Z (signal_437) ) ;
    MUX2_X1 cell_46 ( .S (signal_422), .A (1'b1), .B (signal_416), .Z (signal_439) ) ;
    MUX2_X1 cell_49 ( .S (signal_422), .A (1'b0), .B (signal_421), .Z (signal_441) ) ;
    INV_X1 cell_52 ( .A (signal_418), .ZN (signal_417) ) ;
    INV_X1 cell_64 ( .A (signal_394), .ZN (signal_453) ) ;
    INV_X1 cell_65 ( .A (signal_453), .ZN (signal_455) ) ;
    INV_X1 cell_66 ( .A (signal_393), .ZN (signal_444) ) ;
    INV_X1 cell_67 ( .A (signal_444), .ZN (signal_452) ) ;
    INV_X1 cell_68 ( .A (signal_456), .ZN (signal_464) ) ;
    INV_X1 cell_69 ( .A (signal_453), .ZN (signal_454) ) ;
    INV_X1 cell_70 ( .A (signal_444), .ZN (signal_448) ) ;
    INV_X1 cell_71 ( .A (signal_456), .ZN (signal_460) ) ;
    INV_X1 cell_72 ( .A (signal_444), .ZN (signal_446) ) ;
    INV_X1 cell_73 ( .A (signal_456), .ZN (signal_458) ) ;
    INV_X1 cell_74 ( .A (signal_444), .ZN (signal_450) ) ;
    INV_X1 cell_75 ( .A (signal_456), .ZN (signal_462) ) ;
    INV_X1 cell_76 ( .A (signal_444), .ZN (signal_445) ) ;
    INV_X1 cell_77 ( .A (signal_456), .ZN (signal_457) ) ;
    INV_X1 cell_78 ( .A (signal_444), .ZN (signal_447) ) ;
    INV_X1 cell_79 ( .A (signal_456), .ZN (signal_459) ) ;
    INV_X1 cell_80 ( .A (signal_444), .ZN (signal_449) ) ;
    INV_X1 cell_81 ( .A (signal_456), .ZN (signal_461) ) ;
    INV_X1 cell_82 ( .A (signal_444), .ZN (signal_451) ) ;
    INV_X1 cell_83 ( .A (signal_456), .ZN (signal_463) ) ;
    INV_X1 cell_84 ( .A (signal_395), .ZN (signal_456) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_85 ( .s (signal_457), .b ({signal_2280, signal_1677}), .a ({ciphertext_s1[120], ciphertext_s0[120]}), .c ({signal_3250, signal_465}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_88 ( .s (signal_457), .b ({signal_2283, signal_1676}), .a ({ciphertext_s1[121], ciphertext_s0[121]}), .c ({signal_3251, signal_467}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_91 ( .s (signal_457), .b ({signal_2286, signal_1675}), .a ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({signal_3252, signal_469}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_94 ( .s (signal_457), .b ({signal_2289, signal_1674}), .a ({ciphertext_s1[123], ciphertext_s0[123]}), .c ({signal_3253, signal_471}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_97 ( .s (signal_457), .b ({signal_2292, signal_1673}), .a ({ciphertext_s1[124], ciphertext_s0[124]}), .c ({signal_3254, signal_473}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_100 ( .s (signal_457), .b ({signal_2295, signal_1672}), .a ({ciphertext_s1[125], ciphertext_s0[125]}), .c ({signal_3255, signal_475}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_103 ( .s (signal_457), .b ({signal_2298, signal_1671}), .a ({ciphertext_s1[126], ciphertext_s0[126]}), .c ({signal_3256, signal_477}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_106 ( .s (signal_457), .b ({signal_2301, signal_1670}), .a ({ciphertext_s1[127], ciphertext_s0[127]}), .c ({signal_3257, signal_479}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_109 ( .s (signal_457), .b ({signal_2304, signal_1669}), .a ({ciphertext_s1[112], ciphertext_s0[112]}), .c ({signal_3258, signal_481}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_112 ( .s (signal_457), .b ({signal_2307, signal_1668}), .a ({ciphertext_s1[113], ciphertext_s0[113]}), .c ({signal_3259, signal_483}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_115 ( .s (signal_457), .b ({signal_2310, signal_1667}), .a ({ciphertext_s1[114], ciphertext_s0[114]}), .c ({signal_3260, signal_485}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_118 ( .s (signal_457), .b ({signal_2313, signal_1666}), .a ({ciphertext_s1[115], ciphertext_s0[115]}), .c ({signal_3261, signal_487}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_121 ( .s (signal_457), .b ({signal_2316, signal_1665}), .a ({ciphertext_s1[116], ciphertext_s0[116]}), .c ({signal_3262, signal_489}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_124 ( .s (signal_457), .b ({signal_2319, signal_1664}), .a ({ciphertext_s1[117], ciphertext_s0[117]}), .c ({signal_3263, signal_491}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_127 ( .s (signal_457), .b ({signal_2322, signal_1663}), .a ({ciphertext_s1[118], ciphertext_s0[118]}), .c ({signal_3264, signal_493}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_130 ( .s (signal_457), .b ({signal_2325, signal_1662}), .a ({ciphertext_s1[119], ciphertext_s0[119]}), .c ({signal_3265, signal_495}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_133 ( .s (signal_458), .b ({signal_2328, signal_1661}), .a ({ciphertext_s1[104], ciphertext_s0[104]}), .c ({signal_3266, signal_497}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_136 ( .s (signal_458), .b ({signal_2331, signal_1660}), .a ({ciphertext_s1[105], ciphertext_s0[105]}), .c ({signal_3267, signal_499}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_139 ( .s (signal_458), .b ({signal_2334, signal_1659}), .a ({ciphertext_s1[106], ciphertext_s0[106]}), .c ({signal_3268, signal_501}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_142 ( .s (signal_458), .b ({signal_2337, signal_1658}), .a ({ciphertext_s1[107], ciphertext_s0[107]}), .c ({signal_3269, signal_503}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_145 ( .s (signal_458), .b ({signal_2340, signal_1657}), .a ({ciphertext_s1[108], ciphertext_s0[108]}), .c ({signal_3270, signal_505}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_148 ( .s (signal_458), .b ({signal_2343, signal_1656}), .a ({ciphertext_s1[109], ciphertext_s0[109]}), .c ({signal_3271, signal_507}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_151 ( .s (signal_458), .b ({signal_2346, signal_1655}), .a ({ciphertext_s1[110], ciphertext_s0[110]}), .c ({signal_3272, signal_509}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_154 ( .s (signal_458), .b ({signal_2349, signal_1654}), .a ({ciphertext_s1[111], ciphertext_s0[111]}), .c ({signal_3273, signal_511}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_157 ( .s (signal_458), .b ({signal_3170, signal_1653}), .a ({ciphertext_s1[96], ciphertext_s0[96]}), .c ({signal_3274, signal_513}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_160 ( .s (signal_458), .b ({signal_3172, signal_1652}), .a ({ciphertext_s1[97], ciphertext_s0[97]}), .c ({signal_3275, signal_515}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_163 ( .s (signal_458), .b ({signal_3174, signal_1651}), .a ({ciphertext_s1[98], ciphertext_s0[98]}), .c ({signal_3276, signal_517}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_166 ( .s (signal_458), .b ({signal_3176, signal_1650}), .a ({ciphertext_s1[99], ciphertext_s0[99]}), .c ({signal_3277, signal_519}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_169 ( .s (signal_458), .b ({signal_3178, signal_1649}), .a ({ciphertext_s1[100], ciphertext_s0[100]}), .c ({signal_3278, signal_521}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_172 ( .s (signal_458), .b ({signal_3180, signal_1648}), .a ({ciphertext_s1[101], ciphertext_s0[101]}), .c ({signal_3279, signal_523}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_175 ( .s (signal_458), .b ({signal_3182, signal_1647}), .a ({ciphertext_s1[102], ciphertext_s0[102]}), .c ({signal_3280, signal_525}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_178 ( .s (signal_458), .b ({signal_3184, signal_1646}), .a ({ciphertext_s1[103], ciphertext_s0[103]}), .c ({signal_3281, signal_527}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_181 ( .s (signal_459), .b ({signal_2352, signal_1645}), .a ({ciphertext_s1[80], ciphertext_s0[80]}), .c ({signal_3282, signal_529}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_184 ( .s (signal_459), .b ({signal_2355, signal_1644}), .a ({ciphertext_s1[81], ciphertext_s0[81]}), .c ({signal_3283, signal_531}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_187 ( .s (signal_459), .b ({signal_2358, signal_1643}), .a ({ciphertext_s1[82], ciphertext_s0[82]}), .c ({signal_3284, signal_533}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_190 ( .s (signal_459), .b ({signal_2361, signal_1642}), .a ({ciphertext_s1[83], ciphertext_s0[83]}), .c ({signal_3285, signal_535}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_193 ( .s (signal_459), .b ({signal_2364, signal_1641}), .a ({ciphertext_s1[84], ciphertext_s0[84]}), .c ({signal_3286, signal_537}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_196 ( .s (signal_459), .b ({signal_2367, signal_1640}), .a ({ciphertext_s1[85], ciphertext_s0[85]}), .c ({signal_3287, signal_539}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_199 ( .s (signal_459), .b ({signal_2370, signal_1639}), .a ({ciphertext_s1[86], ciphertext_s0[86]}), .c ({signal_3288, signal_541}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_202 ( .s (signal_459), .b ({signal_2373, signal_1638}), .a ({ciphertext_s1[87], ciphertext_s0[87]}), .c ({signal_3289, signal_543}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_205 ( .s (signal_459), .b ({signal_2376, signal_1637}), .a ({ciphertext_s1[72], ciphertext_s0[72]}), .c ({signal_3290, signal_545}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_208 ( .s (signal_459), .b ({signal_2379, signal_1636}), .a ({ciphertext_s1[73], ciphertext_s0[73]}), .c ({signal_3291, signal_547}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_211 ( .s (signal_459), .b ({signal_2382, signal_1635}), .a ({ciphertext_s1[74], ciphertext_s0[74]}), .c ({signal_3292, signal_549}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_214 ( .s (signal_459), .b ({signal_2385, signal_1634}), .a ({ciphertext_s1[75], ciphertext_s0[75]}), .c ({signal_3293, signal_551}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_217 ( .s (signal_459), .b ({signal_2388, signal_1633}), .a ({ciphertext_s1[76], ciphertext_s0[76]}), .c ({signal_3294, signal_553}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_220 ( .s (signal_459), .b ({signal_2391, signal_1632}), .a ({ciphertext_s1[77], ciphertext_s0[77]}), .c ({signal_3295, signal_555}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_223 ( .s (signal_459), .b ({signal_2394, signal_1631}), .a ({ciphertext_s1[78], ciphertext_s0[78]}), .c ({signal_3296, signal_557}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_226 ( .s (signal_459), .b ({signal_2397, signal_1630}), .a ({ciphertext_s1[79], ciphertext_s0[79]}), .c ({signal_3297, signal_559}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_229 ( .s (signal_460), .b ({signal_2400, signal_1629}), .a ({ciphertext_s1[64], ciphertext_s0[64]}), .c ({signal_3298, signal_561}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_232 ( .s (signal_460), .b ({signal_2403, signal_1628}), .a ({ciphertext_s1[65], ciphertext_s0[65]}), .c ({signal_3299, signal_563}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_235 ( .s (signal_460), .b ({signal_2406, signal_1627}), .a ({ciphertext_s1[66], ciphertext_s0[66]}), .c ({signal_3300, signal_565}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_238 ( .s (signal_460), .b ({signal_2409, signal_1626}), .a ({ciphertext_s1[67], ciphertext_s0[67]}), .c ({signal_3301, signal_567}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_241 ( .s (signal_460), .b ({signal_2412, signal_1625}), .a ({ciphertext_s1[68], ciphertext_s0[68]}), .c ({signal_3302, signal_569}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_244 ( .s (signal_460), .b ({signal_2415, signal_1624}), .a ({ciphertext_s1[69], ciphertext_s0[69]}), .c ({signal_3303, signal_571}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_247 ( .s (signal_460), .b ({signal_2418, signal_1623}), .a ({ciphertext_s1[70], ciphertext_s0[70]}), .c ({signal_3304, signal_573}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_250 ( .s (signal_460), .b ({signal_2421, signal_1622}), .a ({ciphertext_s1[71], ciphertext_s0[71]}), .c ({signal_3305, signal_575}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_253 ( .s (signal_460), .b ({signal_3186, signal_1621}), .a ({ciphertext_s1[88], ciphertext_s0[88]}), .c ({signal_3306, signal_577}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_256 ( .s (signal_460), .b ({signal_3188, signal_1620}), .a ({ciphertext_s1[89], ciphertext_s0[89]}), .c ({signal_3307, signal_579}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_259 ( .s (signal_460), .b ({signal_3190, signal_1619}), .a ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({signal_3308, signal_581}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_262 ( .s (signal_460), .b ({signal_3192, signal_1618}), .a ({ciphertext_s1[91], ciphertext_s0[91]}), .c ({signal_3309, signal_583}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_265 ( .s (signal_460), .b ({signal_3194, signal_1617}), .a ({ciphertext_s1[92], ciphertext_s0[92]}), .c ({signal_3310, signal_585}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_268 ( .s (signal_460), .b ({signal_3196, signal_1616}), .a ({ciphertext_s1[93], ciphertext_s0[93]}), .c ({signal_3311, signal_587}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_271 ( .s (signal_460), .b ({signal_3198, signal_1615}), .a ({ciphertext_s1[94], ciphertext_s0[94]}), .c ({signal_3312, signal_589}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_274 ( .s (signal_460), .b ({signal_3200, signal_1614}), .a ({ciphertext_s1[95], ciphertext_s0[95]}), .c ({signal_3313, signal_591}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_277 ( .s (signal_461), .b ({signal_2424, signal_1613}), .a ({ciphertext_s1[40], ciphertext_s0[40]}), .c ({signal_3314, signal_593}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_280 ( .s (signal_461), .b ({signal_2427, signal_1612}), .a ({ciphertext_s1[41], ciphertext_s0[41]}), .c ({signal_3315, signal_595}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_283 ( .s (signal_461), .b ({signal_2430, signal_1611}), .a ({ciphertext_s1[42], ciphertext_s0[42]}), .c ({signal_3316, signal_597}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_286 ( .s (signal_461), .b ({signal_2433, signal_1610}), .a ({ciphertext_s1[43], ciphertext_s0[43]}), .c ({signal_3317, signal_599}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_289 ( .s (signal_461), .b ({signal_2436, signal_1609}), .a ({ciphertext_s1[44], ciphertext_s0[44]}), .c ({signal_3318, signal_601}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_292 ( .s (signal_461), .b ({signal_2439, signal_1608}), .a ({ciphertext_s1[45], ciphertext_s0[45]}), .c ({signal_3319, signal_603}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_295 ( .s (signal_461), .b ({signal_2442, signal_1607}), .a ({ciphertext_s1[46], ciphertext_s0[46]}), .c ({signal_3320, signal_605}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_298 ( .s (signal_461), .b ({signal_2445, signal_1606}), .a ({ciphertext_s1[47], ciphertext_s0[47]}), .c ({signal_3321, signal_607}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_301 ( .s (signal_461), .b ({signal_2448, signal_1605}), .a ({ciphertext_s1[32], ciphertext_s0[32]}), .c ({signal_3322, signal_609}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_304 ( .s (signal_461), .b ({signal_2451, signal_1604}), .a ({ciphertext_s1[33], ciphertext_s0[33]}), .c ({signal_3323, signal_611}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_307 ( .s (signal_461), .b ({signal_2454, signal_1603}), .a ({ciphertext_s1[34], ciphertext_s0[34]}), .c ({signal_3324, signal_613}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_310 ( .s (signal_461), .b ({signal_2457, signal_1602}), .a ({ciphertext_s1[35], ciphertext_s0[35]}), .c ({signal_3325, signal_615}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_313 ( .s (signal_461), .b ({signal_2460, signal_1601}), .a ({ciphertext_s1[36], ciphertext_s0[36]}), .c ({signal_3326, signal_617}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_316 ( .s (signal_461), .b ({signal_2463, signal_1600}), .a ({ciphertext_s1[37], ciphertext_s0[37]}), .c ({signal_3327, signal_619}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_319 ( .s (signal_461), .b ({signal_2466, signal_1599}), .a ({ciphertext_s1[38], ciphertext_s0[38]}), .c ({signal_3328, signal_621}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_322 ( .s (signal_461), .b ({signal_2469, signal_1598}), .a ({ciphertext_s1[39], ciphertext_s0[39]}), .c ({signal_3329, signal_623}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_325 ( .s (signal_462), .b ({signal_2472, signal_1597}), .a ({ciphertext_s1[56], ciphertext_s0[56]}), .c ({signal_3330, signal_625}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_328 ( .s (signal_462), .b ({signal_2475, signal_1596}), .a ({ciphertext_s1[57], ciphertext_s0[57]}), .c ({signal_3331, signal_627}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_331 ( .s (signal_462), .b ({signal_2478, signal_1595}), .a ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({signal_3332, signal_629}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_334 ( .s (signal_462), .b ({signal_2481, signal_1594}), .a ({ciphertext_s1[59], ciphertext_s0[59]}), .c ({signal_3333, signal_631}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_337 ( .s (signal_462), .b ({signal_2484, signal_1593}), .a ({ciphertext_s1[60], ciphertext_s0[60]}), .c ({signal_3334, signal_633}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_340 ( .s (signal_462), .b ({signal_2487, signal_1592}), .a ({ciphertext_s1[61], ciphertext_s0[61]}), .c ({signal_3335, signal_635}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_343 ( .s (signal_462), .b ({signal_2490, signal_1591}), .a ({ciphertext_s1[62], ciphertext_s0[62]}), .c ({signal_3336, signal_637}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_346 ( .s (signal_462), .b ({signal_2493, signal_1590}), .a ({ciphertext_s1[63], ciphertext_s0[63]}), .c ({signal_3337, signal_639}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_349 ( .s (signal_462), .b ({signal_3202, signal_1589}), .a ({ciphertext_s1[48], ciphertext_s0[48]}), .c ({signal_3338, signal_641}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_352 ( .s (signal_462), .b ({signal_3204, signal_1588}), .a ({ciphertext_s1[49], ciphertext_s0[49]}), .c ({signal_3339, signal_643}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_355 ( .s (signal_462), .b ({signal_3206, signal_1587}), .a ({ciphertext_s1[50], ciphertext_s0[50]}), .c ({signal_3340, signal_645}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_358 ( .s (signal_462), .b ({signal_3208, signal_1586}), .a ({ciphertext_s1[51], ciphertext_s0[51]}), .c ({signal_3341, signal_647}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_361 ( .s (signal_462), .b ({signal_3210, signal_1585}), .a ({ciphertext_s1[52], ciphertext_s0[52]}), .c ({signal_3342, signal_649}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_364 ( .s (signal_462), .b ({signal_3212, signal_1584}), .a ({ciphertext_s1[53], ciphertext_s0[53]}), .c ({signal_3343, signal_651}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_367 ( .s (signal_462), .b ({signal_3214, signal_1583}), .a ({ciphertext_s1[54], ciphertext_s0[54]}), .c ({signal_3344, signal_653}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_370 ( .s (signal_462), .b ({signal_3216, signal_1582}), .a ({ciphertext_s1[55], ciphertext_s0[55]}), .c ({signal_3345, signal_655}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_373 ( .s (signal_463), .b ({signal_2496, signal_1581}), .a ({ciphertext_s1[0], ciphertext_s0[0]}), .c ({signal_3346, signal_657}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_376 ( .s (signal_463), .b ({signal_2499, signal_1580}), .a ({ciphertext_s1[1], ciphertext_s0[1]}), .c ({signal_3347, signal_659}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_379 ( .s (signal_463), .b ({signal_2502, signal_1579}), .a ({ciphertext_s1[2], ciphertext_s0[2]}), .c ({signal_3348, signal_661}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_382 ( .s (signal_463), .b ({signal_2505, signal_1578}), .a ({ciphertext_s1[3], ciphertext_s0[3]}), .c ({signal_3349, signal_663}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_385 ( .s (signal_463), .b ({signal_2508, signal_1577}), .a ({ciphertext_s1[4], ciphertext_s0[4]}), .c ({signal_3350, signal_665}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_388 ( .s (signal_463), .b ({signal_2511, signal_1576}), .a ({ciphertext_s1[5], ciphertext_s0[5]}), .c ({signal_3351, signal_667}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_391 ( .s (signal_463), .b ({signal_2514, signal_1575}), .a ({ciphertext_s1[6], ciphertext_s0[6]}), .c ({signal_3352, signal_669}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_394 ( .s (signal_463), .b ({signal_2517, signal_1574}), .a ({ciphertext_s1[7], ciphertext_s0[7]}), .c ({signal_3353, signal_671}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_397 ( .s (signal_463), .b ({signal_2520, signal_1573}), .a ({ciphertext_s1[24], ciphertext_s0[24]}), .c ({signal_3354, signal_673}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_400 ( .s (signal_463), .b ({signal_2523, signal_1572}), .a ({ciphertext_s1[25], ciphertext_s0[25]}), .c ({signal_3355, signal_675}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_403 ( .s (signal_463), .b ({signal_2526, signal_1571}), .a ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({signal_3356, signal_677}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_406 ( .s (signal_463), .b ({signal_2529, signal_1570}), .a ({ciphertext_s1[27], ciphertext_s0[27]}), .c ({signal_3357, signal_679}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_409 ( .s (signal_463), .b ({signal_2532, signal_1569}), .a ({ciphertext_s1[28], ciphertext_s0[28]}), .c ({signal_3358, signal_681}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_412 ( .s (signal_463), .b ({signal_2535, signal_1568}), .a ({ciphertext_s1[29], ciphertext_s0[29]}), .c ({signal_3359, signal_683}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_415 ( .s (signal_463), .b ({signal_2538, signal_1567}), .a ({ciphertext_s1[30], ciphertext_s0[30]}), .c ({signal_3360, signal_685}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_418 ( .s (signal_463), .b ({signal_2541, signal_1566}), .a ({ciphertext_s1[31], ciphertext_s0[31]}), .c ({signal_3361, signal_687}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_421 ( .s (signal_464), .b ({signal_2544, signal_1565}), .a ({ciphertext_s1[16], ciphertext_s0[16]}), .c ({signal_3362, signal_689}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_424 ( .s (signal_464), .b ({signal_2547, signal_1564}), .a ({ciphertext_s1[17], ciphertext_s0[17]}), .c ({signal_3363, signal_691}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_427 ( .s (signal_464), .b ({signal_2550, signal_1563}), .a ({ciphertext_s1[18], ciphertext_s0[18]}), .c ({signal_3364, signal_693}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_430 ( .s (signal_464), .b ({signal_2553, signal_1562}), .a ({ciphertext_s1[19], ciphertext_s0[19]}), .c ({signal_3365, signal_695}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_433 ( .s (signal_464), .b ({signal_2556, signal_1561}), .a ({ciphertext_s1[20], ciphertext_s0[20]}), .c ({signal_3366, signal_697}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_436 ( .s (signal_464), .b ({signal_2559, signal_1560}), .a ({ciphertext_s1[21], ciphertext_s0[21]}), .c ({signal_3367, signal_699}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_439 ( .s (signal_464), .b ({signal_2562, signal_1559}), .a ({ciphertext_s1[22], ciphertext_s0[22]}), .c ({signal_3368, signal_701}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_442 ( .s (signal_464), .b ({signal_2565, signal_1558}), .a ({ciphertext_s1[23], ciphertext_s0[23]}), .c ({signal_3369, signal_703}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_469 ( .s (signal_445), .b ({plaintext_s1[120], plaintext_s0[120]}), .a ({ciphertext_s1[112], ciphertext_s0[112]}), .c ({signal_2280, signal_1677}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_470 ( .s (signal_445), .b ({plaintext_s1[121], plaintext_s0[121]}), .a ({ciphertext_s1[113], ciphertext_s0[113]}), .c ({signal_2283, signal_1676}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_471 ( .s (signal_445), .b ({plaintext_s1[122], plaintext_s0[122]}), .a ({ciphertext_s1[114], ciphertext_s0[114]}), .c ({signal_2286, signal_1675}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_472 ( .s (signal_445), .b ({plaintext_s1[123], plaintext_s0[123]}), .a ({ciphertext_s1[115], ciphertext_s0[115]}), .c ({signal_2289, signal_1674}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_473 ( .s (signal_445), .b ({plaintext_s1[124], plaintext_s0[124]}), .a ({ciphertext_s1[116], ciphertext_s0[116]}), .c ({signal_2292, signal_1673}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_474 ( .s (signal_445), .b ({plaintext_s1[125], plaintext_s0[125]}), .a ({ciphertext_s1[117], ciphertext_s0[117]}), .c ({signal_2295, signal_1672}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_475 ( .s (signal_445), .b ({plaintext_s1[126], plaintext_s0[126]}), .a ({ciphertext_s1[118], ciphertext_s0[118]}), .c ({signal_2298, signal_1671}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_476 ( .s (signal_445), .b ({plaintext_s1[127], plaintext_s0[127]}), .a ({ciphertext_s1[119], ciphertext_s0[119]}), .c ({signal_2301, signal_1670}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_477 ( .s (signal_445), .b ({plaintext_s1[112], plaintext_s0[112]}), .a ({ciphertext_s1[104], ciphertext_s0[104]}), .c ({signal_2304, signal_1669}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_478 ( .s (signal_445), .b ({plaintext_s1[113], plaintext_s0[113]}), .a ({ciphertext_s1[105], ciphertext_s0[105]}), .c ({signal_2307, signal_1668}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_479 ( .s (signal_445), .b ({plaintext_s1[114], plaintext_s0[114]}), .a ({ciphertext_s1[106], ciphertext_s0[106]}), .c ({signal_2310, signal_1667}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_480 ( .s (signal_445), .b ({plaintext_s1[115], plaintext_s0[115]}), .a ({ciphertext_s1[107], ciphertext_s0[107]}), .c ({signal_2313, signal_1666}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_481 ( .s (signal_445), .b ({plaintext_s1[116], plaintext_s0[116]}), .a ({ciphertext_s1[108], ciphertext_s0[108]}), .c ({signal_2316, signal_1665}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_482 ( .s (signal_445), .b ({plaintext_s1[117], plaintext_s0[117]}), .a ({ciphertext_s1[109], ciphertext_s0[109]}), .c ({signal_2319, signal_1664}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_483 ( .s (signal_445), .b ({plaintext_s1[118], plaintext_s0[118]}), .a ({ciphertext_s1[110], ciphertext_s0[110]}), .c ({signal_2322, signal_1663}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_484 ( .s (signal_445), .b ({plaintext_s1[119], plaintext_s0[119]}), .a ({ciphertext_s1[111], ciphertext_s0[111]}), .c ({signal_2325, signal_1662}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_485 ( .s (signal_446), .b ({plaintext_s1[104], plaintext_s0[104]}), .a ({ciphertext_s1[96], ciphertext_s0[96]}), .c ({signal_2328, signal_1661}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_486 ( .s (signal_446), .b ({plaintext_s1[105], plaintext_s0[105]}), .a ({ciphertext_s1[97], ciphertext_s0[97]}), .c ({signal_2331, signal_1660}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_487 ( .s (signal_446), .b ({plaintext_s1[106], plaintext_s0[106]}), .a ({ciphertext_s1[98], ciphertext_s0[98]}), .c ({signal_2334, signal_1659}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_488 ( .s (signal_446), .b ({plaintext_s1[107], plaintext_s0[107]}), .a ({ciphertext_s1[99], ciphertext_s0[99]}), .c ({signal_2337, signal_1658}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_489 ( .s (signal_446), .b ({plaintext_s1[108], plaintext_s0[108]}), .a ({ciphertext_s1[100], ciphertext_s0[100]}), .c ({signal_2340, signal_1657}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_490 ( .s (signal_446), .b ({plaintext_s1[109], plaintext_s0[109]}), .a ({ciphertext_s1[101], ciphertext_s0[101]}), .c ({signal_2343, signal_1656}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_491 ( .s (signal_446), .b ({plaintext_s1[110], plaintext_s0[110]}), .a ({ciphertext_s1[102], ciphertext_s0[102]}), .c ({signal_2346, signal_1655}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_492 ( .s (signal_446), .b ({plaintext_s1[111], plaintext_s0[111]}), .a ({ciphertext_s1[103], ciphertext_s0[103]}), .c ({signal_2349, signal_1654}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_493 ( .s (signal_454), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .a ({signal_3004, signal_1429}), .c ({signal_3132, signal_1549}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_494 ( .s (signal_454), .b ({ciphertext_s1[89], ciphertext_s0[89]}), .a ({signal_3005, signal_1428}), .c ({signal_3133, signal_1548}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_495 ( .s (signal_454), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .a ({signal_3006, signal_1427}), .c ({signal_3134, signal_1547}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_496 ( .s (signal_454), .b ({ciphertext_s1[91], ciphertext_s0[91]}), .a ({signal_3007, signal_1426}), .c ({signal_3135, signal_1546}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_497 ( .s (signal_454), .b ({ciphertext_s1[92], ciphertext_s0[92]}), .a ({signal_3008, signal_1425}), .c ({signal_3136, signal_1545}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_498 ( .s (signal_454), .b ({ciphertext_s1[93], ciphertext_s0[93]}), .a ({signal_3009, signal_1424}), .c ({signal_3137, signal_1544}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_499 ( .s (signal_454), .b ({ciphertext_s1[94], ciphertext_s0[94]}), .a ({signal_3010, signal_1423}), .c ({signal_3138, signal_1543}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_500 ( .s (signal_454), .b ({ciphertext_s1[95], ciphertext_s0[95]}), .a ({signal_3011, signal_1422}), .c ({signal_3139, signal_1542}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_501 ( .s (signal_446), .b ({plaintext_s1[96], plaintext_s0[96]}), .a ({signal_3132, signal_1549}), .c ({signal_3170, signal_1653}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_502 ( .s (signal_446), .b ({plaintext_s1[97], plaintext_s0[97]}), .a ({signal_3133, signal_1548}), .c ({signal_3172, signal_1652}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_503 ( .s (signal_446), .b ({plaintext_s1[98], plaintext_s0[98]}), .a ({signal_3134, signal_1547}), .c ({signal_3174, signal_1651}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_504 ( .s (signal_446), .b ({plaintext_s1[99], plaintext_s0[99]}), .a ({signal_3135, signal_1546}), .c ({signal_3176, signal_1650}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_505 ( .s (signal_446), .b ({plaintext_s1[100], plaintext_s0[100]}), .a ({signal_3136, signal_1545}), .c ({signal_3178, signal_1649}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_506 ( .s (signal_446), .b ({plaintext_s1[101], plaintext_s0[101]}), .a ({signal_3137, signal_1544}), .c ({signal_3180, signal_1648}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_507 ( .s (signal_446), .b ({plaintext_s1[102], plaintext_s0[102]}), .a ({signal_3138, signal_1543}), .c ({signal_3182, signal_1647}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_508 ( .s (signal_446), .b ({plaintext_s1[103], plaintext_s0[103]}), .a ({signal_3139, signal_1542}), .c ({signal_3184, signal_1646}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_509 ( .s (signal_447), .b ({plaintext_s1[88], plaintext_s0[88]}), .a ({ciphertext_s1[80], ciphertext_s0[80]}), .c ({signal_2352, signal_1645}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_510 ( .s (signal_447), .b ({plaintext_s1[89], plaintext_s0[89]}), .a ({ciphertext_s1[81], ciphertext_s0[81]}), .c ({signal_2355, signal_1644}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_511 ( .s (signal_447), .b ({plaintext_s1[90], plaintext_s0[90]}), .a ({ciphertext_s1[82], ciphertext_s0[82]}), .c ({signal_2358, signal_1643}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_512 ( .s (signal_447), .b ({plaintext_s1[91], plaintext_s0[91]}), .a ({ciphertext_s1[83], ciphertext_s0[83]}), .c ({signal_2361, signal_1642}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_513 ( .s (signal_447), .b ({plaintext_s1[92], plaintext_s0[92]}), .a ({ciphertext_s1[84], ciphertext_s0[84]}), .c ({signal_2364, signal_1641}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_514 ( .s (signal_447), .b ({plaintext_s1[93], plaintext_s0[93]}), .a ({ciphertext_s1[85], ciphertext_s0[85]}), .c ({signal_2367, signal_1640}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_515 ( .s (signal_447), .b ({plaintext_s1[94], plaintext_s0[94]}), .a ({ciphertext_s1[86], ciphertext_s0[86]}), .c ({signal_2370, signal_1639}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_516 ( .s (signal_447), .b ({plaintext_s1[95], plaintext_s0[95]}), .a ({ciphertext_s1[87], ciphertext_s0[87]}), .c ({signal_2373, signal_1638}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_517 ( .s (signal_447), .b ({plaintext_s1[80], plaintext_s0[80]}), .a ({ciphertext_s1[72], ciphertext_s0[72]}), .c ({signal_2376, signal_1637}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_518 ( .s (signal_447), .b ({plaintext_s1[81], plaintext_s0[81]}), .a ({ciphertext_s1[73], ciphertext_s0[73]}), .c ({signal_2379, signal_1636}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_519 ( .s (signal_447), .b ({plaintext_s1[82], plaintext_s0[82]}), .a ({ciphertext_s1[74], ciphertext_s0[74]}), .c ({signal_2382, signal_1635}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_520 ( .s (signal_447), .b ({plaintext_s1[83], plaintext_s0[83]}), .a ({ciphertext_s1[75], ciphertext_s0[75]}), .c ({signal_2385, signal_1634}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_521 ( .s (signal_447), .b ({plaintext_s1[84], plaintext_s0[84]}), .a ({ciphertext_s1[76], ciphertext_s0[76]}), .c ({signal_2388, signal_1633}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_522 ( .s (signal_447), .b ({plaintext_s1[85], plaintext_s0[85]}), .a ({ciphertext_s1[77], ciphertext_s0[77]}), .c ({signal_2391, signal_1632}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_523 ( .s (signal_447), .b ({plaintext_s1[86], plaintext_s0[86]}), .a ({ciphertext_s1[78], ciphertext_s0[78]}), .c ({signal_2394, signal_1631}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_524 ( .s (signal_447), .b ({plaintext_s1[87], plaintext_s0[87]}), .a ({ciphertext_s1[79], ciphertext_s0[79]}), .c ({signal_2397, signal_1630}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_525 ( .s (signal_448), .b ({plaintext_s1[72], plaintext_s0[72]}), .a ({ciphertext_s1[64], ciphertext_s0[64]}), .c ({signal_2400, signal_1629}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_526 ( .s (signal_448), .b ({plaintext_s1[73], plaintext_s0[73]}), .a ({ciphertext_s1[65], ciphertext_s0[65]}), .c ({signal_2403, signal_1628}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_527 ( .s (signal_448), .b ({plaintext_s1[74], plaintext_s0[74]}), .a ({ciphertext_s1[66], ciphertext_s0[66]}), .c ({signal_2406, signal_1627}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_528 ( .s (signal_448), .b ({plaintext_s1[75], plaintext_s0[75]}), .a ({ciphertext_s1[67], ciphertext_s0[67]}), .c ({signal_2409, signal_1626}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_529 ( .s (signal_448), .b ({plaintext_s1[76], plaintext_s0[76]}), .a ({ciphertext_s1[68], ciphertext_s0[68]}), .c ({signal_2412, signal_1625}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_530 ( .s (signal_448), .b ({plaintext_s1[77], plaintext_s0[77]}), .a ({ciphertext_s1[69], ciphertext_s0[69]}), .c ({signal_2415, signal_1624}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_531 ( .s (signal_448), .b ({plaintext_s1[78], plaintext_s0[78]}), .a ({ciphertext_s1[70], ciphertext_s0[70]}), .c ({signal_2418, signal_1623}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_532 ( .s (signal_448), .b ({plaintext_s1[79], plaintext_s0[79]}), .a ({ciphertext_s1[71], ciphertext_s0[71]}), .c ({signal_2421, signal_1622}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_533 ( .s (signal_454), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .a ({signal_2996, signal_1437}), .c ({signal_3140, signal_1541}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_534 ( .s (signal_454), .b ({ciphertext_s1[57], ciphertext_s0[57]}), .a ({signal_2997, signal_1436}), .c ({signal_3141, signal_1540}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_535 ( .s (signal_454), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .a ({signal_2998, signal_1435}), .c ({signal_3142, signal_1539}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_536 ( .s (signal_454), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .a ({signal_2999, signal_1434}), .c ({signal_3143, signal_1538}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_537 ( .s (signal_454), .b ({ciphertext_s1[60], ciphertext_s0[60]}), .a ({signal_3000, signal_1433}), .c ({signal_3144, signal_1537}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_538 ( .s (signal_454), .b ({ciphertext_s1[61], ciphertext_s0[61]}), .a ({signal_3001, signal_1432}), .c ({signal_3145, signal_1536}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_539 ( .s (signal_454), .b ({ciphertext_s1[62], ciphertext_s0[62]}), .a ({signal_3002, signal_1431}), .c ({signal_3146, signal_1535}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_540 ( .s (signal_454), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .a ({signal_3003, signal_1430}), .c ({signal_3147, signal_1534}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_541 ( .s (signal_448), .b ({plaintext_s1[64], plaintext_s0[64]}), .a ({signal_3140, signal_1541}), .c ({signal_3186, signal_1621}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_542 ( .s (signal_448), .b ({plaintext_s1[65], plaintext_s0[65]}), .a ({signal_3141, signal_1540}), .c ({signal_3188, signal_1620}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_543 ( .s (signal_448), .b ({plaintext_s1[66], plaintext_s0[66]}), .a ({signal_3142, signal_1539}), .c ({signal_3190, signal_1619}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_544 ( .s (signal_448), .b ({plaintext_s1[67], plaintext_s0[67]}), .a ({signal_3143, signal_1538}), .c ({signal_3192, signal_1618}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_545 ( .s (signal_448), .b ({plaintext_s1[68], plaintext_s0[68]}), .a ({signal_3144, signal_1537}), .c ({signal_3194, signal_1617}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_546 ( .s (signal_448), .b ({plaintext_s1[69], plaintext_s0[69]}), .a ({signal_3145, signal_1536}), .c ({signal_3196, signal_1616}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_547 ( .s (signal_448), .b ({plaintext_s1[70], plaintext_s0[70]}), .a ({signal_3146, signal_1535}), .c ({signal_3198, signal_1615}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_548 ( .s (signal_448), .b ({plaintext_s1[71], plaintext_s0[71]}), .a ({signal_3147, signal_1534}), .c ({signal_3200, signal_1614}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_549 ( .s (signal_449), .b ({plaintext_s1[56], plaintext_s0[56]}), .a ({ciphertext_s1[48], ciphertext_s0[48]}), .c ({signal_2424, signal_1613}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_550 ( .s (signal_449), .b ({plaintext_s1[57], plaintext_s0[57]}), .a ({ciphertext_s1[49], ciphertext_s0[49]}), .c ({signal_2427, signal_1612}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_551 ( .s (signal_449), .b ({plaintext_s1[58], plaintext_s0[58]}), .a ({ciphertext_s1[50], ciphertext_s0[50]}), .c ({signal_2430, signal_1611}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_552 ( .s (signal_449), .b ({plaintext_s1[59], plaintext_s0[59]}), .a ({ciphertext_s1[51], ciphertext_s0[51]}), .c ({signal_2433, signal_1610}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_553 ( .s (signal_449), .b ({plaintext_s1[60], plaintext_s0[60]}), .a ({ciphertext_s1[52], ciphertext_s0[52]}), .c ({signal_2436, signal_1609}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_554 ( .s (signal_449), .b ({plaintext_s1[61], plaintext_s0[61]}), .a ({ciphertext_s1[53], ciphertext_s0[53]}), .c ({signal_2439, signal_1608}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_555 ( .s (signal_449), .b ({plaintext_s1[62], plaintext_s0[62]}), .a ({ciphertext_s1[54], ciphertext_s0[54]}), .c ({signal_2442, signal_1607}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_556 ( .s (signal_449), .b ({plaintext_s1[63], plaintext_s0[63]}), .a ({ciphertext_s1[55], ciphertext_s0[55]}), .c ({signal_2445, signal_1606}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_557 ( .s (signal_449), .b ({plaintext_s1[48], plaintext_s0[48]}), .a ({ciphertext_s1[40], ciphertext_s0[40]}), .c ({signal_2448, signal_1605}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_558 ( .s (signal_449), .b ({plaintext_s1[49], plaintext_s0[49]}), .a ({ciphertext_s1[41], ciphertext_s0[41]}), .c ({signal_2451, signal_1604}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_559 ( .s (signal_449), .b ({plaintext_s1[50], plaintext_s0[50]}), .a ({ciphertext_s1[42], ciphertext_s0[42]}), .c ({signal_2454, signal_1603}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_560 ( .s (signal_449), .b ({plaintext_s1[51], plaintext_s0[51]}), .a ({ciphertext_s1[43], ciphertext_s0[43]}), .c ({signal_2457, signal_1602}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_561 ( .s (signal_449), .b ({plaintext_s1[52], plaintext_s0[52]}), .a ({ciphertext_s1[44], ciphertext_s0[44]}), .c ({signal_2460, signal_1601}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_562 ( .s (signal_449), .b ({plaintext_s1[53], plaintext_s0[53]}), .a ({ciphertext_s1[45], ciphertext_s0[45]}), .c ({signal_2463, signal_1600}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_563 ( .s (signal_449), .b ({plaintext_s1[54], plaintext_s0[54]}), .a ({ciphertext_s1[46], ciphertext_s0[46]}), .c ({signal_2466, signal_1599}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_564 ( .s (signal_449), .b ({plaintext_s1[55], plaintext_s0[55]}), .a ({ciphertext_s1[47], ciphertext_s0[47]}), .c ({signal_2469, signal_1598}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_565 ( .s (signal_450), .b ({plaintext_s1[40], plaintext_s0[40]}), .a ({ciphertext_s1[32], ciphertext_s0[32]}), .c ({signal_2472, signal_1597}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_566 ( .s (signal_450), .b ({plaintext_s1[41], plaintext_s0[41]}), .a ({ciphertext_s1[33], ciphertext_s0[33]}), .c ({signal_2475, signal_1596}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_567 ( .s (signal_450), .b ({plaintext_s1[42], plaintext_s0[42]}), .a ({ciphertext_s1[34], ciphertext_s0[34]}), .c ({signal_2478, signal_1595}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_568 ( .s (signal_450), .b ({plaintext_s1[43], plaintext_s0[43]}), .a ({ciphertext_s1[35], ciphertext_s0[35]}), .c ({signal_2481, signal_1594}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_569 ( .s (signal_450), .b ({plaintext_s1[44], plaintext_s0[44]}), .a ({ciphertext_s1[36], ciphertext_s0[36]}), .c ({signal_2484, signal_1593}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_570 ( .s (signal_450), .b ({plaintext_s1[45], plaintext_s0[45]}), .a ({ciphertext_s1[37], ciphertext_s0[37]}), .c ({signal_2487, signal_1592}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_571 ( .s (signal_450), .b ({plaintext_s1[46], plaintext_s0[46]}), .a ({ciphertext_s1[38], ciphertext_s0[38]}), .c ({signal_2490, signal_1591}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_572 ( .s (signal_450), .b ({plaintext_s1[47], plaintext_s0[47]}), .a ({ciphertext_s1[39], ciphertext_s0[39]}), .c ({signal_2493, signal_1590}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_573 ( .s (signal_455), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .a ({signal_2988, signal_1445}), .c ({signal_3148, signal_1533}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_574 ( .s (signal_455), .b ({ciphertext_s1[25], ciphertext_s0[25]}), .a ({signal_2989, signal_1444}), .c ({signal_3149, signal_1532}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_575 ( .s (signal_455), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .a ({signal_2990, signal_1443}), .c ({signal_3150, signal_1531}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_576 ( .s (signal_455), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .a ({signal_2991, signal_1442}), .c ({signal_3151, signal_1530}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_577 ( .s (signal_455), .b ({ciphertext_s1[28], ciphertext_s0[28]}), .a ({signal_2992, signal_1441}), .c ({signal_3152, signal_1529}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_578 ( .s (signal_455), .b ({ciphertext_s1[29], ciphertext_s0[29]}), .a ({signal_2993, signal_1440}), .c ({signal_3153, signal_1528}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_579 ( .s (signal_455), .b ({ciphertext_s1[30], ciphertext_s0[30]}), .a ({signal_2994, signal_1439}), .c ({signal_3154, signal_1527}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_580 ( .s (signal_455), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .a ({signal_2995, signal_1438}), .c ({signal_3155, signal_1526}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_581 ( .s (signal_450), .b ({plaintext_s1[32], plaintext_s0[32]}), .a ({signal_3148, signal_1533}), .c ({signal_3202, signal_1589}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_582 ( .s (signal_450), .b ({plaintext_s1[33], plaintext_s0[33]}), .a ({signal_3149, signal_1532}), .c ({signal_3204, signal_1588}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_583 ( .s (signal_450), .b ({plaintext_s1[34], plaintext_s0[34]}), .a ({signal_3150, signal_1531}), .c ({signal_3206, signal_1587}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_584 ( .s (signal_450), .b ({plaintext_s1[35], plaintext_s0[35]}), .a ({signal_3151, signal_1530}), .c ({signal_3208, signal_1586}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_585 ( .s (signal_450), .b ({plaintext_s1[36], plaintext_s0[36]}), .a ({signal_3152, signal_1529}), .c ({signal_3210, signal_1585}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_586 ( .s (signal_450), .b ({plaintext_s1[37], plaintext_s0[37]}), .a ({signal_3153, signal_1528}), .c ({signal_3212, signal_1584}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_587 ( .s (signal_450), .b ({plaintext_s1[38], plaintext_s0[38]}), .a ({signal_3154, signal_1527}), .c ({signal_3214, signal_1583}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_588 ( .s (signal_450), .b ({plaintext_s1[39], plaintext_s0[39]}), .a ({signal_3155, signal_1526}), .c ({signal_3216, signal_1582}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_589 ( .s (signal_451), .b ({plaintext_s1[24], plaintext_s0[24]}), .a ({ciphertext_s1[16], ciphertext_s0[16]}), .c ({signal_2496, signal_1581}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_590 ( .s (signal_451), .b ({plaintext_s1[25], plaintext_s0[25]}), .a ({ciphertext_s1[17], ciphertext_s0[17]}), .c ({signal_2499, signal_1580}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_591 ( .s (signal_451), .b ({plaintext_s1[26], plaintext_s0[26]}), .a ({ciphertext_s1[18], ciphertext_s0[18]}), .c ({signal_2502, signal_1579}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_592 ( .s (signal_451), .b ({plaintext_s1[27], plaintext_s0[27]}), .a ({ciphertext_s1[19], ciphertext_s0[19]}), .c ({signal_2505, signal_1578}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_593 ( .s (signal_451), .b ({plaintext_s1[28], plaintext_s0[28]}), .a ({ciphertext_s1[20], ciphertext_s0[20]}), .c ({signal_2508, signal_1577}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_594 ( .s (signal_451), .b ({plaintext_s1[29], plaintext_s0[29]}), .a ({ciphertext_s1[21], ciphertext_s0[21]}), .c ({signal_2511, signal_1576}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_595 ( .s (signal_451), .b ({plaintext_s1[30], plaintext_s0[30]}), .a ({ciphertext_s1[22], ciphertext_s0[22]}), .c ({signal_2514, signal_1575}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_596 ( .s (signal_451), .b ({plaintext_s1[31], plaintext_s0[31]}), .a ({ciphertext_s1[23], ciphertext_s0[23]}), .c ({signal_2517, signal_1574}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_597 ( .s (signal_451), .b ({plaintext_s1[16], plaintext_s0[16]}), .a ({ciphertext_s1[8], ciphertext_s0[8]}), .c ({signal_2520, signal_1573}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_598 ( .s (signal_451), .b ({plaintext_s1[17], plaintext_s0[17]}), .a ({ciphertext_s1[9], ciphertext_s0[9]}), .c ({signal_2523, signal_1572}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_599 ( .s (signal_451), .b ({plaintext_s1[18], plaintext_s0[18]}), .a ({ciphertext_s1[10], ciphertext_s0[10]}), .c ({signal_2526, signal_1571}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_600 ( .s (signal_451), .b ({plaintext_s1[19], plaintext_s0[19]}), .a ({ciphertext_s1[11], ciphertext_s0[11]}), .c ({signal_2529, signal_1570}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_601 ( .s (signal_451), .b ({plaintext_s1[20], plaintext_s0[20]}), .a ({ciphertext_s1[12], ciphertext_s0[12]}), .c ({signal_2532, signal_1569}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_602 ( .s (signal_451), .b ({plaintext_s1[21], plaintext_s0[21]}), .a ({ciphertext_s1[13], ciphertext_s0[13]}), .c ({signal_2535, signal_1568}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_603 ( .s (signal_451), .b ({plaintext_s1[22], plaintext_s0[22]}), .a ({ciphertext_s1[14], ciphertext_s0[14]}), .c ({signal_2538, signal_1567}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_604 ( .s (signal_451), .b ({plaintext_s1[23], plaintext_s0[23]}), .a ({ciphertext_s1[15], ciphertext_s0[15]}), .c ({signal_2541, signal_1566}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_605 ( .s (signal_452), .b ({plaintext_s1[8], plaintext_s0[8]}), .a ({ciphertext_s1[0], ciphertext_s0[0]}), .c ({signal_2544, signal_1565}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_606 ( .s (signal_452), .b ({plaintext_s1[9], plaintext_s0[9]}), .a ({ciphertext_s1[1], ciphertext_s0[1]}), .c ({signal_2547, signal_1564}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_607 ( .s (signal_452), .b ({plaintext_s1[10], plaintext_s0[10]}), .a ({ciphertext_s1[2], ciphertext_s0[2]}), .c ({signal_2550, signal_1563}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_608 ( .s (signal_452), .b ({plaintext_s1[11], plaintext_s0[11]}), .a ({ciphertext_s1[3], ciphertext_s0[3]}), .c ({signal_2553, signal_1562}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_609 ( .s (signal_452), .b ({plaintext_s1[12], plaintext_s0[12]}), .a ({ciphertext_s1[4], ciphertext_s0[4]}), .c ({signal_2556, signal_1561}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_610 ( .s (signal_452), .b ({plaintext_s1[13], plaintext_s0[13]}), .a ({ciphertext_s1[5], ciphertext_s0[5]}), .c ({signal_2559, signal_1560}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_611 ( .s (signal_452), .b ({plaintext_s1[14], plaintext_s0[14]}), .a ({ciphertext_s1[6], ciphertext_s0[6]}), .c ({signal_2562, signal_1559}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_612 ( .s (signal_452), .b ({plaintext_s1[15], plaintext_s0[15]}), .a ({ciphertext_s1[7], ciphertext_s0[7]}), .c ({signal_2565, signal_1558}) ) ;
    INV_X1 cell_629 ( .A (signal_399), .ZN (signal_721) ) ;
    INV_X1 cell_630 ( .A (signal_721), .ZN (signal_722) ) ;
    INV_X1 cell_631 ( .A (signal_721), .ZN (signal_723) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_632 ( .s (signal_723), .b ({signal_2949, signal_1485}), .a ({ciphertext_s1[24], ciphertext_s0[24]}), .c ({signal_2984, signal_1453}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_633 ( .s (signal_722), .b ({signal_2973, signal_1484}), .a ({ciphertext_s1[25], ciphertext_s0[25]}), .c ({signal_2985, signal_1452}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_634 ( .s (signal_399), .b ({signal_2947, signal_1483}), .a ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({signal_2958, signal_1451}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_635 ( .s (signal_399), .b ({signal_2972, signal_1482}), .a ({ciphertext_s1[27], ciphertext_s0[27]}), .c ({signal_2986, signal_1450}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_636 ( .s (signal_399), .b ({signal_2971, signal_1481}), .a ({ciphertext_s1[28], ciphertext_s0[28]}), .c ({signal_2987, signal_1449}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_637 ( .s (signal_399), .b ({signal_2944, signal_1480}), .a ({ciphertext_s1[29], ciphertext_s0[29]}), .c ({signal_2959, signal_1448}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_638 ( .s (signal_399), .b ({signal_2943, signal_1479}), .a ({ciphertext_s1[30], ciphertext_s0[30]}), .c ({signal_2960, signal_1447}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_639 ( .s (signal_399), .b ({signal_2942, signal_1478}), .a ({ciphertext_s1[31], ciphertext_s0[31]}), .c ({signal_2961, signal_1446}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_640 ( .s (signal_722), .b ({signal_2941, signal_1477}), .a ({ciphertext_s1[56], ciphertext_s0[56]}), .c ({signal_2988, signal_1445}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_641 ( .s (signal_722), .b ({signal_2970, signal_1476}), .a ({ciphertext_s1[57], ciphertext_s0[57]}), .c ({signal_2989, signal_1444}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_642 ( .s (signal_722), .b ({signal_2939, signal_1475}), .a ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({signal_2990, signal_1443}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_643 ( .s (signal_722), .b ({signal_2969, signal_1474}), .a ({ciphertext_s1[59], ciphertext_s0[59]}), .c ({signal_2991, signal_1442}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_644 ( .s (signal_722), .b ({signal_2968, signal_1473}), .a ({ciphertext_s1[60], ciphertext_s0[60]}), .c ({signal_2992, signal_1441}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_645 ( .s (signal_722), .b ({signal_2936, signal_1472}), .a ({ciphertext_s1[61], ciphertext_s0[61]}), .c ({signal_2993, signal_1440}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_646 ( .s (signal_722), .b ({signal_2935, signal_1471}), .a ({ciphertext_s1[62], ciphertext_s0[62]}), .c ({signal_2994, signal_1439}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_647 ( .s (signal_722), .b ({signal_2934, signal_1470}), .a ({ciphertext_s1[63], ciphertext_s0[63]}), .c ({signal_2995, signal_1438}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_648 ( .s (signal_722), .b ({signal_2933, signal_1469}), .a ({ciphertext_s1[88], ciphertext_s0[88]}), .c ({signal_2996, signal_1437}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_649 ( .s (signal_722), .b ({signal_2967, signal_1468}), .a ({ciphertext_s1[89], ciphertext_s0[89]}), .c ({signal_2997, signal_1436}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_650 ( .s (signal_722), .b ({signal_2931, signal_1467}), .a ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({signal_2998, signal_1435}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_651 ( .s (signal_722), .b ({signal_2966, signal_1466}), .a ({ciphertext_s1[91], ciphertext_s0[91]}), .c ({signal_2999, signal_1434}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_652 ( .s (signal_723), .b ({signal_2965, signal_1465}), .a ({ciphertext_s1[92], ciphertext_s0[92]}), .c ({signal_3000, signal_1433}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_653 ( .s (signal_723), .b ({signal_2928, signal_1464}), .a ({ciphertext_s1[93], ciphertext_s0[93]}), .c ({signal_3001, signal_1432}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_654 ( .s (signal_723), .b ({signal_2927, signal_1463}), .a ({ciphertext_s1[94], ciphertext_s0[94]}), .c ({signal_3002, signal_1431}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_655 ( .s (signal_723), .b ({signal_2926, signal_1462}), .a ({ciphertext_s1[95], ciphertext_s0[95]}), .c ({signal_3003, signal_1430}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_656 ( .s (signal_723), .b ({signal_2925, signal_1461}), .a ({ciphertext_s1[120], ciphertext_s0[120]}), .c ({signal_3004, signal_1429}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_657 ( .s (signal_723), .b ({signal_2964, signal_1460}), .a ({ciphertext_s1[121], ciphertext_s0[121]}), .c ({signal_3005, signal_1428}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_658 ( .s (signal_723), .b ({signal_2923, signal_1459}), .a ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({signal_3006, signal_1427}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_659 ( .s (signal_723), .b ({signal_2963, signal_1458}), .a ({ciphertext_s1[123], ciphertext_s0[123]}), .c ({signal_3007, signal_1426}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_660 ( .s (signal_723), .b ({signal_2962, signal_1457}), .a ({ciphertext_s1[124], ciphertext_s0[124]}), .c ({signal_3008, signal_1425}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_661 ( .s (signal_723), .b ({signal_2920, signal_1456}), .a ({ciphertext_s1[125], ciphertext_s0[125]}), .c ({signal_3009, signal_1424}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_662 ( .s (signal_723), .b ({signal_2919, signal_1455}), .a ({ciphertext_s1[126], ciphertext_s0[126]}), .c ({signal_3010, signal_1423}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_663 ( .s (signal_723), .b ({signal_2918, signal_1454}), .a ({ciphertext_s1[127], ciphertext_s0[127]}), .c ({signal_3011, signal_1422}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_664 ( .a ({signal_2130, signal_765}), .b ({signal_2128, signal_1486}), .c ({signal_2131, signal_1686}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_665 ( .a ({signal_2132, signal_764}), .b ({signal_2125, signal_1487}), .c ({signal_2133, signal_1687}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_666 ( .a ({signal_2134, signal_763}), .b ({signal_2122, signal_1488}), .c ({signal_2135, signal_1688}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_667 ( .a ({signal_2136, signal_762}), .b ({signal_2119, signal_1489}), .c ({signal_2137, signal_1689}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_668 ( .a ({signal_2138, signal_761}), .b ({signal_2116, signal_1490}), .c ({signal_2139, signal_1690}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_669 ( .a ({signal_2140, signal_760}), .b ({signal_2113, signal_1491}), .c ({signal_2141, signal_1691}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_670 ( .a ({signal_2142, signal_759}), .b ({signal_2110, signal_1492}), .c ({signal_2143, signal_1692}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_671 ( .a ({signal_2144, signal_758}), .b ({signal_2107, signal_1493}), .c ({signal_2145, signal_1693}) ) ;
    INV_X1 cell_688 ( .A (signal_732), .ZN (signal_733) ) ;
    INV_X1 cell_689 ( .A (signal_732), .ZN (signal_734) ) ;
    INV_X1 cell_690 ( .A (signal_732), .ZN (signal_735) ) ;
    INV_X1 cell_691 ( .A (signal_732), .ZN (signal_736) ) ;
    INV_X1 cell_692 ( .A (signal_732), .ZN (signal_737) ) ;
    INV_X1 cell_693 ( .A (signal_732), .ZN (signal_738) ) ;
    INV_X1 cell_694 ( .A (signal_732), .ZN (signal_739) ) ;
    INV_X1 cell_695 ( .A (signal_732), .ZN (signal_740) ) ;
    INV_X1 cell_696 ( .A (signal_393), .ZN (signal_732) ) ;
    INV_X1 cell_697 ( .A (signal_741), .ZN (signal_748) ) ;
    INV_X1 cell_698 ( .A (signal_750), .ZN (signal_756) ) ;
    INV_X1 cell_699 ( .A (signal_741), .ZN (signal_742) ) ;
    INV_X1 cell_700 ( .A (signal_750), .ZN (signal_751) ) ;
    INV_X1 cell_701 ( .A (signal_741), .ZN (signal_743) ) ;
    INV_X1 cell_702 ( .A (signal_750), .ZN (signal_752) ) ;
    INV_X1 cell_703 ( .A (signal_741), .ZN (signal_744) ) ;
    INV_X1 cell_704 ( .A (signal_750), .ZN (signal_753) ) ;
    INV_X1 cell_705 ( .A (signal_741), .ZN (signal_747) ) ;
    INV_X1 cell_706 ( .A (signal_750), .ZN (signal_755) ) ;
    INV_X1 cell_707 ( .A (signal_741), .ZN (signal_746) ) ;
    INV_X1 cell_708 ( .A (signal_750), .ZN (signal_754) ) ;
    INV_X1 cell_709 ( .A (signal_741), .ZN (signal_749) ) ;
    INV_X1 cell_710 ( .A (signal_750), .ZN (signal_757) ) ;
    INV_X1 cell_711 ( .A (signal_741), .ZN (signal_745) ) ;
    INV_X1 cell_712 ( .A (signal_394), .ZN (signal_741) ) ;
    INV_X1 cell_713 ( .A (signal_404), .ZN (signal_750) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_714 ( .s (signal_751), .b ({signal_2107, signal_1493}), .a ({signal_3391, signal_767}), .c ({signal_3499, signal_766}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_715 ( .s (signal_742), .b ({signal_3371, signal_1933}), .a ({signal_2615, signal_1877}), .c ({signal_3391, signal_767}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_718 ( .s (signal_751), .b ({signal_2110, signal_1492}), .a ({signal_3392, signal_770}), .c ({signal_3500, signal_769}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_719 ( .s (signal_742), .b ({signal_3373, signal_1932}), .a ({signal_2618, signal_1876}), .c ({signal_3392, signal_770}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_722 ( .s (signal_751), .b ({signal_2113, signal_1491}), .a ({signal_3393, signal_773}), .c ({signal_3501, signal_772}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_723 ( .s (signal_742), .b ({signal_3375, signal_1931}), .a ({signal_2621, signal_1875}), .c ({signal_3393, signal_773}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_726 ( .s (signal_751), .b ({signal_2116, signal_1490}), .a ({signal_3394, signal_776}), .c ({signal_3502, signal_775}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_727 ( .s (signal_742), .b ({signal_3377, signal_1930}), .a ({signal_2624, signal_1874}), .c ({signal_3394, signal_776}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_730 ( .s (signal_751), .b ({signal_2119, signal_1489}), .a ({signal_3395, signal_779}), .c ({signal_3503, signal_778}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_731 ( .s (signal_742), .b ({signal_3379, signal_1929}), .a ({signal_2627, signal_1873}), .c ({signal_3395, signal_779}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_734 ( .s (signal_751), .b ({signal_2122, signal_1488}), .a ({signal_3396, signal_782}), .c ({signal_3504, signal_781}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_735 ( .s (signal_742), .b ({signal_3381, signal_1928}), .a ({signal_2630, signal_1872}), .c ({signal_3396, signal_782}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_738 ( .s (signal_751), .b ({signal_2125, signal_1487}), .a ({signal_3397, signal_785}), .c ({signal_3505, signal_784}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_739 ( .s (signal_742), .b ({signal_3383, signal_1927}), .a ({signal_2633, signal_1871}), .c ({signal_3397, signal_785}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_742 ( .s (signal_751), .b ({signal_2128, signal_1486}), .a ({signal_3398, signal_788}), .c ({signal_3506, signal_787}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_743 ( .s (signal_742), .b ({signal_3385, signal_1926}), .a ({signal_2636, signal_1870}), .c ({signal_3398, signal_788}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_746 ( .s (signal_751), .b ({signal_2144, signal_758}), .a ({signal_3012, signal_791}), .c ({signal_3399, signal_790}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_747 ( .s (signal_742), .b ({signal_2568, signal_1925}), .a ({signal_2639, signal_1861}), .c ({signal_3012, signal_791}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_750 ( .s (signal_751), .b ({signal_2142, signal_759}), .a ({signal_3013, signal_794}), .c ({signal_3400, signal_793}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_751 ( .s (signal_742), .b ({signal_2571, signal_1924}), .a ({signal_2642, signal_1860}), .c ({signal_3013, signal_794}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_754 ( .s (signal_751), .b ({signal_2140, signal_760}), .a ({signal_3014, signal_797}), .c ({signal_3401, signal_796}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_755 ( .s (signal_742), .b ({signal_2574, signal_1923}), .a ({signal_2645, signal_1859}), .c ({signal_3014, signal_797}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_758 ( .s (signal_751), .b ({signal_2138, signal_761}), .a ({signal_3015, signal_800}), .c ({signal_3402, signal_799}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_759 ( .s (signal_742), .b ({signal_2577, signal_1922}), .a ({signal_2648, signal_1858}), .c ({signal_3015, signal_800}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_762 ( .s (signal_751), .b ({signal_2136, signal_762}), .a ({signal_3016, signal_803}), .c ({signal_3403, signal_802}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_763 ( .s (signal_742), .b ({signal_2580, signal_1921}), .a ({signal_2651, signal_1857}), .c ({signal_3016, signal_803}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_766 ( .s (signal_751), .b ({signal_2134, signal_763}), .a ({signal_3017, signal_806}), .c ({signal_3404, signal_805}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_767 ( .s (signal_742), .b ({signal_2583, signal_1920}), .a ({signal_2654, signal_1856}), .c ({signal_3017, signal_806}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_770 ( .s (signal_751), .b ({signal_2132, signal_764}), .a ({signal_3018, signal_809}), .c ({signal_3405, signal_808}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_771 ( .s (signal_742), .b ({signal_2586, signal_1919}), .a ({signal_2657, signal_1855}), .c ({signal_3018, signal_809}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_774 ( .s (signal_751), .b ({signal_2130, signal_765}), .a ({signal_3019, signal_812}), .c ({signal_3406, signal_811}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_775 ( .s (signal_742), .b ({signal_2589, signal_1918}), .a ({signal_2660, signal_1854}), .c ({signal_3019, signal_812}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_778 ( .s (signal_752), .b ({signal_2567, signal_1909}), .a ({signal_3020, signal_815}), .c ({signal_3407, signal_814}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_779 ( .s (signal_743), .b ({signal_2592, signal_1917}), .a ({signal_2663, signal_1845}), .c ({signal_3020, signal_815}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_782 ( .s (signal_752), .b ({signal_2570, signal_1908}), .a ({signal_3021, signal_818}), .c ({signal_3408, signal_817}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_783 ( .s (signal_743), .b ({signal_2595, signal_1916}), .a ({signal_2666, signal_1844}), .c ({signal_3021, signal_818}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_786 ( .s (signal_752), .b ({signal_2573, signal_1907}), .a ({signal_3022, signal_821}), .c ({signal_3409, signal_820}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_787 ( .s (signal_743), .b ({signal_2598, signal_1915}), .a ({signal_2669, signal_1843}), .c ({signal_3022, signal_821}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_790 ( .s (signal_752), .b ({signal_2576, signal_1906}), .a ({signal_3023, signal_824}), .c ({signal_3410, signal_823}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_791 ( .s (signal_743), .b ({signal_2601, signal_1914}), .a ({signal_2672, signal_1842}), .c ({signal_3023, signal_824}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_794 ( .s (signal_752), .b ({signal_2579, signal_1905}), .a ({signal_3024, signal_827}), .c ({signal_3411, signal_826}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_795 ( .s (signal_743), .b ({signal_2604, signal_1913}), .a ({signal_2675, signal_1841}), .c ({signal_3024, signal_827}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_798 ( .s (signal_752), .b ({signal_2582, signal_1904}), .a ({signal_3025, signal_830}), .c ({signal_3412, signal_829}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_799 ( .s (signal_743), .b ({signal_2607, signal_1912}), .a ({signal_2678, signal_1840}), .c ({signal_3025, signal_830}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_802 ( .s (signal_752), .b ({signal_2585, signal_1903}), .a ({signal_3026, signal_833}), .c ({signal_3413, signal_832}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_803 ( .s (signal_743), .b ({signal_2610, signal_1911}), .a ({signal_2681, signal_1839}), .c ({signal_3026, signal_833}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_806 ( .s (signal_752), .b ({signal_2588, signal_1902}), .a ({signal_3027, signal_836}), .c ({signal_3414, signal_835}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_807 ( .s (signal_743), .b ({signal_2613, signal_1910}), .a ({signal_2684, signal_1838}), .c ({signal_3027, signal_836}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_810 ( .s (signal_752), .b ({signal_2591, signal_1893}), .a ({signal_3028, signal_839}), .c ({signal_3415, signal_838}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_811 ( .s (signal_743), .b ({signal_2616, signal_1901}), .a ({signal_2687, signal_1509}), .c ({signal_3028, signal_839}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_814 ( .s (signal_752), .b ({signal_2594, signal_1892}), .a ({signal_3029, signal_842}), .c ({signal_3416, signal_841}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_815 ( .s (signal_743), .b ({signal_2619, signal_1900}), .a ({signal_2690, signal_1508}), .c ({signal_3029, signal_842}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_818 ( .s (signal_752), .b ({signal_2597, signal_1891}), .a ({signal_3030, signal_845}), .c ({signal_3417, signal_844}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_819 ( .s (signal_743), .b ({signal_2622, signal_1899}), .a ({signal_2693, signal_1507}), .c ({signal_3030, signal_845}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_822 ( .s (signal_752), .b ({signal_2600, signal_1890}), .a ({signal_3031, signal_848}), .c ({signal_3418, signal_847}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_823 ( .s (signal_743), .b ({signal_2625, signal_1898}), .a ({signal_2696, signal_1506}), .c ({signal_3031, signal_848}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_826 ( .s (signal_752), .b ({signal_2603, signal_1889}), .a ({signal_3032, signal_851}), .c ({signal_3419, signal_850}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_827 ( .s (signal_743), .b ({signal_2628, signal_1897}), .a ({signal_2699, signal_1505}), .c ({signal_3032, signal_851}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_830 ( .s (signal_752), .b ({signal_2606, signal_1888}), .a ({signal_3033, signal_854}), .c ({signal_3420, signal_853}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_831 ( .s (signal_743), .b ({signal_2631, signal_1896}), .a ({signal_2702, signal_1504}), .c ({signal_3033, signal_854}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_834 ( .s (signal_752), .b ({signal_2609, signal_1887}), .a ({signal_3034, signal_857}), .c ({signal_3421, signal_856}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_835 ( .s (signal_743), .b ({signal_2634, signal_1895}), .a ({signal_2705, signal_1503}), .c ({signal_3034, signal_857}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_838 ( .s (signal_752), .b ({signal_2612, signal_1886}), .a ({signal_3035, signal_860}), .c ({signal_3422, signal_859}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_839 ( .s (signal_743), .b ({signal_2637, signal_1894}), .a ({signal_2708, signal_1502}), .c ({signal_3035, signal_860}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_842 ( .s (signal_753), .b ({signal_2615, signal_1877}), .a ({signal_3036, signal_863}), .c ({signal_3423, signal_862}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_843 ( .s (signal_744), .b ({signal_2640, signal_1885}), .a ({signal_2711, signal_1821}), .c ({signal_3036, signal_863}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_846 ( .s (signal_753), .b ({signal_2618, signal_1876}), .a ({signal_3037, signal_866}), .c ({signal_3424, signal_865}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_847 ( .s (signal_744), .b ({signal_2643, signal_1884}), .a ({signal_2714, signal_1820}), .c ({signal_3037, signal_866}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_850 ( .s (signal_753), .b ({signal_2621, signal_1875}), .a ({signal_3038, signal_869}), .c ({signal_3425, signal_868}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_851 ( .s (signal_744), .b ({signal_2646, signal_1883}), .a ({signal_2717, signal_1819}), .c ({signal_3038, signal_869}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_854 ( .s (signal_753), .b ({signal_2624, signal_1874}), .a ({signal_3039, signal_872}), .c ({signal_3426, signal_871}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_855 ( .s (signal_744), .b ({signal_2649, signal_1882}), .a ({signal_2720, signal_1818}), .c ({signal_3039, signal_872}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_858 ( .s (signal_753), .b ({signal_2627, signal_1873}), .a ({signal_3040, signal_875}), .c ({signal_3427, signal_874}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_859 ( .s (signal_744), .b ({signal_2652, signal_1881}), .a ({signal_2723, signal_1817}), .c ({signal_3040, signal_875}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_862 ( .s (signal_753), .b ({signal_2630, signal_1872}), .a ({signal_3041, signal_878}), .c ({signal_3428, signal_877}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_863 ( .s (signal_744), .b ({signal_2655, signal_1880}), .a ({signal_2726, signal_1816}), .c ({signal_3041, signal_878}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_866 ( .s (signal_753), .b ({signal_2633, signal_1871}), .a ({signal_3042, signal_881}), .c ({signal_3429, signal_880}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_867 ( .s (signal_744), .b ({signal_2658, signal_1879}), .a ({signal_2729, signal_1815}), .c ({signal_3042, signal_881}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_870 ( .s (signal_753), .b ({signal_2636, signal_1870}), .a ({signal_3043, signal_884}), .c ({signal_3430, signal_883}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_871 ( .s (signal_744), .b ({signal_2661, signal_1878}), .a ({signal_2732, signal_1814}), .c ({signal_3043, signal_884}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_874 ( .s (signal_753), .b ({signal_2639, signal_1861}), .a ({signal_3044, signal_887}), .c ({signal_3431, signal_886}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_875 ( .s (signal_744), .b ({signal_2664, signal_1869}), .a ({signal_2735, signal_1805}), .c ({signal_3044, signal_887}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_878 ( .s (signal_753), .b ({signal_2642, signal_1860}), .a ({signal_3045, signal_890}), .c ({signal_3432, signal_889}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_879 ( .s (signal_744), .b ({signal_2667, signal_1868}), .a ({signal_2738, signal_1804}), .c ({signal_3045, signal_890}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_882 ( .s (signal_753), .b ({signal_2645, signal_1859}), .a ({signal_3046, signal_893}), .c ({signal_3433, signal_892}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_883 ( .s (signal_744), .b ({signal_2670, signal_1867}), .a ({signal_2741, signal_1803}), .c ({signal_3046, signal_893}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_886 ( .s (signal_753), .b ({signal_2648, signal_1858}), .a ({signal_3047, signal_896}), .c ({signal_3434, signal_895}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_887 ( .s (signal_744), .b ({signal_2673, signal_1866}), .a ({signal_2744, signal_1802}), .c ({signal_3047, signal_896}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_890 ( .s (signal_753), .b ({signal_2651, signal_1857}), .a ({signal_3048, signal_899}), .c ({signal_3435, signal_898}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_891 ( .s (signal_744), .b ({signal_2676, signal_1865}), .a ({signal_2747, signal_1801}), .c ({signal_3048, signal_899}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_894 ( .s (signal_753), .b ({signal_2654, signal_1856}), .a ({signal_3049, signal_902}), .c ({signal_3436, signal_901}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_895 ( .s (signal_744), .b ({signal_2679, signal_1864}), .a ({signal_2750, signal_1800}), .c ({signal_3049, signal_902}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_898 ( .s (signal_753), .b ({signal_2657, signal_1855}), .a ({signal_3050, signal_905}), .c ({signal_3437, signal_904}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_899 ( .s (signal_744), .b ({signal_2682, signal_1863}), .a ({signal_2753, signal_1799}), .c ({signal_3050, signal_905}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_902 ( .s (signal_753), .b ({signal_2660, signal_1854}), .a ({signal_3051, signal_908}), .c ({signal_3438, signal_907}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_903 ( .s (signal_744), .b ({signal_2685, signal_1862}), .a ({signal_2756, signal_1798}), .c ({signal_3051, signal_908}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_906 ( .s (signal_404), .b ({signal_2663, signal_1845}), .a ({signal_3052, signal_911}), .c ({signal_3217, signal_910}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_907 ( .s (signal_745), .b ({signal_2688, signal_1853}), .a ({signal_2759, signal_1789}), .c ({signal_3052, signal_911}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_910 ( .s (signal_404), .b ({signal_2666, signal_1844}), .a ({signal_3053, signal_914}), .c ({signal_3218, signal_913}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_911 ( .s (signal_745), .b ({signal_2691, signal_1852}), .a ({signal_2762, signal_1788}), .c ({signal_3053, signal_914}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_914 ( .s (signal_404), .b ({signal_2669, signal_1843}), .a ({signal_3054, signal_917}), .c ({signal_3219, signal_916}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_915 ( .s (signal_745), .b ({signal_2694, signal_1851}), .a ({signal_2765, signal_1787}), .c ({signal_3054, signal_917}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_918 ( .s (signal_404), .b ({signal_2672, signal_1842}), .a ({signal_3055, signal_920}), .c ({signal_3220, signal_919}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_919 ( .s (signal_745), .b ({signal_2697, signal_1850}), .a ({signal_2768, signal_1786}), .c ({signal_3055, signal_920}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_922 ( .s (signal_404), .b ({signal_2675, signal_1841}), .a ({signal_3056, signal_923}), .c ({signal_3221, signal_922}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_923 ( .s (signal_745), .b ({signal_2700, signal_1849}), .a ({signal_2771, signal_1785}), .c ({signal_3056, signal_923}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_926 ( .s (signal_404), .b ({signal_2678, signal_1840}), .a ({signal_3057, signal_926}), .c ({signal_3222, signal_925}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_927 ( .s (signal_745), .b ({signal_2703, signal_1848}), .a ({signal_2774, signal_1784}), .c ({signal_3057, signal_926}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_930 ( .s (signal_404), .b ({signal_2681, signal_1839}), .a ({signal_3058, signal_929}), .c ({signal_3223, signal_928}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_931 ( .s (signal_745), .b ({signal_2706, signal_1847}), .a ({signal_2777, signal_1783}), .c ({signal_3058, signal_929}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_934 ( .s (signal_404), .b ({signal_2684, signal_1838}), .a ({signal_3059, signal_932}), .c ({signal_3224, signal_931}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_935 ( .s (signal_745), .b ({signal_2709, signal_1846}), .a ({signal_2780, signal_1782}), .c ({signal_3059, signal_932}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_938 ( .s (signal_404), .b ({signal_2687, signal_1509}), .a ({signal_3060, signal_935}), .c ({signal_3225, signal_934}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_939 ( .s (signal_745), .b ({signal_2712, signal_1837}), .a ({signal_2783, signal_1773}), .c ({signal_3060, signal_935}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_942 ( .s (signal_404), .b ({signal_2690, signal_1508}), .a ({signal_3061, signal_938}), .c ({signal_3226, signal_937}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_943 ( .s (signal_745), .b ({signal_2715, signal_1836}), .a ({signal_2786, signal_1772}), .c ({signal_3061, signal_938}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_946 ( .s (signal_404), .b ({signal_2693, signal_1507}), .a ({signal_3062, signal_941}), .c ({signal_3227, signal_940}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_947 ( .s (signal_745), .b ({signal_2718, signal_1835}), .a ({signal_2789, signal_1771}), .c ({signal_3062, signal_941}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_950 ( .s (signal_404), .b ({signal_2696, signal_1506}), .a ({signal_3063, signal_944}), .c ({signal_3228, signal_943}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_951 ( .s (signal_745), .b ({signal_2721, signal_1834}), .a ({signal_2792, signal_1770}), .c ({signal_3063, signal_944}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_954 ( .s (signal_404), .b ({signal_2699, signal_1505}), .a ({signal_3064, signal_947}), .c ({signal_3229, signal_946}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_955 ( .s (signal_745), .b ({signal_2724, signal_1833}), .a ({signal_2795, signal_1769}), .c ({signal_3064, signal_947}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_958 ( .s (signal_404), .b ({signal_2702, signal_1504}), .a ({signal_3065, signal_950}), .c ({signal_3230, signal_949}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_959 ( .s (signal_745), .b ({signal_2727, signal_1832}), .a ({signal_2798, signal_1768}), .c ({signal_3065, signal_950}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_962 ( .s (signal_404), .b ({signal_2705, signal_1503}), .a ({signal_3066, signal_953}), .c ({signal_3231, signal_952}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_963 ( .s (signal_745), .b ({signal_2730, signal_1831}), .a ({signal_2801, signal_1767}), .c ({signal_3066, signal_953}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_966 ( .s (signal_404), .b ({signal_2708, signal_1502}), .a ({signal_3067, signal_956}), .c ({signal_3232, signal_955}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_967 ( .s (signal_745), .b ({signal_2733, signal_1830}), .a ({signal_2804, signal_1766}), .c ({signal_3067, signal_956}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_970 ( .s (signal_754), .b ({signal_2711, signal_1821}), .a ({signal_3068, signal_959}), .c ({signal_3439, signal_958}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_971 ( .s (signal_746), .b ({signal_2736, signal_1829}), .a ({signal_2807, signal_1749}), .c ({signal_3068, signal_959}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_974 ( .s (signal_754), .b ({signal_2714, signal_1820}), .a ({signal_3069, signal_962}), .c ({signal_3440, signal_961}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_975 ( .s (signal_746), .b ({signal_2739, signal_1828}), .a ({signal_2810, signal_1748}), .c ({signal_3069, signal_962}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_978 ( .s (signal_754), .b ({signal_2717, signal_1819}), .a ({signal_3070, signal_965}), .c ({signal_3441, signal_964}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_979 ( .s (signal_746), .b ({signal_2742, signal_1827}), .a ({signal_2813, signal_1747}), .c ({signal_3070, signal_965}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_982 ( .s (signal_754), .b ({signal_2720, signal_1818}), .a ({signal_3071, signal_968}), .c ({signal_3442, signal_967}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_983 ( .s (signal_746), .b ({signal_2745, signal_1826}), .a ({signal_2816, signal_1746}), .c ({signal_3071, signal_968}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_986 ( .s (signal_754), .b ({signal_2723, signal_1817}), .a ({signal_3072, signal_971}), .c ({signal_3443, signal_970}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_987 ( .s (signal_746), .b ({signal_2748, signal_1825}), .a ({signal_2819, signal_1745}), .c ({signal_3072, signal_971}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_990 ( .s (signal_754), .b ({signal_2726, signal_1816}), .a ({signal_3073, signal_974}), .c ({signal_3444, signal_973}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_991 ( .s (signal_746), .b ({signal_2751, signal_1824}), .a ({signal_2822, signal_1744}), .c ({signal_3073, signal_974}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_994 ( .s (signal_754), .b ({signal_2729, signal_1815}), .a ({signal_3074, signal_977}), .c ({signal_3445, signal_976}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_995 ( .s (signal_746), .b ({signal_2754, signal_1823}), .a ({signal_2825, signal_1743}), .c ({signal_3074, signal_977}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_998 ( .s (signal_754), .b ({signal_2732, signal_1814}), .a ({signal_3075, signal_980}), .c ({signal_3446, signal_979}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_999 ( .s (signal_746), .b ({signal_2757, signal_1822}), .a ({signal_2828, signal_1742}), .c ({signal_3075, signal_980}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1002 ( .s (signal_754), .b ({signal_2735, signal_1805}), .a ({signal_3076, signal_983}), .c ({signal_3447, signal_982}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1003 ( .s (signal_746), .b ({signal_2760, signal_1813}), .a ({signal_2831, signal_1733}), .c ({signal_3076, signal_983}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1006 ( .s (signal_754), .b ({signal_2738, signal_1804}), .a ({signal_3077, signal_986}), .c ({signal_3448, signal_985}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1007 ( .s (signal_746), .b ({signal_2763, signal_1812}), .a ({signal_2834, signal_1732}), .c ({signal_3077, signal_986}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1010 ( .s (signal_754), .b ({signal_2741, signal_1803}), .a ({signal_3078, signal_989}), .c ({signal_3449, signal_988}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1011 ( .s (signal_746), .b ({signal_2766, signal_1811}), .a ({signal_2837, signal_1731}), .c ({signal_3078, signal_989}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1014 ( .s (signal_754), .b ({signal_2744, signal_1802}), .a ({signal_3079, signal_992}), .c ({signal_3450, signal_991}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1015 ( .s (signal_746), .b ({signal_2769, signal_1810}), .a ({signal_2840, signal_1730}), .c ({signal_3079, signal_992}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1018 ( .s (signal_754), .b ({signal_2747, signal_1801}), .a ({signal_3080, signal_995}), .c ({signal_3451, signal_994}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1019 ( .s (signal_746), .b ({signal_2772, signal_1809}), .a ({signal_2843, signal_1729}), .c ({signal_3080, signal_995}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1022 ( .s (signal_754), .b ({signal_2750, signal_1800}), .a ({signal_3081, signal_998}), .c ({signal_3452, signal_997}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1023 ( .s (signal_746), .b ({signal_2775, signal_1808}), .a ({signal_2846, signal_1728}), .c ({signal_3081, signal_998}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1026 ( .s (signal_754), .b ({signal_2753, signal_1799}), .a ({signal_3082, signal_1001}), .c ({signal_3453, signal_1000}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1027 ( .s (signal_746), .b ({signal_2778, signal_1807}), .a ({signal_2849, signal_1727}), .c ({signal_3082, signal_1001}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1030 ( .s (signal_754), .b ({signal_2756, signal_1798}), .a ({signal_3083, signal_1004}), .c ({signal_3454, signal_1003}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1031 ( .s (signal_746), .b ({signal_2781, signal_1806}), .a ({signal_2852, signal_1726}), .c ({signal_3083, signal_1004}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1034 ( .s (signal_755), .b ({signal_2759, signal_1789}), .a ({signal_3084, signal_1007}), .c ({signal_3455, signal_1006}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1035 ( .s (signal_747), .b ({signal_2784, signal_1797}), .a ({signal_2855, signal_1717}), .c ({signal_3084, signal_1007}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1038 ( .s (signal_755), .b ({signal_2762, signal_1788}), .a ({signal_3085, signal_1010}), .c ({signal_3456, signal_1009}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1039 ( .s (signal_747), .b ({signal_2787, signal_1796}), .a ({signal_2858, signal_1716}), .c ({signal_3085, signal_1010}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1042 ( .s (signal_755), .b ({signal_2765, signal_1787}), .a ({signal_3086, signal_1013}), .c ({signal_3457, signal_1012}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1043 ( .s (signal_747), .b ({signal_2790, signal_1795}), .a ({signal_2861, signal_1715}), .c ({signal_3086, signal_1013}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1046 ( .s (signal_755), .b ({signal_2768, signal_1786}), .a ({signal_3087, signal_1016}), .c ({signal_3458, signal_1015}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1047 ( .s (signal_747), .b ({signal_2793, signal_1794}), .a ({signal_2864, signal_1714}), .c ({signal_3087, signal_1016}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1050 ( .s (signal_755), .b ({signal_2771, signal_1785}), .a ({signal_3088, signal_1019}), .c ({signal_3459, signal_1018}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1051 ( .s (signal_747), .b ({signal_2796, signal_1793}), .a ({signal_2867, signal_1713}), .c ({signal_3088, signal_1019}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1054 ( .s (signal_755), .b ({signal_2774, signal_1784}), .a ({signal_3089, signal_1022}), .c ({signal_3460, signal_1021}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1055 ( .s (signal_747), .b ({signal_2799, signal_1792}), .a ({signal_2870, signal_1712}), .c ({signal_3089, signal_1022}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1058 ( .s (signal_755), .b ({signal_2777, signal_1783}), .a ({signal_3090, signal_1025}), .c ({signal_3461, signal_1024}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1059 ( .s (signal_747), .b ({signal_2802, signal_1791}), .a ({signal_2873, signal_1711}), .c ({signal_3090, signal_1025}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1062 ( .s (signal_755), .b ({signal_2780, signal_1782}), .a ({signal_3091, signal_1028}), .c ({signal_3462, signal_1027}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1063 ( .s (signal_747), .b ({signal_2805, signal_1790}), .a ({signal_2876, signal_1710}), .c ({signal_3091, signal_1028}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1066 ( .s (signal_755), .b ({signal_2783, signal_1773}), .a ({signal_3092, signal_1031}), .c ({signal_3463, signal_1030}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1067 ( .s (signal_747), .b ({signal_2808, signal_1781}), .a ({signal_2879, signal_1701}), .c ({signal_3092, signal_1031}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1070 ( .s (signal_755), .b ({signal_2786, signal_1772}), .a ({signal_3093, signal_1034}), .c ({signal_3464, signal_1033}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1071 ( .s (signal_747), .b ({signal_2811, signal_1780}), .a ({signal_2882, signal_1700}), .c ({signal_3093, signal_1034}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1074 ( .s (signal_755), .b ({signal_2789, signal_1771}), .a ({signal_3094, signal_1037}), .c ({signal_3465, signal_1036}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1075 ( .s (signal_747), .b ({signal_2814, signal_1779}), .a ({signal_2885, signal_1699}), .c ({signal_3094, signal_1037}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1078 ( .s (signal_755), .b ({signal_2792, signal_1770}), .a ({signal_3095, signal_1040}), .c ({signal_3466, signal_1039}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1079 ( .s (signal_747), .b ({signal_2817, signal_1778}), .a ({signal_2888, signal_1698}), .c ({signal_3095, signal_1040}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1082 ( .s (signal_755), .b ({signal_2795, signal_1769}), .a ({signal_3096, signal_1043}), .c ({signal_3467, signal_1042}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1083 ( .s (signal_747), .b ({signal_2820, signal_1777}), .a ({signal_2891, signal_1697}), .c ({signal_3096, signal_1043}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1086 ( .s (signal_755), .b ({signal_2798, signal_1768}), .a ({signal_3097, signal_1046}), .c ({signal_3468, signal_1045}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1087 ( .s (signal_747), .b ({signal_2823, signal_1776}), .a ({signal_2894, signal_1696}), .c ({signal_3097, signal_1046}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1090 ( .s (signal_755), .b ({signal_2801, signal_1767}), .a ({signal_3098, signal_1049}), .c ({signal_3469, signal_1048}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1091 ( .s (signal_747), .b ({signal_2826, signal_1775}), .a ({signal_2897, signal_1695}), .c ({signal_3098, signal_1049}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1094 ( .s (signal_755), .b ({signal_2804, signal_1766}), .a ({signal_3099, signal_1052}), .c ({signal_3470, signal_1051}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1095 ( .s (signal_747), .b ({signal_2829, signal_1774}), .a ({signal_2900, signal_1694}), .c ({signal_3099, signal_1052}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1130 ( .s (signal_756), .b ({signal_2831, signal_1733}), .a ({signal_3100, signal_1079}), .c ({signal_3471, signal_1078}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1131 ( .s (signal_748), .b ({signal_2856, signal_1741}), .a ({signal_2144, signal_758}), .c ({signal_3100, signal_1079}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1134 ( .s (signal_756), .b ({signal_2834, signal_1732}), .a ({signal_3101, signal_1082}), .c ({signal_3472, signal_1081}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1135 ( .s (signal_748), .b ({signal_2859, signal_1740}), .a ({signal_2142, signal_759}), .c ({signal_3101, signal_1082}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1138 ( .s (signal_756), .b ({signal_2837, signal_1731}), .a ({signal_3102, signal_1085}), .c ({signal_3473, signal_1084}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1139 ( .s (signal_748), .b ({signal_2862, signal_1739}), .a ({signal_2140, signal_760}), .c ({signal_3102, signal_1085}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1142 ( .s (signal_756), .b ({signal_2840, signal_1730}), .a ({signal_3103, signal_1088}), .c ({signal_3474, signal_1087}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1143 ( .s (signal_748), .b ({signal_2865, signal_1738}), .a ({signal_2138, signal_761}), .c ({signal_3103, signal_1088}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1146 ( .s (signal_756), .b ({signal_2843, signal_1729}), .a ({signal_3104, signal_1091}), .c ({signal_3475, signal_1090}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1147 ( .s (signal_748), .b ({signal_2868, signal_1737}), .a ({signal_2136, signal_762}), .c ({signal_3104, signal_1091}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1150 ( .s (signal_756), .b ({signal_2846, signal_1728}), .a ({signal_3105, signal_1094}), .c ({signal_3476, signal_1093}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1151 ( .s (signal_748), .b ({signal_2871, signal_1736}), .a ({signal_2134, signal_763}), .c ({signal_3105, signal_1094}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1154 ( .s (signal_756), .b ({signal_2849, signal_1727}), .a ({signal_3106, signal_1097}), .c ({signal_3477, signal_1096}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1155 ( .s (signal_748), .b ({signal_2874, signal_1735}), .a ({signal_2132, signal_764}), .c ({signal_3106, signal_1097}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1158 ( .s (signal_756), .b ({signal_2852, signal_1726}), .a ({signal_3107, signal_1100}), .c ({signal_3478, signal_1099}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1159 ( .s (signal_748), .b ({signal_2877, signal_1734}), .a ({signal_2130, signal_765}), .c ({signal_3107, signal_1100}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1162 ( .s (signal_757), .b ({signal_2855, signal_1717}), .a ({signal_3108, signal_1103}), .c ({signal_3479, signal_1102}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1163 ( .s (signal_749), .b ({signal_2880, signal_1725}), .a ({signal_2567, signal_1909}), .c ({signal_3108, signal_1103}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1166 ( .s (signal_757), .b ({signal_2858, signal_1716}), .a ({signal_3109, signal_1106}), .c ({signal_3480, signal_1105}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1167 ( .s (signal_749), .b ({signal_2883, signal_1724}), .a ({signal_2570, signal_1908}), .c ({signal_3109, signal_1106}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1170 ( .s (signal_757), .b ({signal_2861, signal_1715}), .a ({signal_3110, signal_1109}), .c ({signal_3481, signal_1108}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1171 ( .s (signal_749), .b ({signal_2886, signal_1723}), .a ({signal_2573, signal_1907}), .c ({signal_3110, signal_1109}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1174 ( .s (signal_757), .b ({signal_2864, signal_1714}), .a ({signal_3111, signal_1112}), .c ({signal_3482, signal_1111}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1175 ( .s (signal_749), .b ({signal_2889, signal_1722}), .a ({signal_2576, signal_1906}), .c ({signal_3111, signal_1112}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1178 ( .s (signal_757), .b ({signal_2867, signal_1713}), .a ({signal_3112, signal_1115}), .c ({signal_3483, signal_1114}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1179 ( .s (signal_749), .b ({signal_2892, signal_1721}), .a ({signal_2579, signal_1905}), .c ({signal_3112, signal_1115}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1182 ( .s (signal_757), .b ({signal_2870, signal_1712}), .a ({signal_3113, signal_1118}), .c ({signal_3484, signal_1117}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1183 ( .s (signal_749), .b ({signal_2895, signal_1720}), .a ({signal_2582, signal_1904}), .c ({signal_3113, signal_1118}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1186 ( .s (signal_757), .b ({signal_2873, signal_1711}), .a ({signal_3114, signal_1121}), .c ({signal_3485, signal_1120}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1187 ( .s (signal_749), .b ({signal_2898, signal_1719}), .a ({signal_2585, signal_1903}), .c ({signal_3114, signal_1121}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1190 ( .s (signal_757), .b ({signal_2876, signal_1710}), .a ({signal_3115, signal_1124}), .c ({signal_3486, signal_1123}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1191 ( .s (signal_749), .b ({signal_2901, signal_1718}), .a ({signal_2588, signal_1902}), .c ({signal_3115, signal_1124}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1194 ( .s (signal_757), .b ({signal_2879, signal_1701}), .a ({signal_3116, signal_1127}), .c ({signal_3487, signal_1126}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1195 ( .s (signal_749), .b ({signal_2903, signal_1709}), .a ({signal_2591, signal_1893}), .c ({signal_3116, signal_1127}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1198 ( .s (signal_757), .b ({signal_2882, signal_1700}), .a ({signal_3117, signal_1130}), .c ({signal_3488, signal_1129}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1199 ( .s (signal_749), .b ({signal_2905, signal_1708}), .a ({signal_2594, signal_1892}), .c ({signal_3117, signal_1130}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1202 ( .s (signal_757), .b ({signal_2885, signal_1699}), .a ({signal_3118, signal_1133}), .c ({signal_3489, signal_1132}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1203 ( .s (signal_749), .b ({signal_2907, signal_1707}), .a ({signal_2597, signal_1891}), .c ({signal_3118, signal_1133}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1206 ( .s (signal_757), .b ({signal_2888, signal_1698}), .a ({signal_3119, signal_1136}), .c ({signal_3490, signal_1135}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1207 ( .s (signal_749), .b ({signal_2909, signal_1706}), .a ({signal_2600, signal_1890}), .c ({signal_3119, signal_1136}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1210 ( .s (signal_757), .b ({signal_2891, signal_1697}), .a ({signal_3120, signal_1139}), .c ({signal_3491, signal_1138}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1211 ( .s (signal_749), .b ({signal_2911, signal_1705}), .a ({signal_2603, signal_1889}), .c ({signal_3120, signal_1139}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1214 ( .s (signal_757), .b ({signal_2894, signal_1696}), .a ({signal_3121, signal_1142}), .c ({signal_3492, signal_1141}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1215 ( .s (signal_749), .b ({signal_2913, signal_1704}), .a ({signal_2606, signal_1888}), .c ({signal_3121, signal_1142}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1218 ( .s (signal_757), .b ({signal_2897, signal_1695}), .a ({signal_3122, signal_1145}), .c ({signal_3493, signal_1144}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1219 ( .s (signal_749), .b ({signal_2915, signal_1703}), .a ({signal_2609, signal_1887}), .c ({signal_3122, signal_1145}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1222 ( .s (signal_757), .b ({signal_2900, signal_1694}), .a ({signal_3123, signal_1148}), .c ({signal_3494, signal_1147}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1223 ( .s (signal_749), .b ({signal_2917, signal_1702}), .a ({signal_2612, signal_1886}), .c ({signal_3123, signal_1148}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1226 ( .s (signal_400), .b ({signal_2144, signal_758}), .a ({signal_2145, signal_1693}), .c ({signal_3233, signal_1685}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1227 ( .s (signal_400), .b ({signal_2142, signal_759}), .a ({signal_2143, signal_1692}), .c ({signal_3234, signal_1684}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1228 ( .s (signal_400), .b ({signal_2140, signal_760}), .a ({signal_2141, signal_1691}), .c ({signal_3235, signal_1683}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1229 ( .s (signal_400), .b ({signal_2138, signal_761}), .a ({signal_2139, signal_1690}), .c ({signal_3236, signal_1682}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1230 ( .s (signal_400), .b ({signal_2136, signal_762}), .a ({signal_2137, signal_1689}), .c ({signal_3237, signal_1681}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1231 ( .s (signal_400), .b ({signal_2134, signal_763}), .a ({signal_2135, signal_1688}), .c ({signal_3238, signal_1680}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1232 ( .s (signal_400), .b ({signal_2132, signal_764}), .a ({signal_2133, signal_1687}), .c ({signal_3239, signal_1679}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1233 ( .s (signal_400), .b ({signal_2130, signal_765}), .a ({signal_2131, signal_1686}), .c ({signal_3240, signal_1678}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1234 ( .s (signal_733), .b ({key_s1[120], key_s0[120]}), .a ({signal_3233, signal_1685}), .c ({signal_3371, signal_1933}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1235 ( .s (signal_733), .b ({key_s1[121], key_s0[121]}), .a ({signal_3234, signal_1684}), .c ({signal_3373, signal_1932}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1236 ( .s (signal_733), .b ({key_s1[122], key_s0[122]}), .a ({signal_3235, signal_1683}), .c ({signal_3375, signal_1931}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1237 ( .s (signal_733), .b ({key_s1[123], key_s0[123]}), .a ({signal_3236, signal_1682}), .c ({signal_3377, signal_1930}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1238 ( .s (signal_733), .b ({key_s1[124], key_s0[124]}), .a ({signal_3237, signal_1681}), .c ({signal_3379, signal_1929}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1239 ( .s (signal_733), .b ({key_s1[125], key_s0[125]}), .a ({signal_3238, signal_1680}), .c ({signal_3381, signal_1928}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1240 ( .s (signal_733), .b ({key_s1[126], key_s0[126]}), .a ({signal_3239, signal_1679}), .c ({signal_3383, signal_1927}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1241 ( .s (signal_733), .b ({key_s1[127], key_s0[127]}), .a ({signal_3240, signal_1678}), .c ({signal_3385, signal_1926}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1242 ( .s (signal_733), .b ({key_s1[112], key_s0[112]}), .a ({signal_2567, signal_1909}), .c ({signal_2568, signal_1925}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1243 ( .s (signal_733), .b ({key_s1[113], key_s0[113]}), .a ({signal_2570, signal_1908}), .c ({signal_2571, signal_1924}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1244 ( .s (signal_733), .b ({key_s1[114], key_s0[114]}), .a ({signal_2573, signal_1907}), .c ({signal_2574, signal_1923}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1245 ( .s (signal_733), .b ({key_s1[115], key_s0[115]}), .a ({signal_2576, signal_1906}), .c ({signal_2577, signal_1922}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1246 ( .s (signal_733), .b ({key_s1[116], key_s0[116]}), .a ({signal_2579, signal_1905}), .c ({signal_2580, signal_1921}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1247 ( .s (signal_733), .b ({key_s1[117], key_s0[117]}), .a ({signal_2582, signal_1904}), .c ({signal_2583, signal_1920}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1248 ( .s (signal_733), .b ({key_s1[118], key_s0[118]}), .a ({signal_2585, signal_1903}), .c ({signal_2586, signal_1919}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1249 ( .s (signal_733), .b ({key_s1[119], key_s0[119]}), .a ({signal_2588, signal_1902}), .c ({signal_2589, signal_1918}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1250 ( .s (signal_734), .b ({key_s1[104], key_s0[104]}), .a ({signal_2591, signal_1893}), .c ({signal_2592, signal_1917}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1251 ( .s (signal_734), .b ({key_s1[105], key_s0[105]}), .a ({signal_2594, signal_1892}), .c ({signal_2595, signal_1916}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1252 ( .s (signal_734), .b ({key_s1[106], key_s0[106]}), .a ({signal_2597, signal_1891}), .c ({signal_2598, signal_1915}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1253 ( .s (signal_734), .b ({key_s1[107], key_s0[107]}), .a ({signal_2600, signal_1890}), .c ({signal_2601, signal_1914}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1254 ( .s (signal_734), .b ({key_s1[108], key_s0[108]}), .a ({signal_2603, signal_1889}), .c ({signal_2604, signal_1913}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1255 ( .s (signal_734), .b ({key_s1[109], key_s0[109]}), .a ({signal_2606, signal_1888}), .c ({signal_2607, signal_1912}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1256 ( .s (signal_734), .b ({key_s1[110], key_s0[110]}), .a ({signal_2609, signal_1887}), .c ({signal_2610, signal_1911}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1257 ( .s (signal_734), .b ({key_s1[111], key_s0[111]}), .a ({signal_2612, signal_1886}), .c ({signal_2613, signal_1910}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1258 ( .s (signal_734), .b ({key_s1[96], key_s0[96]}), .a ({signal_2615, signal_1877}), .c ({signal_2616, signal_1901}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1259 ( .s (signal_734), .b ({key_s1[97], key_s0[97]}), .a ({signal_2618, signal_1876}), .c ({signal_2619, signal_1900}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1260 ( .s (signal_734), .b ({key_s1[98], key_s0[98]}), .a ({signal_2621, signal_1875}), .c ({signal_2622, signal_1899}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1261 ( .s (signal_734), .b ({key_s1[99], key_s0[99]}), .a ({signal_2624, signal_1874}), .c ({signal_2625, signal_1898}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1262 ( .s (signal_734), .b ({key_s1[100], key_s0[100]}), .a ({signal_2627, signal_1873}), .c ({signal_2628, signal_1897}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1263 ( .s (signal_734), .b ({key_s1[101], key_s0[101]}), .a ({signal_2630, signal_1872}), .c ({signal_2631, signal_1896}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1264 ( .s (signal_734), .b ({key_s1[102], key_s0[102]}), .a ({signal_2633, signal_1871}), .c ({signal_2634, signal_1895}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1265 ( .s (signal_734), .b ({key_s1[103], key_s0[103]}), .a ({signal_2636, signal_1870}), .c ({signal_2637, signal_1894}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1266 ( .s (signal_735), .b ({key_s1[88], key_s0[88]}), .a ({signal_2639, signal_1861}), .c ({signal_2640, signal_1885}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1267 ( .s (signal_735), .b ({key_s1[89], key_s0[89]}), .a ({signal_2642, signal_1860}), .c ({signal_2643, signal_1884}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1268 ( .s (signal_735), .b ({key_s1[90], key_s0[90]}), .a ({signal_2645, signal_1859}), .c ({signal_2646, signal_1883}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1269 ( .s (signal_735), .b ({key_s1[91], key_s0[91]}), .a ({signal_2648, signal_1858}), .c ({signal_2649, signal_1882}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1270 ( .s (signal_735), .b ({key_s1[92], key_s0[92]}), .a ({signal_2651, signal_1857}), .c ({signal_2652, signal_1881}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1271 ( .s (signal_735), .b ({key_s1[93], key_s0[93]}), .a ({signal_2654, signal_1856}), .c ({signal_2655, signal_1880}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1272 ( .s (signal_735), .b ({key_s1[94], key_s0[94]}), .a ({signal_2657, signal_1855}), .c ({signal_2658, signal_1879}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1273 ( .s (signal_735), .b ({key_s1[95], key_s0[95]}), .a ({signal_2660, signal_1854}), .c ({signal_2661, signal_1878}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1274 ( .s (signal_735), .b ({key_s1[80], key_s0[80]}), .a ({signal_2663, signal_1845}), .c ({signal_2664, signal_1869}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1275 ( .s (signal_735), .b ({key_s1[81], key_s0[81]}), .a ({signal_2666, signal_1844}), .c ({signal_2667, signal_1868}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1276 ( .s (signal_735), .b ({key_s1[82], key_s0[82]}), .a ({signal_2669, signal_1843}), .c ({signal_2670, signal_1867}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1277 ( .s (signal_735), .b ({key_s1[83], key_s0[83]}), .a ({signal_2672, signal_1842}), .c ({signal_2673, signal_1866}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1278 ( .s (signal_735), .b ({key_s1[84], key_s0[84]}), .a ({signal_2675, signal_1841}), .c ({signal_2676, signal_1865}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1279 ( .s (signal_735), .b ({key_s1[85], key_s0[85]}), .a ({signal_2678, signal_1840}), .c ({signal_2679, signal_1864}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1280 ( .s (signal_735), .b ({key_s1[86], key_s0[86]}), .a ({signal_2681, signal_1839}), .c ({signal_2682, signal_1863}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1281 ( .s (signal_735), .b ({key_s1[87], key_s0[87]}), .a ({signal_2684, signal_1838}), .c ({signal_2685, signal_1862}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1282 ( .s (signal_736), .b ({key_s1[72], key_s0[72]}), .a ({signal_2687, signal_1509}), .c ({signal_2688, signal_1853}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1283 ( .s (signal_736), .b ({key_s1[73], key_s0[73]}), .a ({signal_2690, signal_1508}), .c ({signal_2691, signal_1852}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1284 ( .s (signal_736), .b ({key_s1[74], key_s0[74]}), .a ({signal_2693, signal_1507}), .c ({signal_2694, signal_1851}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1285 ( .s (signal_736), .b ({key_s1[75], key_s0[75]}), .a ({signal_2696, signal_1506}), .c ({signal_2697, signal_1850}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1286 ( .s (signal_736), .b ({key_s1[76], key_s0[76]}), .a ({signal_2699, signal_1505}), .c ({signal_2700, signal_1849}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1287 ( .s (signal_736), .b ({key_s1[77], key_s0[77]}), .a ({signal_2702, signal_1504}), .c ({signal_2703, signal_1848}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1288 ( .s (signal_736), .b ({key_s1[78], key_s0[78]}), .a ({signal_2705, signal_1503}), .c ({signal_2706, signal_1847}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1289 ( .s (signal_736), .b ({key_s1[79], key_s0[79]}), .a ({signal_2708, signal_1502}), .c ({signal_2709, signal_1846}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1290 ( .s (signal_736), .b ({key_s1[64], key_s0[64]}), .a ({signal_2711, signal_1821}), .c ({signal_2712, signal_1837}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1291 ( .s (signal_736), .b ({key_s1[65], key_s0[65]}), .a ({signal_2714, signal_1820}), .c ({signal_2715, signal_1836}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1292 ( .s (signal_736), .b ({key_s1[66], key_s0[66]}), .a ({signal_2717, signal_1819}), .c ({signal_2718, signal_1835}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1293 ( .s (signal_736), .b ({key_s1[67], key_s0[67]}), .a ({signal_2720, signal_1818}), .c ({signal_2721, signal_1834}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1294 ( .s (signal_736), .b ({key_s1[68], key_s0[68]}), .a ({signal_2723, signal_1817}), .c ({signal_2724, signal_1833}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1295 ( .s (signal_736), .b ({key_s1[69], key_s0[69]}), .a ({signal_2726, signal_1816}), .c ({signal_2727, signal_1832}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1296 ( .s (signal_736), .b ({key_s1[70], key_s0[70]}), .a ({signal_2729, signal_1815}), .c ({signal_2730, signal_1831}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1297 ( .s (signal_736), .b ({key_s1[71], key_s0[71]}), .a ({signal_2732, signal_1814}), .c ({signal_2733, signal_1830}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1298 ( .s (signal_737), .b ({key_s1[56], key_s0[56]}), .a ({signal_2735, signal_1805}), .c ({signal_2736, signal_1829}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1299 ( .s (signal_737), .b ({key_s1[57], key_s0[57]}), .a ({signal_2738, signal_1804}), .c ({signal_2739, signal_1828}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1300 ( .s (signal_737), .b ({key_s1[58], key_s0[58]}), .a ({signal_2741, signal_1803}), .c ({signal_2742, signal_1827}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1301 ( .s (signal_737), .b ({key_s1[59], key_s0[59]}), .a ({signal_2744, signal_1802}), .c ({signal_2745, signal_1826}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1302 ( .s (signal_737), .b ({key_s1[60], key_s0[60]}), .a ({signal_2747, signal_1801}), .c ({signal_2748, signal_1825}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1303 ( .s (signal_737), .b ({key_s1[61], key_s0[61]}), .a ({signal_2750, signal_1800}), .c ({signal_2751, signal_1824}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1304 ( .s (signal_737), .b ({key_s1[62], key_s0[62]}), .a ({signal_2753, signal_1799}), .c ({signal_2754, signal_1823}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1305 ( .s (signal_737), .b ({key_s1[63], key_s0[63]}), .a ({signal_2756, signal_1798}), .c ({signal_2757, signal_1822}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1306 ( .s (signal_737), .b ({key_s1[48], key_s0[48]}), .a ({signal_2759, signal_1789}), .c ({signal_2760, signal_1813}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1307 ( .s (signal_737), .b ({key_s1[49], key_s0[49]}), .a ({signal_2762, signal_1788}), .c ({signal_2763, signal_1812}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1308 ( .s (signal_737), .b ({key_s1[50], key_s0[50]}), .a ({signal_2765, signal_1787}), .c ({signal_2766, signal_1811}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1309 ( .s (signal_737), .b ({key_s1[51], key_s0[51]}), .a ({signal_2768, signal_1786}), .c ({signal_2769, signal_1810}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1310 ( .s (signal_737), .b ({key_s1[52], key_s0[52]}), .a ({signal_2771, signal_1785}), .c ({signal_2772, signal_1809}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1311 ( .s (signal_737), .b ({key_s1[53], key_s0[53]}), .a ({signal_2774, signal_1784}), .c ({signal_2775, signal_1808}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1312 ( .s (signal_737), .b ({key_s1[54], key_s0[54]}), .a ({signal_2777, signal_1783}), .c ({signal_2778, signal_1807}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1313 ( .s (signal_737), .b ({key_s1[55], key_s0[55]}), .a ({signal_2780, signal_1782}), .c ({signal_2781, signal_1806}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1314 ( .s (signal_738), .b ({key_s1[40], key_s0[40]}), .a ({signal_2783, signal_1773}), .c ({signal_2784, signal_1797}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1315 ( .s (signal_738), .b ({key_s1[41], key_s0[41]}), .a ({signal_2786, signal_1772}), .c ({signal_2787, signal_1796}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1316 ( .s (signal_738), .b ({key_s1[42], key_s0[42]}), .a ({signal_2789, signal_1771}), .c ({signal_2790, signal_1795}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1317 ( .s (signal_738), .b ({key_s1[43], key_s0[43]}), .a ({signal_2792, signal_1770}), .c ({signal_2793, signal_1794}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1318 ( .s (signal_738), .b ({key_s1[44], key_s0[44]}), .a ({signal_2795, signal_1769}), .c ({signal_2796, signal_1793}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1319 ( .s (signal_738), .b ({key_s1[45], key_s0[45]}), .a ({signal_2798, signal_1768}), .c ({signal_2799, signal_1792}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1320 ( .s (signal_738), .b ({key_s1[46], key_s0[46]}), .a ({signal_2801, signal_1767}), .c ({signal_2802, signal_1791}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1321 ( .s (signal_738), .b ({key_s1[47], key_s0[47]}), .a ({signal_2804, signal_1766}), .c ({signal_2805, signal_1790}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1322 ( .s (signal_738), .b ({key_s1[32], key_s0[32]}), .a ({signal_2807, signal_1749}), .c ({signal_2808, signal_1781}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1323 ( .s (signal_738), .b ({key_s1[33], key_s0[33]}), .a ({signal_2810, signal_1748}), .c ({signal_2811, signal_1780}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1324 ( .s (signal_738), .b ({key_s1[34], key_s0[34]}), .a ({signal_2813, signal_1747}), .c ({signal_2814, signal_1779}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1325 ( .s (signal_738), .b ({key_s1[35], key_s0[35]}), .a ({signal_2816, signal_1746}), .c ({signal_2817, signal_1778}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1326 ( .s (signal_738), .b ({key_s1[36], key_s0[36]}), .a ({signal_2819, signal_1745}), .c ({signal_2820, signal_1777}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1327 ( .s (signal_738), .b ({key_s1[37], key_s0[37]}), .a ({signal_2822, signal_1744}), .c ({signal_2823, signal_1776}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1328 ( .s (signal_738), .b ({key_s1[38], key_s0[38]}), .a ({signal_2825, signal_1743}), .c ({signal_2826, signal_1775}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1329 ( .s (signal_738), .b ({key_s1[39], key_s0[39]}), .a ({signal_2828, signal_1742}), .c ({signal_2829, signal_1774}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1330 ( .s (signal_739), .b ({key_s1[24], key_s0[24]}), .a ({signal_2831, signal_1733}), .c ({signal_2832, signal_1765}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1331 ( .s (signal_739), .b ({key_s1[25], key_s0[25]}), .a ({signal_2834, signal_1732}), .c ({signal_2835, signal_1764}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1332 ( .s (signal_739), .b ({key_s1[26], key_s0[26]}), .a ({signal_2837, signal_1731}), .c ({signal_2838, signal_1763}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1333 ( .s (signal_739), .b ({key_s1[27], key_s0[27]}), .a ({signal_2840, signal_1730}), .c ({signal_2841, signal_1762}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1334 ( .s (signal_739), .b ({key_s1[28], key_s0[28]}), .a ({signal_2843, signal_1729}), .c ({signal_2844, signal_1761}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1335 ( .s (signal_739), .b ({key_s1[29], key_s0[29]}), .a ({signal_2846, signal_1728}), .c ({signal_2847, signal_1760}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1336 ( .s (signal_739), .b ({key_s1[30], key_s0[30]}), .a ({signal_2849, signal_1727}), .c ({signal_2850, signal_1759}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1337 ( .s (signal_739), .b ({key_s1[31], key_s0[31]}), .a ({signal_2852, signal_1726}), .c ({signal_2853, signal_1758}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1338 ( .s (signal_739), .b ({key_s1[16], key_s0[16]}), .a ({signal_2855, signal_1717}), .c ({signal_2856, signal_1741}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1339 ( .s (signal_739), .b ({key_s1[17], key_s0[17]}), .a ({signal_2858, signal_1716}), .c ({signal_2859, signal_1740}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1340 ( .s (signal_739), .b ({key_s1[18], key_s0[18]}), .a ({signal_2861, signal_1715}), .c ({signal_2862, signal_1739}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1341 ( .s (signal_739), .b ({key_s1[19], key_s0[19]}), .a ({signal_2864, signal_1714}), .c ({signal_2865, signal_1738}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1342 ( .s (signal_739), .b ({key_s1[20], key_s0[20]}), .a ({signal_2867, signal_1713}), .c ({signal_2868, signal_1737}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1343 ( .s (signal_739), .b ({key_s1[21], key_s0[21]}), .a ({signal_2870, signal_1712}), .c ({signal_2871, signal_1736}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1344 ( .s (signal_739), .b ({key_s1[22], key_s0[22]}), .a ({signal_2873, signal_1711}), .c ({signal_2874, signal_1735}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1345 ( .s (signal_739), .b ({key_s1[23], key_s0[23]}), .a ({signal_2876, signal_1710}), .c ({signal_2877, signal_1734}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1346 ( .s (signal_740), .b ({key_s1[8], key_s0[8]}), .a ({signal_2879, signal_1701}), .c ({signal_2880, signal_1725}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1347 ( .s (signal_740), .b ({key_s1[9], key_s0[9]}), .a ({signal_2882, signal_1700}), .c ({signal_2883, signal_1724}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1348 ( .s (signal_740), .b ({key_s1[10], key_s0[10]}), .a ({signal_2885, signal_1699}), .c ({signal_2886, signal_1723}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1349 ( .s (signal_740), .b ({key_s1[11], key_s0[11]}), .a ({signal_2888, signal_1698}), .c ({signal_2889, signal_1722}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1350 ( .s (signal_740), .b ({key_s1[12], key_s0[12]}), .a ({signal_2891, signal_1697}), .c ({signal_2892, signal_1721}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1351 ( .s (signal_740), .b ({key_s1[13], key_s0[13]}), .a ({signal_2894, signal_1696}), .c ({signal_2895, signal_1720}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1352 ( .s (signal_740), .b ({key_s1[14], key_s0[14]}), .a ({signal_2897, signal_1695}), .c ({signal_2898, signal_1719}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1353 ( .s (signal_740), .b ({key_s1[15], key_s0[15]}), .a ({signal_2900, signal_1694}), .c ({signal_2901, signal_1718}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1354 ( .s (signal_740), .b ({key_s1[0], key_s0[0]}), .a ({signal_2107, signal_1493}), .c ({signal_2903, signal_1709}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1355 ( .s (signal_740), .b ({key_s1[1], key_s0[1]}), .a ({signal_2110, signal_1492}), .c ({signal_2905, signal_1708}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1356 ( .s (signal_740), .b ({key_s1[2], key_s0[2]}), .a ({signal_2113, signal_1491}), .c ({signal_2907, signal_1707}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1357 ( .s (signal_740), .b ({key_s1[3], key_s0[3]}), .a ({signal_2116, signal_1490}), .c ({signal_2909, signal_1706}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1358 ( .s (signal_740), .b ({key_s1[4], key_s0[4]}), .a ({signal_2119, signal_1489}), .c ({signal_2911, signal_1705}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1359 ( .s (signal_740), .b ({key_s1[5], key_s0[5]}), .a ({signal_2122, signal_1488}), .c ({signal_2913, signal_1704}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1360 ( .s (signal_740), .b ({key_s1[6], key_s0[6]}), .a ({signal_2125, signal_1487}), .c ({signal_2915, signal_1703}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1361 ( .s (signal_740), .b ({key_s1[7], key_s0[7]}), .a ({signal_2128, signal_1486}), .c ({signal_2917, signal_1702}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1362 ( .a ({signal_2246, signal_1150}), .b ({signal_2148, signal_1151}), .c ({signal_2918, signal_1454}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1363 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .c ({signal_2148, signal_1151}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1364 ( .a ({ciphertext_s1[126], ciphertext_s0[126]}), .b ({signal_2175, signal_1934}), .c ({signal_2246, signal_1150}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1365 ( .a ({signal_2247, signal_1152}), .b ({signal_2151, signal_1153}), .c ({signal_2919, signal_1455}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1366 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({ciphertext_s1[30], ciphertext_s0[30]}), .c ({signal_2151, signal_1153}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1367 ( .a ({ciphertext_s1[125], ciphertext_s0[125]}), .b ({signal_2177, signal_1935}), .c ({signal_2247, signal_1152}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1368 ( .a ({signal_2248, signal_1154}), .b ({signal_2154, signal_1155}), .c ({signal_2920, signal_1456}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1369 ( .a ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({ciphertext_s1[29], ciphertext_s0[29]}), .c ({signal_2154, signal_1155}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1370 ( .a ({ciphertext_s1[124], ciphertext_s0[124]}), .b ({signal_2179, signal_1936}), .c ({signal_2248, signal_1154}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1371 ( .a ({signal_2921, signal_1156}), .b ({signal_2157, signal_1157}), .c ({signal_2962, signal_1457}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1372 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({ciphertext_s1[28], ciphertext_s0[28]}), .c ({signal_2157, signal_1157}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1373 ( .a ({signal_2170, signal_1942}), .b ({signal_2251, signal_1937}), .c ({signal_2921, signal_1156}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1374 ( .a ({signal_2922, signal_1158}), .b ({signal_2160, signal_1159}), .c ({signal_2963, signal_1458}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1375 ( .a ({ciphertext_s1[59], ciphertext_s0[59]}), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .c ({signal_2160, signal_1159}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1376 ( .a ({signal_2171, signal_1943}), .b ({signal_2252, signal_1938}), .c ({signal_2922, signal_1158}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1377 ( .a ({signal_2249, signal_1160}), .b ({signal_2163, signal_1161}), .c ({signal_2923, signal_1459}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1378 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({signal_2163, signal_1161}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1379 ( .a ({ciphertext_s1[121], ciphertext_s0[121]}), .b ({signal_2182, signal_1939}), .c ({signal_2249, signal_1160}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1380 ( .a ({signal_2924, signal_1162}), .b ({signal_2166, signal_1163}), .c ({signal_2964, signal_1460}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1381 ( .a ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({ciphertext_s1[57], ciphertext_s0[57]}), .c ({signal_2166, signal_1163}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1382 ( .a ({signal_2172, signal_1945}), .b ({signal_2253, signal_1940}), .c ({signal_2924, signal_1162}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1383 ( .a ({signal_2250, signal_1164}), .b ({signal_2169, signal_1165}), .c ({signal_2925, signal_1461}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1384 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .c ({signal_2169, signal_1165}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1385 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({signal_2184, signal_1941}), .c ({signal_2250, signal_1164}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1386 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[123], ciphertext_s0[123]}), .c ({signal_2170, signal_1942}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1387 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({signal_2171, signal_1943}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1388 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[120], ciphertext_s0[120]}), .c ({signal_2172, signal_1945}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1389 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[94], ciphertext_s0[94]}), .c ({signal_2175, signal_1934}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1390 ( .a ({ciphertext_s1[94], ciphertext_s0[94]}), .b ({ciphertext_s1[93], ciphertext_s0[93]}), .c ({signal_2177, signal_1935}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1391 ( .a ({ciphertext_s1[93], ciphertext_s0[93]}), .b ({ciphertext_s1[92], ciphertext_s0[92]}), .c ({signal_2179, signal_1936}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1392 ( .a ({ciphertext_s1[92], ciphertext_s0[92]}), .b ({signal_2186, signal_1946}), .c ({signal_2251, signal_1937}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1393 ( .a ({ciphertext_s1[91], ciphertext_s0[91]}), .b ({signal_2187, signal_1947}), .c ({signal_2252, signal_1938}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1394 ( .a ({ciphertext_s1[90], ciphertext_s0[90]}), .b ({ciphertext_s1[89], ciphertext_s0[89]}), .c ({signal_2182, signal_1939}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1395 ( .a ({ciphertext_s1[89], ciphertext_s0[89]}), .b ({signal_2188, signal_1949}), .c ({signal_2253, signal_1940}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1396 ( .a ({ciphertext_s1[88], ciphertext_s0[88]}), .b ({ciphertext_s1[95], ciphertext_s0[95]}), .c ({signal_2184, signal_1941}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1397 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[91], ciphertext_s0[91]}), .c ({signal_2186, signal_1946}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1398 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({signal_2187, signal_1947}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1399 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .c ({signal_2188, signal_1949}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1400 ( .a ({signal_2254, signal_1166}), .b ({signal_2189, signal_1167}), .c ({signal_2926, signal_1462}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1401 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[127], ciphertext_s0[127]}), .c ({signal_2189, signal_1167}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1402 ( .a ({ciphertext_s1[94], ciphertext_s0[94]}), .b ({signal_2200, signal_1950}), .c ({signal_2254, signal_1166}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1403 ( .a ({signal_2255, signal_1168}), .b ({signal_2190, signal_1169}), .c ({signal_2927, signal_1463}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1404 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({ciphertext_s1[126], ciphertext_s0[126]}), .c ({signal_2190, signal_1169}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1405 ( .a ({ciphertext_s1[93], ciphertext_s0[93]}), .b ({signal_2201, signal_1951}), .c ({signal_2255, signal_1168}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1406 ( .a ({signal_2256, signal_1170}), .b ({signal_2191, signal_1171}), .c ({signal_2928, signal_1464}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1407 ( .a ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({ciphertext_s1[125], ciphertext_s0[125]}), .c ({signal_2191, signal_1171}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1408 ( .a ({ciphertext_s1[92], ciphertext_s0[92]}), .b ({signal_2202, signal_1952}), .c ({signal_2256, signal_1170}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1409 ( .a ({signal_2929, signal_1172}), .b ({signal_2192, signal_1173}), .c ({signal_2965, signal_1465}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1410 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({ciphertext_s1[124], ciphertext_s0[124]}), .c ({signal_2192, signal_1173}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1411 ( .a ({signal_2197, signal_1184}), .b ({signal_2259, signal_1953}), .c ({signal_2929, signal_1172}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1412 ( .a ({signal_2930, signal_1174}), .b ({signal_2193, signal_1175}), .c ({signal_2966, signal_1466}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1413 ( .a ({ciphertext_s1[27], ciphertext_s0[27]}), .b ({ciphertext_s1[123], ciphertext_s0[123]}), .c ({signal_2193, signal_1175}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1414 ( .a ({signal_2198, signal_1183}), .b ({signal_2260, signal_1954}), .c ({signal_2930, signal_1174}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1415 ( .a ({signal_2257, signal_1176}), .b ({signal_2194, signal_1177}), .c ({signal_2931, signal_1467}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1416 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({signal_2194, signal_1177}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1417 ( .a ({ciphertext_s1[89], ciphertext_s0[89]}), .b ({signal_2203, signal_1955}), .c ({signal_2257, signal_1176}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1418 ( .a ({signal_2932, signal_1178}), .b ({signal_2195, signal_1179}), .c ({signal_2967, signal_1468}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1419 ( .a ({ciphertext_s1[121], ciphertext_s0[121]}), .b ({ciphertext_s1[25], ciphertext_s0[25]}), .c ({signal_2195, signal_1179}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1420 ( .a ({signal_2199, signal_1182}), .b ({signal_2261, signal_1956}), .c ({signal_2932, signal_1178}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1421 ( .a ({signal_2258, signal_1180}), .b ({signal_2196, signal_1181}), .c ({signal_2933, signal_1469}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1422 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .c ({signal_2196, signal_1181}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1423 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({signal_2204, signal_1957}), .c ({signal_2258, signal_1180}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1424 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[91], ciphertext_s0[91]}), .c ({signal_2197, signal_1184}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1425 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({signal_2198, signal_1183}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1426 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .c ({signal_2199, signal_1182}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1427 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[62], ciphertext_s0[62]}), .c ({signal_2200, signal_1950}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1428 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({ciphertext_s1[61], ciphertext_s0[61]}), .c ({signal_2201, signal_1951}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1429 ( .a ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({ciphertext_s1[60], ciphertext_s0[60]}), .c ({signal_2202, signal_1952}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1430 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({signal_2205, signal_1958}), .c ({signal_2259, signal_1953}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1431 ( .a ({ciphertext_s1[59], ciphertext_s0[59]}), .b ({signal_2206, signal_1959}), .c ({signal_2260, signal_1954}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1432 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({ciphertext_s1[57], ciphertext_s0[57]}), .c ({signal_2203, signal_1955}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1433 ( .a ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({signal_2207, signal_1961}), .c ({signal_2261, signal_1956}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1434 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .c ({signal_2204, signal_1957}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1435 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .c ({signal_2205, signal_1958}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1436 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({signal_2206, signal_1959}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1437 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .c ({signal_2207, signal_1961}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1438 ( .a ({signal_2262, signal_1185}), .b ({signal_2208, signal_1186}), .c ({signal_2934, signal_1470}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1439 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[95], ciphertext_s0[95]}), .c ({signal_2208, signal_1186}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1440 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({signal_2219, signal_1962}), .c ({signal_2262, signal_1185}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1441 ( .a ({signal_2263, signal_1187}), .b ({signal_2209, signal_1188}), .c ({signal_2935, signal_1471}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1442 ( .a ({ciphertext_s1[126], ciphertext_s0[126]}), .b ({ciphertext_s1[94], ciphertext_s0[94]}), .c ({signal_2209, signal_1188}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1443 ( .a ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({signal_2220, signal_1963}), .c ({signal_2263, signal_1187}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1444 ( .a ({signal_2264, signal_1189}), .b ({signal_2210, signal_1190}), .c ({signal_2936, signal_1472}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1445 ( .a ({ciphertext_s1[125], ciphertext_s0[125]}), .b ({ciphertext_s1[93], ciphertext_s0[93]}), .c ({signal_2210, signal_1190}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1446 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({signal_2221, signal_1964}), .c ({signal_2264, signal_1189}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1447 ( .a ({signal_2937, signal_1191}), .b ({signal_2211, signal_1192}), .c ({signal_2968, signal_1473}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1448 ( .a ({ciphertext_s1[124], ciphertext_s0[124]}), .b ({ciphertext_s1[92], ciphertext_s0[92]}), .c ({signal_2211, signal_1192}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1449 ( .a ({signal_2216, signal_1203}), .b ({signal_2267, signal_1965}), .c ({signal_2937, signal_1191}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1450 ( .a ({signal_2938, signal_1193}), .b ({signal_2212, signal_1194}), .c ({signal_2969, signal_1474}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1451 ( .a ({ciphertext_s1[123], ciphertext_s0[123]}), .b ({ciphertext_s1[91], ciphertext_s0[91]}), .c ({signal_2212, signal_1194}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1452 ( .a ({signal_2217, signal_1202}), .b ({signal_2268, signal_1966}), .c ({signal_2938, signal_1193}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1453 ( .a ({signal_2265, signal_1195}), .b ({signal_2213, signal_1196}), .c ({signal_2939, signal_1475}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1454 ( .a ({ciphertext_s1[122], ciphertext_s0[122]}), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({signal_2213, signal_1196}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1455 ( .a ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({signal_2222, signal_1967}), .c ({signal_2265, signal_1195}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1456 ( .a ({signal_2940, signal_1197}), .b ({signal_2214, signal_1198}), .c ({signal_2970, signal_1476}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1457 ( .a ({ciphertext_s1[89], ciphertext_s0[89]}), .b ({ciphertext_s1[121], ciphertext_s0[121]}), .c ({signal_2214, signal_1198}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1458 ( .a ({signal_2218, signal_1201}), .b ({signal_2269, signal_1968}), .c ({signal_2940, signal_1197}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1459 ( .a ({signal_2266, signal_1199}), .b ({signal_2215, signal_1200}), .c ({signal_2941, signal_1477}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1460 ( .a ({ciphertext_s1[88], ciphertext_s0[88]}), .b ({ciphertext_s1[120], ciphertext_s0[120]}), .c ({signal_2215, signal_1200}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1461 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({signal_2223, signal_1969}), .c ({signal_2266, signal_1199}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1462 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .c ({signal_2216, signal_1203}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1463 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({signal_2217, signal_1202}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1464 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .c ({signal_2218, signal_1201}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1465 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[30], ciphertext_s0[30]}), .c ({signal_2219, signal_1962}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1466 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({ciphertext_s1[29], ciphertext_s0[29]}), .c ({signal_2220, signal_1963}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1467 ( .a ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({ciphertext_s1[28], ciphertext_s0[28]}), .c ({signal_2221, signal_1964}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1468 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({signal_2224, signal_1970}), .c ({signal_2267, signal_1965}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1469 ( .a ({ciphertext_s1[27], ciphertext_s0[27]}), .b ({signal_2225, signal_1971}), .c ({signal_2268, signal_1966}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1470 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({ciphertext_s1[25], ciphertext_s0[25]}), .c ({signal_2222, signal_1967}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1471 ( .a ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({signal_2226, signal_1973}), .c ({signal_2269, signal_1968}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1472 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .c ({signal_2223, signal_1969}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1473 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .c ({signal_2224, signal_1970}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1474 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({signal_2225, signal_1971}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1475 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .c ({signal_2226, signal_1973}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1476 ( .a ({signal_2270, signal_1204}), .b ({signal_2227, signal_1205}), .c ({signal_2942, signal_1478}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1477 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .c ({signal_2227, signal_1205}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1478 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({signal_2238, signal_1974}), .c ({signal_2270, signal_1204}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1479 ( .a ({signal_2271, signal_1206}), .b ({signal_2228, signal_1207}), .c ({signal_2943, signal_1479}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1480 ( .a ({ciphertext_s1[94], ciphertext_s0[94]}), .b ({ciphertext_s1[62], ciphertext_s0[62]}), .c ({signal_2228, signal_1207}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1481 ( .a ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({signal_2239, signal_1975}), .c ({signal_2271, signal_1206}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1482 ( .a ({signal_2272, signal_1208}), .b ({signal_2229, signal_1209}), .c ({signal_2944, signal_1480}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1483 ( .a ({ciphertext_s1[93], ciphertext_s0[93]}), .b ({ciphertext_s1[61], ciphertext_s0[61]}), .c ({signal_2229, signal_1209}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1484 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({signal_2240, signal_1976}), .c ({signal_2272, signal_1208}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1485 ( .a ({signal_2945, signal_1210}), .b ({signal_2230, signal_1211}), .c ({signal_2971, signal_1481}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1486 ( .a ({ciphertext_s1[92], ciphertext_s0[92]}), .b ({ciphertext_s1[60], ciphertext_s0[60]}), .c ({signal_2230, signal_1211}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1487 ( .a ({signal_2235, signal_1222}), .b ({signal_2275, signal_1977}), .c ({signal_2945, signal_1210}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1488 ( .a ({signal_2946, signal_1212}), .b ({signal_2231, signal_1213}), .c ({signal_2972, signal_1482}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1489 ( .a ({ciphertext_s1[91], ciphertext_s0[91]}), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .c ({signal_2231, signal_1213}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1490 ( .a ({signal_2236, signal_1221}), .b ({signal_2276, signal_1978}), .c ({signal_2946, signal_1212}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1491 ( .a ({signal_2273, signal_1214}), .b ({signal_2232, signal_1215}), .c ({signal_2947, signal_1483}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1492 ( .a ({ciphertext_s1[90], ciphertext_s0[90]}), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({signal_2232, signal_1215}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1493 ( .a ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({signal_2241, signal_1979}), .c ({signal_2273, signal_1214}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1494 ( .a ({signal_2948, signal_1216}), .b ({signal_2233, signal_1217}), .c ({signal_2973, signal_1484}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1495 ( .a ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({ciphertext_s1[89], ciphertext_s0[89]}), .c ({signal_2233, signal_1217}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1496 ( .a ({signal_2237, signal_1220}), .b ({signal_2277, signal_1980}), .c ({signal_2948, signal_1216}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1497 ( .a ({signal_2274, signal_1218}), .b ({signal_2234, signal_1219}), .c ({signal_2949, signal_1485}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1498 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .c ({signal_2234, signal_1219}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1499 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({signal_2242, signal_1981}), .c ({signal_2274, signal_1218}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1500 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .c ({signal_2235, signal_1222}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1501 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({signal_2236, signal_1221}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1502 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .c ({signal_2237, signal_1220}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1503 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[126], ciphertext_s0[126]}), .c ({signal_2238, signal_1974}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1504 ( .a ({ciphertext_s1[126], ciphertext_s0[126]}), .b ({ciphertext_s1[125], ciphertext_s0[125]}), .c ({signal_2239, signal_1975}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1505 ( .a ({ciphertext_s1[125], ciphertext_s0[125]}), .b ({ciphertext_s1[124], ciphertext_s0[124]}), .c ({signal_2240, signal_1976}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1506 ( .a ({ciphertext_s1[124], ciphertext_s0[124]}), .b ({signal_2243, signal_1225}), .c ({signal_2275, signal_1977}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1507 ( .a ({ciphertext_s1[123], ciphertext_s0[123]}), .b ({signal_2244, signal_1224}), .c ({signal_2276, signal_1978}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1508 ( .a ({ciphertext_s1[122], ciphertext_s0[122]}), .b ({ciphertext_s1[121], ciphertext_s0[121]}), .c ({signal_2241, signal_1979}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1509 ( .a ({ciphertext_s1[121], ciphertext_s0[121]}), .b ({signal_2245, signal_1223}), .c ({signal_2277, signal_1980}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1510 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({ciphertext_s1[127], ciphertext_s0[127]}), .c ({signal_2242, signal_1981}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1511 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[123], ciphertext_s0[123]}), .c ({signal_2243, signal_1225}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1512 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({signal_2244, signal_1224}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1513 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[120], ciphertext_s0[120]}), .c ({signal_2245, signal_1223}) ) ;
    NOR2_X1 cell_1514 ( .A1 (signal_1255), .A2 (signal_1226), .ZN (signal_1494) ) ;
    NOR2_X1 cell_1515 ( .A1 (signal_1257), .A2 (signal_1226), .ZN (signal_1495) ) ;
    AND2_X1 cell_1516 ( .A1 (signal_1273), .A2 (signal_397), .ZN (signal_1496) ) ;
    AND2_X1 cell_1517 ( .A1 (signal_1272), .A2 (signal_397), .ZN (signal_1497) ) ;
    NOR2_X1 cell_1518 ( .A1 (signal_1261), .A2 (signal_1226), .ZN (signal_1498) ) ;
    NOR2_X1 cell_1519 ( .A1 (signal_1263), .A2 (signal_1226), .ZN (signal_1499) ) ;
    NOR2_X1 cell_1520 ( .A1 (signal_1265), .A2 (signal_1226), .ZN (signal_1500) ) ;
    NOR2_X1 cell_1521 ( .A1 (signal_1267), .A2 (signal_1226), .ZN (signal_1501) ) ;
    INV_X1 cell_1522 ( .A (signal_397), .ZN (signal_1226) ) ;
    NAND2_X1 cell_1523 ( .A1 (signal_1227), .A2 (signal_1228), .ZN (signal_401) ) ;
    NOR2_X1 cell_1524 ( .A1 (signal_1229), .A2 (signal_1230), .ZN (signal_1228) ) ;
    NAND2_X1 cell_1525 ( .A1 (signal_1231), .A2 (signal_1232), .ZN (signal_1230) ) ;
    NOR2_X1 cell_1526 ( .A1 (signal_1269), .A2 (signal_1261), .ZN (signal_1232) ) ;
    NOR2_X1 cell_1527 ( .A1 (signal_1274), .A2 (signal_1267), .ZN (signal_1231) ) ;
    NAND2_X1 cell_1528 ( .A1 (signal_1270), .A2 (signal_1254), .ZN (signal_1229) ) ;
    NOR2_X1 cell_1529 ( .A1 (signal_1272), .A2 (signal_1273), .ZN (signal_1227) ) ;
    NAND2_X1 cell_1530 ( .A1 (signal_393), .A2 (signal_1233), .ZN (signal_1275) ) ;
    MUX2_X1 cell_1531 ( .S (signal_1253), .A (signal_1255), .B (signal_1267), .Z (signal_1233) ) ;
    NAND2_X1 cell_1532 ( .A1 (signal_1234), .A2 (signal_1235), .ZN (signal_1266) ) ;
    NAND2_X1 cell_1533 ( .A1 (signal_1236), .A2 (signal_1269), .ZN (signal_1235) ) ;
    NAND2_X1 cell_1534 ( .A1 (signal_1237), .A2 (signal_1238), .ZN (signal_1234) ) ;
    XOR2_X1 cell_1535 ( .A (signal_1268), .B (signal_1254), .Z (signal_1237) ) ;
    NAND2_X1 cell_1536 ( .A1 (signal_393), .A2 (signal_1239), .ZN (signal_1264) ) ;
    MUX2_X1 cell_1537 ( .S (signal_1253), .A (signal_1265), .B (signal_1263), .Z (signal_1239) ) ;
    NAND2_X1 cell_1538 ( .A1 (signal_393), .A2 (signal_1240), .ZN (signal_1262) ) ;
    MUX2_X1 cell_1539 ( .S (signal_1253), .A (signal_1241), .B (signal_1261), .Z (signal_1240) ) ;
    XNOR2_X1 cell_1540 ( .A (signal_1254), .B (signal_1270), .ZN (signal_1241) ) ;
    NAND2_X1 cell_1541 ( .A1 (signal_1242), .A2 (signal_1243), .ZN (signal_1260) ) ;
    NAND2_X1 cell_1542 ( .A1 (signal_1272), .A2 (signal_1236), .ZN (signal_1243) ) ;
    NAND2_X1 cell_1543 ( .A1 (signal_1244), .A2 (signal_1238), .ZN (signal_1242) ) ;
    XOR2_X1 cell_1544 ( .A (signal_1261), .B (signal_1255), .Z (signal_1244) ) ;
    NAND2_X1 cell_1545 ( .A1 (signal_1245), .A2 (signal_1246), .ZN (signal_1259) ) ;
    NAND2_X1 cell_1546 ( .A1 (signal_1272), .A2 (signal_1238), .ZN (signal_1246) ) ;
    NAND2_X1 cell_1547 ( .A1 (signal_1273), .A2 (signal_1236), .ZN (signal_1245) ) ;
    NAND2_X1 cell_1548 ( .A1 (signal_1247), .A2 (signal_1248), .ZN (signal_1258) ) ;
    NAND2_X1 cell_1549 ( .A1 (signal_1273), .A2 (signal_1238), .ZN (signal_1248) ) ;
    NOR2_X1 cell_1550 ( .A1 (signal_1253), .A2 (signal_1252), .ZN (signal_1238) ) ;
    NAND2_X1 cell_1551 ( .A1 (signal_1274), .A2 (signal_1236), .ZN (signal_1247) ) ;
    NOR2_X1 cell_1552 ( .A1 (signal_395), .A2 (signal_1252), .ZN (signal_1236) ) ;
    NAND2_X1 cell_1553 ( .A1 (signal_393), .A2 (signal_1249), .ZN (signal_1256) ) ;
    MUX2_X1 cell_1554 ( .S (signal_1253), .A (signal_1257), .B (signal_1255), .Z (signal_1249) ) ;
    NAND2_X1 cell_1555 ( .A1 (signal_1272), .A2 (signal_1270), .ZN (signal_1251) ) ;
    NAND2_X1 cell_1556 ( .A1 (signal_1269), .A2 (signal_1273), .ZN (signal_1250) ) ;
    INV_X1 cell_1557 ( .A (signal_393), .ZN (signal_1252) ) ;
    INV_X1 cell_1558 ( .A (signal_395), .ZN (signal_1253) ) ;
    NOR2_X1 cell_1559 ( .A1 (signal_1250), .A2 (signal_1251), .ZN (signal_399) ) ;
    INV_X1 cell_1560 ( .A (signal_1268), .ZN (signal_1267) ) ;
    INV_X1 cell_1562 ( .A (signal_1269), .ZN (signal_1265) ) ;
    INV_X1 cell_1564 ( .A (signal_1270), .ZN (signal_1263) ) ;
    INV_X1 cell_1566 ( .A (signal_1271), .ZN (signal_1261) ) ;
    INV_X1 cell_1572 ( .A (signal_1274), .ZN (signal_1257) ) ;
    INV_X1 cell_1574 ( .A (signal_1254), .ZN (signal_1255) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1576 ( .s (signal_394), .b ({signal_2108, signal_1413}), .a ({signal_2687, signal_1509}), .c ({signal_2950, signal_1517}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1577 ( .s (signal_394), .b ({signal_2111, signal_1412}), .a ({signal_2690, signal_1508}), .c ({signal_2951, signal_1516}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1578 ( .s (signal_394), .b ({signal_2114, signal_1411}), .a ({signal_2693, signal_1507}), .c ({signal_2952, signal_1515}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1579 ( .s (signal_394), .b ({signal_2117, signal_1410}), .a ({signal_2696, signal_1506}), .c ({signal_2953, signal_1514}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1580 ( .s (signal_394), .b ({signal_2120, signal_1409}), .a ({signal_2699, signal_1505}), .c ({signal_2954, signal_1513}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1581 ( .s (signal_394), .b ({signal_2123, signal_1408}), .a ({signal_2702, signal_1504}), .c ({signal_2955, signal_1512}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1582 ( .s (signal_394), .b ({signal_2126, signal_1407}), .a ({signal_2705, signal_1503}), .c ({signal_2956, signal_1511}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1583 ( .s (signal_394), .b ({signal_2129, signal_1406}), .a ({signal_2708, signal_1502}), .c ({signal_2957, signal_1510}) ) ;
    INV_X1 cell_1712 ( .A (signal_393), .ZN (signal_402) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1714 ( .a ({signal_2954, signal_1513}), .b ({signal_2957, signal_1510}), .c ({signal_2974, signal_1982}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1715 ( .a ({signal_2952, signal_1515}), .b ({signal_2957, signal_1510}), .c ({signal_2975, signal_1983}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1716 ( .a ({signal_2951, signal_1516}), .b ({signal_2957, signal_1510}), .c ({signal_2976, signal_1984}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1717 ( .a ({signal_2952, signal_1515}), .b ({signal_2954, signal_1513}), .c ({signal_2977, signal_1985}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1718 ( .a ({signal_2951, signal_1516}), .b ({signal_2953, signal_1514}), .c ({signal_2978, signal_1986}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1719 ( .a ({signal_2955, signal_1512}), .b ({signal_2956, signal_1511}), .c ({signal_2979, signal_1987}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1720 ( .a ({signal_2952, signal_1515}), .b ({signal_2956, signal_1511}), .c ({signal_2980, signal_1988}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1721 ( .a ({signal_2952, signal_1515}), .b ({signal_2955, signal_1512}), .c ({signal_2981, signal_1989}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1722 ( .a ({signal_2950, signal_1517}), .b ({signal_2954, signal_1513}), .c ({signal_2982, signal_1990}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1723 ( .a ({signal_2950, signal_1517}), .b ({signal_2951, signal_1516}), .c ({signal_2983, signal_1991}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1724 ( .a ({signal_2974, signal_1982}), .b ({signal_2978, signal_1986}), .c ({signal_3124, signal_1992}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1725 ( .a ({signal_2950, signal_1517}), .b ({signal_2979, signal_1987}), .c ({signal_3125, signal_1993}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1726 ( .a ({signal_2976, signal_1984}), .b ({signal_2977, signal_1985}), .c ({signal_3126, signal_1994}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1727 ( .a ({signal_2978, signal_1986}), .b ({signal_2980, signal_1988}), .c ({signal_3127, signal_1995}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1728 ( .a ({signal_2978, signal_1986}), .b ({signal_2981, signal_1989}), .c ({signal_3128, signal_1996}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1729 ( .a ({signal_2979, signal_1987}), .b ({signal_2982, signal_1990}), .c ({signal_3129, signal_1997}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1730 ( .a ({signal_2979, signal_1987}), .b ({signal_2983, signal_1991}), .c ({signal_3130, signal_1998}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1731 ( .a ({signal_2974, signal_1982}), .b ({signal_2981, signal_1989}), .c ({signal_3131, signal_1999}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1738 ( .a ({signal_2950, signal_1517}), .b ({signal_3124, signal_1992}), .c ({signal_3162, signal_2006}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1739 ( .a ({signal_2979, signal_1987}), .b ({signal_3124, signal_1992}), .c ({signal_3163, signal_2007}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1740 ( .a ({signal_2980, signal_1988}), .b ({signal_3124, signal_1992}), .c ({signal_3164, signal_2008}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1741 ( .a ({signal_3125, signal_1993}), .b ({signal_3128, signal_1996}), .c ({signal_3165, signal_2009}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1742 ( .a ({signal_2974, signal_1982}), .b ({signal_3129, signal_1997}), .c ({signal_3166, signal_2010}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1743 ( .a ({signal_2975, signal_1983}), .b ({signal_3130, signal_1998}), .c ({signal_3167, signal_2011}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1744 ( .a ({signal_2976, signal_1984}), .b ({signal_3128, signal_1996}), .c ({signal_3168, signal_2012}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1748 ( .a ({signal_2975, signal_1983}), .b ({signal_3163, signal_2007}), .c ({signal_3244, signal_2016}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1749 ( .a ({signal_3165, signal_2009}), .b ({signal_3166, signal_2010}), .c ({signal_3245, signal_2017}) ) ;

    /* cells in depth 1 */
    buf_clk cell_1846 ( .C (clk), .D (signal_2008), .Q (signal_3696) ) ;
    buf_clk cell_1848 ( .C (clk), .D (signal_3164), .Q (signal_3698) ) ;
    buf_clk cell_1850 ( .C (clk), .D (signal_2012), .Q (signal_3700) ) ;
    buf_clk cell_1852 ( .C (clk), .D (signal_3168), .Q (signal_3702) ) ;
    buf_clk cell_1854 ( .C (clk), .D (signal_2016), .Q (signal_3704) ) ;
    buf_clk cell_1856 ( .C (clk), .D (signal_3244), .Q (signal_3706) ) ;
    buf_clk cell_1858 ( .C (clk), .D (signal_2017), .Q (signal_3708) ) ;
    buf_clk cell_1860 ( .C (clk), .D (signal_3245), .Q (signal_3710) ) ;
    buf_clk cell_1894 ( .C (clk), .D (signal_399), .Q (signal_3744) ) ;
    buf_clk cell_1902 ( .C (clk), .D (signal_1413), .Q (signal_3752) ) ;
    buf_clk cell_1910 ( .C (clk), .D (signal_2108), .Q (signal_3760) ) ;
    buf_clk cell_1918 ( .C (clk), .D (signal_1412), .Q (signal_3768) ) ;
    buf_clk cell_1926 ( .C (clk), .D (signal_2111), .Q (signal_3776) ) ;
    buf_clk cell_1934 ( .C (clk), .D (signal_1411), .Q (signal_3784) ) ;
    buf_clk cell_1942 ( .C (clk), .D (signal_2114), .Q (signal_3792) ) ;
    buf_clk cell_1950 ( .C (clk), .D (signal_1410), .Q (signal_3800) ) ;
    buf_clk cell_1958 ( .C (clk), .D (signal_2117), .Q (signal_3808) ) ;
    buf_clk cell_1966 ( .C (clk), .D (signal_1409), .Q (signal_3816) ) ;
    buf_clk cell_1974 ( .C (clk), .D (signal_2120), .Q (signal_3824) ) ;
    buf_clk cell_1982 ( .C (clk), .D (signal_1408), .Q (signal_3832) ) ;
    buf_clk cell_1990 ( .C (clk), .D (signal_2123), .Q (signal_3840) ) ;
    buf_clk cell_1998 ( .C (clk), .D (signal_1407), .Q (signal_3848) ) ;
    buf_clk cell_2006 ( .C (clk), .D (signal_2126), .Q (signal_3856) ) ;
    buf_clk cell_2014 ( .C (clk), .D (signal_1406), .Q (signal_3864) ) ;
    buf_clk cell_2022 ( .C (clk), .D (signal_2129), .Q (signal_3872) ) ;
    buf_clk cell_2030 ( .C (clk), .D (signal_464), .Q (signal_3880) ) ;
    buf_clk cell_2038 ( .C (clk), .D (ciphertext_s0[8]), .Q (signal_3888) ) ;
    buf_clk cell_2046 ( .C (clk), .D (ciphertext_s1[8]), .Q (signal_3896) ) ;
    buf_clk cell_2054 ( .C (clk), .D (ciphertext_s0[9]), .Q (signal_3904) ) ;
    buf_clk cell_2062 ( .C (clk), .D (ciphertext_s1[9]), .Q (signal_3912) ) ;
    buf_clk cell_2070 ( .C (clk), .D (ciphertext_s0[10]), .Q (signal_3920) ) ;
    buf_clk cell_2078 ( .C (clk), .D (ciphertext_s1[10]), .Q (signal_3928) ) ;
    buf_clk cell_2086 ( .C (clk), .D (ciphertext_s0[11]), .Q (signal_3936) ) ;
    buf_clk cell_2094 ( .C (clk), .D (ciphertext_s1[11]), .Q (signal_3944) ) ;
    buf_clk cell_2102 ( .C (clk), .D (ciphertext_s0[12]), .Q (signal_3952) ) ;
    buf_clk cell_2110 ( .C (clk), .D (ciphertext_s1[12]), .Q (signal_3960) ) ;
    buf_clk cell_2118 ( .C (clk), .D (ciphertext_s0[13]), .Q (signal_3968) ) ;
    buf_clk cell_2126 ( .C (clk), .D (ciphertext_s1[13]), .Q (signal_3976) ) ;
    buf_clk cell_2134 ( .C (clk), .D (ciphertext_s0[14]), .Q (signal_3984) ) ;
    buf_clk cell_2142 ( .C (clk), .D (ciphertext_s1[14]), .Q (signal_3992) ) ;
    buf_clk cell_2150 ( .C (clk), .D (ciphertext_s0[15]), .Q (signal_4000) ) ;
    buf_clk cell_2158 ( .C (clk), .D (ciphertext_s1[15]), .Q (signal_4008) ) ;
    buf_clk cell_2166 ( .C (clk), .D (signal_455), .Q (signal_4016) ) ;
    buf_clk cell_2174 ( .C (clk), .D (signal_1453), .Q (signal_4024) ) ;
    buf_clk cell_2182 ( .C (clk), .D (signal_2984), .Q (signal_4032) ) ;
    buf_clk cell_2190 ( .C (clk), .D (signal_1452), .Q (signal_4040) ) ;
    buf_clk cell_2198 ( .C (clk), .D (signal_2985), .Q (signal_4048) ) ;
    buf_clk cell_2206 ( .C (clk), .D (signal_1451), .Q (signal_4056) ) ;
    buf_clk cell_2214 ( .C (clk), .D (signal_2958), .Q (signal_4064) ) ;
    buf_clk cell_2222 ( .C (clk), .D (signal_1450), .Q (signal_4072) ) ;
    buf_clk cell_2230 ( .C (clk), .D (signal_2986), .Q (signal_4080) ) ;
    buf_clk cell_2238 ( .C (clk), .D (signal_1449), .Q (signal_4088) ) ;
    buf_clk cell_2246 ( .C (clk), .D (signal_2987), .Q (signal_4096) ) ;
    buf_clk cell_2254 ( .C (clk), .D (signal_1448), .Q (signal_4104) ) ;
    buf_clk cell_2262 ( .C (clk), .D (signal_2959), .Q (signal_4112) ) ;
    buf_clk cell_2270 ( .C (clk), .D (signal_1447), .Q (signal_4120) ) ;
    buf_clk cell_2278 ( .C (clk), .D (signal_2960), .Q (signal_4128) ) ;
    buf_clk cell_2286 ( .C (clk), .D (signal_1446), .Q (signal_4136) ) ;
    buf_clk cell_2294 ( .C (clk), .D (signal_2961), .Q (signal_4144) ) ;
    buf_clk cell_2302 ( .C (clk), .D (signal_452), .Q (signal_4152) ) ;
    buf_clk cell_2310 ( .C (clk), .D (plaintext_s0[0]), .Q (signal_4160) ) ;
    buf_clk cell_2318 ( .C (clk), .D (plaintext_s1[0]), .Q (signal_4168) ) ;
    buf_clk cell_2326 ( .C (clk), .D (plaintext_s0[1]), .Q (signal_4176) ) ;
    buf_clk cell_2334 ( .C (clk), .D (plaintext_s1[1]), .Q (signal_4184) ) ;
    buf_clk cell_2342 ( .C (clk), .D (plaintext_s0[2]), .Q (signal_4192) ) ;
    buf_clk cell_2350 ( .C (clk), .D (plaintext_s1[2]), .Q (signal_4200) ) ;
    buf_clk cell_2358 ( .C (clk), .D (plaintext_s0[3]), .Q (signal_4208) ) ;
    buf_clk cell_2366 ( .C (clk), .D (plaintext_s1[3]), .Q (signal_4216) ) ;
    buf_clk cell_2374 ( .C (clk), .D (plaintext_s0[4]), .Q (signal_4224) ) ;
    buf_clk cell_2382 ( .C (clk), .D (plaintext_s1[4]), .Q (signal_4232) ) ;
    buf_clk cell_2390 ( .C (clk), .D (plaintext_s0[5]), .Q (signal_4240) ) ;
    buf_clk cell_2398 ( .C (clk), .D (plaintext_s1[5]), .Q (signal_4248) ) ;
    buf_clk cell_2406 ( .C (clk), .D (plaintext_s0[6]), .Q (signal_4256) ) ;
    buf_clk cell_2414 ( .C (clk), .D (plaintext_s1[6]), .Q (signal_4264) ) ;
    buf_clk cell_2422 ( .C (clk), .D (plaintext_s0[7]), .Q (signal_4272) ) ;
    buf_clk cell_2430 ( .C (clk), .D (plaintext_s1[7]), .Q (signal_4280) ) ;
    buf_clk cell_2438 ( .C (clk), .D (signal_1486), .Q (signal_4288) ) ;
    buf_clk cell_2446 ( .C (clk), .D (signal_2128), .Q (signal_4296) ) ;
    buf_clk cell_2454 ( .C (clk), .D (signal_1494), .Q (signal_4304) ) ;
    buf_clk cell_2462 ( .C (clk), .D (signal_1487), .Q (signal_4312) ) ;
    buf_clk cell_2470 ( .C (clk), .D (signal_2125), .Q (signal_4320) ) ;
    buf_clk cell_2478 ( .C (clk), .D (signal_1495), .Q (signal_4328) ) ;
    buf_clk cell_2486 ( .C (clk), .D (signal_1488), .Q (signal_4336) ) ;
    buf_clk cell_2494 ( .C (clk), .D (signal_2122), .Q (signal_4344) ) ;
    buf_clk cell_2502 ( .C (clk), .D (signal_1496), .Q (signal_4352) ) ;
    buf_clk cell_2510 ( .C (clk), .D (signal_1489), .Q (signal_4360) ) ;
    buf_clk cell_2518 ( .C (clk), .D (signal_2119), .Q (signal_4368) ) ;
    buf_clk cell_2526 ( .C (clk), .D (signal_1497), .Q (signal_4376) ) ;
    buf_clk cell_2534 ( .C (clk), .D (signal_1490), .Q (signal_4384) ) ;
    buf_clk cell_2542 ( .C (clk), .D (signal_2116), .Q (signal_4392) ) ;
    buf_clk cell_2550 ( .C (clk), .D (signal_1498), .Q (signal_4400) ) ;
    buf_clk cell_2558 ( .C (clk), .D (signal_1491), .Q (signal_4408) ) ;
    buf_clk cell_2566 ( .C (clk), .D (signal_2113), .Q (signal_4416) ) ;
    buf_clk cell_2574 ( .C (clk), .D (signal_1499), .Q (signal_4424) ) ;
    buf_clk cell_2582 ( .C (clk), .D (signal_1492), .Q (signal_4432) ) ;
    buf_clk cell_2590 ( .C (clk), .D (signal_2110), .Q (signal_4440) ) ;
    buf_clk cell_2598 ( .C (clk), .D (signal_1500), .Q (signal_4448) ) ;
    buf_clk cell_2606 ( .C (clk), .D (signal_1493), .Q (signal_4456) ) ;
    buf_clk cell_2614 ( .C (clk), .D (signal_2107), .Q (signal_4464) ) ;
    buf_clk cell_2622 ( .C (clk), .D (signal_1501), .Q (signal_4472) ) ;
    buf_clk cell_2630 ( .C (clk), .D (signal_756), .Q (signal_4480) ) ;
    buf_clk cell_2638 ( .C (clk), .D (signal_1749), .Q (signal_4488) ) ;
    buf_clk cell_2646 ( .C (clk), .D (signal_2807), .Q (signal_4496) ) ;
    buf_clk cell_2654 ( .C (clk), .D (signal_748), .Q (signal_4504) ) ;
    buf_clk cell_2662 ( .C (clk), .D (signal_1765), .Q (signal_4512) ) ;
    buf_clk cell_2670 ( .C (clk), .D (signal_2832), .Q (signal_4520) ) ;
    buf_clk cell_2678 ( .C (clk), .D (signal_1748), .Q (signal_4528) ) ;
    buf_clk cell_2686 ( .C (clk), .D (signal_2810), .Q (signal_4536) ) ;
    buf_clk cell_2694 ( .C (clk), .D (signal_1764), .Q (signal_4544) ) ;
    buf_clk cell_2702 ( .C (clk), .D (signal_2835), .Q (signal_4552) ) ;
    buf_clk cell_2710 ( .C (clk), .D (signal_1747), .Q (signal_4560) ) ;
    buf_clk cell_2718 ( .C (clk), .D (signal_2813), .Q (signal_4568) ) ;
    buf_clk cell_2726 ( .C (clk), .D (signal_1763), .Q (signal_4576) ) ;
    buf_clk cell_2734 ( .C (clk), .D (signal_2838), .Q (signal_4584) ) ;
    buf_clk cell_2742 ( .C (clk), .D (signal_1746), .Q (signal_4592) ) ;
    buf_clk cell_2750 ( .C (clk), .D (signal_2816), .Q (signal_4600) ) ;
    buf_clk cell_2758 ( .C (clk), .D (signal_1762), .Q (signal_4608) ) ;
    buf_clk cell_2766 ( .C (clk), .D (signal_2841), .Q (signal_4616) ) ;
    buf_clk cell_2774 ( .C (clk), .D (signal_1745), .Q (signal_4624) ) ;
    buf_clk cell_2782 ( .C (clk), .D (signal_2819), .Q (signal_4632) ) ;
    buf_clk cell_2790 ( .C (clk), .D (signal_1761), .Q (signal_4640) ) ;
    buf_clk cell_2798 ( .C (clk), .D (signal_2844), .Q (signal_4648) ) ;
    buf_clk cell_2806 ( .C (clk), .D (signal_1744), .Q (signal_4656) ) ;
    buf_clk cell_2814 ( .C (clk), .D (signal_2822), .Q (signal_4664) ) ;
    buf_clk cell_2822 ( .C (clk), .D (signal_1760), .Q (signal_4672) ) ;
    buf_clk cell_2830 ( .C (clk), .D (signal_2847), .Q (signal_4680) ) ;
    buf_clk cell_2838 ( .C (clk), .D (signal_1743), .Q (signal_4688) ) ;
    buf_clk cell_2846 ( .C (clk), .D (signal_2825), .Q (signal_4696) ) ;
    buf_clk cell_2854 ( .C (clk), .D (signal_1759), .Q (signal_4704) ) ;
    buf_clk cell_2862 ( .C (clk), .D (signal_2850), .Q (signal_4712) ) ;
    buf_clk cell_2870 ( .C (clk), .D (signal_1742), .Q (signal_4720) ) ;
    buf_clk cell_2878 ( .C (clk), .D (signal_2828), .Q (signal_4728) ) ;
    buf_clk cell_2886 ( .C (clk), .D (signal_1758), .Q (signal_4736) ) ;
    buf_clk cell_2894 ( .C (clk), .D (signal_2853), .Q (signal_4744) ) ;
    buf_clk cell_2902 ( .C (clk), .D (signal_2006), .Q (signal_4752) ) ;
    buf_clk cell_2908 ( .C (clk), .D (signal_3162), .Q (signal_4758) ) ;
    buf_clk cell_2914 ( .C (clk), .D (signal_1517), .Q (signal_4764) ) ;
    buf_clk cell_2920 ( .C (clk), .D (signal_2950), .Q (signal_4770) ) ;
    buf_clk cell_2926 ( .C (clk), .D (signal_1993), .Q (signal_4776) ) ;
    buf_clk cell_2932 ( .C (clk), .D (signal_3125), .Q (signal_4782) ) ;
    buf_clk cell_2938 ( .C (clk), .D (signal_2009), .Q (signal_4788) ) ;
    buf_clk cell_2944 ( .C (clk), .D (signal_3165), .Q (signal_4794) ) ;
    buf_clk cell_2950 ( .C (clk), .D (signal_2011), .Q (signal_4800) ) ;
    buf_clk cell_2956 ( .C (clk), .D (signal_3167), .Q (signal_4806) ) ;
    buf_clk cell_2962 ( .C (clk), .D (signal_1997), .Q (signal_4812) ) ;
    buf_clk cell_2968 ( .C (clk), .D (signal_3129), .Q (signal_4818) ) ;
    buf_clk cell_2974 ( .C (clk), .D (signal_1998), .Q (signal_4824) ) ;
    buf_clk cell_2980 ( .C (clk), .D (signal_3130), .Q (signal_4830) ) ;
    buf_clk cell_2986 ( .C (clk), .D (signal_2010), .Q (signal_4836) ) ;
    buf_clk cell_2992 ( .C (clk), .D (signal_3166), .Q (signal_4842) ) ;
    buf_clk cell_2998 ( .C (clk), .D (signal_1992), .Q (signal_4848) ) ;
    buf_clk cell_3004 ( .C (clk), .D (signal_3124), .Q (signal_4854) ) ;
    buf_clk cell_3010 ( .C (clk), .D (signal_1996), .Q (signal_4860) ) ;
    buf_clk cell_3016 ( .C (clk), .D (signal_3128), .Q (signal_4866) ) ;
    buf_clk cell_3022 ( .C (clk), .D (signal_1995), .Q (signal_4872) ) ;
    buf_clk cell_3028 ( .C (clk), .D (signal_3127), .Q (signal_4878) ) ;
    buf_clk cell_3034 ( .C (clk), .D (signal_2007), .Q (signal_4884) ) ;
    buf_clk cell_3040 ( .C (clk), .D (signal_3163), .Q (signal_4890) ) ;
    buf_clk cell_3046 ( .C (clk), .D (signal_1994), .Q (signal_4896) ) ;
    buf_clk cell_3052 ( .C (clk), .D (signal_3126), .Q (signal_4902) ) ;
    buf_clk cell_3058 ( .C (clk), .D (signal_1984), .Q (signal_4908) ) ;
    buf_clk cell_3064 ( .C (clk), .D (signal_2976), .Q (signal_4914) ) ;
    buf_clk cell_3070 ( .C (clk), .D (signal_1982), .Q (signal_4920) ) ;
    buf_clk cell_3076 ( .C (clk), .D (signal_2974), .Q (signal_4926) ) ;
    buf_clk cell_3082 ( .C (clk), .D (signal_1983), .Q (signal_4932) ) ;
    buf_clk cell_3088 ( .C (clk), .D (signal_2975), .Q (signal_4938) ) ;
    buf_clk cell_3094 ( .C (clk), .D (signal_1999), .Q (signal_4944) ) ;
    buf_clk cell_3100 ( .C (clk), .D (signal_3131), .Q (signal_4950) ) ;
    buf_clk cell_3106 ( .C (clk), .D (signal_1985), .Q (signal_4956) ) ;
    buf_clk cell_3112 ( .C (clk), .D (signal_2977), .Q (signal_4962) ) ;
    buf_clk cell_3118 ( .C (clk), .D (signal_429), .Q (signal_4968) ) ;
    buf_clk cell_3126 ( .C (clk), .D (signal_431), .Q (signal_4976) ) ;
    buf_clk cell_3134 ( .C (clk), .D (signal_433), .Q (signal_4984) ) ;
    buf_clk cell_3142 ( .C (clk), .D (signal_435), .Q (signal_4992) ) ;
    buf_clk cell_3150 ( .C (clk), .D (signal_437), .Q (signal_5000) ) ;
    buf_clk cell_3158 ( .C (clk), .D (signal_439), .Q (signal_5008) ) ;
    buf_clk cell_3166 ( .C (clk), .D (signal_441), .Q (signal_5016) ) ;
    buf_clk cell_3174 ( .C (clk), .D (signal_419), .Q (signal_5024) ) ;
    buf_clk cell_3182 ( .C (clk), .D (signal_395), .Q (signal_5032) ) ;
    buf_clk cell_3190 ( .C (clk), .D (signal_465), .Q (signal_5040) ) ;
    buf_clk cell_3198 ( .C (clk), .D (signal_3250), .Q (signal_5048) ) ;
    buf_clk cell_3206 ( .C (clk), .D (signal_467), .Q (signal_5056) ) ;
    buf_clk cell_3214 ( .C (clk), .D (signal_3251), .Q (signal_5064) ) ;
    buf_clk cell_3222 ( .C (clk), .D (signal_469), .Q (signal_5072) ) ;
    buf_clk cell_3230 ( .C (clk), .D (signal_3252), .Q (signal_5080) ) ;
    buf_clk cell_3238 ( .C (clk), .D (signal_471), .Q (signal_5088) ) ;
    buf_clk cell_3246 ( .C (clk), .D (signal_3253), .Q (signal_5096) ) ;
    buf_clk cell_3254 ( .C (clk), .D (signal_473), .Q (signal_5104) ) ;
    buf_clk cell_3262 ( .C (clk), .D (signal_3254), .Q (signal_5112) ) ;
    buf_clk cell_3270 ( .C (clk), .D (signal_475), .Q (signal_5120) ) ;
    buf_clk cell_3278 ( .C (clk), .D (signal_3255), .Q (signal_5128) ) ;
    buf_clk cell_3286 ( .C (clk), .D (signal_477), .Q (signal_5136) ) ;
    buf_clk cell_3294 ( .C (clk), .D (signal_3256), .Q (signal_5144) ) ;
    buf_clk cell_3302 ( .C (clk), .D (signal_479), .Q (signal_5152) ) ;
    buf_clk cell_3310 ( .C (clk), .D (signal_3257), .Q (signal_5160) ) ;
    buf_clk cell_3318 ( .C (clk), .D (signal_481), .Q (signal_5168) ) ;
    buf_clk cell_3326 ( .C (clk), .D (signal_3258), .Q (signal_5176) ) ;
    buf_clk cell_3334 ( .C (clk), .D (signal_483), .Q (signal_5184) ) ;
    buf_clk cell_3342 ( .C (clk), .D (signal_3259), .Q (signal_5192) ) ;
    buf_clk cell_3350 ( .C (clk), .D (signal_485), .Q (signal_5200) ) ;
    buf_clk cell_3358 ( .C (clk), .D (signal_3260), .Q (signal_5208) ) ;
    buf_clk cell_3366 ( .C (clk), .D (signal_487), .Q (signal_5216) ) ;
    buf_clk cell_3374 ( .C (clk), .D (signal_3261), .Q (signal_5224) ) ;
    buf_clk cell_3382 ( .C (clk), .D (signal_489), .Q (signal_5232) ) ;
    buf_clk cell_3390 ( .C (clk), .D (signal_3262), .Q (signal_5240) ) ;
    buf_clk cell_3398 ( .C (clk), .D (signal_491), .Q (signal_5248) ) ;
    buf_clk cell_3406 ( .C (clk), .D (signal_3263), .Q (signal_5256) ) ;
    buf_clk cell_3414 ( .C (clk), .D (signal_493), .Q (signal_5264) ) ;
    buf_clk cell_3422 ( .C (clk), .D (signal_3264), .Q (signal_5272) ) ;
    buf_clk cell_3430 ( .C (clk), .D (signal_495), .Q (signal_5280) ) ;
    buf_clk cell_3438 ( .C (clk), .D (signal_3265), .Q (signal_5288) ) ;
    buf_clk cell_3446 ( .C (clk), .D (signal_497), .Q (signal_5296) ) ;
    buf_clk cell_3454 ( .C (clk), .D (signal_3266), .Q (signal_5304) ) ;
    buf_clk cell_3462 ( .C (clk), .D (signal_499), .Q (signal_5312) ) ;
    buf_clk cell_3470 ( .C (clk), .D (signal_3267), .Q (signal_5320) ) ;
    buf_clk cell_3478 ( .C (clk), .D (signal_501), .Q (signal_5328) ) ;
    buf_clk cell_3486 ( .C (clk), .D (signal_3268), .Q (signal_5336) ) ;
    buf_clk cell_3494 ( .C (clk), .D (signal_503), .Q (signal_5344) ) ;
    buf_clk cell_3502 ( .C (clk), .D (signal_3269), .Q (signal_5352) ) ;
    buf_clk cell_3510 ( .C (clk), .D (signal_505), .Q (signal_5360) ) ;
    buf_clk cell_3518 ( .C (clk), .D (signal_3270), .Q (signal_5368) ) ;
    buf_clk cell_3526 ( .C (clk), .D (signal_507), .Q (signal_5376) ) ;
    buf_clk cell_3534 ( .C (clk), .D (signal_3271), .Q (signal_5384) ) ;
    buf_clk cell_3542 ( .C (clk), .D (signal_509), .Q (signal_5392) ) ;
    buf_clk cell_3550 ( .C (clk), .D (signal_3272), .Q (signal_5400) ) ;
    buf_clk cell_3558 ( .C (clk), .D (signal_511), .Q (signal_5408) ) ;
    buf_clk cell_3566 ( .C (clk), .D (signal_3273), .Q (signal_5416) ) ;
    buf_clk cell_3574 ( .C (clk), .D (signal_513), .Q (signal_5424) ) ;
    buf_clk cell_3582 ( .C (clk), .D (signal_3274), .Q (signal_5432) ) ;
    buf_clk cell_3590 ( .C (clk), .D (signal_515), .Q (signal_5440) ) ;
    buf_clk cell_3598 ( .C (clk), .D (signal_3275), .Q (signal_5448) ) ;
    buf_clk cell_3606 ( .C (clk), .D (signal_517), .Q (signal_5456) ) ;
    buf_clk cell_3614 ( .C (clk), .D (signal_3276), .Q (signal_5464) ) ;
    buf_clk cell_3622 ( .C (clk), .D (signal_519), .Q (signal_5472) ) ;
    buf_clk cell_3630 ( .C (clk), .D (signal_3277), .Q (signal_5480) ) ;
    buf_clk cell_3638 ( .C (clk), .D (signal_521), .Q (signal_5488) ) ;
    buf_clk cell_3646 ( .C (clk), .D (signal_3278), .Q (signal_5496) ) ;
    buf_clk cell_3654 ( .C (clk), .D (signal_523), .Q (signal_5504) ) ;
    buf_clk cell_3662 ( .C (clk), .D (signal_3279), .Q (signal_5512) ) ;
    buf_clk cell_3670 ( .C (clk), .D (signal_525), .Q (signal_5520) ) ;
    buf_clk cell_3678 ( .C (clk), .D (signal_3280), .Q (signal_5528) ) ;
    buf_clk cell_3686 ( .C (clk), .D (signal_527), .Q (signal_5536) ) ;
    buf_clk cell_3694 ( .C (clk), .D (signal_3281), .Q (signal_5544) ) ;
    buf_clk cell_3702 ( .C (clk), .D (signal_529), .Q (signal_5552) ) ;
    buf_clk cell_3710 ( .C (clk), .D (signal_3282), .Q (signal_5560) ) ;
    buf_clk cell_3718 ( .C (clk), .D (signal_531), .Q (signal_5568) ) ;
    buf_clk cell_3726 ( .C (clk), .D (signal_3283), .Q (signal_5576) ) ;
    buf_clk cell_3734 ( .C (clk), .D (signal_533), .Q (signal_5584) ) ;
    buf_clk cell_3742 ( .C (clk), .D (signal_3284), .Q (signal_5592) ) ;
    buf_clk cell_3750 ( .C (clk), .D (signal_535), .Q (signal_5600) ) ;
    buf_clk cell_3758 ( .C (clk), .D (signal_3285), .Q (signal_5608) ) ;
    buf_clk cell_3766 ( .C (clk), .D (signal_537), .Q (signal_5616) ) ;
    buf_clk cell_3774 ( .C (clk), .D (signal_3286), .Q (signal_5624) ) ;
    buf_clk cell_3782 ( .C (clk), .D (signal_539), .Q (signal_5632) ) ;
    buf_clk cell_3790 ( .C (clk), .D (signal_3287), .Q (signal_5640) ) ;
    buf_clk cell_3798 ( .C (clk), .D (signal_541), .Q (signal_5648) ) ;
    buf_clk cell_3806 ( .C (clk), .D (signal_3288), .Q (signal_5656) ) ;
    buf_clk cell_3814 ( .C (clk), .D (signal_543), .Q (signal_5664) ) ;
    buf_clk cell_3822 ( .C (clk), .D (signal_3289), .Q (signal_5672) ) ;
    buf_clk cell_3830 ( .C (clk), .D (signal_545), .Q (signal_5680) ) ;
    buf_clk cell_3838 ( .C (clk), .D (signal_3290), .Q (signal_5688) ) ;
    buf_clk cell_3846 ( .C (clk), .D (signal_547), .Q (signal_5696) ) ;
    buf_clk cell_3854 ( .C (clk), .D (signal_3291), .Q (signal_5704) ) ;
    buf_clk cell_3862 ( .C (clk), .D (signal_549), .Q (signal_5712) ) ;
    buf_clk cell_3870 ( .C (clk), .D (signal_3292), .Q (signal_5720) ) ;
    buf_clk cell_3878 ( .C (clk), .D (signal_551), .Q (signal_5728) ) ;
    buf_clk cell_3886 ( .C (clk), .D (signal_3293), .Q (signal_5736) ) ;
    buf_clk cell_3894 ( .C (clk), .D (signal_553), .Q (signal_5744) ) ;
    buf_clk cell_3902 ( .C (clk), .D (signal_3294), .Q (signal_5752) ) ;
    buf_clk cell_3910 ( .C (clk), .D (signal_555), .Q (signal_5760) ) ;
    buf_clk cell_3918 ( .C (clk), .D (signal_3295), .Q (signal_5768) ) ;
    buf_clk cell_3926 ( .C (clk), .D (signal_557), .Q (signal_5776) ) ;
    buf_clk cell_3934 ( .C (clk), .D (signal_3296), .Q (signal_5784) ) ;
    buf_clk cell_3942 ( .C (clk), .D (signal_559), .Q (signal_5792) ) ;
    buf_clk cell_3950 ( .C (clk), .D (signal_3297), .Q (signal_5800) ) ;
    buf_clk cell_3958 ( .C (clk), .D (signal_561), .Q (signal_5808) ) ;
    buf_clk cell_3966 ( .C (clk), .D (signal_3298), .Q (signal_5816) ) ;
    buf_clk cell_3974 ( .C (clk), .D (signal_563), .Q (signal_5824) ) ;
    buf_clk cell_3982 ( .C (clk), .D (signal_3299), .Q (signal_5832) ) ;
    buf_clk cell_3990 ( .C (clk), .D (signal_565), .Q (signal_5840) ) ;
    buf_clk cell_3998 ( .C (clk), .D (signal_3300), .Q (signal_5848) ) ;
    buf_clk cell_4006 ( .C (clk), .D (signal_567), .Q (signal_5856) ) ;
    buf_clk cell_4014 ( .C (clk), .D (signal_3301), .Q (signal_5864) ) ;
    buf_clk cell_4022 ( .C (clk), .D (signal_569), .Q (signal_5872) ) ;
    buf_clk cell_4030 ( .C (clk), .D (signal_3302), .Q (signal_5880) ) ;
    buf_clk cell_4038 ( .C (clk), .D (signal_571), .Q (signal_5888) ) ;
    buf_clk cell_4046 ( .C (clk), .D (signal_3303), .Q (signal_5896) ) ;
    buf_clk cell_4054 ( .C (clk), .D (signal_573), .Q (signal_5904) ) ;
    buf_clk cell_4062 ( .C (clk), .D (signal_3304), .Q (signal_5912) ) ;
    buf_clk cell_4070 ( .C (clk), .D (signal_575), .Q (signal_5920) ) ;
    buf_clk cell_4078 ( .C (clk), .D (signal_3305), .Q (signal_5928) ) ;
    buf_clk cell_4086 ( .C (clk), .D (signal_577), .Q (signal_5936) ) ;
    buf_clk cell_4094 ( .C (clk), .D (signal_3306), .Q (signal_5944) ) ;
    buf_clk cell_4102 ( .C (clk), .D (signal_579), .Q (signal_5952) ) ;
    buf_clk cell_4110 ( .C (clk), .D (signal_3307), .Q (signal_5960) ) ;
    buf_clk cell_4118 ( .C (clk), .D (signal_581), .Q (signal_5968) ) ;
    buf_clk cell_4126 ( .C (clk), .D (signal_3308), .Q (signal_5976) ) ;
    buf_clk cell_4134 ( .C (clk), .D (signal_583), .Q (signal_5984) ) ;
    buf_clk cell_4142 ( .C (clk), .D (signal_3309), .Q (signal_5992) ) ;
    buf_clk cell_4150 ( .C (clk), .D (signal_585), .Q (signal_6000) ) ;
    buf_clk cell_4158 ( .C (clk), .D (signal_3310), .Q (signal_6008) ) ;
    buf_clk cell_4166 ( .C (clk), .D (signal_587), .Q (signal_6016) ) ;
    buf_clk cell_4174 ( .C (clk), .D (signal_3311), .Q (signal_6024) ) ;
    buf_clk cell_4182 ( .C (clk), .D (signal_589), .Q (signal_6032) ) ;
    buf_clk cell_4190 ( .C (clk), .D (signal_3312), .Q (signal_6040) ) ;
    buf_clk cell_4198 ( .C (clk), .D (signal_591), .Q (signal_6048) ) ;
    buf_clk cell_4206 ( .C (clk), .D (signal_3313), .Q (signal_6056) ) ;
    buf_clk cell_4214 ( .C (clk), .D (signal_593), .Q (signal_6064) ) ;
    buf_clk cell_4222 ( .C (clk), .D (signal_3314), .Q (signal_6072) ) ;
    buf_clk cell_4230 ( .C (clk), .D (signal_595), .Q (signal_6080) ) ;
    buf_clk cell_4238 ( .C (clk), .D (signal_3315), .Q (signal_6088) ) ;
    buf_clk cell_4246 ( .C (clk), .D (signal_597), .Q (signal_6096) ) ;
    buf_clk cell_4254 ( .C (clk), .D (signal_3316), .Q (signal_6104) ) ;
    buf_clk cell_4262 ( .C (clk), .D (signal_599), .Q (signal_6112) ) ;
    buf_clk cell_4270 ( .C (clk), .D (signal_3317), .Q (signal_6120) ) ;
    buf_clk cell_4278 ( .C (clk), .D (signal_601), .Q (signal_6128) ) ;
    buf_clk cell_4286 ( .C (clk), .D (signal_3318), .Q (signal_6136) ) ;
    buf_clk cell_4294 ( .C (clk), .D (signal_603), .Q (signal_6144) ) ;
    buf_clk cell_4302 ( .C (clk), .D (signal_3319), .Q (signal_6152) ) ;
    buf_clk cell_4310 ( .C (clk), .D (signal_605), .Q (signal_6160) ) ;
    buf_clk cell_4318 ( .C (clk), .D (signal_3320), .Q (signal_6168) ) ;
    buf_clk cell_4326 ( .C (clk), .D (signal_607), .Q (signal_6176) ) ;
    buf_clk cell_4334 ( .C (clk), .D (signal_3321), .Q (signal_6184) ) ;
    buf_clk cell_4342 ( .C (clk), .D (signal_609), .Q (signal_6192) ) ;
    buf_clk cell_4350 ( .C (clk), .D (signal_3322), .Q (signal_6200) ) ;
    buf_clk cell_4358 ( .C (clk), .D (signal_611), .Q (signal_6208) ) ;
    buf_clk cell_4366 ( .C (clk), .D (signal_3323), .Q (signal_6216) ) ;
    buf_clk cell_4374 ( .C (clk), .D (signal_613), .Q (signal_6224) ) ;
    buf_clk cell_4382 ( .C (clk), .D (signal_3324), .Q (signal_6232) ) ;
    buf_clk cell_4390 ( .C (clk), .D (signal_615), .Q (signal_6240) ) ;
    buf_clk cell_4398 ( .C (clk), .D (signal_3325), .Q (signal_6248) ) ;
    buf_clk cell_4406 ( .C (clk), .D (signal_617), .Q (signal_6256) ) ;
    buf_clk cell_4414 ( .C (clk), .D (signal_3326), .Q (signal_6264) ) ;
    buf_clk cell_4422 ( .C (clk), .D (signal_619), .Q (signal_6272) ) ;
    buf_clk cell_4430 ( .C (clk), .D (signal_3327), .Q (signal_6280) ) ;
    buf_clk cell_4438 ( .C (clk), .D (signal_621), .Q (signal_6288) ) ;
    buf_clk cell_4446 ( .C (clk), .D (signal_3328), .Q (signal_6296) ) ;
    buf_clk cell_4454 ( .C (clk), .D (signal_623), .Q (signal_6304) ) ;
    buf_clk cell_4462 ( .C (clk), .D (signal_3329), .Q (signal_6312) ) ;
    buf_clk cell_4470 ( .C (clk), .D (signal_625), .Q (signal_6320) ) ;
    buf_clk cell_4478 ( .C (clk), .D (signal_3330), .Q (signal_6328) ) ;
    buf_clk cell_4486 ( .C (clk), .D (signal_627), .Q (signal_6336) ) ;
    buf_clk cell_4494 ( .C (clk), .D (signal_3331), .Q (signal_6344) ) ;
    buf_clk cell_4502 ( .C (clk), .D (signal_629), .Q (signal_6352) ) ;
    buf_clk cell_4510 ( .C (clk), .D (signal_3332), .Q (signal_6360) ) ;
    buf_clk cell_4518 ( .C (clk), .D (signal_631), .Q (signal_6368) ) ;
    buf_clk cell_4526 ( .C (clk), .D (signal_3333), .Q (signal_6376) ) ;
    buf_clk cell_4534 ( .C (clk), .D (signal_633), .Q (signal_6384) ) ;
    buf_clk cell_4542 ( .C (clk), .D (signal_3334), .Q (signal_6392) ) ;
    buf_clk cell_4550 ( .C (clk), .D (signal_635), .Q (signal_6400) ) ;
    buf_clk cell_4558 ( .C (clk), .D (signal_3335), .Q (signal_6408) ) ;
    buf_clk cell_4566 ( .C (clk), .D (signal_637), .Q (signal_6416) ) ;
    buf_clk cell_4574 ( .C (clk), .D (signal_3336), .Q (signal_6424) ) ;
    buf_clk cell_4582 ( .C (clk), .D (signal_639), .Q (signal_6432) ) ;
    buf_clk cell_4590 ( .C (clk), .D (signal_3337), .Q (signal_6440) ) ;
    buf_clk cell_4598 ( .C (clk), .D (signal_641), .Q (signal_6448) ) ;
    buf_clk cell_4606 ( .C (clk), .D (signal_3338), .Q (signal_6456) ) ;
    buf_clk cell_4614 ( .C (clk), .D (signal_643), .Q (signal_6464) ) ;
    buf_clk cell_4622 ( .C (clk), .D (signal_3339), .Q (signal_6472) ) ;
    buf_clk cell_4630 ( .C (clk), .D (signal_645), .Q (signal_6480) ) ;
    buf_clk cell_4638 ( .C (clk), .D (signal_3340), .Q (signal_6488) ) ;
    buf_clk cell_4646 ( .C (clk), .D (signal_647), .Q (signal_6496) ) ;
    buf_clk cell_4654 ( .C (clk), .D (signal_3341), .Q (signal_6504) ) ;
    buf_clk cell_4662 ( .C (clk), .D (signal_649), .Q (signal_6512) ) ;
    buf_clk cell_4670 ( .C (clk), .D (signal_3342), .Q (signal_6520) ) ;
    buf_clk cell_4678 ( .C (clk), .D (signal_651), .Q (signal_6528) ) ;
    buf_clk cell_4686 ( .C (clk), .D (signal_3343), .Q (signal_6536) ) ;
    buf_clk cell_4694 ( .C (clk), .D (signal_653), .Q (signal_6544) ) ;
    buf_clk cell_4702 ( .C (clk), .D (signal_3344), .Q (signal_6552) ) ;
    buf_clk cell_4710 ( .C (clk), .D (signal_655), .Q (signal_6560) ) ;
    buf_clk cell_4718 ( .C (clk), .D (signal_3345), .Q (signal_6568) ) ;
    buf_clk cell_4726 ( .C (clk), .D (signal_657), .Q (signal_6576) ) ;
    buf_clk cell_4734 ( .C (clk), .D (signal_3346), .Q (signal_6584) ) ;
    buf_clk cell_4742 ( .C (clk), .D (signal_659), .Q (signal_6592) ) ;
    buf_clk cell_4750 ( .C (clk), .D (signal_3347), .Q (signal_6600) ) ;
    buf_clk cell_4758 ( .C (clk), .D (signal_661), .Q (signal_6608) ) ;
    buf_clk cell_4766 ( .C (clk), .D (signal_3348), .Q (signal_6616) ) ;
    buf_clk cell_4774 ( .C (clk), .D (signal_663), .Q (signal_6624) ) ;
    buf_clk cell_4782 ( .C (clk), .D (signal_3349), .Q (signal_6632) ) ;
    buf_clk cell_4790 ( .C (clk), .D (signal_665), .Q (signal_6640) ) ;
    buf_clk cell_4798 ( .C (clk), .D (signal_3350), .Q (signal_6648) ) ;
    buf_clk cell_4806 ( .C (clk), .D (signal_667), .Q (signal_6656) ) ;
    buf_clk cell_4814 ( .C (clk), .D (signal_3351), .Q (signal_6664) ) ;
    buf_clk cell_4822 ( .C (clk), .D (signal_669), .Q (signal_6672) ) ;
    buf_clk cell_4830 ( .C (clk), .D (signal_3352), .Q (signal_6680) ) ;
    buf_clk cell_4838 ( .C (clk), .D (signal_671), .Q (signal_6688) ) ;
    buf_clk cell_4846 ( .C (clk), .D (signal_3353), .Q (signal_6696) ) ;
    buf_clk cell_4854 ( .C (clk), .D (signal_673), .Q (signal_6704) ) ;
    buf_clk cell_4862 ( .C (clk), .D (signal_3354), .Q (signal_6712) ) ;
    buf_clk cell_4870 ( .C (clk), .D (signal_675), .Q (signal_6720) ) ;
    buf_clk cell_4878 ( .C (clk), .D (signal_3355), .Q (signal_6728) ) ;
    buf_clk cell_4886 ( .C (clk), .D (signal_677), .Q (signal_6736) ) ;
    buf_clk cell_4894 ( .C (clk), .D (signal_3356), .Q (signal_6744) ) ;
    buf_clk cell_4902 ( .C (clk), .D (signal_679), .Q (signal_6752) ) ;
    buf_clk cell_4910 ( .C (clk), .D (signal_3357), .Q (signal_6760) ) ;
    buf_clk cell_4918 ( .C (clk), .D (signal_681), .Q (signal_6768) ) ;
    buf_clk cell_4926 ( .C (clk), .D (signal_3358), .Q (signal_6776) ) ;
    buf_clk cell_4934 ( .C (clk), .D (signal_683), .Q (signal_6784) ) ;
    buf_clk cell_4942 ( .C (clk), .D (signal_3359), .Q (signal_6792) ) ;
    buf_clk cell_4950 ( .C (clk), .D (signal_685), .Q (signal_6800) ) ;
    buf_clk cell_4958 ( .C (clk), .D (signal_3360), .Q (signal_6808) ) ;
    buf_clk cell_4966 ( .C (clk), .D (signal_687), .Q (signal_6816) ) ;
    buf_clk cell_4974 ( .C (clk), .D (signal_3361), .Q (signal_6824) ) ;
    buf_clk cell_4982 ( .C (clk), .D (signal_689), .Q (signal_6832) ) ;
    buf_clk cell_4990 ( .C (clk), .D (signal_3362), .Q (signal_6840) ) ;
    buf_clk cell_4998 ( .C (clk), .D (signal_691), .Q (signal_6848) ) ;
    buf_clk cell_5006 ( .C (clk), .D (signal_3363), .Q (signal_6856) ) ;
    buf_clk cell_5014 ( .C (clk), .D (signal_693), .Q (signal_6864) ) ;
    buf_clk cell_5022 ( .C (clk), .D (signal_3364), .Q (signal_6872) ) ;
    buf_clk cell_5030 ( .C (clk), .D (signal_695), .Q (signal_6880) ) ;
    buf_clk cell_5038 ( .C (clk), .D (signal_3365), .Q (signal_6888) ) ;
    buf_clk cell_5046 ( .C (clk), .D (signal_697), .Q (signal_6896) ) ;
    buf_clk cell_5054 ( .C (clk), .D (signal_3366), .Q (signal_6904) ) ;
    buf_clk cell_5062 ( .C (clk), .D (signal_699), .Q (signal_6912) ) ;
    buf_clk cell_5070 ( .C (clk), .D (signal_3367), .Q (signal_6920) ) ;
    buf_clk cell_5078 ( .C (clk), .D (signal_701), .Q (signal_6928) ) ;
    buf_clk cell_5086 ( .C (clk), .D (signal_3368), .Q (signal_6936) ) ;
    buf_clk cell_5094 ( .C (clk), .D (signal_703), .Q (signal_6944) ) ;
    buf_clk cell_5102 ( .C (clk), .D (signal_3369), .Q (signal_6952) ) ;
    buf_clk cell_5110 ( .C (clk), .D (signal_766), .Q (signal_6960) ) ;
    buf_clk cell_5118 ( .C (clk), .D (signal_3499), .Q (signal_6968) ) ;
    buf_clk cell_5126 ( .C (clk), .D (signal_769), .Q (signal_6976) ) ;
    buf_clk cell_5134 ( .C (clk), .D (signal_3500), .Q (signal_6984) ) ;
    buf_clk cell_5142 ( .C (clk), .D (signal_772), .Q (signal_6992) ) ;
    buf_clk cell_5150 ( .C (clk), .D (signal_3501), .Q (signal_7000) ) ;
    buf_clk cell_5158 ( .C (clk), .D (signal_775), .Q (signal_7008) ) ;
    buf_clk cell_5166 ( .C (clk), .D (signal_3502), .Q (signal_7016) ) ;
    buf_clk cell_5174 ( .C (clk), .D (signal_778), .Q (signal_7024) ) ;
    buf_clk cell_5182 ( .C (clk), .D (signal_3503), .Q (signal_7032) ) ;
    buf_clk cell_5190 ( .C (clk), .D (signal_781), .Q (signal_7040) ) ;
    buf_clk cell_5198 ( .C (clk), .D (signal_3504), .Q (signal_7048) ) ;
    buf_clk cell_5206 ( .C (clk), .D (signal_784), .Q (signal_7056) ) ;
    buf_clk cell_5214 ( .C (clk), .D (signal_3505), .Q (signal_7064) ) ;
    buf_clk cell_5222 ( .C (clk), .D (signal_787), .Q (signal_7072) ) ;
    buf_clk cell_5230 ( .C (clk), .D (signal_3506), .Q (signal_7080) ) ;
    buf_clk cell_5238 ( .C (clk), .D (signal_790), .Q (signal_7088) ) ;
    buf_clk cell_5246 ( .C (clk), .D (signal_3399), .Q (signal_7096) ) ;
    buf_clk cell_5254 ( .C (clk), .D (signal_793), .Q (signal_7104) ) ;
    buf_clk cell_5262 ( .C (clk), .D (signal_3400), .Q (signal_7112) ) ;
    buf_clk cell_5270 ( .C (clk), .D (signal_796), .Q (signal_7120) ) ;
    buf_clk cell_5278 ( .C (clk), .D (signal_3401), .Q (signal_7128) ) ;
    buf_clk cell_5286 ( .C (clk), .D (signal_799), .Q (signal_7136) ) ;
    buf_clk cell_5294 ( .C (clk), .D (signal_3402), .Q (signal_7144) ) ;
    buf_clk cell_5302 ( .C (clk), .D (signal_802), .Q (signal_7152) ) ;
    buf_clk cell_5310 ( .C (clk), .D (signal_3403), .Q (signal_7160) ) ;
    buf_clk cell_5318 ( .C (clk), .D (signal_805), .Q (signal_7168) ) ;
    buf_clk cell_5326 ( .C (clk), .D (signal_3404), .Q (signal_7176) ) ;
    buf_clk cell_5334 ( .C (clk), .D (signal_808), .Q (signal_7184) ) ;
    buf_clk cell_5342 ( .C (clk), .D (signal_3405), .Q (signal_7192) ) ;
    buf_clk cell_5350 ( .C (clk), .D (signal_811), .Q (signal_7200) ) ;
    buf_clk cell_5358 ( .C (clk), .D (signal_3406), .Q (signal_7208) ) ;
    buf_clk cell_5366 ( .C (clk), .D (signal_814), .Q (signal_7216) ) ;
    buf_clk cell_5374 ( .C (clk), .D (signal_3407), .Q (signal_7224) ) ;
    buf_clk cell_5382 ( .C (clk), .D (signal_817), .Q (signal_7232) ) ;
    buf_clk cell_5390 ( .C (clk), .D (signal_3408), .Q (signal_7240) ) ;
    buf_clk cell_5398 ( .C (clk), .D (signal_820), .Q (signal_7248) ) ;
    buf_clk cell_5406 ( .C (clk), .D (signal_3409), .Q (signal_7256) ) ;
    buf_clk cell_5414 ( .C (clk), .D (signal_823), .Q (signal_7264) ) ;
    buf_clk cell_5422 ( .C (clk), .D (signal_3410), .Q (signal_7272) ) ;
    buf_clk cell_5430 ( .C (clk), .D (signal_826), .Q (signal_7280) ) ;
    buf_clk cell_5438 ( .C (clk), .D (signal_3411), .Q (signal_7288) ) ;
    buf_clk cell_5446 ( .C (clk), .D (signal_829), .Q (signal_7296) ) ;
    buf_clk cell_5454 ( .C (clk), .D (signal_3412), .Q (signal_7304) ) ;
    buf_clk cell_5462 ( .C (clk), .D (signal_832), .Q (signal_7312) ) ;
    buf_clk cell_5470 ( .C (clk), .D (signal_3413), .Q (signal_7320) ) ;
    buf_clk cell_5478 ( .C (clk), .D (signal_835), .Q (signal_7328) ) ;
    buf_clk cell_5486 ( .C (clk), .D (signal_3414), .Q (signal_7336) ) ;
    buf_clk cell_5494 ( .C (clk), .D (signal_838), .Q (signal_7344) ) ;
    buf_clk cell_5502 ( .C (clk), .D (signal_3415), .Q (signal_7352) ) ;
    buf_clk cell_5510 ( .C (clk), .D (signal_841), .Q (signal_7360) ) ;
    buf_clk cell_5518 ( .C (clk), .D (signal_3416), .Q (signal_7368) ) ;
    buf_clk cell_5526 ( .C (clk), .D (signal_844), .Q (signal_7376) ) ;
    buf_clk cell_5534 ( .C (clk), .D (signal_3417), .Q (signal_7384) ) ;
    buf_clk cell_5542 ( .C (clk), .D (signal_847), .Q (signal_7392) ) ;
    buf_clk cell_5550 ( .C (clk), .D (signal_3418), .Q (signal_7400) ) ;
    buf_clk cell_5558 ( .C (clk), .D (signal_850), .Q (signal_7408) ) ;
    buf_clk cell_5566 ( .C (clk), .D (signal_3419), .Q (signal_7416) ) ;
    buf_clk cell_5574 ( .C (clk), .D (signal_853), .Q (signal_7424) ) ;
    buf_clk cell_5582 ( .C (clk), .D (signal_3420), .Q (signal_7432) ) ;
    buf_clk cell_5590 ( .C (clk), .D (signal_856), .Q (signal_7440) ) ;
    buf_clk cell_5598 ( .C (clk), .D (signal_3421), .Q (signal_7448) ) ;
    buf_clk cell_5606 ( .C (clk), .D (signal_859), .Q (signal_7456) ) ;
    buf_clk cell_5614 ( .C (clk), .D (signal_3422), .Q (signal_7464) ) ;
    buf_clk cell_5622 ( .C (clk), .D (signal_862), .Q (signal_7472) ) ;
    buf_clk cell_5630 ( .C (clk), .D (signal_3423), .Q (signal_7480) ) ;
    buf_clk cell_5638 ( .C (clk), .D (signal_865), .Q (signal_7488) ) ;
    buf_clk cell_5646 ( .C (clk), .D (signal_3424), .Q (signal_7496) ) ;
    buf_clk cell_5654 ( .C (clk), .D (signal_868), .Q (signal_7504) ) ;
    buf_clk cell_5662 ( .C (clk), .D (signal_3425), .Q (signal_7512) ) ;
    buf_clk cell_5670 ( .C (clk), .D (signal_871), .Q (signal_7520) ) ;
    buf_clk cell_5678 ( .C (clk), .D (signal_3426), .Q (signal_7528) ) ;
    buf_clk cell_5686 ( .C (clk), .D (signal_874), .Q (signal_7536) ) ;
    buf_clk cell_5694 ( .C (clk), .D (signal_3427), .Q (signal_7544) ) ;
    buf_clk cell_5702 ( .C (clk), .D (signal_877), .Q (signal_7552) ) ;
    buf_clk cell_5710 ( .C (clk), .D (signal_3428), .Q (signal_7560) ) ;
    buf_clk cell_5718 ( .C (clk), .D (signal_880), .Q (signal_7568) ) ;
    buf_clk cell_5726 ( .C (clk), .D (signal_3429), .Q (signal_7576) ) ;
    buf_clk cell_5734 ( .C (clk), .D (signal_883), .Q (signal_7584) ) ;
    buf_clk cell_5742 ( .C (clk), .D (signal_3430), .Q (signal_7592) ) ;
    buf_clk cell_5750 ( .C (clk), .D (signal_886), .Q (signal_7600) ) ;
    buf_clk cell_5758 ( .C (clk), .D (signal_3431), .Q (signal_7608) ) ;
    buf_clk cell_5766 ( .C (clk), .D (signal_889), .Q (signal_7616) ) ;
    buf_clk cell_5774 ( .C (clk), .D (signal_3432), .Q (signal_7624) ) ;
    buf_clk cell_5782 ( .C (clk), .D (signal_892), .Q (signal_7632) ) ;
    buf_clk cell_5790 ( .C (clk), .D (signal_3433), .Q (signal_7640) ) ;
    buf_clk cell_5798 ( .C (clk), .D (signal_895), .Q (signal_7648) ) ;
    buf_clk cell_5806 ( .C (clk), .D (signal_3434), .Q (signal_7656) ) ;
    buf_clk cell_5814 ( .C (clk), .D (signal_898), .Q (signal_7664) ) ;
    buf_clk cell_5822 ( .C (clk), .D (signal_3435), .Q (signal_7672) ) ;
    buf_clk cell_5830 ( .C (clk), .D (signal_901), .Q (signal_7680) ) ;
    buf_clk cell_5838 ( .C (clk), .D (signal_3436), .Q (signal_7688) ) ;
    buf_clk cell_5846 ( .C (clk), .D (signal_904), .Q (signal_7696) ) ;
    buf_clk cell_5854 ( .C (clk), .D (signal_3437), .Q (signal_7704) ) ;
    buf_clk cell_5862 ( .C (clk), .D (signal_907), .Q (signal_7712) ) ;
    buf_clk cell_5870 ( .C (clk), .D (signal_3438), .Q (signal_7720) ) ;
    buf_clk cell_5878 ( .C (clk), .D (signal_910), .Q (signal_7728) ) ;
    buf_clk cell_5886 ( .C (clk), .D (signal_3217), .Q (signal_7736) ) ;
    buf_clk cell_5894 ( .C (clk), .D (signal_913), .Q (signal_7744) ) ;
    buf_clk cell_5902 ( .C (clk), .D (signal_3218), .Q (signal_7752) ) ;
    buf_clk cell_5910 ( .C (clk), .D (signal_916), .Q (signal_7760) ) ;
    buf_clk cell_5918 ( .C (clk), .D (signal_3219), .Q (signal_7768) ) ;
    buf_clk cell_5926 ( .C (clk), .D (signal_919), .Q (signal_7776) ) ;
    buf_clk cell_5934 ( .C (clk), .D (signal_3220), .Q (signal_7784) ) ;
    buf_clk cell_5942 ( .C (clk), .D (signal_922), .Q (signal_7792) ) ;
    buf_clk cell_5950 ( .C (clk), .D (signal_3221), .Q (signal_7800) ) ;
    buf_clk cell_5958 ( .C (clk), .D (signal_925), .Q (signal_7808) ) ;
    buf_clk cell_5966 ( .C (clk), .D (signal_3222), .Q (signal_7816) ) ;
    buf_clk cell_5974 ( .C (clk), .D (signal_928), .Q (signal_7824) ) ;
    buf_clk cell_5982 ( .C (clk), .D (signal_3223), .Q (signal_7832) ) ;
    buf_clk cell_5990 ( .C (clk), .D (signal_931), .Q (signal_7840) ) ;
    buf_clk cell_5998 ( .C (clk), .D (signal_3224), .Q (signal_7848) ) ;
    buf_clk cell_6006 ( .C (clk), .D (signal_934), .Q (signal_7856) ) ;
    buf_clk cell_6014 ( .C (clk), .D (signal_3225), .Q (signal_7864) ) ;
    buf_clk cell_6022 ( .C (clk), .D (signal_937), .Q (signal_7872) ) ;
    buf_clk cell_6030 ( .C (clk), .D (signal_3226), .Q (signal_7880) ) ;
    buf_clk cell_6038 ( .C (clk), .D (signal_940), .Q (signal_7888) ) ;
    buf_clk cell_6046 ( .C (clk), .D (signal_3227), .Q (signal_7896) ) ;
    buf_clk cell_6054 ( .C (clk), .D (signal_943), .Q (signal_7904) ) ;
    buf_clk cell_6062 ( .C (clk), .D (signal_3228), .Q (signal_7912) ) ;
    buf_clk cell_6070 ( .C (clk), .D (signal_946), .Q (signal_7920) ) ;
    buf_clk cell_6078 ( .C (clk), .D (signal_3229), .Q (signal_7928) ) ;
    buf_clk cell_6086 ( .C (clk), .D (signal_949), .Q (signal_7936) ) ;
    buf_clk cell_6094 ( .C (clk), .D (signal_3230), .Q (signal_7944) ) ;
    buf_clk cell_6102 ( .C (clk), .D (signal_952), .Q (signal_7952) ) ;
    buf_clk cell_6110 ( .C (clk), .D (signal_3231), .Q (signal_7960) ) ;
    buf_clk cell_6118 ( .C (clk), .D (signal_955), .Q (signal_7968) ) ;
    buf_clk cell_6126 ( .C (clk), .D (signal_3232), .Q (signal_7976) ) ;
    buf_clk cell_6134 ( .C (clk), .D (signal_958), .Q (signal_7984) ) ;
    buf_clk cell_6142 ( .C (clk), .D (signal_3439), .Q (signal_7992) ) ;
    buf_clk cell_6150 ( .C (clk), .D (signal_961), .Q (signal_8000) ) ;
    buf_clk cell_6158 ( .C (clk), .D (signal_3440), .Q (signal_8008) ) ;
    buf_clk cell_6166 ( .C (clk), .D (signal_964), .Q (signal_8016) ) ;
    buf_clk cell_6174 ( .C (clk), .D (signal_3441), .Q (signal_8024) ) ;
    buf_clk cell_6182 ( .C (clk), .D (signal_967), .Q (signal_8032) ) ;
    buf_clk cell_6190 ( .C (clk), .D (signal_3442), .Q (signal_8040) ) ;
    buf_clk cell_6198 ( .C (clk), .D (signal_970), .Q (signal_8048) ) ;
    buf_clk cell_6206 ( .C (clk), .D (signal_3443), .Q (signal_8056) ) ;
    buf_clk cell_6214 ( .C (clk), .D (signal_973), .Q (signal_8064) ) ;
    buf_clk cell_6222 ( .C (clk), .D (signal_3444), .Q (signal_8072) ) ;
    buf_clk cell_6230 ( .C (clk), .D (signal_976), .Q (signal_8080) ) ;
    buf_clk cell_6238 ( .C (clk), .D (signal_3445), .Q (signal_8088) ) ;
    buf_clk cell_6246 ( .C (clk), .D (signal_979), .Q (signal_8096) ) ;
    buf_clk cell_6254 ( .C (clk), .D (signal_3446), .Q (signal_8104) ) ;
    buf_clk cell_6262 ( .C (clk), .D (signal_982), .Q (signal_8112) ) ;
    buf_clk cell_6270 ( .C (clk), .D (signal_3447), .Q (signal_8120) ) ;
    buf_clk cell_6278 ( .C (clk), .D (signal_985), .Q (signal_8128) ) ;
    buf_clk cell_6286 ( .C (clk), .D (signal_3448), .Q (signal_8136) ) ;
    buf_clk cell_6294 ( .C (clk), .D (signal_988), .Q (signal_8144) ) ;
    buf_clk cell_6302 ( .C (clk), .D (signal_3449), .Q (signal_8152) ) ;
    buf_clk cell_6310 ( .C (clk), .D (signal_991), .Q (signal_8160) ) ;
    buf_clk cell_6318 ( .C (clk), .D (signal_3450), .Q (signal_8168) ) ;
    buf_clk cell_6326 ( .C (clk), .D (signal_994), .Q (signal_8176) ) ;
    buf_clk cell_6334 ( .C (clk), .D (signal_3451), .Q (signal_8184) ) ;
    buf_clk cell_6342 ( .C (clk), .D (signal_997), .Q (signal_8192) ) ;
    buf_clk cell_6350 ( .C (clk), .D (signal_3452), .Q (signal_8200) ) ;
    buf_clk cell_6358 ( .C (clk), .D (signal_1000), .Q (signal_8208) ) ;
    buf_clk cell_6366 ( .C (clk), .D (signal_3453), .Q (signal_8216) ) ;
    buf_clk cell_6374 ( .C (clk), .D (signal_1003), .Q (signal_8224) ) ;
    buf_clk cell_6382 ( .C (clk), .D (signal_3454), .Q (signal_8232) ) ;
    buf_clk cell_6390 ( .C (clk), .D (signal_1006), .Q (signal_8240) ) ;
    buf_clk cell_6398 ( .C (clk), .D (signal_3455), .Q (signal_8248) ) ;
    buf_clk cell_6406 ( .C (clk), .D (signal_1009), .Q (signal_8256) ) ;
    buf_clk cell_6414 ( .C (clk), .D (signal_3456), .Q (signal_8264) ) ;
    buf_clk cell_6422 ( .C (clk), .D (signal_1012), .Q (signal_8272) ) ;
    buf_clk cell_6430 ( .C (clk), .D (signal_3457), .Q (signal_8280) ) ;
    buf_clk cell_6438 ( .C (clk), .D (signal_1015), .Q (signal_8288) ) ;
    buf_clk cell_6446 ( .C (clk), .D (signal_3458), .Q (signal_8296) ) ;
    buf_clk cell_6454 ( .C (clk), .D (signal_1018), .Q (signal_8304) ) ;
    buf_clk cell_6462 ( .C (clk), .D (signal_3459), .Q (signal_8312) ) ;
    buf_clk cell_6470 ( .C (clk), .D (signal_1021), .Q (signal_8320) ) ;
    buf_clk cell_6478 ( .C (clk), .D (signal_3460), .Q (signal_8328) ) ;
    buf_clk cell_6486 ( .C (clk), .D (signal_1024), .Q (signal_8336) ) ;
    buf_clk cell_6494 ( .C (clk), .D (signal_3461), .Q (signal_8344) ) ;
    buf_clk cell_6502 ( .C (clk), .D (signal_1027), .Q (signal_8352) ) ;
    buf_clk cell_6510 ( .C (clk), .D (signal_3462), .Q (signal_8360) ) ;
    buf_clk cell_6518 ( .C (clk), .D (signal_1030), .Q (signal_8368) ) ;
    buf_clk cell_6526 ( .C (clk), .D (signal_3463), .Q (signal_8376) ) ;
    buf_clk cell_6534 ( .C (clk), .D (signal_1033), .Q (signal_8384) ) ;
    buf_clk cell_6542 ( .C (clk), .D (signal_3464), .Q (signal_8392) ) ;
    buf_clk cell_6550 ( .C (clk), .D (signal_1036), .Q (signal_8400) ) ;
    buf_clk cell_6558 ( .C (clk), .D (signal_3465), .Q (signal_8408) ) ;
    buf_clk cell_6566 ( .C (clk), .D (signal_1039), .Q (signal_8416) ) ;
    buf_clk cell_6574 ( .C (clk), .D (signal_3466), .Q (signal_8424) ) ;
    buf_clk cell_6582 ( .C (clk), .D (signal_1042), .Q (signal_8432) ) ;
    buf_clk cell_6590 ( .C (clk), .D (signal_3467), .Q (signal_8440) ) ;
    buf_clk cell_6598 ( .C (clk), .D (signal_1045), .Q (signal_8448) ) ;
    buf_clk cell_6606 ( .C (clk), .D (signal_3468), .Q (signal_8456) ) ;
    buf_clk cell_6614 ( .C (clk), .D (signal_1048), .Q (signal_8464) ) ;
    buf_clk cell_6622 ( .C (clk), .D (signal_3469), .Q (signal_8472) ) ;
    buf_clk cell_6630 ( .C (clk), .D (signal_1051), .Q (signal_8480) ) ;
    buf_clk cell_6638 ( .C (clk), .D (signal_3470), .Q (signal_8488) ) ;
    buf_clk cell_6646 ( .C (clk), .D (signal_1078), .Q (signal_8496) ) ;
    buf_clk cell_6654 ( .C (clk), .D (signal_3471), .Q (signal_8504) ) ;
    buf_clk cell_6662 ( .C (clk), .D (signal_1081), .Q (signal_8512) ) ;
    buf_clk cell_6670 ( .C (clk), .D (signal_3472), .Q (signal_8520) ) ;
    buf_clk cell_6678 ( .C (clk), .D (signal_1084), .Q (signal_8528) ) ;
    buf_clk cell_6686 ( .C (clk), .D (signal_3473), .Q (signal_8536) ) ;
    buf_clk cell_6694 ( .C (clk), .D (signal_1087), .Q (signal_8544) ) ;
    buf_clk cell_6702 ( .C (clk), .D (signal_3474), .Q (signal_8552) ) ;
    buf_clk cell_6710 ( .C (clk), .D (signal_1090), .Q (signal_8560) ) ;
    buf_clk cell_6718 ( .C (clk), .D (signal_3475), .Q (signal_8568) ) ;
    buf_clk cell_6726 ( .C (clk), .D (signal_1093), .Q (signal_8576) ) ;
    buf_clk cell_6734 ( .C (clk), .D (signal_3476), .Q (signal_8584) ) ;
    buf_clk cell_6742 ( .C (clk), .D (signal_1096), .Q (signal_8592) ) ;
    buf_clk cell_6750 ( .C (clk), .D (signal_3477), .Q (signal_8600) ) ;
    buf_clk cell_6758 ( .C (clk), .D (signal_1099), .Q (signal_8608) ) ;
    buf_clk cell_6766 ( .C (clk), .D (signal_3478), .Q (signal_8616) ) ;
    buf_clk cell_6774 ( .C (clk), .D (signal_1102), .Q (signal_8624) ) ;
    buf_clk cell_6782 ( .C (clk), .D (signal_3479), .Q (signal_8632) ) ;
    buf_clk cell_6790 ( .C (clk), .D (signal_1105), .Q (signal_8640) ) ;
    buf_clk cell_6798 ( .C (clk), .D (signal_3480), .Q (signal_8648) ) ;
    buf_clk cell_6806 ( .C (clk), .D (signal_1108), .Q (signal_8656) ) ;
    buf_clk cell_6814 ( .C (clk), .D (signal_3481), .Q (signal_8664) ) ;
    buf_clk cell_6822 ( .C (clk), .D (signal_1111), .Q (signal_8672) ) ;
    buf_clk cell_6830 ( .C (clk), .D (signal_3482), .Q (signal_8680) ) ;
    buf_clk cell_6838 ( .C (clk), .D (signal_1114), .Q (signal_8688) ) ;
    buf_clk cell_6846 ( .C (clk), .D (signal_3483), .Q (signal_8696) ) ;
    buf_clk cell_6854 ( .C (clk), .D (signal_1117), .Q (signal_8704) ) ;
    buf_clk cell_6862 ( .C (clk), .D (signal_3484), .Q (signal_8712) ) ;
    buf_clk cell_6870 ( .C (clk), .D (signal_1120), .Q (signal_8720) ) ;
    buf_clk cell_6878 ( .C (clk), .D (signal_3485), .Q (signal_8728) ) ;
    buf_clk cell_6886 ( .C (clk), .D (signal_1123), .Q (signal_8736) ) ;
    buf_clk cell_6894 ( .C (clk), .D (signal_3486), .Q (signal_8744) ) ;
    buf_clk cell_6902 ( .C (clk), .D (signal_1126), .Q (signal_8752) ) ;
    buf_clk cell_6910 ( .C (clk), .D (signal_3487), .Q (signal_8760) ) ;
    buf_clk cell_6918 ( .C (clk), .D (signal_1129), .Q (signal_8768) ) ;
    buf_clk cell_6926 ( .C (clk), .D (signal_3488), .Q (signal_8776) ) ;
    buf_clk cell_6934 ( .C (clk), .D (signal_1132), .Q (signal_8784) ) ;
    buf_clk cell_6942 ( .C (clk), .D (signal_3489), .Q (signal_8792) ) ;
    buf_clk cell_6950 ( .C (clk), .D (signal_1135), .Q (signal_8800) ) ;
    buf_clk cell_6958 ( .C (clk), .D (signal_3490), .Q (signal_8808) ) ;
    buf_clk cell_6966 ( .C (clk), .D (signal_1138), .Q (signal_8816) ) ;
    buf_clk cell_6974 ( .C (clk), .D (signal_3491), .Q (signal_8824) ) ;
    buf_clk cell_6982 ( .C (clk), .D (signal_1141), .Q (signal_8832) ) ;
    buf_clk cell_6990 ( .C (clk), .D (signal_3492), .Q (signal_8840) ) ;
    buf_clk cell_6998 ( .C (clk), .D (signal_1144), .Q (signal_8848) ) ;
    buf_clk cell_7006 ( .C (clk), .D (signal_3493), .Q (signal_8856) ) ;
    buf_clk cell_7014 ( .C (clk), .D (signal_1147), .Q (signal_8864) ) ;
    buf_clk cell_7022 ( .C (clk), .D (signal_3494), .Q (signal_8872) ) ;
    buf_clk cell_7030 ( .C (clk), .D (signal_1275), .Q (signal_8880) ) ;
    buf_clk cell_7038 ( .C (clk), .D (signal_1266), .Q (signal_8888) ) ;
    buf_clk cell_7046 ( .C (clk), .D (signal_1264), .Q (signal_8896) ) ;
    buf_clk cell_7054 ( .C (clk), .D (signal_1262), .Q (signal_8904) ) ;
    buf_clk cell_7062 ( .C (clk), .D (signal_1260), .Q (signal_8912) ) ;
    buf_clk cell_7070 ( .C (clk), .D (signal_1259), .Q (signal_8920) ) ;
    buf_clk cell_7078 ( .C (clk), .D (signal_1258), .Q (signal_8928) ) ;
    buf_clk cell_7086 ( .C (clk), .D (signal_1256), .Q (signal_8936) ) ;
    buf_clk cell_7094 ( .C (clk), .D (signal_403), .Q (signal_8944) ) ;

    /* cells in depth 2 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1732 ( .a ({signal_3124, signal_1992}), .b ({signal_3126, signal_1994}), .clk (clk), .r (Fresh[0]), .c ({signal_3156, signal_2000}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1733 ( .a ({signal_2950, signal_1517}), .b ({signal_3129, signal_1997}), .clk (clk), .r (Fresh[1]), .c ({signal_3157, signal_2001}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1734 ( .a ({signal_2976, signal_1984}), .b ({signal_3128, signal_1996}), .clk (clk), .r (Fresh[2]), .c ({signal_3158, signal_2002}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1735 ( .a ({signal_3125, signal_1993}), .b ({signal_3130, signal_1998}), .clk (clk), .r (Fresh[3]), .c ({signal_3159, signal_2003}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1736 ( .a ({signal_2974, signal_1982}), .b ({signal_3127, signal_1995}), .clk (clk), .r (Fresh[4]), .c ({signal_3160, signal_2004}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1737 ( .a ({signal_2977, signal_1985}), .b ({signal_3131, signal_1999}), .clk (clk), .r (Fresh[5]), .c ({signal_3161, signal_2005}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1745 ( .a ({signal_3162, signal_2006}), .b ({signal_3167, signal_2011}), .clk (clk), .r (Fresh[6]), .c ({signal_3241, signal_2013}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1746 ( .a ({signal_3165, signal_2009}), .b ({signal_3166, signal_2010}), .clk (clk), .r (Fresh[7]), .c ({signal_3242, signal_2014}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1747 ( .a ({signal_2975, signal_1983}), .b ({signal_3163, signal_2007}), .clk (clk), .r (Fresh[8]), .c ({signal_3243, signal_2015}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1750 ( .a ({signal_3699, signal_3697}), .b ({signal_3156, signal_2000}), .c ({signal_3246, signal_2018}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1751 ( .a ({signal_3156, signal_2000}), .b ({signal_3157, signal_2001}), .c ({signal_3247, signal_2019}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1752 ( .a ({signal_3703, signal_3701}), .b ({signal_3158, signal_2002}), .c ({signal_3248, signal_2020}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1753 ( .a ({signal_3160, signal_2004}), .b ({signal_3161, signal_2005}), .c ({signal_3249, signal_2021}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1754 ( .a ({signal_3158, signal_2002}), .b ({signal_3242, signal_2014}), .c ({signal_3386, signal_2022}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1755 ( .a ({signal_3160, signal_2004}), .b ({signal_3243, signal_2015}), .c ({signal_3387, signal_2023}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1756 ( .a ({signal_3241, signal_2013}), .b ({signal_3246, signal_2018}), .c ({signal_3388, signal_2024}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1757 ( .a ({signal_3707, signal_3705}), .b ({signal_3247, signal_2019}), .c ({signal_3389, signal_2025}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1758 ( .a ({signal_3159, signal_2003}), .b ({signal_3248, signal_2020}), .c ({signal_3390, signal_2026}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1759 ( .a ({signal_3386, signal_2022}), .b ({signal_3387, signal_2023}), .c ({signal_3495, signal_2027}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1760 ( .a ({signal_3249, signal_2021}), .b ({signal_3388, signal_2024}), .c ({signal_3496, signal_2028}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1761 ( .a ({signal_3387, signal_2023}), .b ({signal_3389, signal_2025}), .c ({signal_3497, signal_2029}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1762 ( .a ({signal_3249, signal_2021}), .b ({signal_3390, signal_2026}), .c ({signal_3498, signal_2030}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1765 ( .a ({signal_3711, signal_3709}), .b ({signal_3495, signal_2027}), .c ({signal_3509, signal_2033}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1766 ( .a ({signal_3496, signal_2028}), .b ({signal_3497, signal_2029}), .c ({signal_3510, signal_2034}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1768 ( .a ({signal_3498, signal_2030}), .b ({signal_3509, signal_2033}), .c ({signal_3512, signal_2036}) ) ;
    buf_clk cell_1847 ( .C (clk), .D (signal_3696), .Q (signal_3697) ) ;
    buf_clk cell_1849 ( .C (clk), .D (signal_3698), .Q (signal_3699) ) ;
    buf_clk cell_1851 ( .C (clk), .D (signal_3700), .Q (signal_3701) ) ;
    buf_clk cell_1853 ( .C (clk), .D (signal_3702), .Q (signal_3703) ) ;
    buf_clk cell_1855 ( .C (clk), .D (signal_3704), .Q (signal_3705) ) ;
    buf_clk cell_1857 ( .C (clk), .D (signal_3706), .Q (signal_3707) ) ;
    buf_clk cell_1859 ( .C (clk), .D (signal_3708), .Q (signal_3709) ) ;
    buf_clk cell_1861 ( .C (clk), .D (signal_3710), .Q (signal_3711) ) ;
    buf_clk cell_1895 ( .C (clk), .D (signal_3744), .Q (signal_3745) ) ;
    buf_clk cell_1903 ( .C (clk), .D (signal_3752), .Q (signal_3753) ) ;
    buf_clk cell_1911 ( .C (clk), .D (signal_3760), .Q (signal_3761) ) ;
    buf_clk cell_1919 ( .C (clk), .D (signal_3768), .Q (signal_3769) ) ;
    buf_clk cell_1927 ( .C (clk), .D (signal_3776), .Q (signal_3777) ) ;
    buf_clk cell_1935 ( .C (clk), .D (signal_3784), .Q (signal_3785) ) ;
    buf_clk cell_1943 ( .C (clk), .D (signal_3792), .Q (signal_3793) ) ;
    buf_clk cell_1951 ( .C (clk), .D (signal_3800), .Q (signal_3801) ) ;
    buf_clk cell_1959 ( .C (clk), .D (signal_3808), .Q (signal_3809) ) ;
    buf_clk cell_1967 ( .C (clk), .D (signal_3816), .Q (signal_3817) ) ;
    buf_clk cell_1975 ( .C (clk), .D (signal_3824), .Q (signal_3825) ) ;
    buf_clk cell_1983 ( .C (clk), .D (signal_3832), .Q (signal_3833) ) ;
    buf_clk cell_1991 ( .C (clk), .D (signal_3840), .Q (signal_3841) ) ;
    buf_clk cell_1999 ( .C (clk), .D (signal_3848), .Q (signal_3849) ) ;
    buf_clk cell_2007 ( .C (clk), .D (signal_3856), .Q (signal_3857) ) ;
    buf_clk cell_2015 ( .C (clk), .D (signal_3864), .Q (signal_3865) ) ;
    buf_clk cell_2023 ( .C (clk), .D (signal_3872), .Q (signal_3873) ) ;
    buf_clk cell_2031 ( .C (clk), .D (signal_3880), .Q (signal_3881) ) ;
    buf_clk cell_2039 ( .C (clk), .D (signal_3888), .Q (signal_3889) ) ;
    buf_clk cell_2047 ( .C (clk), .D (signal_3896), .Q (signal_3897) ) ;
    buf_clk cell_2055 ( .C (clk), .D (signal_3904), .Q (signal_3905) ) ;
    buf_clk cell_2063 ( .C (clk), .D (signal_3912), .Q (signal_3913) ) ;
    buf_clk cell_2071 ( .C (clk), .D (signal_3920), .Q (signal_3921) ) ;
    buf_clk cell_2079 ( .C (clk), .D (signal_3928), .Q (signal_3929) ) ;
    buf_clk cell_2087 ( .C (clk), .D (signal_3936), .Q (signal_3937) ) ;
    buf_clk cell_2095 ( .C (clk), .D (signal_3944), .Q (signal_3945) ) ;
    buf_clk cell_2103 ( .C (clk), .D (signal_3952), .Q (signal_3953) ) ;
    buf_clk cell_2111 ( .C (clk), .D (signal_3960), .Q (signal_3961) ) ;
    buf_clk cell_2119 ( .C (clk), .D (signal_3968), .Q (signal_3969) ) ;
    buf_clk cell_2127 ( .C (clk), .D (signal_3976), .Q (signal_3977) ) ;
    buf_clk cell_2135 ( .C (clk), .D (signal_3984), .Q (signal_3985) ) ;
    buf_clk cell_2143 ( .C (clk), .D (signal_3992), .Q (signal_3993) ) ;
    buf_clk cell_2151 ( .C (clk), .D (signal_4000), .Q (signal_4001) ) ;
    buf_clk cell_2159 ( .C (clk), .D (signal_4008), .Q (signal_4009) ) ;
    buf_clk cell_2167 ( .C (clk), .D (signal_4016), .Q (signal_4017) ) ;
    buf_clk cell_2175 ( .C (clk), .D (signal_4024), .Q (signal_4025) ) ;
    buf_clk cell_2183 ( .C (clk), .D (signal_4032), .Q (signal_4033) ) ;
    buf_clk cell_2191 ( .C (clk), .D (signal_4040), .Q (signal_4041) ) ;
    buf_clk cell_2199 ( .C (clk), .D (signal_4048), .Q (signal_4049) ) ;
    buf_clk cell_2207 ( .C (clk), .D (signal_4056), .Q (signal_4057) ) ;
    buf_clk cell_2215 ( .C (clk), .D (signal_4064), .Q (signal_4065) ) ;
    buf_clk cell_2223 ( .C (clk), .D (signal_4072), .Q (signal_4073) ) ;
    buf_clk cell_2231 ( .C (clk), .D (signal_4080), .Q (signal_4081) ) ;
    buf_clk cell_2239 ( .C (clk), .D (signal_4088), .Q (signal_4089) ) ;
    buf_clk cell_2247 ( .C (clk), .D (signal_4096), .Q (signal_4097) ) ;
    buf_clk cell_2255 ( .C (clk), .D (signal_4104), .Q (signal_4105) ) ;
    buf_clk cell_2263 ( .C (clk), .D (signal_4112), .Q (signal_4113) ) ;
    buf_clk cell_2271 ( .C (clk), .D (signal_4120), .Q (signal_4121) ) ;
    buf_clk cell_2279 ( .C (clk), .D (signal_4128), .Q (signal_4129) ) ;
    buf_clk cell_2287 ( .C (clk), .D (signal_4136), .Q (signal_4137) ) ;
    buf_clk cell_2295 ( .C (clk), .D (signal_4144), .Q (signal_4145) ) ;
    buf_clk cell_2303 ( .C (clk), .D (signal_4152), .Q (signal_4153) ) ;
    buf_clk cell_2311 ( .C (clk), .D (signal_4160), .Q (signal_4161) ) ;
    buf_clk cell_2319 ( .C (clk), .D (signal_4168), .Q (signal_4169) ) ;
    buf_clk cell_2327 ( .C (clk), .D (signal_4176), .Q (signal_4177) ) ;
    buf_clk cell_2335 ( .C (clk), .D (signal_4184), .Q (signal_4185) ) ;
    buf_clk cell_2343 ( .C (clk), .D (signal_4192), .Q (signal_4193) ) ;
    buf_clk cell_2351 ( .C (clk), .D (signal_4200), .Q (signal_4201) ) ;
    buf_clk cell_2359 ( .C (clk), .D (signal_4208), .Q (signal_4209) ) ;
    buf_clk cell_2367 ( .C (clk), .D (signal_4216), .Q (signal_4217) ) ;
    buf_clk cell_2375 ( .C (clk), .D (signal_4224), .Q (signal_4225) ) ;
    buf_clk cell_2383 ( .C (clk), .D (signal_4232), .Q (signal_4233) ) ;
    buf_clk cell_2391 ( .C (clk), .D (signal_4240), .Q (signal_4241) ) ;
    buf_clk cell_2399 ( .C (clk), .D (signal_4248), .Q (signal_4249) ) ;
    buf_clk cell_2407 ( .C (clk), .D (signal_4256), .Q (signal_4257) ) ;
    buf_clk cell_2415 ( .C (clk), .D (signal_4264), .Q (signal_4265) ) ;
    buf_clk cell_2423 ( .C (clk), .D (signal_4272), .Q (signal_4273) ) ;
    buf_clk cell_2431 ( .C (clk), .D (signal_4280), .Q (signal_4281) ) ;
    buf_clk cell_2439 ( .C (clk), .D (signal_4288), .Q (signal_4289) ) ;
    buf_clk cell_2447 ( .C (clk), .D (signal_4296), .Q (signal_4297) ) ;
    buf_clk cell_2455 ( .C (clk), .D (signal_4304), .Q (signal_4305) ) ;
    buf_clk cell_2463 ( .C (clk), .D (signal_4312), .Q (signal_4313) ) ;
    buf_clk cell_2471 ( .C (clk), .D (signal_4320), .Q (signal_4321) ) ;
    buf_clk cell_2479 ( .C (clk), .D (signal_4328), .Q (signal_4329) ) ;
    buf_clk cell_2487 ( .C (clk), .D (signal_4336), .Q (signal_4337) ) ;
    buf_clk cell_2495 ( .C (clk), .D (signal_4344), .Q (signal_4345) ) ;
    buf_clk cell_2503 ( .C (clk), .D (signal_4352), .Q (signal_4353) ) ;
    buf_clk cell_2511 ( .C (clk), .D (signal_4360), .Q (signal_4361) ) ;
    buf_clk cell_2519 ( .C (clk), .D (signal_4368), .Q (signal_4369) ) ;
    buf_clk cell_2527 ( .C (clk), .D (signal_4376), .Q (signal_4377) ) ;
    buf_clk cell_2535 ( .C (clk), .D (signal_4384), .Q (signal_4385) ) ;
    buf_clk cell_2543 ( .C (clk), .D (signal_4392), .Q (signal_4393) ) ;
    buf_clk cell_2551 ( .C (clk), .D (signal_4400), .Q (signal_4401) ) ;
    buf_clk cell_2559 ( .C (clk), .D (signal_4408), .Q (signal_4409) ) ;
    buf_clk cell_2567 ( .C (clk), .D (signal_4416), .Q (signal_4417) ) ;
    buf_clk cell_2575 ( .C (clk), .D (signal_4424), .Q (signal_4425) ) ;
    buf_clk cell_2583 ( .C (clk), .D (signal_4432), .Q (signal_4433) ) ;
    buf_clk cell_2591 ( .C (clk), .D (signal_4440), .Q (signal_4441) ) ;
    buf_clk cell_2599 ( .C (clk), .D (signal_4448), .Q (signal_4449) ) ;
    buf_clk cell_2607 ( .C (clk), .D (signal_4456), .Q (signal_4457) ) ;
    buf_clk cell_2615 ( .C (clk), .D (signal_4464), .Q (signal_4465) ) ;
    buf_clk cell_2623 ( .C (clk), .D (signal_4472), .Q (signal_4473) ) ;
    buf_clk cell_2631 ( .C (clk), .D (signal_4480), .Q (signal_4481) ) ;
    buf_clk cell_2639 ( .C (clk), .D (signal_4488), .Q (signal_4489) ) ;
    buf_clk cell_2647 ( .C (clk), .D (signal_4496), .Q (signal_4497) ) ;
    buf_clk cell_2655 ( .C (clk), .D (signal_4504), .Q (signal_4505) ) ;
    buf_clk cell_2663 ( .C (clk), .D (signal_4512), .Q (signal_4513) ) ;
    buf_clk cell_2671 ( .C (clk), .D (signal_4520), .Q (signal_4521) ) ;
    buf_clk cell_2679 ( .C (clk), .D (signal_4528), .Q (signal_4529) ) ;
    buf_clk cell_2687 ( .C (clk), .D (signal_4536), .Q (signal_4537) ) ;
    buf_clk cell_2695 ( .C (clk), .D (signal_4544), .Q (signal_4545) ) ;
    buf_clk cell_2703 ( .C (clk), .D (signal_4552), .Q (signal_4553) ) ;
    buf_clk cell_2711 ( .C (clk), .D (signal_4560), .Q (signal_4561) ) ;
    buf_clk cell_2719 ( .C (clk), .D (signal_4568), .Q (signal_4569) ) ;
    buf_clk cell_2727 ( .C (clk), .D (signal_4576), .Q (signal_4577) ) ;
    buf_clk cell_2735 ( .C (clk), .D (signal_4584), .Q (signal_4585) ) ;
    buf_clk cell_2743 ( .C (clk), .D (signal_4592), .Q (signal_4593) ) ;
    buf_clk cell_2751 ( .C (clk), .D (signal_4600), .Q (signal_4601) ) ;
    buf_clk cell_2759 ( .C (clk), .D (signal_4608), .Q (signal_4609) ) ;
    buf_clk cell_2767 ( .C (clk), .D (signal_4616), .Q (signal_4617) ) ;
    buf_clk cell_2775 ( .C (clk), .D (signal_4624), .Q (signal_4625) ) ;
    buf_clk cell_2783 ( .C (clk), .D (signal_4632), .Q (signal_4633) ) ;
    buf_clk cell_2791 ( .C (clk), .D (signal_4640), .Q (signal_4641) ) ;
    buf_clk cell_2799 ( .C (clk), .D (signal_4648), .Q (signal_4649) ) ;
    buf_clk cell_2807 ( .C (clk), .D (signal_4656), .Q (signal_4657) ) ;
    buf_clk cell_2815 ( .C (clk), .D (signal_4664), .Q (signal_4665) ) ;
    buf_clk cell_2823 ( .C (clk), .D (signal_4672), .Q (signal_4673) ) ;
    buf_clk cell_2831 ( .C (clk), .D (signal_4680), .Q (signal_4681) ) ;
    buf_clk cell_2839 ( .C (clk), .D (signal_4688), .Q (signal_4689) ) ;
    buf_clk cell_2847 ( .C (clk), .D (signal_4696), .Q (signal_4697) ) ;
    buf_clk cell_2855 ( .C (clk), .D (signal_4704), .Q (signal_4705) ) ;
    buf_clk cell_2863 ( .C (clk), .D (signal_4712), .Q (signal_4713) ) ;
    buf_clk cell_2871 ( .C (clk), .D (signal_4720), .Q (signal_4721) ) ;
    buf_clk cell_2879 ( .C (clk), .D (signal_4728), .Q (signal_4729) ) ;
    buf_clk cell_2887 ( .C (clk), .D (signal_4736), .Q (signal_4737) ) ;
    buf_clk cell_2895 ( .C (clk), .D (signal_4744), .Q (signal_4745) ) ;
    buf_clk cell_2903 ( .C (clk), .D (signal_4752), .Q (signal_4753) ) ;
    buf_clk cell_2909 ( .C (clk), .D (signal_4758), .Q (signal_4759) ) ;
    buf_clk cell_2915 ( .C (clk), .D (signal_4764), .Q (signal_4765) ) ;
    buf_clk cell_2921 ( .C (clk), .D (signal_4770), .Q (signal_4771) ) ;
    buf_clk cell_2927 ( .C (clk), .D (signal_4776), .Q (signal_4777) ) ;
    buf_clk cell_2933 ( .C (clk), .D (signal_4782), .Q (signal_4783) ) ;
    buf_clk cell_2939 ( .C (clk), .D (signal_4788), .Q (signal_4789) ) ;
    buf_clk cell_2945 ( .C (clk), .D (signal_4794), .Q (signal_4795) ) ;
    buf_clk cell_2951 ( .C (clk), .D (signal_4800), .Q (signal_4801) ) ;
    buf_clk cell_2957 ( .C (clk), .D (signal_4806), .Q (signal_4807) ) ;
    buf_clk cell_2963 ( .C (clk), .D (signal_4812), .Q (signal_4813) ) ;
    buf_clk cell_2969 ( .C (clk), .D (signal_4818), .Q (signal_4819) ) ;
    buf_clk cell_2975 ( .C (clk), .D (signal_4824), .Q (signal_4825) ) ;
    buf_clk cell_2981 ( .C (clk), .D (signal_4830), .Q (signal_4831) ) ;
    buf_clk cell_2987 ( .C (clk), .D (signal_4836), .Q (signal_4837) ) ;
    buf_clk cell_2993 ( .C (clk), .D (signal_4842), .Q (signal_4843) ) ;
    buf_clk cell_2999 ( .C (clk), .D (signal_4848), .Q (signal_4849) ) ;
    buf_clk cell_3005 ( .C (clk), .D (signal_4854), .Q (signal_4855) ) ;
    buf_clk cell_3011 ( .C (clk), .D (signal_4860), .Q (signal_4861) ) ;
    buf_clk cell_3017 ( .C (clk), .D (signal_4866), .Q (signal_4867) ) ;
    buf_clk cell_3023 ( .C (clk), .D (signal_4872), .Q (signal_4873) ) ;
    buf_clk cell_3029 ( .C (clk), .D (signal_4878), .Q (signal_4879) ) ;
    buf_clk cell_3035 ( .C (clk), .D (signal_4884), .Q (signal_4885) ) ;
    buf_clk cell_3041 ( .C (clk), .D (signal_4890), .Q (signal_4891) ) ;
    buf_clk cell_3047 ( .C (clk), .D (signal_4896), .Q (signal_4897) ) ;
    buf_clk cell_3053 ( .C (clk), .D (signal_4902), .Q (signal_4903) ) ;
    buf_clk cell_3059 ( .C (clk), .D (signal_4908), .Q (signal_4909) ) ;
    buf_clk cell_3065 ( .C (clk), .D (signal_4914), .Q (signal_4915) ) ;
    buf_clk cell_3071 ( .C (clk), .D (signal_4920), .Q (signal_4921) ) ;
    buf_clk cell_3077 ( .C (clk), .D (signal_4926), .Q (signal_4927) ) ;
    buf_clk cell_3083 ( .C (clk), .D (signal_4932), .Q (signal_4933) ) ;
    buf_clk cell_3089 ( .C (clk), .D (signal_4938), .Q (signal_4939) ) ;
    buf_clk cell_3095 ( .C (clk), .D (signal_4944), .Q (signal_4945) ) ;
    buf_clk cell_3101 ( .C (clk), .D (signal_4950), .Q (signal_4951) ) ;
    buf_clk cell_3107 ( .C (clk), .D (signal_4956), .Q (signal_4957) ) ;
    buf_clk cell_3113 ( .C (clk), .D (signal_4962), .Q (signal_4963) ) ;
    buf_clk cell_3119 ( .C (clk), .D (signal_4968), .Q (signal_4969) ) ;
    buf_clk cell_3127 ( .C (clk), .D (signal_4976), .Q (signal_4977) ) ;
    buf_clk cell_3135 ( .C (clk), .D (signal_4984), .Q (signal_4985) ) ;
    buf_clk cell_3143 ( .C (clk), .D (signal_4992), .Q (signal_4993) ) ;
    buf_clk cell_3151 ( .C (clk), .D (signal_5000), .Q (signal_5001) ) ;
    buf_clk cell_3159 ( .C (clk), .D (signal_5008), .Q (signal_5009) ) ;
    buf_clk cell_3167 ( .C (clk), .D (signal_5016), .Q (signal_5017) ) ;
    buf_clk cell_3175 ( .C (clk), .D (signal_5024), .Q (signal_5025) ) ;
    buf_clk cell_3183 ( .C (clk), .D (signal_5032), .Q (signal_5033) ) ;
    buf_clk cell_3191 ( .C (clk), .D (signal_5040), .Q (signal_5041) ) ;
    buf_clk cell_3199 ( .C (clk), .D (signal_5048), .Q (signal_5049) ) ;
    buf_clk cell_3207 ( .C (clk), .D (signal_5056), .Q (signal_5057) ) ;
    buf_clk cell_3215 ( .C (clk), .D (signal_5064), .Q (signal_5065) ) ;
    buf_clk cell_3223 ( .C (clk), .D (signal_5072), .Q (signal_5073) ) ;
    buf_clk cell_3231 ( .C (clk), .D (signal_5080), .Q (signal_5081) ) ;
    buf_clk cell_3239 ( .C (clk), .D (signal_5088), .Q (signal_5089) ) ;
    buf_clk cell_3247 ( .C (clk), .D (signal_5096), .Q (signal_5097) ) ;
    buf_clk cell_3255 ( .C (clk), .D (signal_5104), .Q (signal_5105) ) ;
    buf_clk cell_3263 ( .C (clk), .D (signal_5112), .Q (signal_5113) ) ;
    buf_clk cell_3271 ( .C (clk), .D (signal_5120), .Q (signal_5121) ) ;
    buf_clk cell_3279 ( .C (clk), .D (signal_5128), .Q (signal_5129) ) ;
    buf_clk cell_3287 ( .C (clk), .D (signal_5136), .Q (signal_5137) ) ;
    buf_clk cell_3295 ( .C (clk), .D (signal_5144), .Q (signal_5145) ) ;
    buf_clk cell_3303 ( .C (clk), .D (signal_5152), .Q (signal_5153) ) ;
    buf_clk cell_3311 ( .C (clk), .D (signal_5160), .Q (signal_5161) ) ;
    buf_clk cell_3319 ( .C (clk), .D (signal_5168), .Q (signal_5169) ) ;
    buf_clk cell_3327 ( .C (clk), .D (signal_5176), .Q (signal_5177) ) ;
    buf_clk cell_3335 ( .C (clk), .D (signal_5184), .Q (signal_5185) ) ;
    buf_clk cell_3343 ( .C (clk), .D (signal_5192), .Q (signal_5193) ) ;
    buf_clk cell_3351 ( .C (clk), .D (signal_5200), .Q (signal_5201) ) ;
    buf_clk cell_3359 ( .C (clk), .D (signal_5208), .Q (signal_5209) ) ;
    buf_clk cell_3367 ( .C (clk), .D (signal_5216), .Q (signal_5217) ) ;
    buf_clk cell_3375 ( .C (clk), .D (signal_5224), .Q (signal_5225) ) ;
    buf_clk cell_3383 ( .C (clk), .D (signal_5232), .Q (signal_5233) ) ;
    buf_clk cell_3391 ( .C (clk), .D (signal_5240), .Q (signal_5241) ) ;
    buf_clk cell_3399 ( .C (clk), .D (signal_5248), .Q (signal_5249) ) ;
    buf_clk cell_3407 ( .C (clk), .D (signal_5256), .Q (signal_5257) ) ;
    buf_clk cell_3415 ( .C (clk), .D (signal_5264), .Q (signal_5265) ) ;
    buf_clk cell_3423 ( .C (clk), .D (signal_5272), .Q (signal_5273) ) ;
    buf_clk cell_3431 ( .C (clk), .D (signal_5280), .Q (signal_5281) ) ;
    buf_clk cell_3439 ( .C (clk), .D (signal_5288), .Q (signal_5289) ) ;
    buf_clk cell_3447 ( .C (clk), .D (signal_5296), .Q (signal_5297) ) ;
    buf_clk cell_3455 ( .C (clk), .D (signal_5304), .Q (signal_5305) ) ;
    buf_clk cell_3463 ( .C (clk), .D (signal_5312), .Q (signal_5313) ) ;
    buf_clk cell_3471 ( .C (clk), .D (signal_5320), .Q (signal_5321) ) ;
    buf_clk cell_3479 ( .C (clk), .D (signal_5328), .Q (signal_5329) ) ;
    buf_clk cell_3487 ( .C (clk), .D (signal_5336), .Q (signal_5337) ) ;
    buf_clk cell_3495 ( .C (clk), .D (signal_5344), .Q (signal_5345) ) ;
    buf_clk cell_3503 ( .C (clk), .D (signal_5352), .Q (signal_5353) ) ;
    buf_clk cell_3511 ( .C (clk), .D (signal_5360), .Q (signal_5361) ) ;
    buf_clk cell_3519 ( .C (clk), .D (signal_5368), .Q (signal_5369) ) ;
    buf_clk cell_3527 ( .C (clk), .D (signal_5376), .Q (signal_5377) ) ;
    buf_clk cell_3535 ( .C (clk), .D (signal_5384), .Q (signal_5385) ) ;
    buf_clk cell_3543 ( .C (clk), .D (signal_5392), .Q (signal_5393) ) ;
    buf_clk cell_3551 ( .C (clk), .D (signal_5400), .Q (signal_5401) ) ;
    buf_clk cell_3559 ( .C (clk), .D (signal_5408), .Q (signal_5409) ) ;
    buf_clk cell_3567 ( .C (clk), .D (signal_5416), .Q (signal_5417) ) ;
    buf_clk cell_3575 ( .C (clk), .D (signal_5424), .Q (signal_5425) ) ;
    buf_clk cell_3583 ( .C (clk), .D (signal_5432), .Q (signal_5433) ) ;
    buf_clk cell_3591 ( .C (clk), .D (signal_5440), .Q (signal_5441) ) ;
    buf_clk cell_3599 ( .C (clk), .D (signal_5448), .Q (signal_5449) ) ;
    buf_clk cell_3607 ( .C (clk), .D (signal_5456), .Q (signal_5457) ) ;
    buf_clk cell_3615 ( .C (clk), .D (signal_5464), .Q (signal_5465) ) ;
    buf_clk cell_3623 ( .C (clk), .D (signal_5472), .Q (signal_5473) ) ;
    buf_clk cell_3631 ( .C (clk), .D (signal_5480), .Q (signal_5481) ) ;
    buf_clk cell_3639 ( .C (clk), .D (signal_5488), .Q (signal_5489) ) ;
    buf_clk cell_3647 ( .C (clk), .D (signal_5496), .Q (signal_5497) ) ;
    buf_clk cell_3655 ( .C (clk), .D (signal_5504), .Q (signal_5505) ) ;
    buf_clk cell_3663 ( .C (clk), .D (signal_5512), .Q (signal_5513) ) ;
    buf_clk cell_3671 ( .C (clk), .D (signal_5520), .Q (signal_5521) ) ;
    buf_clk cell_3679 ( .C (clk), .D (signal_5528), .Q (signal_5529) ) ;
    buf_clk cell_3687 ( .C (clk), .D (signal_5536), .Q (signal_5537) ) ;
    buf_clk cell_3695 ( .C (clk), .D (signal_5544), .Q (signal_5545) ) ;
    buf_clk cell_3703 ( .C (clk), .D (signal_5552), .Q (signal_5553) ) ;
    buf_clk cell_3711 ( .C (clk), .D (signal_5560), .Q (signal_5561) ) ;
    buf_clk cell_3719 ( .C (clk), .D (signal_5568), .Q (signal_5569) ) ;
    buf_clk cell_3727 ( .C (clk), .D (signal_5576), .Q (signal_5577) ) ;
    buf_clk cell_3735 ( .C (clk), .D (signal_5584), .Q (signal_5585) ) ;
    buf_clk cell_3743 ( .C (clk), .D (signal_5592), .Q (signal_5593) ) ;
    buf_clk cell_3751 ( .C (clk), .D (signal_5600), .Q (signal_5601) ) ;
    buf_clk cell_3759 ( .C (clk), .D (signal_5608), .Q (signal_5609) ) ;
    buf_clk cell_3767 ( .C (clk), .D (signal_5616), .Q (signal_5617) ) ;
    buf_clk cell_3775 ( .C (clk), .D (signal_5624), .Q (signal_5625) ) ;
    buf_clk cell_3783 ( .C (clk), .D (signal_5632), .Q (signal_5633) ) ;
    buf_clk cell_3791 ( .C (clk), .D (signal_5640), .Q (signal_5641) ) ;
    buf_clk cell_3799 ( .C (clk), .D (signal_5648), .Q (signal_5649) ) ;
    buf_clk cell_3807 ( .C (clk), .D (signal_5656), .Q (signal_5657) ) ;
    buf_clk cell_3815 ( .C (clk), .D (signal_5664), .Q (signal_5665) ) ;
    buf_clk cell_3823 ( .C (clk), .D (signal_5672), .Q (signal_5673) ) ;
    buf_clk cell_3831 ( .C (clk), .D (signal_5680), .Q (signal_5681) ) ;
    buf_clk cell_3839 ( .C (clk), .D (signal_5688), .Q (signal_5689) ) ;
    buf_clk cell_3847 ( .C (clk), .D (signal_5696), .Q (signal_5697) ) ;
    buf_clk cell_3855 ( .C (clk), .D (signal_5704), .Q (signal_5705) ) ;
    buf_clk cell_3863 ( .C (clk), .D (signal_5712), .Q (signal_5713) ) ;
    buf_clk cell_3871 ( .C (clk), .D (signal_5720), .Q (signal_5721) ) ;
    buf_clk cell_3879 ( .C (clk), .D (signal_5728), .Q (signal_5729) ) ;
    buf_clk cell_3887 ( .C (clk), .D (signal_5736), .Q (signal_5737) ) ;
    buf_clk cell_3895 ( .C (clk), .D (signal_5744), .Q (signal_5745) ) ;
    buf_clk cell_3903 ( .C (clk), .D (signal_5752), .Q (signal_5753) ) ;
    buf_clk cell_3911 ( .C (clk), .D (signal_5760), .Q (signal_5761) ) ;
    buf_clk cell_3919 ( .C (clk), .D (signal_5768), .Q (signal_5769) ) ;
    buf_clk cell_3927 ( .C (clk), .D (signal_5776), .Q (signal_5777) ) ;
    buf_clk cell_3935 ( .C (clk), .D (signal_5784), .Q (signal_5785) ) ;
    buf_clk cell_3943 ( .C (clk), .D (signal_5792), .Q (signal_5793) ) ;
    buf_clk cell_3951 ( .C (clk), .D (signal_5800), .Q (signal_5801) ) ;
    buf_clk cell_3959 ( .C (clk), .D (signal_5808), .Q (signal_5809) ) ;
    buf_clk cell_3967 ( .C (clk), .D (signal_5816), .Q (signal_5817) ) ;
    buf_clk cell_3975 ( .C (clk), .D (signal_5824), .Q (signal_5825) ) ;
    buf_clk cell_3983 ( .C (clk), .D (signal_5832), .Q (signal_5833) ) ;
    buf_clk cell_3991 ( .C (clk), .D (signal_5840), .Q (signal_5841) ) ;
    buf_clk cell_3999 ( .C (clk), .D (signal_5848), .Q (signal_5849) ) ;
    buf_clk cell_4007 ( .C (clk), .D (signal_5856), .Q (signal_5857) ) ;
    buf_clk cell_4015 ( .C (clk), .D (signal_5864), .Q (signal_5865) ) ;
    buf_clk cell_4023 ( .C (clk), .D (signal_5872), .Q (signal_5873) ) ;
    buf_clk cell_4031 ( .C (clk), .D (signal_5880), .Q (signal_5881) ) ;
    buf_clk cell_4039 ( .C (clk), .D (signal_5888), .Q (signal_5889) ) ;
    buf_clk cell_4047 ( .C (clk), .D (signal_5896), .Q (signal_5897) ) ;
    buf_clk cell_4055 ( .C (clk), .D (signal_5904), .Q (signal_5905) ) ;
    buf_clk cell_4063 ( .C (clk), .D (signal_5912), .Q (signal_5913) ) ;
    buf_clk cell_4071 ( .C (clk), .D (signal_5920), .Q (signal_5921) ) ;
    buf_clk cell_4079 ( .C (clk), .D (signal_5928), .Q (signal_5929) ) ;
    buf_clk cell_4087 ( .C (clk), .D (signal_5936), .Q (signal_5937) ) ;
    buf_clk cell_4095 ( .C (clk), .D (signal_5944), .Q (signal_5945) ) ;
    buf_clk cell_4103 ( .C (clk), .D (signal_5952), .Q (signal_5953) ) ;
    buf_clk cell_4111 ( .C (clk), .D (signal_5960), .Q (signal_5961) ) ;
    buf_clk cell_4119 ( .C (clk), .D (signal_5968), .Q (signal_5969) ) ;
    buf_clk cell_4127 ( .C (clk), .D (signal_5976), .Q (signal_5977) ) ;
    buf_clk cell_4135 ( .C (clk), .D (signal_5984), .Q (signal_5985) ) ;
    buf_clk cell_4143 ( .C (clk), .D (signal_5992), .Q (signal_5993) ) ;
    buf_clk cell_4151 ( .C (clk), .D (signal_6000), .Q (signal_6001) ) ;
    buf_clk cell_4159 ( .C (clk), .D (signal_6008), .Q (signal_6009) ) ;
    buf_clk cell_4167 ( .C (clk), .D (signal_6016), .Q (signal_6017) ) ;
    buf_clk cell_4175 ( .C (clk), .D (signal_6024), .Q (signal_6025) ) ;
    buf_clk cell_4183 ( .C (clk), .D (signal_6032), .Q (signal_6033) ) ;
    buf_clk cell_4191 ( .C (clk), .D (signal_6040), .Q (signal_6041) ) ;
    buf_clk cell_4199 ( .C (clk), .D (signal_6048), .Q (signal_6049) ) ;
    buf_clk cell_4207 ( .C (clk), .D (signal_6056), .Q (signal_6057) ) ;
    buf_clk cell_4215 ( .C (clk), .D (signal_6064), .Q (signal_6065) ) ;
    buf_clk cell_4223 ( .C (clk), .D (signal_6072), .Q (signal_6073) ) ;
    buf_clk cell_4231 ( .C (clk), .D (signal_6080), .Q (signal_6081) ) ;
    buf_clk cell_4239 ( .C (clk), .D (signal_6088), .Q (signal_6089) ) ;
    buf_clk cell_4247 ( .C (clk), .D (signal_6096), .Q (signal_6097) ) ;
    buf_clk cell_4255 ( .C (clk), .D (signal_6104), .Q (signal_6105) ) ;
    buf_clk cell_4263 ( .C (clk), .D (signal_6112), .Q (signal_6113) ) ;
    buf_clk cell_4271 ( .C (clk), .D (signal_6120), .Q (signal_6121) ) ;
    buf_clk cell_4279 ( .C (clk), .D (signal_6128), .Q (signal_6129) ) ;
    buf_clk cell_4287 ( .C (clk), .D (signal_6136), .Q (signal_6137) ) ;
    buf_clk cell_4295 ( .C (clk), .D (signal_6144), .Q (signal_6145) ) ;
    buf_clk cell_4303 ( .C (clk), .D (signal_6152), .Q (signal_6153) ) ;
    buf_clk cell_4311 ( .C (clk), .D (signal_6160), .Q (signal_6161) ) ;
    buf_clk cell_4319 ( .C (clk), .D (signal_6168), .Q (signal_6169) ) ;
    buf_clk cell_4327 ( .C (clk), .D (signal_6176), .Q (signal_6177) ) ;
    buf_clk cell_4335 ( .C (clk), .D (signal_6184), .Q (signal_6185) ) ;
    buf_clk cell_4343 ( .C (clk), .D (signal_6192), .Q (signal_6193) ) ;
    buf_clk cell_4351 ( .C (clk), .D (signal_6200), .Q (signal_6201) ) ;
    buf_clk cell_4359 ( .C (clk), .D (signal_6208), .Q (signal_6209) ) ;
    buf_clk cell_4367 ( .C (clk), .D (signal_6216), .Q (signal_6217) ) ;
    buf_clk cell_4375 ( .C (clk), .D (signal_6224), .Q (signal_6225) ) ;
    buf_clk cell_4383 ( .C (clk), .D (signal_6232), .Q (signal_6233) ) ;
    buf_clk cell_4391 ( .C (clk), .D (signal_6240), .Q (signal_6241) ) ;
    buf_clk cell_4399 ( .C (clk), .D (signal_6248), .Q (signal_6249) ) ;
    buf_clk cell_4407 ( .C (clk), .D (signal_6256), .Q (signal_6257) ) ;
    buf_clk cell_4415 ( .C (clk), .D (signal_6264), .Q (signal_6265) ) ;
    buf_clk cell_4423 ( .C (clk), .D (signal_6272), .Q (signal_6273) ) ;
    buf_clk cell_4431 ( .C (clk), .D (signal_6280), .Q (signal_6281) ) ;
    buf_clk cell_4439 ( .C (clk), .D (signal_6288), .Q (signal_6289) ) ;
    buf_clk cell_4447 ( .C (clk), .D (signal_6296), .Q (signal_6297) ) ;
    buf_clk cell_4455 ( .C (clk), .D (signal_6304), .Q (signal_6305) ) ;
    buf_clk cell_4463 ( .C (clk), .D (signal_6312), .Q (signal_6313) ) ;
    buf_clk cell_4471 ( .C (clk), .D (signal_6320), .Q (signal_6321) ) ;
    buf_clk cell_4479 ( .C (clk), .D (signal_6328), .Q (signal_6329) ) ;
    buf_clk cell_4487 ( .C (clk), .D (signal_6336), .Q (signal_6337) ) ;
    buf_clk cell_4495 ( .C (clk), .D (signal_6344), .Q (signal_6345) ) ;
    buf_clk cell_4503 ( .C (clk), .D (signal_6352), .Q (signal_6353) ) ;
    buf_clk cell_4511 ( .C (clk), .D (signal_6360), .Q (signal_6361) ) ;
    buf_clk cell_4519 ( .C (clk), .D (signal_6368), .Q (signal_6369) ) ;
    buf_clk cell_4527 ( .C (clk), .D (signal_6376), .Q (signal_6377) ) ;
    buf_clk cell_4535 ( .C (clk), .D (signal_6384), .Q (signal_6385) ) ;
    buf_clk cell_4543 ( .C (clk), .D (signal_6392), .Q (signal_6393) ) ;
    buf_clk cell_4551 ( .C (clk), .D (signal_6400), .Q (signal_6401) ) ;
    buf_clk cell_4559 ( .C (clk), .D (signal_6408), .Q (signal_6409) ) ;
    buf_clk cell_4567 ( .C (clk), .D (signal_6416), .Q (signal_6417) ) ;
    buf_clk cell_4575 ( .C (clk), .D (signal_6424), .Q (signal_6425) ) ;
    buf_clk cell_4583 ( .C (clk), .D (signal_6432), .Q (signal_6433) ) ;
    buf_clk cell_4591 ( .C (clk), .D (signal_6440), .Q (signal_6441) ) ;
    buf_clk cell_4599 ( .C (clk), .D (signal_6448), .Q (signal_6449) ) ;
    buf_clk cell_4607 ( .C (clk), .D (signal_6456), .Q (signal_6457) ) ;
    buf_clk cell_4615 ( .C (clk), .D (signal_6464), .Q (signal_6465) ) ;
    buf_clk cell_4623 ( .C (clk), .D (signal_6472), .Q (signal_6473) ) ;
    buf_clk cell_4631 ( .C (clk), .D (signal_6480), .Q (signal_6481) ) ;
    buf_clk cell_4639 ( .C (clk), .D (signal_6488), .Q (signal_6489) ) ;
    buf_clk cell_4647 ( .C (clk), .D (signal_6496), .Q (signal_6497) ) ;
    buf_clk cell_4655 ( .C (clk), .D (signal_6504), .Q (signal_6505) ) ;
    buf_clk cell_4663 ( .C (clk), .D (signal_6512), .Q (signal_6513) ) ;
    buf_clk cell_4671 ( .C (clk), .D (signal_6520), .Q (signal_6521) ) ;
    buf_clk cell_4679 ( .C (clk), .D (signal_6528), .Q (signal_6529) ) ;
    buf_clk cell_4687 ( .C (clk), .D (signal_6536), .Q (signal_6537) ) ;
    buf_clk cell_4695 ( .C (clk), .D (signal_6544), .Q (signal_6545) ) ;
    buf_clk cell_4703 ( .C (clk), .D (signal_6552), .Q (signal_6553) ) ;
    buf_clk cell_4711 ( .C (clk), .D (signal_6560), .Q (signal_6561) ) ;
    buf_clk cell_4719 ( .C (clk), .D (signal_6568), .Q (signal_6569) ) ;
    buf_clk cell_4727 ( .C (clk), .D (signal_6576), .Q (signal_6577) ) ;
    buf_clk cell_4735 ( .C (clk), .D (signal_6584), .Q (signal_6585) ) ;
    buf_clk cell_4743 ( .C (clk), .D (signal_6592), .Q (signal_6593) ) ;
    buf_clk cell_4751 ( .C (clk), .D (signal_6600), .Q (signal_6601) ) ;
    buf_clk cell_4759 ( .C (clk), .D (signal_6608), .Q (signal_6609) ) ;
    buf_clk cell_4767 ( .C (clk), .D (signal_6616), .Q (signal_6617) ) ;
    buf_clk cell_4775 ( .C (clk), .D (signal_6624), .Q (signal_6625) ) ;
    buf_clk cell_4783 ( .C (clk), .D (signal_6632), .Q (signal_6633) ) ;
    buf_clk cell_4791 ( .C (clk), .D (signal_6640), .Q (signal_6641) ) ;
    buf_clk cell_4799 ( .C (clk), .D (signal_6648), .Q (signal_6649) ) ;
    buf_clk cell_4807 ( .C (clk), .D (signal_6656), .Q (signal_6657) ) ;
    buf_clk cell_4815 ( .C (clk), .D (signal_6664), .Q (signal_6665) ) ;
    buf_clk cell_4823 ( .C (clk), .D (signal_6672), .Q (signal_6673) ) ;
    buf_clk cell_4831 ( .C (clk), .D (signal_6680), .Q (signal_6681) ) ;
    buf_clk cell_4839 ( .C (clk), .D (signal_6688), .Q (signal_6689) ) ;
    buf_clk cell_4847 ( .C (clk), .D (signal_6696), .Q (signal_6697) ) ;
    buf_clk cell_4855 ( .C (clk), .D (signal_6704), .Q (signal_6705) ) ;
    buf_clk cell_4863 ( .C (clk), .D (signal_6712), .Q (signal_6713) ) ;
    buf_clk cell_4871 ( .C (clk), .D (signal_6720), .Q (signal_6721) ) ;
    buf_clk cell_4879 ( .C (clk), .D (signal_6728), .Q (signal_6729) ) ;
    buf_clk cell_4887 ( .C (clk), .D (signal_6736), .Q (signal_6737) ) ;
    buf_clk cell_4895 ( .C (clk), .D (signal_6744), .Q (signal_6745) ) ;
    buf_clk cell_4903 ( .C (clk), .D (signal_6752), .Q (signal_6753) ) ;
    buf_clk cell_4911 ( .C (clk), .D (signal_6760), .Q (signal_6761) ) ;
    buf_clk cell_4919 ( .C (clk), .D (signal_6768), .Q (signal_6769) ) ;
    buf_clk cell_4927 ( .C (clk), .D (signal_6776), .Q (signal_6777) ) ;
    buf_clk cell_4935 ( .C (clk), .D (signal_6784), .Q (signal_6785) ) ;
    buf_clk cell_4943 ( .C (clk), .D (signal_6792), .Q (signal_6793) ) ;
    buf_clk cell_4951 ( .C (clk), .D (signal_6800), .Q (signal_6801) ) ;
    buf_clk cell_4959 ( .C (clk), .D (signal_6808), .Q (signal_6809) ) ;
    buf_clk cell_4967 ( .C (clk), .D (signal_6816), .Q (signal_6817) ) ;
    buf_clk cell_4975 ( .C (clk), .D (signal_6824), .Q (signal_6825) ) ;
    buf_clk cell_4983 ( .C (clk), .D (signal_6832), .Q (signal_6833) ) ;
    buf_clk cell_4991 ( .C (clk), .D (signal_6840), .Q (signal_6841) ) ;
    buf_clk cell_4999 ( .C (clk), .D (signal_6848), .Q (signal_6849) ) ;
    buf_clk cell_5007 ( .C (clk), .D (signal_6856), .Q (signal_6857) ) ;
    buf_clk cell_5015 ( .C (clk), .D (signal_6864), .Q (signal_6865) ) ;
    buf_clk cell_5023 ( .C (clk), .D (signal_6872), .Q (signal_6873) ) ;
    buf_clk cell_5031 ( .C (clk), .D (signal_6880), .Q (signal_6881) ) ;
    buf_clk cell_5039 ( .C (clk), .D (signal_6888), .Q (signal_6889) ) ;
    buf_clk cell_5047 ( .C (clk), .D (signal_6896), .Q (signal_6897) ) ;
    buf_clk cell_5055 ( .C (clk), .D (signal_6904), .Q (signal_6905) ) ;
    buf_clk cell_5063 ( .C (clk), .D (signal_6912), .Q (signal_6913) ) ;
    buf_clk cell_5071 ( .C (clk), .D (signal_6920), .Q (signal_6921) ) ;
    buf_clk cell_5079 ( .C (clk), .D (signal_6928), .Q (signal_6929) ) ;
    buf_clk cell_5087 ( .C (clk), .D (signal_6936), .Q (signal_6937) ) ;
    buf_clk cell_5095 ( .C (clk), .D (signal_6944), .Q (signal_6945) ) ;
    buf_clk cell_5103 ( .C (clk), .D (signal_6952), .Q (signal_6953) ) ;
    buf_clk cell_5111 ( .C (clk), .D (signal_6960), .Q (signal_6961) ) ;
    buf_clk cell_5119 ( .C (clk), .D (signal_6968), .Q (signal_6969) ) ;
    buf_clk cell_5127 ( .C (clk), .D (signal_6976), .Q (signal_6977) ) ;
    buf_clk cell_5135 ( .C (clk), .D (signal_6984), .Q (signal_6985) ) ;
    buf_clk cell_5143 ( .C (clk), .D (signal_6992), .Q (signal_6993) ) ;
    buf_clk cell_5151 ( .C (clk), .D (signal_7000), .Q (signal_7001) ) ;
    buf_clk cell_5159 ( .C (clk), .D (signal_7008), .Q (signal_7009) ) ;
    buf_clk cell_5167 ( .C (clk), .D (signal_7016), .Q (signal_7017) ) ;
    buf_clk cell_5175 ( .C (clk), .D (signal_7024), .Q (signal_7025) ) ;
    buf_clk cell_5183 ( .C (clk), .D (signal_7032), .Q (signal_7033) ) ;
    buf_clk cell_5191 ( .C (clk), .D (signal_7040), .Q (signal_7041) ) ;
    buf_clk cell_5199 ( .C (clk), .D (signal_7048), .Q (signal_7049) ) ;
    buf_clk cell_5207 ( .C (clk), .D (signal_7056), .Q (signal_7057) ) ;
    buf_clk cell_5215 ( .C (clk), .D (signal_7064), .Q (signal_7065) ) ;
    buf_clk cell_5223 ( .C (clk), .D (signal_7072), .Q (signal_7073) ) ;
    buf_clk cell_5231 ( .C (clk), .D (signal_7080), .Q (signal_7081) ) ;
    buf_clk cell_5239 ( .C (clk), .D (signal_7088), .Q (signal_7089) ) ;
    buf_clk cell_5247 ( .C (clk), .D (signal_7096), .Q (signal_7097) ) ;
    buf_clk cell_5255 ( .C (clk), .D (signal_7104), .Q (signal_7105) ) ;
    buf_clk cell_5263 ( .C (clk), .D (signal_7112), .Q (signal_7113) ) ;
    buf_clk cell_5271 ( .C (clk), .D (signal_7120), .Q (signal_7121) ) ;
    buf_clk cell_5279 ( .C (clk), .D (signal_7128), .Q (signal_7129) ) ;
    buf_clk cell_5287 ( .C (clk), .D (signal_7136), .Q (signal_7137) ) ;
    buf_clk cell_5295 ( .C (clk), .D (signal_7144), .Q (signal_7145) ) ;
    buf_clk cell_5303 ( .C (clk), .D (signal_7152), .Q (signal_7153) ) ;
    buf_clk cell_5311 ( .C (clk), .D (signal_7160), .Q (signal_7161) ) ;
    buf_clk cell_5319 ( .C (clk), .D (signal_7168), .Q (signal_7169) ) ;
    buf_clk cell_5327 ( .C (clk), .D (signal_7176), .Q (signal_7177) ) ;
    buf_clk cell_5335 ( .C (clk), .D (signal_7184), .Q (signal_7185) ) ;
    buf_clk cell_5343 ( .C (clk), .D (signal_7192), .Q (signal_7193) ) ;
    buf_clk cell_5351 ( .C (clk), .D (signal_7200), .Q (signal_7201) ) ;
    buf_clk cell_5359 ( .C (clk), .D (signal_7208), .Q (signal_7209) ) ;
    buf_clk cell_5367 ( .C (clk), .D (signal_7216), .Q (signal_7217) ) ;
    buf_clk cell_5375 ( .C (clk), .D (signal_7224), .Q (signal_7225) ) ;
    buf_clk cell_5383 ( .C (clk), .D (signal_7232), .Q (signal_7233) ) ;
    buf_clk cell_5391 ( .C (clk), .D (signal_7240), .Q (signal_7241) ) ;
    buf_clk cell_5399 ( .C (clk), .D (signal_7248), .Q (signal_7249) ) ;
    buf_clk cell_5407 ( .C (clk), .D (signal_7256), .Q (signal_7257) ) ;
    buf_clk cell_5415 ( .C (clk), .D (signal_7264), .Q (signal_7265) ) ;
    buf_clk cell_5423 ( .C (clk), .D (signal_7272), .Q (signal_7273) ) ;
    buf_clk cell_5431 ( .C (clk), .D (signal_7280), .Q (signal_7281) ) ;
    buf_clk cell_5439 ( .C (clk), .D (signal_7288), .Q (signal_7289) ) ;
    buf_clk cell_5447 ( .C (clk), .D (signal_7296), .Q (signal_7297) ) ;
    buf_clk cell_5455 ( .C (clk), .D (signal_7304), .Q (signal_7305) ) ;
    buf_clk cell_5463 ( .C (clk), .D (signal_7312), .Q (signal_7313) ) ;
    buf_clk cell_5471 ( .C (clk), .D (signal_7320), .Q (signal_7321) ) ;
    buf_clk cell_5479 ( .C (clk), .D (signal_7328), .Q (signal_7329) ) ;
    buf_clk cell_5487 ( .C (clk), .D (signal_7336), .Q (signal_7337) ) ;
    buf_clk cell_5495 ( .C (clk), .D (signal_7344), .Q (signal_7345) ) ;
    buf_clk cell_5503 ( .C (clk), .D (signal_7352), .Q (signal_7353) ) ;
    buf_clk cell_5511 ( .C (clk), .D (signal_7360), .Q (signal_7361) ) ;
    buf_clk cell_5519 ( .C (clk), .D (signal_7368), .Q (signal_7369) ) ;
    buf_clk cell_5527 ( .C (clk), .D (signal_7376), .Q (signal_7377) ) ;
    buf_clk cell_5535 ( .C (clk), .D (signal_7384), .Q (signal_7385) ) ;
    buf_clk cell_5543 ( .C (clk), .D (signal_7392), .Q (signal_7393) ) ;
    buf_clk cell_5551 ( .C (clk), .D (signal_7400), .Q (signal_7401) ) ;
    buf_clk cell_5559 ( .C (clk), .D (signal_7408), .Q (signal_7409) ) ;
    buf_clk cell_5567 ( .C (clk), .D (signal_7416), .Q (signal_7417) ) ;
    buf_clk cell_5575 ( .C (clk), .D (signal_7424), .Q (signal_7425) ) ;
    buf_clk cell_5583 ( .C (clk), .D (signal_7432), .Q (signal_7433) ) ;
    buf_clk cell_5591 ( .C (clk), .D (signal_7440), .Q (signal_7441) ) ;
    buf_clk cell_5599 ( .C (clk), .D (signal_7448), .Q (signal_7449) ) ;
    buf_clk cell_5607 ( .C (clk), .D (signal_7456), .Q (signal_7457) ) ;
    buf_clk cell_5615 ( .C (clk), .D (signal_7464), .Q (signal_7465) ) ;
    buf_clk cell_5623 ( .C (clk), .D (signal_7472), .Q (signal_7473) ) ;
    buf_clk cell_5631 ( .C (clk), .D (signal_7480), .Q (signal_7481) ) ;
    buf_clk cell_5639 ( .C (clk), .D (signal_7488), .Q (signal_7489) ) ;
    buf_clk cell_5647 ( .C (clk), .D (signal_7496), .Q (signal_7497) ) ;
    buf_clk cell_5655 ( .C (clk), .D (signal_7504), .Q (signal_7505) ) ;
    buf_clk cell_5663 ( .C (clk), .D (signal_7512), .Q (signal_7513) ) ;
    buf_clk cell_5671 ( .C (clk), .D (signal_7520), .Q (signal_7521) ) ;
    buf_clk cell_5679 ( .C (clk), .D (signal_7528), .Q (signal_7529) ) ;
    buf_clk cell_5687 ( .C (clk), .D (signal_7536), .Q (signal_7537) ) ;
    buf_clk cell_5695 ( .C (clk), .D (signal_7544), .Q (signal_7545) ) ;
    buf_clk cell_5703 ( .C (clk), .D (signal_7552), .Q (signal_7553) ) ;
    buf_clk cell_5711 ( .C (clk), .D (signal_7560), .Q (signal_7561) ) ;
    buf_clk cell_5719 ( .C (clk), .D (signal_7568), .Q (signal_7569) ) ;
    buf_clk cell_5727 ( .C (clk), .D (signal_7576), .Q (signal_7577) ) ;
    buf_clk cell_5735 ( .C (clk), .D (signal_7584), .Q (signal_7585) ) ;
    buf_clk cell_5743 ( .C (clk), .D (signal_7592), .Q (signal_7593) ) ;
    buf_clk cell_5751 ( .C (clk), .D (signal_7600), .Q (signal_7601) ) ;
    buf_clk cell_5759 ( .C (clk), .D (signal_7608), .Q (signal_7609) ) ;
    buf_clk cell_5767 ( .C (clk), .D (signal_7616), .Q (signal_7617) ) ;
    buf_clk cell_5775 ( .C (clk), .D (signal_7624), .Q (signal_7625) ) ;
    buf_clk cell_5783 ( .C (clk), .D (signal_7632), .Q (signal_7633) ) ;
    buf_clk cell_5791 ( .C (clk), .D (signal_7640), .Q (signal_7641) ) ;
    buf_clk cell_5799 ( .C (clk), .D (signal_7648), .Q (signal_7649) ) ;
    buf_clk cell_5807 ( .C (clk), .D (signal_7656), .Q (signal_7657) ) ;
    buf_clk cell_5815 ( .C (clk), .D (signal_7664), .Q (signal_7665) ) ;
    buf_clk cell_5823 ( .C (clk), .D (signal_7672), .Q (signal_7673) ) ;
    buf_clk cell_5831 ( .C (clk), .D (signal_7680), .Q (signal_7681) ) ;
    buf_clk cell_5839 ( .C (clk), .D (signal_7688), .Q (signal_7689) ) ;
    buf_clk cell_5847 ( .C (clk), .D (signal_7696), .Q (signal_7697) ) ;
    buf_clk cell_5855 ( .C (clk), .D (signal_7704), .Q (signal_7705) ) ;
    buf_clk cell_5863 ( .C (clk), .D (signal_7712), .Q (signal_7713) ) ;
    buf_clk cell_5871 ( .C (clk), .D (signal_7720), .Q (signal_7721) ) ;
    buf_clk cell_5879 ( .C (clk), .D (signal_7728), .Q (signal_7729) ) ;
    buf_clk cell_5887 ( .C (clk), .D (signal_7736), .Q (signal_7737) ) ;
    buf_clk cell_5895 ( .C (clk), .D (signal_7744), .Q (signal_7745) ) ;
    buf_clk cell_5903 ( .C (clk), .D (signal_7752), .Q (signal_7753) ) ;
    buf_clk cell_5911 ( .C (clk), .D (signal_7760), .Q (signal_7761) ) ;
    buf_clk cell_5919 ( .C (clk), .D (signal_7768), .Q (signal_7769) ) ;
    buf_clk cell_5927 ( .C (clk), .D (signal_7776), .Q (signal_7777) ) ;
    buf_clk cell_5935 ( .C (clk), .D (signal_7784), .Q (signal_7785) ) ;
    buf_clk cell_5943 ( .C (clk), .D (signal_7792), .Q (signal_7793) ) ;
    buf_clk cell_5951 ( .C (clk), .D (signal_7800), .Q (signal_7801) ) ;
    buf_clk cell_5959 ( .C (clk), .D (signal_7808), .Q (signal_7809) ) ;
    buf_clk cell_5967 ( .C (clk), .D (signal_7816), .Q (signal_7817) ) ;
    buf_clk cell_5975 ( .C (clk), .D (signal_7824), .Q (signal_7825) ) ;
    buf_clk cell_5983 ( .C (clk), .D (signal_7832), .Q (signal_7833) ) ;
    buf_clk cell_5991 ( .C (clk), .D (signal_7840), .Q (signal_7841) ) ;
    buf_clk cell_5999 ( .C (clk), .D (signal_7848), .Q (signal_7849) ) ;
    buf_clk cell_6007 ( .C (clk), .D (signal_7856), .Q (signal_7857) ) ;
    buf_clk cell_6015 ( .C (clk), .D (signal_7864), .Q (signal_7865) ) ;
    buf_clk cell_6023 ( .C (clk), .D (signal_7872), .Q (signal_7873) ) ;
    buf_clk cell_6031 ( .C (clk), .D (signal_7880), .Q (signal_7881) ) ;
    buf_clk cell_6039 ( .C (clk), .D (signal_7888), .Q (signal_7889) ) ;
    buf_clk cell_6047 ( .C (clk), .D (signal_7896), .Q (signal_7897) ) ;
    buf_clk cell_6055 ( .C (clk), .D (signal_7904), .Q (signal_7905) ) ;
    buf_clk cell_6063 ( .C (clk), .D (signal_7912), .Q (signal_7913) ) ;
    buf_clk cell_6071 ( .C (clk), .D (signal_7920), .Q (signal_7921) ) ;
    buf_clk cell_6079 ( .C (clk), .D (signal_7928), .Q (signal_7929) ) ;
    buf_clk cell_6087 ( .C (clk), .D (signal_7936), .Q (signal_7937) ) ;
    buf_clk cell_6095 ( .C (clk), .D (signal_7944), .Q (signal_7945) ) ;
    buf_clk cell_6103 ( .C (clk), .D (signal_7952), .Q (signal_7953) ) ;
    buf_clk cell_6111 ( .C (clk), .D (signal_7960), .Q (signal_7961) ) ;
    buf_clk cell_6119 ( .C (clk), .D (signal_7968), .Q (signal_7969) ) ;
    buf_clk cell_6127 ( .C (clk), .D (signal_7976), .Q (signal_7977) ) ;
    buf_clk cell_6135 ( .C (clk), .D (signal_7984), .Q (signal_7985) ) ;
    buf_clk cell_6143 ( .C (clk), .D (signal_7992), .Q (signal_7993) ) ;
    buf_clk cell_6151 ( .C (clk), .D (signal_8000), .Q (signal_8001) ) ;
    buf_clk cell_6159 ( .C (clk), .D (signal_8008), .Q (signal_8009) ) ;
    buf_clk cell_6167 ( .C (clk), .D (signal_8016), .Q (signal_8017) ) ;
    buf_clk cell_6175 ( .C (clk), .D (signal_8024), .Q (signal_8025) ) ;
    buf_clk cell_6183 ( .C (clk), .D (signal_8032), .Q (signal_8033) ) ;
    buf_clk cell_6191 ( .C (clk), .D (signal_8040), .Q (signal_8041) ) ;
    buf_clk cell_6199 ( .C (clk), .D (signal_8048), .Q (signal_8049) ) ;
    buf_clk cell_6207 ( .C (clk), .D (signal_8056), .Q (signal_8057) ) ;
    buf_clk cell_6215 ( .C (clk), .D (signal_8064), .Q (signal_8065) ) ;
    buf_clk cell_6223 ( .C (clk), .D (signal_8072), .Q (signal_8073) ) ;
    buf_clk cell_6231 ( .C (clk), .D (signal_8080), .Q (signal_8081) ) ;
    buf_clk cell_6239 ( .C (clk), .D (signal_8088), .Q (signal_8089) ) ;
    buf_clk cell_6247 ( .C (clk), .D (signal_8096), .Q (signal_8097) ) ;
    buf_clk cell_6255 ( .C (clk), .D (signal_8104), .Q (signal_8105) ) ;
    buf_clk cell_6263 ( .C (clk), .D (signal_8112), .Q (signal_8113) ) ;
    buf_clk cell_6271 ( .C (clk), .D (signal_8120), .Q (signal_8121) ) ;
    buf_clk cell_6279 ( .C (clk), .D (signal_8128), .Q (signal_8129) ) ;
    buf_clk cell_6287 ( .C (clk), .D (signal_8136), .Q (signal_8137) ) ;
    buf_clk cell_6295 ( .C (clk), .D (signal_8144), .Q (signal_8145) ) ;
    buf_clk cell_6303 ( .C (clk), .D (signal_8152), .Q (signal_8153) ) ;
    buf_clk cell_6311 ( .C (clk), .D (signal_8160), .Q (signal_8161) ) ;
    buf_clk cell_6319 ( .C (clk), .D (signal_8168), .Q (signal_8169) ) ;
    buf_clk cell_6327 ( .C (clk), .D (signal_8176), .Q (signal_8177) ) ;
    buf_clk cell_6335 ( .C (clk), .D (signal_8184), .Q (signal_8185) ) ;
    buf_clk cell_6343 ( .C (clk), .D (signal_8192), .Q (signal_8193) ) ;
    buf_clk cell_6351 ( .C (clk), .D (signal_8200), .Q (signal_8201) ) ;
    buf_clk cell_6359 ( .C (clk), .D (signal_8208), .Q (signal_8209) ) ;
    buf_clk cell_6367 ( .C (clk), .D (signal_8216), .Q (signal_8217) ) ;
    buf_clk cell_6375 ( .C (clk), .D (signal_8224), .Q (signal_8225) ) ;
    buf_clk cell_6383 ( .C (clk), .D (signal_8232), .Q (signal_8233) ) ;
    buf_clk cell_6391 ( .C (clk), .D (signal_8240), .Q (signal_8241) ) ;
    buf_clk cell_6399 ( .C (clk), .D (signal_8248), .Q (signal_8249) ) ;
    buf_clk cell_6407 ( .C (clk), .D (signal_8256), .Q (signal_8257) ) ;
    buf_clk cell_6415 ( .C (clk), .D (signal_8264), .Q (signal_8265) ) ;
    buf_clk cell_6423 ( .C (clk), .D (signal_8272), .Q (signal_8273) ) ;
    buf_clk cell_6431 ( .C (clk), .D (signal_8280), .Q (signal_8281) ) ;
    buf_clk cell_6439 ( .C (clk), .D (signal_8288), .Q (signal_8289) ) ;
    buf_clk cell_6447 ( .C (clk), .D (signal_8296), .Q (signal_8297) ) ;
    buf_clk cell_6455 ( .C (clk), .D (signal_8304), .Q (signal_8305) ) ;
    buf_clk cell_6463 ( .C (clk), .D (signal_8312), .Q (signal_8313) ) ;
    buf_clk cell_6471 ( .C (clk), .D (signal_8320), .Q (signal_8321) ) ;
    buf_clk cell_6479 ( .C (clk), .D (signal_8328), .Q (signal_8329) ) ;
    buf_clk cell_6487 ( .C (clk), .D (signal_8336), .Q (signal_8337) ) ;
    buf_clk cell_6495 ( .C (clk), .D (signal_8344), .Q (signal_8345) ) ;
    buf_clk cell_6503 ( .C (clk), .D (signal_8352), .Q (signal_8353) ) ;
    buf_clk cell_6511 ( .C (clk), .D (signal_8360), .Q (signal_8361) ) ;
    buf_clk cell_6519 ( .C (clk), .D (signal_8368), .Q (signal_8369) ) ;
    buf_clk cell_6527 ( .C (clk), .D (signal_8376), .Q (signal_8377) ) ;
    buf_clk cell_6535 ( .C (clk), .D (signal_8384), .Q (signal_8385) ) ;
    buf_clk cell_6543 ( .C (clk), .D (signal_8392), .Q (signal_8393) ) ;
    buf_clk cell_6551 ( .C (clk), .D (signal_8400), .Q (signal_8401) ) ;
    buf_clk cell_6559 ( .C (clk), .D (signal_8408), .Q (signal_8409) ) ;
    buf_clk cell_6567 ( .C (clk), .D (signal_8416), .Q (signal_8417) ) ;
    buf_clk cell_6575 ( .C (clk), .D (signal_8424), .Q (signal_8425) ) ;
    buf_clk cell_6583 ( .C (clk), .D (signal_8432), .Q (signal_8433) ) ;
    buf_clk cell_6591 ( .C (clk), .D (signal_8440), .Q (signal_8441) ) ;
    buf_clk cell_6599 ( .C (clk), .D (signal_8448), .Q (signal_8449) ) ;
    buf_clk cell_6607 ( .C (clk), .D (signal_8456), .Q (signal_8457) ) ;
    buf_clk cell_6615 ( .C (clk), .D (signal_8464), .Q (signal_8465) ) ;
    buf_clk cell_6623 ( .C (clk), .D (signal_8472), .Q (signal_8473) ) ;
    buf_clk cell_6631 ( .C (clk), .D (signal_8480), .Q (signal_8481) ) ;
    buf_clk cell_6639 ( .C (clk), .D (signal_8488), .Q (signal_8489) ) ;
    buf_clk cell_6647 ( .C (clk), .D (signal_8496), .Q (signal_8497) ) ;
    buf_clk cell_6655 ( .C (clk), .D (signal_8504), .Q (signal_8505) ) ;
    buf_clk cell_6663 ( .C (clk), .D (signal_8512), .Q (signal_8513) ) ;
    buf_clk cell_6671 ( .C (clk), .D (signal_8520), .Q (signal_8521) ) ;
    buf_clk cell_6679 ( .C (clk), .D (signal_8528), .Q (signal_8529) ) ;
    buf_clk cell_6687 ( .C (clk), .D (signal_8536), .Q (signal_8537) ) ;
    buf_clk cell_6695 ( .C (clk), .D (signal_8544), .Q (signal_8545) ) ;
    buf_clk cell_6703 ( .C (clk), .D (signal_8552), .Q (signal_8553) ) ;
    buf_clk cell_6711 ( .C (clk), .D (signal_8560), .Q (signal_8561) ) ;
    buf_clk cell_6719 ( .C (clk), .D (signal_8568), .Q (signal_8569) ) ;
    buf_clk cell_6727 ( .C (clk), .D (signal_8576), .Q (signal_8577) ) ;
    buf_clk cell_6735 ( .C (clk), .D (signal_8584), .Q (signal_8585) ) ;
    buf_clk cell_6743 ( .C (clk), .D (signal_8592), .Q (signal_8593) ) ;
    buf_clk cell_6751 ( .C (clk), .D (signal_8600), .Q (signal_8601) ) ;
    buf_clk cell_6759 ( .C (clk), .D (signal_8608), .Q (signal_8609) ) ;
    buf_clk cell_6767 ( .C (clk), .D (signal_8616), .Q (signal_8617) ) ;
    buf_clk cell_6775 ( .C (clk), .D (signal_8624), .Q (signal_8625) ) ;
    buf_clk cell_6783 ( .C (clk), .D (signal_8632), .Q (signal_8633) ) ;
    buf_clk cell_6791 ( .C (clk), .D (signal_8640), .Q (signal_8641) ) ;
    buf_clk cell_6799 ( .C (clk), .D (signal_8648), .Q (signal_8649) ) ;
    buf_clk cell_6807 ( .C (clk), .D (signal_8656), .Q (signal_8657) ) ;
    buf_clk cell_6815 ( .C (clk), .D (signal_8664), .Q (signal_8665) ) ;
    buf_clk cell_6823 ( .C (clk), .D (signal_8672), .Q (signal_8673) ) ;
    buf_clk cell_6831 ( .C (clk), .D (signal_8680), .Q (signal_8681) ) ;
    buf_clk cell_6839 ( .C (clk), .D (signal_8688), .Q (signal_8689) ) ;
    buf_clk cell_6847 ( .C (clk), .D (signal_8696), .Q (signal_8697) ) ;
    buf_clk cell_6855 ( .C (clk), .D (signal_8704), .Q (signal_8705) ) ;
    buf_clk cell_6863 ( .C (clk), .D (signal_8712), .Q (signal_8713) ) ;
    buf_clk cell_6871 ( .C (clk), .D (signal_8720), .Q (signal_8721) ) ;
    buf_clk cell_6879 ( .C (clk), .D (signal_8728), .Q (signal_8729) ) ;
    buf_clk cell_6887 ( .C (clk), .D (signal_8736), .Q (signal_8737) ) ;
    buf_clk cell_6895 ( .C (clk), .D (signal_8744), .Q (signal_8745) ) ;
    buf_clk cell_6903 ( .C (clk), .D (signal_8752), .Q (signal_8753) ) ;
    buf_clk cell_6911 ( .C (clk), .D (signal_8760), .Q (signal_8761) ) ;
    buf_clk cell_6919 ( .C (clk), .D (signal_8768), .Q (signal_8769) ) ;
    buf_clk cell_6927 ( .C (clk), .D (signal_8776), .Q (signal_8777) ) ;
    buf_clk cell_6935 ( .C (clk), .D (signal_8784), .Q (signal_8785) ) ;
    buf_clk cell_6943 ( .C (clk), .D (signal_8792), .Q (signal_8793) ) ;
    buf_clk cell_6951 ( .C (clk), .D (signal_8800), .Q (signal_8801) ) ;
    buf_clk cell_6959 ( .C (clk), .D (signal_8808), .Q (signal_8809) ) ;
    buf_clk cell_6967 ( .C (clk), .D (signal_8816), .Q (signal_8817) ) ;
    buf_clk cell_6975 ( .C (clk), .D (signal_8824), .Q (signal_8825) ) ;
    buf_clk cell_6983 ( .C (clk), .D (signal_8832), .Q (signal_8833) ) ;
    buf_clk cell_6991 ( .C (clk), .D (signal_8840), .Q (signal_8841) ) ;
    buf_clk cell_6999 ( .C (clk), .D (signal_8848), .Q (signal_8849) ) ;
    buf_clk cell_7007 ( .C (clk), .D (signal_8856), .Q (signal_8857) ) ;
    buf_clk cell_7015 ( .C (clk), .D (signal_8864), .Q (signal_8865) ) ;
    buf_clk cell_7023 ( .C (clk), .D (signal_8872), .Q (signal_8873) ) ;
    buf_clk cell_7031 ( .C (clk), .D (signal_8880), .Q (signal_8881) ) ;
    buf_clk cell_7039 ( .C (clk), .D (signal_8888), .Q (signal_8889) ) ;
    buf_clk cell_7047 ( .C (clk), .D (signal_8896), .Q (signal_8897) ) ;
    buf_clk cell_7055 ( .C (clk), .D (signal_8904), .Q (signal_8905) ) ;
    buf_clk cell_7063 ( .C (clk), .D (signal_8912), .Q (signal_8913) ) ;
    buf_clk cell_7071 ( .C (clk), .D (signal_8920), .Q (signal_8921) ) ;
    buf_clk cell_7079 ( .C (clk), .D (signal_8928), .Q (signal_8929) ) ;
    buf_clk cell_7087 ( .C (clk), .D (signal_8936), .Q (signal_8937) ) ;
    buf_clk cell_7095 ( .C (clk), .D (signal_8944), .Q (signal_8945) ) ;

    /* cells in depth 3 */
    buf_clk cell_1862 ( .C (clk), .D (signal_2029), .Q (signal_3712) ) ;
    buf_clk cell_1864 ( .C (clk), .D (signal_3497), .Q (signal_3714) ) ;
    buf_clk cell_1866 ( .C (clk), .D (signal_2033), .Q (signal_3716) ) ;
    buf_clk cell_1868 ( .C (clk), .D (signal_3509), .Q (signal_3718) ) ;
    buf_clk cell_1870 ( .C (clk), .D (signal_2034), .Q (signal_3720) ) ;
    buf_clk cell_1872 ( .C (clk), .D (signal_3510), .Q (signal_3722) ) ;
    buf_clk cell_1874 ( .C (clk), .D (signal_2036), .Q (signal_3724) ) ;
    buf_clk cell_1876 ( .C (clk), .D (signal_3512), .Q (signal_3726) ) ;
    buf_clk cell_1896 ( .C (clk), .D (signal_3745), .Q (signal_3746) ) ;
    buf_clk cell_1904 ( .C (clk), .D (signal_3753), .Q (signal_3754) ) ;
    buf_clk cell_1912 ( .C (clk), .D (signal_3761), .Q (signal_3762) ) ;
    buf_clk cell_1920 ( .C (clk), .D (signal_3769), .Q (signal_3770) ) ;
    buf_clk cell_1928 ( .C (clk), .D (signal_3777), .Q (signal_3778) ) ;
    buf_clk cell_1936 ( .C (clk), .D (signal_3785), .Q (signal_3786) ) ;
    buf_clk cell_1944 ( .C (clk), .D (signal_3793), .Q (signal_3794) ) ;
    buf_clk cell_1952 ( .C (clk), .D (signal_3801), .Q (signal_3802) ) ;
    buf_clk cell_1960 ( .C (clk), .D (signal_3809), .Q (signal_3810) ) ;
    buf_clk cell_1968 ( .C (clk), .D (signal_3817), .Q (signal_3818) ) ;
    buf_clk cell_1976 ( .C (clk), .D (signal_3825), .Q (signal_3826) ) ;
    buf_clk cell_1984 ( .C (clk), .D (signal_3833), .Q (signal_3834) ) ;
    buf_clk cell_1992 ( .C (clk), .D (signal_3841), .Q (signal_3842) ) ;
    buf_clk cell_2000 ( .C (clk), .D (signal_3849), .Q (signal_3850) ) ;
    buf_clk cell_2008 ( .C (clk), .D (signal_3857), .Q (signal_3858) ) ;
    buf_clk cell_2016 ( .C (clk), .D (signal_3865), .Q (signal_3866) ) ;
    buf_clk cell_2024 ( .C (clk), .D (signal_3873), .Q (signal_3874) ) ;
    buf_clk cell_2032 ( .C (clk), .D (signal_3881), .Q (signal_3882) ) ;
    buf_clk cell_2040 ( .C (clk), .D (signal_3889), .Q (signal_3890) ) ;
    buf_clk cell_2048 ( .C (clk), .D (signal_3897), .Q (signal_3898) ) ;
    buf_clk cell_2056 ( .C (clk), .D (signal_3905), .Q (signal_3906) ) ;
    buf_clk cell_2064 ( .C (clk), .D (signal_3913), .Q (signal_3914) ) ;
    buf_clk cell_2072 ( .C (clk), .D (signal_3921), .Q (signal_3922) ) ;
    buf_clk cell_2080 ( .C (clk), .D (signal_3929), .Q (signal_3930) ) ;
    buf_clk cell_2088 ( .C (clk), .D (signal_3937), .Q (signal_3938) ) ;
    buf_clk cell_2096 ( .C (clk), .D (signal_3945), .Q (signal_3946) ) ;
    buf_clk cell_2104 ( .C (clk), .D (signal_3953), .Q (signal_3954) ) ;
    buf_clk cell_2112 ( .C (clk), .D (signal_3961), .Q (signal_3962) ) ;
    buf_clk cell_2120 ( .C (clk), .D (signal_3969), .Q (signal_3970) ) ;
    buf_clk cell_2128 ( .C (clk), .D (signal_3977), .Q (signal_3978) ) ;
    buf_clk cell_2136 ( .C (clk), .D (signal_3985), .Q (signal_3986) ) ;
    buf_clk cell_2144 ( .C (clk), .D (signal_3993), .Q (signal_3994) ) ;
    buf_clk cell_2152 ( .C (clk), .D (signal_4001), .Q (signal_4002) ) ;
    buf_clk cell_2160 ( .C (clk), .D (signal_4009), .Q (signal_4010) ) ;
    buf_clk cell_2168 ( .C (clk), .D (signal_4017), .Q (signal_4018) ) ;
    buf_clk cell_2176 ( .C (clk), .D (signal_4025), .Q (signal_4026) ) ;
    buf_clk cell_2184 ( .C (clk), .D (signal_4033), .Q (signal_4034) ) ;
    buf_clk cell_2192 ( .C (clk), .D (signal_4041), .Q (signal_4042) ) ;
    buf_clk cell_2200 ( .C (clk), .D (signal_4049), .Q (signal_4050) ) ;
    buf_clk cell_2208 ( .C (clk), .D (signal_4057), .Q (signal_4058) ) ;
    buf_clk cell_2216 ( .C (clk), .D (signal_4065), .Q (signal_4066) ) ;
    buf_clk cell_2224 ( .C (clk), .D (signal_4073), .Q (signal_4074) ) ;
    buf_clk cell_2232 ( .C (clk), .D (signal_4081), .Q (signal_4082) ) ;
    buf_clk cell_2240 ( .C (clk), .D (signal_4089), .Q (signal_4090) ) ;
    buf_clk cell_2248 ( .C (clk), .D (signal_4097), .Q (signal_4098) ) ;
    buf_clk cell_2256 ( .C (clk), .D (signal_4105), .Q (signal_4106) ) ;
    buf_clk cell_2264 ( .C (clk), .D (signal_4113), .Q (signal_4114) ) ;
    buf_clk cell_2272 ( .C (clk), .D (signal_4121), .Q (signal_4122) ) ;
    buf_clk cell_2280 ( .C (clk), .D (signal_4129), .Q (signal_4130) ) ;
    buf_clk cell_2288 ( .C (clk), .D (signal_4137), .Q (signal_4138) ) ;
    buf_clk cell_2296 ( .C (clk), .D (signal_4145), .Q (signal_4146) ) ;
    buf_clk cell_2304 ( .C (clk), .D (signal_4153), .Q (signal_4154) ) ;
    buf_clk cell_2312 ( .C (clk), .D (signal_4161), .Q (signal_4162) ) ;
    buf_clk cell_2320 ( .C (clk), .D (signal_4169), .Q (signal_4170) ) ;
    buf_clk cell_2328 ( .C (clk), .D (signal_4177), .Q (signal_4178) ) ;
    buf_clk cell_2336 ( .C (clk), .D (signal_4185), .Q (signal_4186) ) ;
    buf_clk cell_2344 ( .C (clk), .D (signal_4193), .Q (signal_4194) ) ;
    buf_clk cell_2352 ( .C (clk), .D (signal_4201), .Q (signal_4202) ) ;
    buf_clk cell_2360 ( .C (clk), .D (signal_4209), .Q (signal_4210) ) ;
    buf_clk cell_2368 ( .C (clk), .D (signal_4217), .Q (signal_4218) ) ;
    buf_clk cell_2376 ( .C (clk), .D (signal_4225), .Q (signal_4226) ) ;
    buf_clk cell_2384 ( .C (clk), .D (signal_4233), .Q (signal_4234) ) ;
    buf_clk cell_2392 ( .C (clk), .D (signal_4241), .Q (signal_4242) ) ;
    buf_clk cell_2400 ( .C (clk), .D (signal_4249), .Q (signal_4250) ) ;
    buf_clk cell_2408 ( .C (clk), .D (signal_4257), .Q (signal_4258) ) ;
    buf_clk cell_2416 ( .C (clk), .D (signal_4265), .Q (signal_4266) ) ;
    buf_clk cell_2424 ( .C (clk), .D (signal_4273), .Q (signal_4274) ) ;
    buf_clk cell_2432 ( .C (clk), .D (signal_4281), .Q (signal_4282) ) ;
    buf_clk cell_2440 ( .C (clk), .D (signal_4289), .Q (signal_4290) ) ;
    buf_clk cell_2448 ( .C (clk), .D (signal_4297), .Q (signal_4298) ) ;
    buf_clk cell_2456 ( .C (clk), .D (signal_4305), .Q (signal_4306) ) ;
    buf_clk cell_2464 ( .C (clk), .D (signal_4313), .Q (signal_4314) ) ;
    buf_clk cell_2472 ( .C (clk), .D (signal_4321), .Q (signal_4322) ) ;
    buf_clk cell_2480 ( .C (clk), .D (signal_4329), .Q (signal_4330) ) ;
    buf_clk cell_2488 ( .C (clk), .D (signal_4337), .Q (signal_4338) ) ;
    buf_clk cell_2496 ( .C (clk), .D (signal_4345), .Q (signal_4346) ) ;
    buf_clk cell_2504 ( .C (clk), .D (signal_4353), .Q (signal_4354) ) ;
    buf_clk cell_2512 ( .C (clk), .D (signal_4361), .Q (signal_4362) ) ;
    buf_clk cell_2520 ( .C (clk), .D (signal_4369), .Q (signal_4370) ) ;
    buf_clk cell_2528 ( .C (clk), .D (signal_4377), .Q (signal_4378) ) ;
    buf_clk cell_2536 ( .C (clk), .D (signal_4385), .Q (signal_4386) ) ;
    buf_clk cell_2544 ( .C (clk), .D (signal_4393), .Q (signal_4394) ) ;
    buf_clk cell_2552 ( .C (clk), .D (signal_4401), .Q (signal_4402) ) ;
    buf_clk cell_2560 ( .C (clk), .D (signal_4409), .Q (signal_4410) ) ;
    buf_clk cell_2568 ( .C (clk), .D (signal_4417), .Q (signal_4418) ) ;
    buf_clk cell_2576 ( .C (clk), .D (signal_4425), .Q (signal_4426) ) ;
    buf_clk cell_2584 ( .C (clk), .D (signal_4433), .Q (signal_4434) ) ;
    buf_clk cell_2592 ( .C (clk), .D (signal_4441), .Q (signal_4442) ) ;
    buf_clk cell_2600 ( .C (clk), .D (signal_4449), .Q (signal_4450) ) ;
    buf_clk cell_2608 ( .C (clk), .D (signal_4457), .Q (signal_4458) ) ;
    buf_clk cell_2616 ( .C (clk), .D (signal_4465), .Q (signal_4466) ) ;
    buf_clk cell_2624 ( .C (clk), .D (signal_4473), .Q (signal_4474) ) ;
    buf_clk cell_2632 ( .C (clk), .D (signal_4481), .Q (signal_4482) ) ;
    buf_clk cell_2640 ( .C (clk), .D (signal_4489), .Q (signal_4490) ) ;
    buf_clk cell_2648 ( .C (clk), .D (signal_4497), .Q (signal_4498) ) ;
    buf_clk cell_2656 ( .C (clk), .D (signal_4505), .Q (signal_4506) ) ;
    buf_clk cell_2664 ( .C (clk), .D (signal_4513), .Q (signal_4514) ) ;
    buf_clk cell_2672 ( .C (clk), .D (signal_4521), .Q (signal_4522) ) ;
    buf_clk cell_2680 ( .C (clk), .D (signal_4529), .Q (signal_4530) ) ;
    buf_clk cell_2688 ( .C (clk), .D (signal_4537), .Q (signal_4538) ) ;
    buf_clk cell_2696 ( .C (clk), .D (signal_4545), .Q (signal_4546) ) ;
    buf_clk cell_2704 ( .C (clk), .D (signal_4553), .Q (signal_4554) ) ;
    buf_clk cell_2712 ( .C (clk), .D (signal_4561), .Q (signal_4562) ) ;
    buf_clk cell_2720 ( .C (clk), .D (signal_4569), .Q (signal_4570) ) ;
    buf_clk cell_2728 ( .C (clk), .D (signal_4577), .Q (signal_4578) ) ;
    buf_clk cell_2736 ( .C (clk), .D (signal_4585), .Q (signal_4586) ) ;
    buf_clk cell_2744 ( .C (clk), .D (signal_4593), .Q (signal_4594) ) ;
    buf_clk cell_2752 ( .C (clk), .D (signal_4601), .Q (signal_4602) ) ;
    buf_clk cell_2760 ( .C (clk), .D (signal_4609), .Q (signal_4610) ) ;
    buf_clk cell_2768 ( .C (clk), .D (signal_4617), .Q (signal_4618) ) ;
    buf_clk cell_2776 ( .C (clk), .D (signal_4625), .Q (signal_4626) ) ;
    buf_clk cell_2784 ( .C (clk), .D (signal_4633), .Q (signal_4634) ) ;
    buf_clk cell_2792 ( .C (clk), .D (signal_4641), .Q (signal_4642) ) ;
    buf_clk cell_2800 ( .C (clk), .D (signal_4649), .Q (signal_4650) ) ;
    buf_clk cell_2808 ( .C (clk), .D (signal_4657), .Q (signal_4658) ) ;
    buf_clk cell_2816 ( .C (clk), .D (signal_4665), .Q (signal_4666) ) ;
    buf_clk cell_2824 ( .C (clk), .D (signal_4673), .Q (signal_4674) ) ;
    buf_clk cell_2832 ( .C (clk), .D (signal_4681), .Q (signal_4682) ) ;
    buf_clk cell_2840 ( .C (clk), .D (signal_4689), .Q (signal_4690) ) ;
    buf_clk cell_2848 ( .C (clk), .D (signal_4697), .Q (signal_4698) ) ;
    buf_clk cell_2856 ( .C (clk), .D (signal_4705), .Q (signal_4706) ) ;
    buf_clk cell_2864 ( .C (clk), .D (signal_4713), .Q (signal_4714) ) ;
    buf_clk cell_2872 ( .C (clk), .D (signal_4721), .Q (signal_4722) ) ;
    buf_clk cell_2880 ( .C (clk), .D (signal_4729), .Q (signal_4730) ) ;
    buf_clk cell_2888 ( .C (clk), .D (signal_4737), .Q (signal_4738) ) ;
    buf_clk cell_2896 ( .C (clk), .D (signal_4745), .Q (signal_4746) ) ;
    buf_clk cell_2904 ( .C (clk), .D (signal_4753), .Q (signal_4754) ) ;
    buf_clk cell_2910 ( .C (clk), .D (signal_4759), .Q (signal_4760) ) ;
    buf_clk cell_2916 ( .C (clk), .D (signal_4765), .Q (signal_4766) ) ;
    buf_clk cell_2922 ( .C (clk), .D (signal_4771), .Q (signal_4772) ) ;
    buf_clk cell_2928 ( .C (clk), .D (signal_4777), .Q (signal_4778) ) ;
    buf_clk cell_2934 ( .C (clk), .D (signal_4783), .Q (signal_4784) ) ;
    buf_clk cell_2940 ( .C (clk), .D (signal_4789), .Q (signal_4790) ) ;
    buf_clk cell_2946 ( .C (clk), .D (signal_4795), .Q (signal_4796) ) ;
    buf_clk cell_2952 ( .C (clk), .D (signal_4801), .Q (signal_4802) ) ;
    buf_clk cell_2958 ( .C (clk), .D (signal_4807), .Q (signal_4808) ) ;
    buf_clk cell_2964 ( .C (clk), .D (signal_4813), .Q (signal_4814) ) ;
    buf_clk cell_2970 ( .C (clk), .D (signal_4819), .Q (signal_4820) ) ;
    buf_clk cell_2976 ( .C (clk), .D (signal_4825), .Q (signal_4826) ) ;
    buf_clk cell_2982 ( .C (clk), .D (signal_4831), .Q (signal_4832) ) ;
    buf_clk cell_2988 ( .C (clk), .D (signal_4837), .Q (signal_4838) ) ;
    buf_clk cell_2994 ( .C (clk), .D (signal_4843), .Q (signal_4844) ) ;
    buf_clk cell_3000 ( .C (clk), .D (signal_4849), .Q (signal_4850) ) ;
    buf_clk cell_3006 ( .C (clk), .D (signal_4855), .Q (signal_4856) ) ;
    buf_clk cell_3012 ( .C (clk), .D (signal_4861), .Q (signal_4862) ) ;
    buf_clk cell_3018 ( .C (clk), .D (signal_4867), .Q (signal_4868) ) ;
    buf_clk cell_3024 ( .C (clk), .D (signal_4873), .Q (signal_4874) ) ;
    buf_clk cell_3030 ( .C (clk), .D (signal_4879), .Q (signal_4880) ) ;
    buf_clk cell_3036 ( .C (clk), .D (signal_4885), .Q (signal_4886) ) ;
    buf_clk cell_3042 ( .C (clk), .D (signal_4891), .Q (signal_4892) ) ;
    buf_clk cell_3048 ( .C (clk), .D (signal_4897), .Q (signal_4898) ) ;
    buf_clk cell_3054 ( .C (clk), .D (signal_4903), .Q (signal_4904) ) ;
    buf_clk cell_3060 ( .C (clk), .D (signal_4909), .Q (signal_4910) ) ;
    buf_clk cell_3066 ( .C (clk), .D (signal_4915), .Q (signal_4916) ) ;
    buf_clk cell_3072 ( .C (clk), .D (signal_4921), .Q (signal_4922) ) ;
    buf_clk cell_3078 ( .C (clk), .D (signal_4927), .Q (signal_4928) ) ;
    buf_clk cell_3084 ( .C (clk), .D (signal_4933), .Q (signal_4934) ) ;
    buf_clk cell_3090 ( .C (clk), .D (signal_4939), .Q (signal_4940) ) ;
    buf_clk cell_3096 ( .C (clk), .D (signal_4945), .Q (signal_4946) ) ;
    buf_clk cell_3102 ( .C (clk), .D (signal_4951), .Q (signal_4952) ) ;
    buf_clk cell_3108 ( .C (clk), .D (signal_4957), .Q (signal_4958) ) ;
    buf_clk cell_3114 ( .C (clk), .D (signal_4963), .Q (signal_4964) ) ;
    buf_clk cell_3120 ( .C (clk), .D (signal_4969), .Q (signal_4970) ) ;
    buf_clk cell_3128 ( .C (clk), .D (signal_4977), .Q (signal_4978) ) ;
    buf_clk cell_3136 ( .C (clk), .D (signal_4985), .Q (signal_4986) ) ;
    buf_clk cell_3144 ( .C (clk), .D (signal_4993), .Q (signal_4994) ) ;
    buf_clk cell_3152 ( .C (clk), .D (signal_5001), .Q (signal_5002) ) ;
    buf_clk cell_3160 ( .C (clk), .D (signal_5009), .Q (signal_5010) ) ;
    buf_clk cell_3168 ( .C (clk), .D (signal_5017), .Q (signal_5018) ) ;
    buf_clk cell_3176 ( .C (clk), .D (signal_5025), .Q (signal_5026) ) ;
    buf_clk cell_3184 ( .C (clk), .D (signal_5033), .Q (signal_5034) ) ;
    buf_clk cell_3192 ( .C (clk), .D (signal_5041), .Q (signal_5042) ) ;
    buf_clk cell_3200 ( .C (clk), .D (signal_5049), .Q (signal_5050) ) ;
    buf_clk cell_3208 ( .C (clk), .D (signal_5057), .Q (signal_5058) ) ;
    buf_clk cell_3216 ( .C (clk), .D (signal_5065), .Q (signal_5066) ) ;
    buf_clk cell_3224 ( .C (clk), .D (signal_5073), .Q (signal_5074) ) ;
    buf_clk cell_3232 ( .C (clk), .D (signal_5081), .Q (signal_5082) ) ;
    buf_clk cell_3240 ( .C (clk), .D (signal_5089), .Q (signal_5090) ) ;
    buf_clk cell_3248 ( .C (clk), .D (signal_5097), .Q (signal_5098) ) ;
    buf_clk cell_3256 ( .C (clk), .D (signal_5105), .Q (signal_5106) ) ;
    buf_clk cell_3264 ( .C (clk), .D (signal_5113), .Q (signal_5114) ) ;
    buf_clk cell_3272 ( .C (clk), .D (signal_5121), .Q (signal_5122) ) ;
    buf_clk cell_3280 ( .C (clk), .D (signal_5129), .Q (signal_5130) ) ;
    buf_clk cell_3288 ( .C (clk), .D (signal_5137), .Q (signal_5138) ) ;
    buf_clk cell_3296 ( .C (clk), .D (signal_5145), .Q (signal_5146) ) ;
    buf_clk cell_3304 ( .C (clk), .D (signal_5153), .Q (signal_5154) ) ;
    buf_clk cell_3312 ( .C (clk), .D (signal_5161), .Q (signal_5162) ) ;
    buf_clk cell_3320 ( .C (clk), .D (signal_5169), .Q (signal_5170) ) ;
    buf_clk cell_3328 ( .C (clk), .D (signal_5177), .Q (signal_5178) ) ;
    buf_clk cell_3336 ( .C (clk), .D (signal_5185), .Q (signal_5186) ) ;
    buf_clk cell_3344 ( .C (clk), .D (signal_5193), .Q (signal_5194) ) ;
    buf_clk cell_3352 ( .C (clk), .D (signal_5201), .Q (signal_5202) ) ;
    buf_clk cell_3360 ( .C (clk), .D (signal_5209), .Q (signal_5210) ) ;
    buf_clk cell_3368 ( .C (clk), .D (signal_5217), .Q (signal_5218) ) ;
    buf_clk cell_3376 ( .C (clk), .D (signal_5225), .Q (signal_5226) ) ;
    buf_clk cell_3384 ( .C (clk), .D (signal_5233), .Q (signal_5234) ) ;
    buf_clk cell_3392 ( .C (clk), .D (signal_5241), .Q (signal_5242) ) ;
    buf_clk cell_3400 ( .C (clk), .D (signal_5249), .Q (signal_5250) ) ;
    buf_clk cell_3408 ( .C (clk), .D (signal_5257), .Q (signal_5258) ) ;
    buf_clk cell_3416 ( .C (clk), .D (signal_5265), .Q (signal_5266) ) ;
    buf_clk cell_3424 ( .C (clk), .D (signal_5273), .Q (signal_5274) ) ;
    buf_clk cell_3432 ( .C (clk), .D (signal_5281), .Q (signal_5282) ) ;
    buf_clk cell_3440 ( .C (clk), .D (signal_5289), .Q (signal_5290) ) ;
    buf_clk cell_3448 ( .C (clk), .D (signal_5297), .Q (signal_5298) ) ;
    buf_clk cell_3456 ( .C (clk), .D (signal_5305), .Q (signal_5306) ) ;
    buf_clk cell_3464 ( .C (clk), .D (signal_5313), .Q (signal_5314) ) ;
    buf_clk cell_3472 ( .C (clk), .D (signal_5321), .Q (signal_5322) ) ;
    buf_clk cell_3480 ( .C (clk), .D (signal_5329), .Q (signal_5330) ) ;
    buf_clk cell_3488 ( .C (clk), .D (signal_5337), .Q (signal_5338) ) ;
    buf_clk cell_3496 ( .C (clk), .D (signal_5345), .Q (signal_5346) ) ;
    buf_clk cell_3504 ( .C (clk), .D (signal_5353), .Q (signal_5354) ) ;
    buf_clk cell_3512 ( .C (clk), .D (signal_5361), .Q (signal_5362) ) ;
    buf_clk cell_3520 ( .C (clk), .D (signal_5369), .Q (signal_5370) ) ;
    buf_clk cell_3528 ( .C (clk), .D (signal_5377), .Q (signal_5378) ) ;
    buf_clk cell_3536 ( .C (clk), .D (signal_5385), .Q (signal_5386) ) ;
    buf_clk cell_3544 ( .C (clk), .D (signal_5393), .Q (signal_5394) ) ;
    buf_clk cell_3552 ( .C (clk), .D (signal_5401), .Q (signal_5402) ) ;
    buf_clk cell_3560 ( .C (clk), .D (signal_5409), .Q (signal_5410) ) ;
    buf_clk cell_3568 ( .C (clk), .D (signal_5417), .Q (signal_5418) ) ;
    buf_clk cell_3576 ( .C (clk), .D (signal_5425), .Q (signal_5426) ) ;
    buf_clk cell_3584 ( .C (clk), .D (signal_5433), .Q (signal_5434) ) ;
    buf_clk cell_3592 ( .C (clk), .D (signal_5441), .Q (signal_5442) ) ;
    buf_clk cell_3600 ( .C (clk), .D (signal_5449), .Q (signal_5450) ) ;
    buf_clk cell_3608 ( .C (clk), .D (signal_5457), .Q (signal_5458) ) ;
    buf_clk cell_3616 ( .C (clk), .D (signal_5465), .Q (signal_5466) ) ;
    buf_clk cell_3624 ( .C (clk), .D (signal_5473), .Q (signal_5474) ) ;
    buf_clk cell_3632 ( .C (clk), .D (signal_5481), .Q (signal_5482) ) ;
    buf_clk cell_3640 ( .C (clk), .D (signal_5489), .Q (signal_5490) ) ;
    buf_clk cell_3648 ( .C (clk), .D (signal_5497), .Q (signal_5498) ) ;
    buf_clk cell_3656 ( .C (clk), .D (signal_5505), .Q (signal_5506) ) ;
    buf_clk cell_3664 ( .C (clk), .D (signal_5513), .Q (signal_5514) ) ;
    buf_clk cell_3672 ( .C (clk), .D (signal_5521), .Q (signal_5522) ) ;
    buf_clk cell_3680 ( .C (clk), .D (signal_5529), .Q (signal_5530) ) ;
    buf_clk cell_3688 ( .C (clk), .D (signal_5537), .Q (signal_5538) ) ;
    buf_clk cell_3696 ( .C (clk), .D (signal_5545), .Q (signal_5546) ) ;
    buf_clk cell_3704 ( .C (clk), .D (signal_5553), .Q (signal_5554) ) ;
    buf_clk cell_3712 ( .C (clk), .D (signal_5561), .Q (signal_5562) ) ;
    buf_clk cell_3720 ( .C (clk), .D (signal_5569), .Q (signal_5570) ) ;
    buf_clk cell_3728 ( .C (clk), .D (signal_5577), .Q (signal_5578) ) ;
    buf_clk cell_3736 ( .C (clk), .D (signal_5585), .Q (signal_5586) ) ;
    buf_clk cell_3744 ( .C (clk), .D (signal_5593), .Q (signal_5594) ) ;
    buf_clk cell_3752 ( .C (clk), .D (signal_5601), .Q (signal_5602) ) ;
    buf_clk cell_3760 ( .C (clk), .D (signal_5609), .Q (signal_5610) ) ;
    buf_clk cell_3768 ( .C (clk), .D (signal_5617), .Q (signal_5618) ) ;
    buf_clk cell_3776 ( .C (clk), .D (signal_5625), .Q (signal_5626) ) ;
    buf_clk cell_3784 ( .C (clk), .D (signal_5633), .Q (signal_5634) ) ;
    buf_clk cell_3792 ( .C (clk), .D (signal_5641), .Q (signal_5642) ) ;
    buf_clk cell_3800 ( .C (clk), .D (signal_5649), .Q (signal_5650) ) ;
    buf_clk cell_3808 ( .C (clk), .D (signal_5657), .Q (signal_5658) ) ;
    buf_clk cell_3816 ( .C (clk), .D (signal_5665), .Q (signal_5666) ) ;
    buf_clk cell_3824 ( .C (clk), .D (signal_5673), .Q (signal_5674) ) ;
    buf_clk cell_3832 ( .C (clk), .D (signal_5681), .Q (signal_5682) ) ;
    buf_clk cell_3840 ( .C (clk), .D (signal_5689), .Q (signal_5690) ) ;
    buf_clk cell_3848 ( .C (clk), .D (signal_5697), .Q (signal_5698) ) ;
    buf_clk cell_3856 ( .C (clk), .D (signal_5705), .Q (signal_5706) ) ;
    buf_clk cell_3864 ( .C (clk), .D (signal_5713), .Q (signal_5714) ) ;
    buf_clk cell_3872 ( .C (clk), .D (signal_5721), .Q (signal_5722) ) ;
    buf_clk cell_3880 ( .C (clk), .D (signal_5729), .Q (signal_5730) ) ;
    buf_clk cell_3888 ( .C (clk), .D (signal_5737), .Q (signal_5738) ) ;
    buf_clk cell_3896 ( .C (clk), .D (signal_5745), .Q (signal_5746) ) ;
    buf_clk cell_3904 ( .C (clk), .D (signal_5753), .Q (signal_5754) ) ;
    buf_clk cell_3912 ( .C (clk), .D (signal_5761), .Q (signal_5762) ) ;
    buf_clk cell_3920 ( .C (clk), .D (signal_5769), .Q (signal_5770) ) ;
    buf_clk cell_3928 ( .C (clk), .D (signal_5777), .Q (signal_5778) ) ;
    buf_clk cell_3936 ( .C (clk), .D (signal_5785), .Q (signal_5786) ) ;
    buf_clk cell_3944 ( .C (clk), .D (signal_5793), .Q (signal_5794) ) ;
    buf_clk cell_3952 ( .C (clk), .D (signal_5801), .Q (signal_5802) ) ;
    buf_clk cell_3960 ( .C (clk), .D (signal_5809), .Q (signal_5810) ) ;
    buf_clk cell_3968 ( .C (clk), .D (signal_5817), .Q (signal_5818) ) ;
    buf_clk cell_3976 ( .C (clk), .D (signal_5825), .Q (signal_5826) ) ;
    buf_clk cell_3984 ( .C (clk), .D (signal_5833), .Q (signal_5834) ) ;
    buf_clk cell_3992 ( .C (clk), .D (signal_5841), .Q (signal_5842) ) ;
    buf_clk cell_4000 ( .C (clk), .D (signal_5849), .Q (signal_5850) ) ;
    buf_clk cell_4008 ( .C (clk), .D (signal_5857), .Q (signal_5858) ) ;
    buf_clk cell_4016 ( .C (clk), .D (signal_5865), .Q (signal_5866) ) ;
    buf_clk cell_4024 ( .C (clk), .D (signal_5873), .Q (signal_5874) ) ;
    buf_clk cell_4032 ( .C (clk), .D (signal_5881), .Q (signal_5882) ) ;
    buf_clk cell_4040 ( .C (clk), .D (signal_5889), .Q (signal_5890) ) ;
    buf_clk cell_4048 ( .C (clk), .D (signal_5897), .Q (signal_5898) ) ;
    buf_clk cell_4056 ( .C (clk), .D (signal_5905), .Q (signal_5906) ) ;
    buf_clk cell_4064 ( .C (clk), .D (signal_5913), .Q (signal_5914) ) ;
    buf_clk cell_4072 ( .C (clk), .D (signal_5921), .Q (signal_5922) ) ;
    buf_clk cell_4080 ( .C (clk), .D (signal_5929), .Q (signal_5930) ) ;
    buf_clk cell_4088 ( .C (clk), .D (signal_5937), .Q (signal_5938) ) ;
    buf_clk cell_4096 ( .C (clk), .D (signal_5945), .Q (signal_5946) ) ;
    buf_clk cell_4104 ( .C (clk), .D (signal_5953), .Q (signal_5954) ) ;
    buf_clk cell_4112 ( .C (clk), .D (signal_5961), .Q (signal_5962) ) ;
    buf_clk cell_4120 ( .C (clk), .D (signal_5969), .Q (signal_5970) ) ;
    buf_clk cell_4128 ( .C (clk), .D (signal_5977), .Q (signal_5978) ) ;
    buf_clk cell_4136 ( .C (clk), .D (signal_5985), .Q (signal_5986) ) ;
    buf_clk cell_4144 ( .C (clk), .D (signal_5993), .Q (signal_5994) ) ;
    buf_clk cell_4152 ( .C (clk), .D (signal_6001), .Q (signal_6002) ) ;
    buf_clk cell_4160 ( .C (clk), .D (signal_6009), .Q (signal_6010) ) ;
    buf_clk cell_4168 ( .C (clk), .D (signal_6017), .Q (signal_6018) ) ;
    buf_clk cell_4176 ( .C (clk), .D (signal_6025), .Q (signal_6026) ) ;
    buf_clk cell_4184 ( .C (clk), .D (signal_6033), .Q (signal_6034) ) ;
    buf_clk cell_4192 ( .C (clk), .D (signal_6041), .Q (signal_6042) ) ;
    buf_clk cell_4200 ( .C (clk), .D (signal_6049), .Q (signal_6050) ) ;
    buf_clk cell_4208 ( .C (clk), .D (signal_6057), .Q (signal_6058) ) ;
    buf_clk cell_4216 ( .C (clk), .D (signal_6065), .Q (signal_6066) ) ;
    buf_clk cell_4224 ( .C (clk), .D (signal_6073), .Q (signal_6074) ) ;
    buf_clk cell_4232 ( .C (clk), .D (signal_6081), .Q (signal_6082) ) ;
    buf_clk cell_4240 ( .C (clk), .D (signal_6089), .Q (signal_6090) ) ;
    buf_clk cell_4248 ( .C (clk), .D (signal_6097), .Q (signal_6098) ) ;
    buf_clk cell_4256 ( .C (clk), .D (signal_6105), .Q (signal_6106) ) ;
    buf_clk cell_4264 ( .C (clk), .D (signal_6113), .Q (signal_6114) ) ;
    buf_clk cell_4272 ( .C (clk), .D (signal_6121), .Q (signal_6122) ) ;
    buf_clk cell_4280 ( .C (clk), .D (signal_6129), .Q (signal_6130) ) ;
    buf_clk cell_4288 ( .C (clk), .D (signal_6137), .Q (signal_6138) ) ;
    buf_clk cell_4296 ( .C (clk), .D (signal_6145), .Q (signal_6146) ) ;
    buf_clk cell_4304 ( .C (clk), .D (signal_6153), .Q (signal_6154) ) ;
    buf_clk cell_4312 ( .C (clk), .D (signal_6161), .Q (signal_6162) ) ;
    buf_clk cell_4320 ( .C (clk), .D (signal_6169), .Q (signal_6170) ) ;
    buf_clk cell_4328 ( .C (clk), .D (signal_6177), .Q (signal_6178) ) ;
    buf_clk cell_4336 ( .C (clk), .D (signal_6185), .Q (signal_6186) ) ;
    buf_clk cell_4344 ( .C (clk), .D (signal_6193), .Q (signal_6194) ) ;
    buf_clk cell_4352 ( .C (clk), .D (signal_6201), .Q (signal_6202) ) ;
    buf_clk cell_4360 ( .C (clk), .D (signal_6209), .Q (signal_6210) ) ;
    buf_clk cell_4368 ( .C (clk), .D (signal_6217), .Q (signal_6218) ) ;
    buf_clk cell_4376 ( .C (clk), .D (signal_6225), .Q (signal_6226) ) ;
    buf_clk cell_4384 ( .C (clk), .D (signal_6233), .Q (signal_6234) ) ;
    buf_clk cell_4392 ( .C (clk), .D (signal_6241), .Q (signal_6242) ) ;
    buf_clk cell_4400 ( .C (clk), .D (signal_6249), .Q (signal_6250) ) ;
    buf_clk cell_4408 ( .C (clk), .D (signal_6257), .Q (signal_6258) ) ;
    buf_clk cell_4416 ( .C (clk), .D (signal_6265), .Q (signal_6266) ) ;
    buf_clk cell_4424 ( .C (clk), .D (signal_6273), .Q (signal_6274) ) ;
    buf_clk cell_4432 ( .C (clk), .D (signal_6281), .Q (signal_6282) ) ;
    buf_clk cell_4440 ( .C (clk), .D (signal_6289), .Q (signal_6290) ) ;
    buf_clk cell_4448 ( .C (clk), .D (signal_6297), .Q (signal_6298) ) ;
    buf_clk cell_4456 ( .C (clk), .D (signal_6305), .Q (signal_6306) ) ;
    buf_clk cell_4464 ( .C (clk), .D (signal_6313), .Q (signal_6314) ) ;
    buf_clk cell_4472 ( .C (clk), .D (signal_6321), .Q (signal_6322) ) ;
    buf_clk cell_4480 ( .C (clk), .D (signal_6329), .Q (signal_6330) ) ;
    buf_clk cell_4488 ( .C (clk), .D (signal_6337), .Q (signal_6338) ) ;
    buf_clk cell_4496 ( .C (clk), .D (signal_6345), .Q (signal_6346) ) ;
    buf_clk cell_4504 ( .C (clk), .D (signal_6353), .Q (signal_6354) ) ;
    buf_clk cell_4512 ( .C (clk), .D (signal_6361), .Q (signal_6362) ) ;
    buf_clk cell_4520 ( .C (clk), .D (signal_6369), .Q (signal_6370) ) ;
    buf_clk cell_4528 ( .C (clk), .D (signal_6377), .Q (signal_6378) ) ;
    buf_clk cell_4536 ( .C (clk), .D (signal_6385), .Q (signal_6386) ) ;
    buf_clk cell_4544 ( .C (clk), .D (signal_6393), .Q (signal_6394) ) ;
    buf_clk cell_4552 ( .C (clk), .D (signal_6401), .Q (signal_6402) ) ;
    buf_clk cell_4560 ( .C (clk), .D (signal_6409), .Q (signal_6410) ) ;
    buf_clk cell_4568 ( .C (clk), .D (signal_6417), .Q (signal_6418) ) ;
    buf_clk cell_4576 ( .C (clk), .D (signal_6425), .Q (signal_6426) ) ;
    buf_clk cell_4584 ( .C (clk), .D (signal_6433), .Q (signal_6434) ) ;
    buf_clk cell_4592 ( .C (clk), .D (signal_6441), .Q (signal_6442) ) ;
    buf_clk cell_4600 ( .C (clk), .D (signal_6449), .Q (signal_6450) ) ;
    buf_clk cell_4608 ( .C (clk), .D (signal_6457), .Q (signal_6458) ) ;
    buf_clk cell_4616 ( .C (clk), .D (signal_6465), .Q (signal_6466) ) ;
    buf_clk cell_4624 ( .C (clk), .D (signal_6473), .Q (signal_6474) ) ;
    buf_clk cell_4632 ( .C (clk), .D (signal_6481), .Q (signal_6482) ) ;
    buf_clk cell_4640 ( .C (clk), .D (signal_6489), .Q (signal_6490) ) ;
    buf_clk cell_4648 ( .C (clk), .D (signal_6497), .Q (signal_6498) ) ;
    buf_clk cell_4656 ( .C (clk), .D (signal_6505), .Q (signal_6506) ) ;
    buf_clk cell_4664 ( .C (clk), .D (signal_6513), .Q (signal_6514) ) ;
    buf_clk cell_4672 ( .C (clk), .D (signal_6521), .Q (signal_6522) ) ;
    buf_clk cell_4680 ( .C (clk), .D (signal_6529), .Q (signal_6530) ) ;
    buf_clk cell_4688 ( .C (clk), .D (signal_6537), .Q (signal_6538) ) ;
    buf_clk cell_4696 ( .C (clk), .D (signal_6545), .Q (signal_6546) ) ;
    buf_clk cell_4704 ( .C (clk), .D (signal_6553), .Q (signal_6554) ) ;
    buf_clk cell_4712 ( .C (clk), .D (signal_6561), .Q (signal_6562) ) ;
    buf_clk cell_4720 ( .C (clk), .D (signal_6569), .Q (signal_6570) ) ;
    buf_clk cell_4728 ( .C (clk), .D (signal_6577), .Q (signal_6578) ) ;
    buf_clk cell_4736 ( .C (clk), .D (signal_6585), .Q (signal_6586) ) ;
    buf_clk cell_4744 ( .C (clk), .D (signal_6593), .Q (signal_6594) ) ;
    buf_clk cell_4752 ( .C (clk), .D (signal_6601), .Q (signal_6602) ) ;
    buf_clk cell_4760 ( .C (clk), .D (signal_6609), .Q (signal_6610) ) ;
    buf_clk cell_4768 ( .C (clk), .D (signal_6617), .Q (signal_6618) ) ;
    buf_clk cell_4776 ( .C (clk), .D (signal_6625), .Q (signal_6626) ) ;
    buf_clk cell_4784 ( .C (clk), .D (signal_6633), .Q (signal_6634) ) ;
    buf_clk cell_4792 ( .C (clk), .D (signal_6641), .Q (signal_6642) ) ;
    buf_clk cell_4800 ( .C (clk), .D (signal_6649), .Q (signal_6650) ) ;
    buf_clk cell_4808 ( .C (clk), .D (signal_6657), .Q (signal_6658) ) ;
    buf_clk cell_4816 ( .C (clk), .D (signal_6665), .Q (signal_6666) ) ;
    buf_clk cell_4824 ( .C (clk), .D (signal_6673), .Q (signal_6674) ) ;
    buf_clk cell_4832 ( .C (clk), .D (signal_6681), .Q (signal_6682) ) ;
    buf_clk cell_4840 ( .C (clk), .D (signal_6689), .Q (signal_6690) ) ;
    buf_clk cell_4848 ( .C (clk), .D (signal_6697), .Q (signal_6698) ) ;
    buf_clk cell_4856 ( .C (clk), .D (signal_6705), .Q (signal_6706) ) ;
    buf_clk cell_4864 ( .C (clk), .D (signal_6713), .Q (signal_6714) ) ;
    buf_clk cell_4872 ( .C (clk), .D (signal_6721), .Q (signal_6722) ) ;
    buf_clk cell_4880 ( .C (clk), .D (signal_6729), .Q (signal_6730) ) ;
    buf_clk cell_4888 ( .C (clk), .D (signal_6737), .Q (signal_6738) ) ;
    buf_clk cell_4896 ( .C (clk), .D (signal_6745), .Q (signal_6746) ) ;
    buf_clk cell_4904 ( .C (clk), .D (signal_6753), .Q (signal_6754) ) ;
    buf_clk cell_4912 ( .C (clk), .D (signal_6761), .Q (signal_6762) ) ;
    buf_clk cell_4920 ( .C (clk), .D (signal_6769), .Q (signal_6770) ) ;
    buf_clk cell_4928 ( .C (clk), .D (signal_6777), .Q (signal_6778) ) ;
    buf_clk cell_4936 ( .C (clk), .D (signal_6785), .Q (signal_6786) ) ;
    buf_clk cell_4944 ( .C (clk), .D (signal_6793), .Q (signal_6794) ) ;
    buf_clk cell_4952 ( .C (clk), .D (signal_6801), .Q (signal_6802) ) ;
    buf_clk cell_4960 ( .C (clk), .D (signal_6809), .Q (signal_6810) ) ;
    buf_clk cell_4968 ( .C (clk), .D (signal_6817), .Q (signal_6818) ) ;
    buf_clk cell_4976 ( .C (clk), .D (signal_6825), .Q (signal_6826) ) ;
    buf_clk cell_4984 ( .C (clk), .D (signal_6833), .Q (signal_6834) ) ;
    buf_clk cell_4992 ( .C (clk), .D (signal_6841), .Q (signal_6842) ) ;
    buf_clk cell_5000 ( .C (clk), .D (signal_6849), .Q (signal_6850) ) ;
    buf_clk cell_5008 ( .C (clk), .D (signal_6857), .Q (signal_6858) ) ;
    buf_clk cell_5016 ( .C (clk), .D (signal_6865), .Q (signal_6866) ) ;
    buf_clk cell_5024 ( .C (clk), .D (signal_6873), .Q (signal_6874) ) ;
    buf_clk cell_5032 ( .C (clk), .D (signal_6881), .Q (signal_6882) ) ;
    buf_clk cell_5040 ( .C (clk), .D (signal_6889), .Q (signal_6890) ) ;
    buf_clk cell_5048 ( .C (clk), .D (signal_6897), .Q (signal_6898) ) ;
    buf_clk cell_5056 ( .C (clk), .D (signal_6905), .Q (signal_6906) ) ;
    buf_clk cell_5064 ( .C (clk), .D (signal_6913), .Q (signal_6914) ) ;
    buf_clk cell_5072 ( .C (clk), .D (signal_6921), .Q (signal_6922) ) ;
    buf_clk cell_5080 ( .C (clk), .D (signal_6929), .Q (signal_6930) ) ;
    buf_clk cell_5088 ( .C (clk), .D (signal_6937), .Q (signal_6938) ) ;
    buf_clk cell_5096 ( .C (clk), .D (signal_6945), .Q (signal_6946) ) ;
    buf_clk cell_5104 ( .C (clk), .D (signal_6953), .Q (signal_6954) ) ;
    buf_clk cell_5112 ( .C (clk), .D (signal_6961), .Q (signal_6962) ) ;
    buf_clk cell_5120 ( .C (clk), .D (signal_6969), .Q (signal_6970) ) ;
    buf_clk cell_5128 ( .C (clk), .D (signal_6977), .Q (signal_6978) ) ;
    buf_clk cell_5136 ( .C (clk), .D (signal_6985), .Q (signal_6986) ) ;
    buf_clk cell_5144 ( .C (clk), .D (signal_6993), .Q (signal_6994) ) ;
    buf_clk cell_5152 ( .C (clk), .D (signal_7001), .Q (signal_7002) ) ;
    buf_clk cell_5160 ( .C (clk), .D (signal_7009), .Q (signal_7010) ) ;
    buf_clk cell_5168 ( .C (clk), .D (signal_7017), .Q (signal_7018) ) ;
    buf_clk cell_5176 ( .C (clk), .D (signal_7025), .Q (signal_7026) ) ;
    buf_clk cell_5184 ( .C (clk), .D (signal_7033), .Q (signal_7034) ) ;
    buf_clk cell_5192 ( .C (clk), .D (signal_7041), .Q (signal_7042) ) ;
    buf_clk cell_5200 ( .C (clk), .D (signal_7049), .Q (signal_7050) ) ;
    buf_clk cell_5208 ( .C (clk), .D (signal_7057), .Q (signal_7058) ) ;
    buf_clk cell_5216 ( .C (clk), .D (signal_7065), .Q (signal_7066) ) ;
    buf_clk cell_5224 ( .C (clk), .D (signal_7073), .Q (signal_7074) ) ;
    buf_clk cell_5232 ( .C (clk), .D (signal_7081), .Q (signal_7082) ) ;
    buf_clk cell_5240 ( .C (clk), .D (signal_7089), .Q (signal_7090) ) ;
    buf_clk cell_5248 ( .C (clk), .D (signal_7097), .Q (signal_7098) ) ;
    buf_clk cell_5256 ( .C (clk), .D (signal_7105), .Q (signal_7106) ) ;
    buf_clk cell_5264 ( .C (clk), .D (signal_7113), .Q (signal_7114) ) ;
    buf_clk cell_5272 ( .C (clk), .D (signal_7121), .Q (signal_7122) ) ;
    buf_clk cell_5280 ( .C (clk), .D (signal_7129), .Q (signal_7130) ) ;
    buf_clk cell_5288 ( .C (clk), .D (signal_7137), .Q (signal_7138) ) ;
    buf_clk cell_5296 ( .C (clk), .D (signal_7145), .Q (signal_7146) ) ;
    buf_clk cell_5304 ( .C (clk), .D (signal_7153), .Q (signal_7154) ) ;
    buf_clk cell_5312 ( .C (clk), .D (signal_7161), .Q (signal_7162) ) ;
    buf_clk cell_5320 ( .C (clk), .D (signal_7169), .Q (signal_7170) ) ;
    buf_clk cell_5328 ( .C (clk), .D (signal_7177), .Q (signal_7178) ) ;
    buf_clk cell_5336 ( .C (clk), .D (signal_7185), .Q (signal_7186) ) ;
    buf_clk cell_5344 ( .C (clk), .D (signal_7193), .Q (signal_7194) ) ;
    buf_clk cell_5352 ( .C (clk), .D (signal_7201), .Q (signal_7202) ) ;
    buf_clk cell_5360 ( .C (clk), .D (signal_7209), .Q (signal_7210) ) ;
    buf_clk cell_5368 ( .C (clk), .D (signal_7217), .Q (signal_7218) ) ;
    buf_clk cell_5376 ( .C (clk), .D (signal_7225), .Q (signal_7226) ) ;
    buf_clk cell_5384 ( .C (clk), .D (signal_7233), .Q (signal_7234) ) ;
    buf_clk cell_5392 ( .C (clk), .D (signal_7241), .Q (signal_7242) ) ;
    buf_clk cell_5400 ( .C (clk), .D (signal_7249), .Q (signal_7250) ) ;
    buf_clk cell_5408 ( .C (clk), .D (signal_7257), .Q (signal_7258) ) ;
    buf_clk cell_5416 ( .C (clk), .D (signal_7265), .Q (signal_7266) ) ;
    buf_clk cell_5424 ( .C (clk), .D (signal_7273), .Q (signal_7274) ) ;
    buf_clk cell_5432 ( .C (clk), .D (signal_7281), .Q (signal_7282) ) ;
    buf_clk cell_5440 ( .C (clk), .D (signal_7289), .Q (signal_7290) ) ;
    buf_clk cell_5448 ( .C (clk), .D (signal_7297), .Q (signal_7298) ) ;
    buf_clk cell_5456 ( .C (clk), .D (signal_7305), .Q (signal_7306) ) ;
    buf_clk cell_5464 ( .C (clk), .D (signal_7313), .Q (signal_7314) ) ;
    buf_clk cell_5472 ( .C (clk), .D (signal_7321), .Q (signal_7322) ) ;
    buf_clk cell_5480 ( .C (clk), .D (signal_7329), .Q (signal_7330) ) ;
    buf_clk cell_5488 ( .C (clk), .D (signal_7337), .Q (signal_7338) ) ;
    buf_clk cell_5496 ( .C (clk), .D (signal_7345), .Q (signal_7346) ) ;
    buf_clk cell_5504 ( .C (clk), .D (signal_7353), .Q (signal_7354) ) ;
    buf_clk cell_5512 ( .C (clk), .D (signal_7361), .Q (signal_7362) ) ;
    buf_clk cell_5520 ( .C (clk), .D (signal_7369), .Q (signal_7370) ) ;
    buf_clk cell_5528 ( .C (clk), .D (signal_7377), .Q (signal_7378) ) ;
    buf_clk cell_5536 ( .C (clk), .D (signal_7385), .Q (signal_7386) ) ;
    buf_clk cell_5544 ( .C (clk), .D (signal_7393), .Q (signal_7394) ) ;
    buf_clk cell_5552 ( .C (clk), .D (signal_7401), .Q (signal_7402) ) ;
    buf_clk cell_5560 ( .C (clk), .D (signal_7409), .Q (signal_7410) ) ;
    buf_clk cell_5568 ( .C (clk), .D (signal_7417), .Q (signal_7418) ) ;
    buf_clk cell_5576 ( .C (clk), .D (signal_7425), .Q (signal_7426) ) ;
    buf_clk cell_5584 ( .C (clk), .D (signal_7433), .Q (signal_7434) ) ;
    buf_clk cell_5592 ( .C (clk), .D (signal_7441), .Q (signal_7442) ) ;
    buf_clk cell_5600 ( .C (clk), .D (signal_7449), .Q (signal_7450) ) ;
    buf_clk cell_5608 ( .C (clk), .D (signal_7457), .Q (signal_7458) ) ;
    buf_clk cell_5616 ( .C (clk), .D (signal_7465), .Q (signal_7466) ) ;
    buf_clk cell_5624 ( .C (clk), .D (signal_7473), .Q (signal_7474) ) ;
    buf_clk cell_5632 ( .C (clk), .D (signal_7481), .Q (signal_7482) ) ;
    buf_clk cell_5640 ( .C (clk), .D (signal_7489), .Q (signal_7490) ) ;
    buf_clk cell_5648 ( .C (clk), .D (signal_7497), .Q (signal_7498) ) ;
    buf_clk cell_5656 ( .C (clk), .D (signal_7505), .Q (signal_7506) ) ;
    buf_clk cell_5664 ( .C (clk), .D (signal_7513), .Q (signal_7514) ) ;
    buf_clk cell_5672 ( .C (clk), .D (signal_7521), .Q (signal_7522) ) ;
    buf_clk cell_5680 ( .C (clk), .D (signal_7529), .Q (signal_7530) ) ;
    buf_clk cell_5688 ( .C (clk), .D (signal_7537), .Q (signal_7538) ) ;
    buf_clk cell_5696 ( .C (clk), .D (signal_7545), .Q (signal_7546) ) ;
    buf_clk cell_5704 ( .C (clk), .D (signal_7553), .Q (signal_7554) ) ;
    buf_clk cell_5712 ( .C (clk), .D (signal_7561), .Q (signal_7562) ) ;
    buf_clk cell_5720 ( .C (clk), .D (signal_7569), .Q (signal_7570) ) ;
    buf_clk cell_5728 ( .C (clk), .D (signal_7577), .Q (signal_7578) ) ;
    buf_clk cell_5736 ( .C (clk), .D (signal_7585), .Q (signal_7586) ) ;
    buf_clk cell_5744 ( .C (clk), .D (signal_7593), .Q (signal_7594) ) ;
    buf_clk cell_5752 ( .C (clk), .D (signal_7601), .Q (signal_7602) ) ;
    buf_clk cell_5760 ( .C (clk), .D (signal_7609), .Q (signal_7610) ) ;
    buf_clk cell_5768 ( .C (clk), .D (signal_7617), .Q (signal_7618) ) ;
    buf_clk cell_5776 ( .C (clk), .D (signal_7625), .Q (signal_7626) ) ;
    buf_clk cell_5784 ( .C (clk), .D (signal_7633), .Q (signal_7634) ) ;
    buf_clk cell_5792 ( .C (clk), .D (signal_7641), .Q (signal_7642) ) ;
    buf_clk cell_5800 ( .C (clk), .D (signal_7649), .Q (signal_7650) ) ;
    buf_clk cell_5808 ( .C (clk), .D (signal_7657), .Q (signal_7658) ) ;
    buf_clk cell_5816 ( .C (clk), .D (signal_7665), .Q (signal_7666) ) ;
    buf_clk cell_5824 ( .C (clk), .D (signal_7673), .Q (signal_7674) ) ;
    buf_clk cell_5832 ( .C (clk), .D (signal_7681), .Q (signal_7682) ) ;
    buf_clk cell_5840 ( .C (clk), .D (signal_7689), .Q (signal_7690) ) ;
    buf_clk cell_5848 ( .C (clk), .D (signal_7697), .Q (signal_7698) ) ;
    buf_clk cell_5856 ( .C (clk), .D (signal_7705), .Q (signal_7706) ) ;
    buf_clk cell_5864 ( .C (clk), .D (signal_7713), .Q (signal_7714) ) ;
    buf_clk cell_5872 ( .C (clk), .D (signal_7721), .Q (signal_7722) ) ;
    buf_clk cell_5880 ( .C (clk), .D (signal_7729), .Q (signal_7730) ) ;
    buf_clk cell_5888 ( .C (clk), .D (signal_7737), .Q (signal_7738) ) ;
    buf_clk cell_5896 ( .C (clk), .D (signal_7745), .Q (signal_7746) ) ;
    buf_clk cell_5904 ( .C (clk), .D (signal_7753), .Q (signal_7754) ) ;
    buf_clk cell_5912 ( .C (clk), .D (signal_7761), .Q (signal_7762) ) ;
    buf_clk cell_5920 ( .C (clk), .D (signal_7769), .Q (signal_7770) ) ;
    buf_clk cell_5928 ( .C (clk), .D (signal_7777), .Q (signal_7778) ) ;
    buf_clk cell_5936 ( .C (clk), .D (signal_7785), .Q (signal_7786) ) ;
    buf_clk cell_5944 ( .C (clk), .D (signal_7793), .Q (signal_7794) ) ;
    buf_clk cell_5952 ( .C (clk), .D (signal_7801), .Q (signal_7802) ) ;
    buf_clk cell_5960 ( .C (clk), .D (signal_7809), .Q (signal_7810) ) ;
    buf_clk cell_5968 ( .C (clk), .D (signal_7817), .Q (signal_7818) ) ;
    buf_clk cell_5976 ( .C (clk), .D (signal_7825), .Q (signal_7826) ) ;
    buf_clk cell_5984 ( .C (clk), .D (signal_7833), .Q (signal_7834) ) ;
    buf_clk cell_5992 ( .C (clk), .D (signal_7841), .Q (signal_7842) ) ;
    buf_clk cell_6000 ( .C (clk), .D (signal_7849), .Q (signal_7850) ) ;
    buf_clk cell_6008 ( .C (clk), .D (signal_7857), .Q (signal_7858) ) ;
    buf_clk cell_6016 ( .C (clk), .D (signal_7865), .Q (signal_7866) ) ;
    buf_clk cell_6024 ( .C (clk), .D (signal_7873), .Q (signal_7874) ) ;
    buf_clk cell_6032 ( .C (clk), .D (signal_7881), .Q (signal_7882) ) ;
    buf_clk cell_6040 ( .C (clk), .D (signal_7889), .Q (signal_7890) ) ;
    buf_clk cell_6048 ( .C (clk), .D (signal_7897), .Q (signal_7898) ) ;
    buf_clk cell_6056 ( .C (clk), .D (signal_7905), .Q (signal_7906) ) ;
    buf_clk cell_6064 ( .C (clk), .D (signal_7913), .Q (signal_7914) ) ;
    buf_clk cell_6072 ( .C (clk), .D (signal_7921), .Q (signal_7922) ) ;
    buf_clk cell_6080 ( .C (clk), .D (signal_7929), .Q (signal_7930) ) ;
    buf_clk cell_6088 ( .C (clk), .D (signal_7937), .Q (signal_7938) ) ;
    buf_clk cell_6096 ( .C (clk), .D (signal_7945), .Q (signal_7946) ) ;
    buf_clk cell_6104 ( .C (clk), .D (signal_7953), .Q (signal_7954) ) ;
    buf_clk cell_6112 ( .C (clk), .D (signal_7961), .Q (signal_7962) ) ;
    buf_clk cell_6120 ( .C (clk), .D (signal_7969), .Q (signal_7970) ) ;
    buf_clk cell_6128 ( .C (clk), .D (signal_7977), .Q (signal_7978) ) ;
    buf_clk cell_6136 ( .C (clk), .D (signal_7985), .Q (signal_7986) ) ;
    buf_clk cell_6144 ( .C (clk), .D (signal_7993), .Q (signal_7994) ) ;
    buf_clk cell_6152 ( .C (clk), .D (signal_8001), .Q (signal_8002) ) ;
    buf_clk cell_6160 ( .C (clk), .D (signal_8009), .Q (signal_8010) ) ;
    buf_clk cell_6168 ( .C (clk), .D (signal_8017), .Q (signal_8018) ) ;
    buf_clk cell_6176 ( .C (clk), .D (signal_8025), .Q (signal_8026) ) ;
    buf_clk cell_6184 ( .C (clk), .D (signal_8033), .Q (signal_8034) ) ;
    buf_clk cell_6192 ( .C (clk), .D (signal_8041), .Q (signal_8042) ) ;
    buf_clk cell_6200 ( .C (clk), .D (signal_8049), .Q (signal_8050) ) ;
    buf_clk cell_6208 ( .C (clk), .D (signal_8057), .Q (signal_8058) ) ;
    buf_clk cell_6216 ( .C (clk), .D (signal_8065), .Q (signal_8066) ) ;
    buf_clk cell_6224 ( .C (clk), .D (signal_8073), .Q (signal_8074) ) ;
    buf_clk cell_6232 ( .C (clk), .D (signal_8081), .Q (signal_8082) ) ;
    buf_clk cell_6240 ( .C (clk), .D (signal_8089), .Q (signal_8090) ) ;
    buf_clk cell_6248 ( .C (clk), .D (signal_8097), .Q (signal_8098) ) ;
    buf_clk cell_6256 ( .C (clk), .D (signal_8105), .Q (signal_8106) ) ;
    buf_clk cell_6264 ( .C (clk), .D (signal_8113), .Q (signal_8114) ) ;
    buf_clk cell_6272 ( .C (clk), .D (signal_8121), .Q (signal_8122) ) ;
    buf_clk cell_6280 ( .C (clk), .D (signal_8129), .Q (signal_8130) ) ;
    buf_clk cell_6288 ( .C (clk), .D (signal_8137), .Q (signal_8138) ) ;
    buf_clk cell_6296 ( .C (clk), .D (signal_8145), .Q (signal_8146) ) ;
    buf_clk cell_6304 ( .C (clk), .D (signal_8153), .Q (signal_8154) ) ;
    buf_clk cell_6312 ( .C (clk), .D (signal_8161), .Q (signal_8162) ) ;
    buf_clk cell_6320 ( .C (clk), .D (signal_8169), .Q (signal_8170) ) ;
    buf_clk cell_6328 ( .C (clk), .D (signal_8177), .Q (signal_8178) ) ;
    buf_clk cell_6336 ( .C (clk), .D (signal_8185), .Q (signal_8186) ) ;
    buf_clk cell_6344 ( .C (clk), .D (signal_8193), .Q (signal_8194) ) ;
    buf_clk cell_6352 ( .C (clk), .D (signal_8201), .Q (signal_8202) ) ;
    buf_clk cell_6360 ( .C (clk), .D (signal_8209), .Q (signal_8210) ) ;
    buf_clk cell_6368 ( .C (clk), .D (signal_8217), .Q (signal_8218) ) ;
    buf_clk cell_6376 ( .C (clk), .D (signal_8225), .Q (signal_8226) ) ;
    buf_clk cell_6384 ( .C (clk), .D (signal_8233), .Q (signal_8234) ) ;
    buf_clk cell_6392 ( .C (clk), .D (signal_8241), .Q (signal_8242) ) ;
    buf_clk cell_6400 ( .C (clk), .D (signal_8249), .Q (signal_8250) ) ;
    buf_clk cell_6408 ( .C (clk), .D (signal_8257), .Q (signal_8258) ) ;
    buf_clk cell_6416 ( .C (clk), .D (signal_8265), .Q (signal_8266) ) ;
    buf_clk cell_6424 ( .C (clk), .D (signal_8273), .Q (signal_8274) ) ;
    buf_clk cell_6432 ( .C (clk), .D (signal_8281), .Q (signal_8282) ) ;
    buf_clk cell_6440 ( .C (clk), .D (signal_8289), .Q (signal_8290) ) ;
    buf_clk cell_6448 ( .C (clk), .D (signal_8297), .Q (signal_8298) ) ;
    buf_clk cell_6456 ( .C (clk), .D (signal_8305), .Q (signal_8306) ) ;
    buf_clk cell_6464 ( .C (clk), .D (signal_8313), .Q (signal_8314) ) ;
    buf_clk cell_6472 ( .C (clk), .D (signal_8321), .Q (signal_8322) ) ;
    buf_clk cell_6480 ( .C (clk), .D (signal_8329), .Q (signal_8330) ) ;
    buf_clk cell_6488 ( .C (clk), .D (signal_8337), .Q (signal_8338) ) ;
    buf_clk cell_6496 ( .C (clk), .D (signal_8345), .Q (signal_8346) ) ;
    buf_clk cell_6504 ( .C (clk), .D (signal_8353), .Q (signal_8354) ) ;
    buf_clk cell_6512 ( .C (clk), .D (signal_8361), .Q (signal_8362) ) ;
    buf_clk cell_6520 ( .C (clk), .D (signal_8369), .Q (signal_8370) ) ;
    buf_clk cell_6528 ( .C (clk), .D (signal_8377), .Q (signal_8378) ) ;
    buf_clk cell_6536 ( .C (clk), .D (signal_8385), .Q (signal_8386) ) ;
    buf_clk cell_6544 ( .C (clk), .D (signal_8393), .Q (signal_8394) ) ;
    buf_clk cell_6552 ( .C (clk), .D (signal_8401), .Q (signal_8402) ) ;
    buf_clk cell_6560 ( .C (clk), .D (signal_8409), .Q (signal_8410) ) ;
    buf_clk cell_6568 ( .C (clk), .D (signal_8417), .Q (signal_8418) ) ;
    buf_clk cell_6576 ( .C (clk), .D (signal_8425), .Q (signal_8426) ) ;
    buf_clk cell_6584 ( .C (clk), .D (signal_8433), .Q (signal_8434) ) ;
    buf_clk cell_6592 ( .C (clk), .D (signal_8441), .Q (signal_8442) ) ;
    buf_clk cell_6600 ( .C (clk), .D (signal_8449), .Q (signal_8450) ) ;
    buf_clk cell_6608 ( .C (clk), .D (signal_8457), .Q (signal_8458) ) ;
    buf_clk cell_6616 ( .C (clk), .D (signal_8465), .Q (signal_8466) ) ;
    buf_clk cell_6624 ( .C (clk), .D (signal_8473), .Q (signal_8474) ) ;
    buf_clk cell_6632 ( .C (clk), .D (signal_8481), .Q (signal_8482) ) ;
    buf_clk cell_6640 ( .C (clk), .D (signal_8489), .Q (signal_8490) ) ;
    buf_clk cell_6648 ( .C (clk), .D (signal_8497), .Q (signal_8498) ) ;
    buf_clk cell_6656 ( .C (clk), .D (signal_8505), .Q (signal_8506) ) ;
    buf_clk cell_6664 ( .C (clk), .D (signal_8513), .Q (signal_8514) ) ;
    buf_clk cell_6672 ( .C (clk), .D (signal_8521), .Q (signal_8522) ) ;
    buf_clk cell_6680 ( .C (clk), .D (signal_8529), .Q (signal_8530) ) ;
    buf_clk cell_6688 ( .C (clk), .D (signal_8537), .Q (signal_8538) ) ;
    buf_clk cell_6696 ( .C (clk), .D (signal_8545), .Q (signal_8546) ) ;
    buf_clk cell_6704 ( .C (clk), .D (signal_8553), .Q (signal_8554) ) ;
    buf_clk cell_6712 ( .C (clk), .D (signal_8561), .Q (signal_8562) ) ;
    buf_clk cell_6720 ( .C (clk), .D (signal_8569), .Q (signal_8570) ) ;
    buf_clk cell_6728 ( .C (clk), .D (signal_8577), .Q (signal_8578) ) ;
    buf_clk cell_6736 ( .C (clk), .D (signal_8585), .Q (signal_8586) ) ;
    buf_clk cell_6744 ( .C (clk), .D (signal_8593), .Q (signal_8594) ) ;
    buf_clk cell_6752 ( .C (clk), .D (signal_8601), .Q (signal_8602) ) ;
    buf_clk cell_6760 ( .C (clk), .D (signal_8609), .Q (signal_8610) ) ;
    buf_clk cell_6768 ( .C (clk), .D (signal_8617), .Q (signal_8618) ) ;
    buf_clk cell_6776 ( .C (clk), .D (signal_8625), .Q (signal_8626) ) ;
    buf_clk cell_6784 ( .C (clk), .D (signal_8633), .Q (signal_8634) ) ;
    buf_clk cell_6792 ( .C (clk), .D (signal_8641), .Q (signal_8642) ) ;
    buf_clk cell_6800 ( .C (clk), .D (signal_8649), .Q (signal_8650) ) ;
    buf_clk cell_6808 ( .C (clk), .D (signal_8657), .Q (signal_8658) ) ;
    buf_clk cell_6816 ( .C (clk), .D (signal_8665), .Q (signal_8666) ) ;
    buf_clk cell_6824 ( .C (clk), .D (signal_8673), .Q (signal_8674) ) ;
    buf_clk cell_6832 ( .C (clk), .D (signal_8681), .Q (signal_8682) ) ;
    buf_clk cell_6840 ( .C (clk), .D (signal_8689), .Q (signal_8690) ) ;
    buf_clk cell_6848 ( .C (clk), .D (signal_8697), .Q (signal_8698) ) ;
    buf_clk cell_6856 ( .C (clk), .D (signal_8705), .Q (signal_8706) ) ;
    buf_clk cell_6864 ( .C (clk), .D (signal_8713), .Q (signal_8714) ) ;
    buf_clk cell_6872 ( .C (clk), .D (signal_8721), .Q (signal_8722) ) ;
    buf_clk cell_6880 ( .C (clk), .D (signal_8729), .Q (signal_8730) ) ;
    buf_clk cell_6888 ( .C (clk), .D (signal_8737), .Q (signal_8738) ) ;
    buf_clk cell_6896 ( .C (clk), .D (signal_8745), .Q (signal_8746) ) ;
    buf_clk cell_6904 ( .C (clk), .D (signal_8753), .Q (signal_8754) ) ;
    buf_clk cell_6912 ( .C (clk), .D (signal_8761), .Q (signal_8762) ) ;
    buf_clk cell_6920 ( .C (clk), .D (signal_8769), .Q (signal_8770) ) ;
    buf_clk cell_6928 ( .C (clk), .D (signal_8777), .Q (signal_8778) ) ;
    buf_clk cell_6936 ( .C (clk), .D (signal_8785), .Q (signal_8786) ) ;
    buf_clk cell_6944 ( .C (clk), .D (signal_8793), .Q (signal_8794) ) ;
    buf_clk cell_6952 ( .C (clk), .D (signal_8801), .Q (signal_8802) ) ;
    buf_clk cell_6960 ( .C (clk), .D (signal_8809), .Q (signal_8810) ) ;
    buf_clk cell_6968 ( .C (clk), .D (signal_8817), .Q (signal_8818) ) ;
    buf_clk cell_6976 ( .C (clk), .D (signal_8825), .Q (signal_8826) ) ;
    buf_clk cell_6984 ( .C (clk), .D (signal_8833), .Q (signal_8834) ) ;
    buf_clk cell_6992 ( .C (clk), .D (signal_8841), .Q (signal_8842) ) ;
    buf_clk cell_7000 ( .C (clk), .D (signal_8849), .Q (signal_8850) ) ;
    buf_clk cell_7008 ( .C (clk), .D (signal_8857), .Q (signal_8858) ) ;
    buf_clk cell_7016 ( .C (clk), .D (signal_8865), .Q (signal_8866) ) ;
    buf_clk cell_7024 ( .C (clk), .D (signal_8873), .Q (signal_8874) ) ;
    buf_clk cell_7032 ( .C (clk), .D (signal_8881), .Q (signal_8882) ) ;
    buf_clk cell_7040 ( .C (clk), .D (signal_8889), .Q (signal_8890) ) ;
    buf_clk cell_7048 ( .C (clk), .D (signal_8897), .Q (signal_8898) ) ;
    buf_clk cell_7056 ( .C (clk), .D (signal_8905), .Q (signal_8906) ) ;
    buf_clk cell_7064 ( .C (clk), .D (signal_8913), .Q (signal_8914) ) ;
    buf_clk cell_7072 ( .C (clk), .D (signal_8921), .Q (signal_8922) ) ;
    buf_clk cell_7080 ( .C (clk), .D (signal_8929), .Q (signal_8930) ) ;
    buf_clk cell_7088 ( .C (clk), .D (signal_8937), .Q (signal_8938) ) ;
    buf_clk cell_7096 ( .C (clk), .D (signal_8945), .Q (signal_8946) ) ;

    /* cells in depth 4 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1763 ( .a ({signal_3496, signal_2028}), .b ({signal_3498, signal_2030}), .clk (clk), .r (Fresh[9]), .c ({signal_3507, signal_2031}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1764 ( .a ({signal_3497, signal_2029}), .b ({signal_3498, signal_2030}), .clk (clk), .r (Fresh[10]), .c ({signal_3508, signal_2032}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1767 ( .a ({signal_3496, signal_2028}), .b ({signal_3509, signal_2033}), .clk (clk), .r (Fresh[11]), .c ({signal_3511, signal_2035}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1769 ( .a ({signal_3715, signal_3713}), .b ({signal_3507, signal_2031}), .c ({signal_3513, signal_2037}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1770 ( .a ({signal_3719, signal_3717}), .b ({signal_3507, signal_2031}), .c ({signal_3514, signal_2038}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1771 ( .a ({signal_3507, signal_2031}), .b ({signal_3723, signal_3721}), .c ({signal_3515, signal_2039}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1776 ( .a ({signal_3507, signal_2031}), .b ({signal_3727, signal_3725}), .c ({signal_3520, signal_2044}) ) ;
    buf_clk cell_1863 ( .C (clk), .D (signal_3712), .Q (signal_3713) ) ;
    buf_clk cell_1865 ( .C (clk), .D (signal_3714), .Q (signal_3715) ) ;
    buf_clk cell_1867 ( .C (clk), .D (signal_3716), .Q (signal_3717) ) ;
    buf_clk cell_1869 ( .C (clk), .D (signal_3718), .Q (signal_3719) ) ;
    buf_clk cell_1871 ( .C (clk), .D (signal_3720), .Q (signal_3721) ) ;
    buf_clk cell_1873 ( .C (clk), .D (signal_3722), .Q (signal_3723) ) ;
    buf_clk cell_1875 ( .C (clk), .D (signal_3724), .Q (signal_3725) ) ;
    buf_clk cell_1877 ( .C (clk), .D (signal_3726), .Q (signal_3727) ) ;
    buf_clk cell_1897 ( .C (clk), .D (signal_3746), .Q (signal_3747) ) ;
    buf_clk cell_1905 ( .C (clk), .D (signal_3754), .Q (signal_3755) ) ;
    buf_clk cell_1913 ( .C (clk), .D (signal_3762), .Q (signal_3763) ) ;
    buf_clk cell_1921 ( .C (clk), .D (signal_3770), .Q (signal_3771) ) ;
    buf_clk cell_1929 ( .C (clk), .D (signal_3778), .Q (signal_3779) ) ;
    buf_clk cell_1937 ( .C (clk), .D (signal_3786), .Q (signal_3787) ) ;
    buf_clk cell_1945 ( .C (clk), .D (signal_3794), .Q (signal_3795) ) ;
    buf_clk cell_1953 ( .C (clk), .D (signal_3802), .Q (signal_3803) ) ;
    buf_clk cell_1961 ( .C (clk), .D (signal_3810), .Q (signal_3811) ) ;
    buf_clk cell_1969 ( .C (clk), .D (signal_3818), .Q (signal_3819) ) ;
    buf_clk cell_1977 ( .C (clk), .D (signal_3826), .Q (signal_3827) ) ;
    buf_clk cell_1985 ( .C (clk), .D (signal_3834), .Q (signal_3835) ) ;
    buf_clk cell_1993 ( .C (clk), .D (signal_3842), .Q (signal_3843) ) ;
    buf_clk cell_2001 ( .C (clk), .D (signal_3850), .Q (signal_3851) ) ;
    buf_clk cell_2009 ( .C (clk), .D (signal_3858), .Q (signal_3859) ) ;
    buf_clk cell_2017 ( .C (clk), .D (signal_3866), .Q (signal_3867) ) ;
    buf_clk cell_2025 ( .C (clk), .D (signal_3874), .Q (signal_3875) ) ;
    buf_clk cell_2033 ( .C (clk), .D (signal_3882), .Q (signal_3883) ) ;
    buf_clk cell_2041 ( .C (clk), .D (signal_3890), .Q (signal_3891) ) ;
    buf_clk cell_2049 ( .C (clk), .D (signal_3898), .Q (signal_3899) ) ;
    buf_clk cell_2057 ( .C (clk), .D (signal_3906), .Q (signal_3907) ) ;
    buf_clk cell_2065 ( .C (clk), .D (signal_3914), .Q (signal_3915) ) ;
    buf_clk cell_2073 ( .C (clk), .D (signal_3922), .Q (signal_3923) ) ;
    buf_clk cell_2081 ( .C (clk), .D (signal_3930), .Q (signal_3931) ) ;
    buf_clk cell_2089 ( .C (clk), .D (signal_3938), .Q (signal_3939) ) ;
    buf_clk cell_2097 ( .C (clk), .D (signal_3946), .Q (signal_3947) ) ;
    buf_clk cell_2105 ( .C (clk), .D (signal_3954), .Q (signal_3955) ) ;
    buf_clk cell_2113 ( .C (clk), .D (signal_3962), .Q (signal_3963) ) ;
    buf_clk cell_2121 ( .C (clk), .D (signal_3970), .Q (signal_3971) ) ;
    buf_clk cell_2129 ( .C (clk), .D (signal_3978), .Q (signal_3979) ) ;
    buf_clk cell_2137 ( .C (clk), .D (signal_3986), .Q (signal_3987) ) ;
    buf_clk cell_2145 ( .C (clk), .D (signal_3994), .Q (signal_3995) ) ;
    buf_clk cell_2153 ( .C (clk), .D (signal_4002), .Q (signal_4003) ) ;
    buf_clk cell_2161 ( .C (clk), .D (signal_4010), .Q (signal_4011) ) ;
    buf_clk cell_2169 ( .C (clk), .D (signal_4018), .Q (signal_4019) ) ;
    buf_clk cell_2177 ( .C (clk), .D (signal_4026), .Q (signal_4027) ) ;
    buf_clk cell_2185 ( .C (clk), .D (signal_4034), .Q (signal_4035) ) ;
    buf_clk cell_2193 ( .C (clk), .D (signal_4042), .Q (signal_4043) ) ;
    buf_clk cell_2201 ( .C (clk), .D (signal_4050), .Q (signal_4051) ) ;
    buf_clk cell_2209 ( .C (clk), .D (signal_4058), .Q (signal_4059) ) ;
    buf_clk cell_2217 ( .C (clk), .D (signal_4066), .Q (signal_4067) ) ;
    buf_clk cell_2225 ( .C (clk), .D (signal_4074), .Q (signal_4075) ) ;
    buf_clk cell_2233 ( .C (clk), .D (signal_4082), .Q (signal_4083) ) ;
    buf_clk cell_2241 ( .C (clk), .D (signal_4090), .Q (signal_4091) ) ;
    buf_clk cell_2249 ( .C (clk), .D (signal_4098), .Q (signal_4099) ) ;
    buf_clk cell_2257 ( .C (clk), .D (signal_4106), .Q (signal_4107) ) ;
    buf_clk cell_2265 ( .C (clk), .D (signal_4114), .Q (signal_4115) ) ;
    buf_clk cell_2273 ( .C (clk), .D (signal_4122), .Q (signal_4123) ) ;
    buf_clk cell_2281 ( .C (clk), .D (signal_4130), .Q (signal_4131) ) ;
    buf_clk cell_2289 ( .C (clk), .D (signal_4138), .Q (signal_4139) ) ;
    buf_clk cell_2297 ( .C (clk), .D (signal_4146), .Q (signal_4147) ) ;
    buf_clk cell_2305 ( .C (clk), .D (signal_4154), .Q (signal_4155) ) ;
    buf_clk cell_2313 ( .C (clk), .D (signal_4162), .Q (signal_4163) ) ;
    buf_clk cell_2321 ( .C (clk), .D (signal_4170), .Q (signal_4171) ) ;
    buf_clk cell_2329 ( .C (clk), .D (signal_4178), .Q (signal_4179) ) ;
    buf_clk cell_2337 ( .C (clk), .D (signal_4186), .Q (signal_4187) ) ;
    buf_clk cell_2345 ( .C (clk), .D (signal_4194), .Q (signal_4195) ) ;
    buf_clk cell_2353 ( .C (clk), .D (signal_4202), .Q (signal_4203) ) ;
    buf_clk cell_2361 ( .C (clk), .D (signal_4210), .Q (signal_4211) ) ;
    buf_clk cell_2369 ( .C (clk), .D (signal_4218), .Q (signal_4219) ) ;
    buf_clk cell_2377 ( .C (clk), .D (signal_4226), .Q (signal_4227) ) ;
    buf_clk cell_2385 ( .C (clk), .D (signal_4234), .Q (signal_4235) ) ;
    buf_clk cell_2393 ( .C (clk), .D (signal_4242), .Q (signal_4243) ) ;
    buf_clk cell_2401 ( .C (clk), .D (signal_4250), .Q (signal_4251) ) ;
    buf_clk cell_2409 ( .C (clk), .D (signal_4258), .Q (signal_4259) ) ;
    buf_clk cell_2417 ( .C (clk), .D (signal_4266), .Q (signal_4267) ) ;
    buf_clk cell_2425 ( .C (clk), .D (signal_4274), .Q (signal_4275) ) ;
    buf_clk cell_2433 ( .C (clk), .D (signal_4282), .Q (signal_4283) ) ;
    buf_clk cell_2441 ( .C (clk), .D (signal_4290), .Q (signal_4291) ) ;
    buf_clk cell_2449 ( .C (clk), .D (signal_4298), .Q (signal_4299) ) ;
    buf_clk cell_2457 ( .C (clk), .D (signal_4306), .Q (signal_4307) ) ;
    buf_clk cell_2465 ( .C (clk), .D (signal_4314), .Q (signal_4315) ) ;
    buf_clk cell_2473 ( .C (clk), .D (signal_4322), .Q (signal_4323) ) ;
    buf_clk cell_2481 ( .C (clk), .D (signal_4330), .Q (signal_4331) ) ;
    buf_clk cell_2489 ( .C (clk), .D (signal_4338), .Q (signal_4339) ) ;
    buf_clk cell_2497 ( .C (clk), .D (signal_4346), .Q (signal_4347) ) ;
    buf_clk cell_2505 ( .C (clk), .D (signal_4354), .Q (signal_4355) ) ;
    buf_clk cell_2513 ( .C (clk), .D (signal_4362), .Q (signal_4363) ) ;
    buf_clk cell_2521 ( .C (clk), .D (signal_4370), .Q (signal_4371) ) ;
    buf_clk cell_2529 ( .C (clk), .D (signal_4378), .Q (signal_4379) ) ;
    buf_clk cell_2537 ( .C (clk), .D (signal_4386), .Q (signal_4387) ) ;
    buf_clk cell_2545 ( .C (clk), .D (signal_4394), .Q (signal_4395) ) ;
    buf_clk cell_2553 ( .C (clk), .D (signal_4402), .Q (signal_4403) ) ;
    buf_clk cell_2561 ( .C (clk), .D (signal_4410), .Q (signal_4411) ) ;
    buf_clk cell_2569 ( .C (clk), .D (signal_4418), .Q (signal_4419) ) ;
    buf_clk cell_2577 ( .C (clk), .D (signal_4426), .Q (signal_4427) ) ;
    buf_clk cell_2585 ( .C (clk), .D (signal_4434), .Q (signal_4435) ) ;
    buf_clk cell_2593 ( .C (clk), .D (signal_4442), .Q (signal_4443) ) ;
    buf_clk cell_2601 ( .C (clk), .D (signal_4450), .Q (signal_4451) ) ;
    buf_clk cell_2609 ( .C (clk), .D (signal_4458), .Q (signal_4459) ) ;
    buf_clk cell_2617 ( .C (clk), .D (signal_4466), .Q (signal_4467) ) ;
    buf_clk cell_2625 ( .C (clk), .D (signal_4474), .Q (signal_4475) ) ;
    buf_clk cell_2633 ( .C (clk), .D (signal_4482), .Q (signal_4483) ) ;
    buf_clk cell_2641 ( .C (clk), .D (signal_4490), .Q (signal_4491) ) ;
    buf_clk cell_2649 ( .C (clk), .D (signal_4498), .Q (signal_4499) ) ;
    buf_clk cell_2657 ( .C (clk), .D (signal_4506), .Q (signal_4507) ) ;
    buf_clk cell_2665 ( .C (clk), .D (signal_4514), .Q (signal_4515) ) ;
    buf_clk cell_2673 ( .C (clk), .D (signal_4522), .Q (signal_4523) ) ;
    buf_clk cell_2681 ( .C (clk), .D (signal_4530), .Q (signal_4531) ) ;
    buf_clk cell_2689 ( .C (clk), .D (signal_4538), .Q (signal_4539) ) ;
    buf_clk cell_2697 ( .C (clk), .D (signal_4546), .Q (signal_4547) ) ;
    buf_clk cell_2705 ( .C (clk), .D (signal_4554), .Q (signal_4555) ) ;
    buf_clk cell_2713 ( .C (clk), .D (signal_4562), .Q (signal_4563) ) ;
    buf_clk cell_2721 ( .C (clk), .D (signal_4570), .Q (signal_4571) ) ;
    buf_clk cell_2729 ( .C (clk), .D (signal_4578), .Q (signal_4579) ) ;
    buf_clk cell_2737 ( .C (clk), .D (signal_4586), .Q (signal_4587) ) ;
    buf_clk cell_2745 ( .C (clk), .D (signal_4594), .Q (signal_4595) ) ;
    buf_clk cell_2753 ( .C (clk), .D (signal_4602), .Q (signal_4603) ) ;
    buf_clk cell_2761 ( .C (clk), .D (signal_4610), .Q (signal_4611) ) ;
    buf_clk cell_2769 ( .C (clk), .D (signal_4618), .Q (signal_4619) ) ;
    buf_clk cell_2777 ( .C (clk), .D (signal_4626), .Q (signal_4627) ) ;
    buf_clk cell_2785 ( .C (clk), .D (signal_4634), .Q (signal_4635) ) ;
    buf_clk cell_2793 ( .C (clk), .D (signal_4642), .Q (signal_4643) ) ;
    buf_clk cell_2801 ( .C (clk), .D (signal_4650), .Q (signal_4651) ) ;
    buf_clk cell_2809 ( .C (clk), .D (signal_4658), .Q (signal_4659) ) ;
    buf_clk cell_2817 ( .C (clk), .D (signal_4666), .Q (signal_4667) ) ;
    buf_clk cell_2825 ( .C (clk), .D (signal_4674), .Q (signal_4675) ) ;
    buf_clk cell_2833 ( .C (clk), .D (signal_4682), .Q (signal_4683) ) ;
    buf_clk cell_2841 ( .C (clk), .D (signal_4690), .Q (signal_4691) ) ;
    buf_clk cell_2849 ( .C (clk), .D (signal_4698), .Q (signal_4699) ) ;
    buf_clk cell_2857 ( .C (clk), .D (signal_4706), .Q (signal_4707) ) ;
    buf_clk cell_2865 ( .C (clk), .D (signal_4714), .Q (signal_4715) ) ;
    buf_clk cell_2873 ( .C (clk), .D (signal_4722), .Q (signal_4723) ) ;
    buf_clk cell_2881 ( .C (clk), .D (signal_4730), .Q (signal_4731) ) ;
    buf_clk cell_2889 ( .C (clk), .D (signal_4738), .Q (signal_4739) ) ;
    buf_clk cell_2897 ( .C (clk), .D (signal_4746), .Q (signal_4747) ) ;
    buf_clk cell_2905 ( .C (clk), .D (signal_4754), .Q (signal_4755) ) ;
    buf_clk cell_2911 ( .C (clk), .D (signal_4760), .Q (signal_4761) ) ;
    buf_clk cell_2917 ( .C (clk), .D (signal_4766), .Q (signal_4767) ) ;
    buf_clk cell_2923 ( .C (clk), .D (signal_4772), .Q (signal_4773) ) ;
    buf_clk cell_2929 ( .C (clk), .D (signal_4778), .Q (signal_4779) ) ;
    buf_clk cell_2935 ( .C (clk), .D (signal_4784), .Q (signal_4785) ) ;
    buf_clk cell_2941 ( .C (clk), .D (signal_4790), .Q (signal_4791) ) ;
    buf_clk cell_2947 ( .C (clk), .D (signal_4796), .Q (signal_4797) ) ;
    buf_clk cell_2953 ( .C (clk), .D (signal_4802), .Q (signal_4803) ) ;
    buf_clk cell_2959 ( .C (clk), .D (signal_4808), .Q (signal_4809) ) ;
    buf_clk cell_2965 ( .C (clk), .D (signal_4814), .Q (signal_4815) ) ;
    buf_clk cell_2971 ( .C (clk), .D (signal_4820), .Q (signal_4821) ) ;
    buf_clk cell_2977 ( .C (clk), .D (signal_4826), .Q (signal_4827) ) ;
    buf_clk cell_2983 ( .C (clk), .D (signal_4832), .Q (signal_4833) ) ;
    buf_clk cell_2989 ( .C (clk), .D (signal_4838), .Q (signal_4839) ) ;
    buf_clk cell_2995 ( .C (clk), .D (signal_4844), .Q (signal_4845) ) ;
    buf_clk cell_3001 ( .C (clk), .D (signal_4850), .Q (signal_4851) ) ;
    buf_clk cell_3007 ( .C (clk), .D (signal_4856), .Q (signal_4857) ) ;
    buf_clk cell_3013 ( .C (clk), .D (signal_4862), .Q (signal_4863) ) ;
    buf_clk cell_3019 ( .C (clk), .D (signal_4868), .Q (signal_4869) ) ;
    buf_clk cell_3025 ( .C (clk), .D (signal_4874), .Q (signal_4875) ) ;
    buf_clk cell_3031 ( .C (clk), .D (signal_4880), .Q (signal_4881) ) ;
    buf_clk cell_3037 ( .C (clk), .D (signal_4886), .Q (signal_4887) ) ;
    buf_clk cell_3043 ( .C (clk), .D (signal_4892), .Q (signal_4893) ) ;
    buf_clk cell_3049 ( .C (clk), .D (signal_4898), .Q (signal_4899) ) ;
    buf_clk cell_3055 ( .C (clk), .D (signal_4904), .Q (signal_4905) ) ;
    buf_clk cell_3061 ( .C (clk), .D (signal_4910), .Q (signal_4911) ) ;
    buf_clk cell_3067 ( .C (clk), .D (signal_4916), .Q (signal_4917) ) ;
    buf_clk cell_3073 ( .C (clk), .D (signal_4922), .Q (signal_4923) ) ;
    buf_clk cell_3079 ( .C (clk), .D (signal_4928), .Q (signal_4929) ) ;
    buf_clk cell_3085 ( .C (clk), .D (signal_4934), .Q (signal_4935) ) ;
    buf_clk cell_3091 ( .C (clk), .D (signal_4940), .Q (signal_4941) ) ;
    buf_clk cell_3097 ( .C (clk), .D (signal_4946), .Q (signal_4947) ) ;
    buf_clk cell_3103 ( .C (clk), .D (signal_4952), .Q (signal_4953) ) ;
    buf_clk cell_3109 ( .C (clk), .D (signal_4958), .Q (signal_4959) ) ;
    buf_clk cell_3115 ( .C (clk), .D (signal_4964), .Q (signal_4965) ) ;
    buf_clk cell_3121 ( .C (clk), .D (signal_4970), .Q (signal_4971) ) ;
    buf_clk cell_3129 ( .C (clk), .D (signal_4978), .Q (signal_4979) ) ;
    buf_clk cell_3137 ( .C (clk), .D (signal_4986), .Q (signal_4987) ) ;
    buf_clk cell_3145 ( .C (clk), .D (signal_4994), .Q (signal_4995) ) ;
    buf_clk cell_3153 ( .C (clk), .D (signal_5002), .Q (signal_5003) ) ;
    buf_clk cell_3161 ( .C (clk), .D (signal_5010), .Q (signal_5011) ) ;
    buf_clk cell_3169 ( .C (clk), .D (signal_5018), .Q (signal_5019) ) ;
    buf_clk cell_3177 ( .C (clk), .D (signal_5026), .Q (signal_5027) ) ;
    buf_clk cell_3185 ( .C (clk), .D (signal_5034), .Q (signal_5035) ) ;
    buf_clk cell_3193 ( .C (clk), .D (signal_5042), .Q (signal_5043) ) ;
    buf_clk cell_3201 ( .C (clk), .D (signal_5050), .Q (signal_5051) ) ;
    buf_clk cell_3209 ( .C (clk), .D (signal_5058), .Q (signal_5059) ) ;
    buf_clk cell_3217 ( .C (clk), .D (signal_5066), .Q (signal_5067) ) ;
    buf_clk cell_3225 ( .C (clk), .D (signal_5074), .Q (signal_5075) ) ;
    buf_clk cell_3233 ( .C (clk), .D (signal_5082), .Q (signal_5083) ) ;
    buf_clk cell_3241 ( .C (clk), .D (signal_5090), .Q (signal_5091) ) ;
    buf_clk cell_3249 ( .C (clk), .D (signal_5098), .Q (signal_5099) ) ;
    buf_clk cell_3257 ( .C (clk), .D (signal_5106), .Q (signal_5107) ) ;
    buf_clk cell_3265 ( .C (clk), .D (signal_5114), .Q (signal_5115) ) ;
    buf_clk cell_3273 ( .C (clk), .D (signal_5122), .Q (signal_5123) ) ;
    buf_clk cell_3281 ( .C (clk), .D (signal_5130), .Q (signal_5131) ) ;
    buf_clk cell_3289 ( .C (clk), .D (signal_5138), .Q (signal_5139) ) ;
    buf_clk cell_3297 ( .C (clk), .D (signal_5146), .Q (signal_5147) ) ;
    buf_clk cell_3305 ( .C (clk), .D (signal_5154), .Q (signal_5155) ) ;
    buf_clk cell_3313 ( .C (clk), .D (signal_5162), .Q (signal_5163) ) ;
    buf_clk cell_3321 ( .C (clk), .D (signal_5170), .Q (signal_5171) ) ;
    buf_clk cell_3329 ( .C (clk), .D (signal_5178), .Q (signal_5179) ) ;
    buf_clk cell_3337 ( .C (clk), .D (signal_5186), .Q (signal_5187) ) ;
    buf_clk cell_3345 ( .C (clk), .D (signal_5194), .Q (signal_5195) ) ;
    buf_clk cell_3353 ( .C (clk), .D (signal_5202), .Q (signal_5203) ) ;
    buf_clk cell_3361 ( .C (clk), .D (signal_5210), .Q (signal_5211) ) ;
    buf_clk cell_3369 ( .C (clk), .D (signal_5218), .Q (signal_5219) ) ;
    buf_clk cell_3377 ( .C (clk), .D (signal_5226), .Q (signal_5227) ) ;
    buf_clk cell_3385 ( .C (clk), .D (signal_5234), .Q (signal_5235) ) ;
    buf_clk cell_3393 ( .C (clk), .D (signal_5242), .Q (signal_5243) ) ;
    buf_clk cell_3401 ( .C (clk), .D (signal_5250), .Q (signal_5251) ) ;
    buf_clk cell_3409 ( .C (clk), .D (signal_5258), .Q (signal_5259) ) ;
    buf_clk cell_3417 ( .C (clk), .D (signal_5266), .Q (signal_5267) ) ;
    buf_clk cell_3425 ( .C (clk), .D (signal_5274), .Q (signal_5275) ) ;
    buf_clk cell_3433 ( .C (clk), .D (signal_5282), .Q (signal_5283) ) ;
    buf_clk cell_3441 ( .C (clk), .D (signal_5290), .Q (signal_5291) ) ;
    buf_clk cell_3449 ( .C (clk), .D (signal_5298), .Q (signal_5299) ) ;
    buf_clk cell_3457 ( .C (clk), .D (signal_5306), .Q (signal_5307) ) ;
    buf_clk cell_3465 ( .C (clk), .D (signal_5314), .Q (signal_5315) ) ;
    buf_clk cell_3473 ( .C (clk), .D (signal_5322), .Q (signal_5323) ) ;
    buf_clk cell_3481 ( .C (clk), .D (signal_5330), .Q (signal_5331) ) ;
    buf_clk cell_3489 ( .C (clk), .D (signal_5338), .Q (signal_5339) ) ;
    buf_clk cell_3497 ( .C (clk), .D (signal_5346), .Q (signal_5347) ) ;
    buf_clk cell_3505 ( .C (clk), .D (signal_5354), .Q (signal_5355) ) ;
    buf_clk cell_3513 ( .C (clk), .D (signal_5362), .Q (signal_5363) ) ;
    buf_clk cell_3521 ( .C (clk), .D (signal_5370), .Q (signal_5371) ) ;
    buf_clk cell_3529 ( .C (clk), .D (signal_5378), .Q (signal_5379) ) ;
    buf_clk cell_3537 ( .C (clk), .D (signal_5386), .Q (signal_5387) ) ;
    buf_clk cell_3545 ( .C (clk), .D (signal_5394), .Q (signal_5395) ) ;
    buf_clk cell_3553 ( .C (clk), .D (signal_5402), .Q (signal_5403) ) ;
    buf_clk cell_3561 ( .C (clk), .D (signal_5410), .Q (signal_5411) ) ;
    buf_clk cell_3569 ( .C (clk), .D (signal_5418), .Q (signal_5419) ) ;
    buf_clk cell_3577 ( .C (clk), .D (signal_5426), .Q (signal_5427) ) ;
    buf_clk cell_3585 ( .C (clk), .D (signal_5434), .Q (signal_5435) ) ;
    buf_clk cell_3593 ( .C (clk), .D (signal_5442), .Q (signal_5443) ) ;
    buf_clk cell_3601 ( .C (clk), .D (signal_5450), .Q (signal_5451) ) ;
    buf_clk cell_3609 ( .C (clk), .D (signal_5458), .Q (signal_5459) ) ;
    buf_clk cell_3617 ( .C (clk), .D (signal_5466), .Q (signal_5467) ) ;
    buf_clk cell_3625 ( .C (clk), .D (signal_5474), .Q (signal_5475) ) ;
    buf_clk cell_3633 ( .C (clk), .D (signal_5482), .Q (signal_5483) ) ;
    buf_clk cell_3641 ( .C (clk), .D (signal_5490), .Q (signal_5491) ) ;
    buf_clk cell_3649 ( .C (clk), .D (signal_5498), .Q (signal_5499) ) ;
    buf_clk cell_3657 ( .C (clk), .D (signal_5506), .Q (signal_5507) ) ;
    buf_clk cell_3665 ( .C (clk), .D (signal_5514), .Q (signal_5515) ) ;
    buf_clk cell_3673 ( .C (clk), .D (signal_5522), .Q (signal_5523) ) ;
    buf_clk cell_3681 ( .C (clk), .D (signal_5530), .Q (signal_5531) ) ;
    buf_clk cell_3689 ( .C (clk), .D (signal_5538), .Q (signal_5539) ) ;
    buf_clk cell_3697 ( .C (clk), .D (signal_5546), .Q (signal_5547) ) ;
    buf_clk cell_3705 ( .C (clk), .D (signal_5554), .Q (signal_5555) ) ;
    buf_clk cell_3713 ( .C (clk), .D (signal_5562), .Q (signal_5563) ) ;
    buf_clk cell_3721 ( .C (clk), .D (signal_5570), .Q (signal_5571) ) ;
    buf_clk cell_3729 ( .C (clk), .D (signal_5578), .Q (signal_5579) ) ;
    buf_clk cell_3737 ( .C (clk), .D (signal_5586), .Q (signal_5587) ) ;
    buf_clk cell_3745 ( .C (clk), .D (signal_5594), .Q (signal_5595) ) ;
    buf_clk cell_3753 ( .C (clk), .D (signal_5602), .Q (signal_5603) ) ;
    buf_clk cell_3761 ( .C (clk), .D (signal_5610), .Q (signal_5611) ) ;
    buf_clk cell_3769 ( .C (clk), .D (signal_5618), .Q (signal_5619) ) ;
    buf_clk cell_3777 ( .C (clk), .D (signal_5626), .Q (signal_5627) ) ;
    buf_clk cell_3785 ( .C (clk), .D (signal_5634), .Q (signal_5635) ) ;
    buf_clk cell_3793 ( .C (clk), .D (signal_5642), .Q (signal_5643) ) ;
    buf_clk cell_3801 ( .C (clk), .D (signal_5650), .Q (signal_5651) ) ;
    buf_clk cell_3809 ( .C (clk), .D (signal_5658), .Q (signal_5659) ) ;
    buf_clk cell_3817 ( .C (clk), .D (signal_5666), .Q (signal_5667) ) ;
    buf_clk cell_3825 ( .C (clk), .D (signal_5674), .Q (signal_5675) ) ;
    buf_clk cell_3833 ( .C (clk), .D (signal_5682), .Q (signal_5683) ) ;
    buf_clk cell_3841 ( .C (clk), .D (signal_5690), .Q (signal_5691) ) ;
    buf_clk cell_3849 ( .C (clk), .D (signal_5698), .Q (signal_5699) ) ;
    buf_clk cell_3857 ( .C (clk), .D (signal_5706), .Q (signal_5707) ) ;
    buf_clk cell_3865 ( .C (clk), .D (signal_5714), .Q (signal_5715) ) ;
    buf_clk cell_3873 ( .C (clk), .D (signal_5722), .Q (signal_5723) ) ;
    buf_clk cell_3881 ( .C (clk), .D (signal_5730), .Q (signal_5731) ) ;
    buf_clk cell_3889 ( .C (clk), .D (signal_5738), .Q (signal_5739) ) ;
    buf_clk cell_3897 ( .C (clk), .D (signal_5746), .Q (signal_5747) ) ;
    buf_clk cell_3905 ( .C (clk), .D (signal_5754), .Q (signal_5755) ) ;
    buf_clk cell_3913 ( .C (clk), .D (signal_5762), .Q (signal_5763) ) ;
    buf_clk cell_3921 ( .C (clk), .D (signal_5770), .Q (signal_5771) ) ;
    buf_clk cell_3929 ( .C (clk), .D (signal_5778), .Q (signal_5779) ) ;
    buf_clk cell_3937 ( .C (clk), .D (signal_5786), .Q (signal_5787) ) ;
    buf_clk cell_3945 ( .C (clk), .D (signal_5794), .Q (signal_5795) ) ;
    buf_clk cell_3953 ( .C (clk), .D (signal_5802), .Q (signal_5803) ) ;
    buf_clk cell_3961 ( .C (clk), .D (signal_5810), .Q (signal_5811) ) ;
    buf_clk cell_3969 ( .C (clk), .D (signal_5818), .Q (signal_5819) ) ;
    buf_clk cell_3977 ( .C (clk), .D (signal_5826), .Q (signal_5827) ) ;
    buf_clk cell_3985 ( .C (clk), .D (signal_5834), .Q (signal_5835) ) ;
    buf_clk cell_3993 ( .C (clk), .D (signal_5842), .Q (signal_5843) ) ;
    buf_clk cell_4001 ( .C (clk), .D (signal_5850), .Q (signal_5851) ) ;
    buf_clk cell_4009 ( .C (clk), .D (signal_5858), .Q (signal_5859) ) ;
    buf_clk cell_4017 ( .C (clk), .D (signal_5866), .Q (signal_5867) ) ;
    buf_clk cell_4025 ( .C (clk), .D (signal_5874), .Q (signal_5875) ) ;
    buf_clk cell_4033 ( .C (clk), .D (signal_5882), .Q (signal_5883) ) ;
    buf_clk cell_4041 ( .C (clk), .D (signal_5890), .Q (signal_5891) ) ;
    buf_clk cell_4049 ( .C (clk), .D (signal_5898), .Q (signal_5899) ) ;
    buf_clk cell_4057 ( .C (clk), .D (signal_5906), .Q (signal_5907) ) ;
    buf_clk cell_4065 ( .C (clk), .D (signal_5914), .Q (signal_5915) ) ;
    buf_clk cell_4073 ( .C (clk), .D (signal_5922), .Q (signal_5923) ) ;
    buf_clk cell_4081 ( .C (clk), .D (signal_5930), .Q (signal_5931) ) ;
    buf_clk cell_4089 ( .C (clk), .D (signal_5938), .Q (signal_5939) ) ;
    buf_clk cell_4097 ( .C (clk), .D (signal_5946), .Q (signal_5947) ) ;
    buf_clk cell_4105 ( .C (clk), .D (signal_5954), .Q (signal_5955) ) ;
    buf_clk cell_4113 ( .C (clk), .D (signal_5962), .Q (signal_5963) ) ;
    buf_clk cell_4121 ( .C (clk), .D (signal_5970), .Q (signal_5971) ) ;
    buf_clk cell_4129 ( .C (clk), .D (signal_5978), .Q (signal_5979) ) ;
    buf_clk cell_4137 ( .C (clk), .D (signal_5986), .Q (signal_5987) ) ;
    buf_clk cell_4145 ( .C (clk), .D (signal_5994), .Q (signal_5995) ) ;
    buf_clk cell_4153 ( .C (clk), .D (signal_6002), .Q (signal_6003) ) ;
    buf_clk cell_4161 ( .C (clk), .D (signal_6010), .Q (signal_6011) ) ;
    buf_clk cell_4169 ( .C (clk), .D (signal_6018), .Q (signal_6019) ) ;
    buf_clk cell_4177 ( .C (clk), .D (signal_6026), .Q (signal_6027) ) ;
    buf_clk cell_4185 ( .C (clk), .D (signal_6034), .Q (signal_6035) ) ;
    buf_clk cell_4193 ( .C (clk), .D (signal_6042), .Q (signal_6043) ) ;
    buf_clk cell_4201 ( .C (clk), .D (signal_6050), .Q (signal_6051) ) ;
    buf_clk cell_4209 ( .C (clk), .D (signal_6058), .Q (signal_6059) ) ;
    buf_clk cell_4217 ( .C (clk), .D (signal_6066), .Q (signal_6067) ) ;
    buf_clk cell_4225 ( .C (clk), .D (signal_6074), .Q (signal_6075) ) ;
    buf_clk cell_4233 ( .C (clk), .D (signal_6082), .Q (signal_6083) ) ;
    buf_clk cell_4241 ( .C (clk), .D (signal_6090), .Q (signal_6091) ) ;
    buf_clk cell_4249 ( .C (clk), .D (signal_6098), .Q (signal_6099) ) ;
    buf_clk cell_4257 ( .C (clk), .D (signal_6106), .Q (signal_6107) ) ;
    buf_clk cell_4265 ( .C (clk), .D (signal_6114), .Q (signal_6115) ) ;
    buf_clk cell_4273 ( .C (clk), .D (signal_6122), .Q (signal_6123) ) ;
    buf_clk cell_4281 ( .C (clk), .D (signal_6130), .Q (signal_6131) ) ;
    buf_clk cell_4289 ( .C (clk), .D (signal_6138), .Q (signal_6139) ) ;
    buf_clk cell_4297 ( .C (clk), .D (signal_6146), .Q (signal_6147) ) ;
    buf_clk cell_4305 ( .C (clk), .D (signal_6154), .Q (signal_6155) ) ;
    buf_clk cell_4313 ( .C (clk), .D (signal_6162), .Q (signal_6163) ) ;
    buf_clk cell_4321 ( .C (clk), .D (signal_6170), .Q (signal_6171) ) ;
    buf_clk cell_4329 ( .C (clk), .D (signal_6178), .Q (signal_6179) ) ;
    buf_clk cell_4337 ( .C (clk), .D (signal_6186), .Q (signal_6187) ) ;
    buf_clk cell_4345 ( .C (clk), .D (signal_6194), .Q (signal_6195) ) ;
    buf_clk cell_4353 ( .C (clk), .D (signal_6202), .Q (signal_6203) ) ;
    buf_clk cell_4361 ( .C (clk), .D (signal_6210), .Q (signal_6211) ) ;
    buf_clk cell_4369 ( .C (clk), .D (signal_6218), .Q (signal_6219) ) ;
    buf_clk cell_4377 ( .C (clk), .D (signal_6226), .Q (signal_6227) ) ;
    buf_clk cell_4385 ( .C (clk), .D (signal_6234), .Q (signal_6235) ) ;
    buf_clk cell_4393 ( .C (clk), .D (signal_6242), .Q (signal_6243) ) ;
    buf_clk cell_4401 ( .C (clk), .D (signal_6250), .Q (signal_6251) ) ;
    buf_clk cell_4409 ( .C (clk), .D (signal_6258), .Q (signal_6259) ) ;
    buf_clk cell_4417 ( .C (clk), .D (signal_6266), .Q (signal_6267) ) ;
    buf_clk cell_4425 ( .C (clk), .D (signal_6274), .Q (signal_6275) ) ;
    buf_clk cell_4433 ( .C (clk), .D (signal_6282), .Q (signal_6283) ) ;
    buf_clk cell_4441 ( .C (clk), .D (signal_6290), .Q (signal_6291) ) ;
    buf_clk cell_4449 ( .C (clk), .D (signal_6298), .Q (signal_6299) ) ;
    buf_clk cell_4457 ( .C (clk), .D (signal_6306), .Q (signal_6307) ) ;
    buf_clk cell_4465 ( .C (clk), .D (signal_6314), .Q (signal_6315) ) ;
    buf_clk cell_4473 ( .C (clk), .D (signal_6322), .Q (signal_6323) ) ;
    buf_clk cell_4481 ( .C (clk), .D (signal_6330), .Q (signal_6331) ) ;
    buf_clk cell_4489 ( .C (clk), .D (signal_6338), .Q (signal_6339) ) ;
    buf_clk cell_4497 ( .C (clk), .D (signal_6346), .Q (signal_6347) ) ;
    buf_clk cell_4505 ( .C (clk), .D (signal_6354), .Q (signal_6355) ) ;
    buf_clk cell_4513 ( .C (clk), .D (signal_6362), .Q (signal_6363) ) ;
    buf_clk cell_4521 ( .C (clk), .D (signal_6370), .Q (signal_6371) ) ;
    buf_clk cell_4529 ( .C (clk), .D (signal_6378), .Q (signal_6379) ) ;
    buf_clk cell_4537 ( .C (clk), .D (signal_6386), .Q (signal_6387) ) ;
    buf_clk cell_4545 ( .C (clk), .D (signal_6394), .Q (signal_6395) ) ;
    buf_clk cell_4553 ( .C (clk), .D (signal_6402), .Q (signal_6403) ) ;
    buf_clk cell_4561 ( .C (clk), .D (signal_6410), .Q (signal_6411) ) ;
    buf_clk cell_4569 ( .C (clk), .D (signal_6418), .Q (signal_6419) ) ;
    buf_clk cell_4577 ( .C (clk), .D (signal_6426), .Q (signal_6427) ) ;
    buf_clk cell_4585 ( .C (clk), .D (signal_6434), .Q (signal_6435) ) ;
    buf_clk cell_4593 ( .C (clk), .D (signal_6442), .Q (signal_6443) ) ;
    buf_clk cell_4601 ( .C (clk), .D (signal_6450), .Q (signal_6451) ) ;
    buf_clk cell_4609 ( .C (clk), .D (signal_6458), .Q (signal_6459) ) ;
    buf_clk cell_4617 ( .C (clk), .D (signal_6466), .Q (signal_6467) ) ;
    buf_clk cell_4625 ( .C (clk), .D (signal_6474), .Q (signal_6475) ) ;
    buf_clk cell_4633 ( .C (clk), .D (signal_6482), .Q (signal_6483) ) ;
    buf_clk cell_4641 ( .C (clk), .D (signal_6490), .Q (signal_6491) ) ;
    buf_clk cell_4649 ( .C (clk), .D (signal_6498), .Q (signal_6499) ) ;
    buf_clk cell_4657 ( .C (clk), .D (signal_6506), .Q (signal_6507) ) ;
    buf_clk cell_4665 ( .C (clk), .D (signal_6514), .Q (signal_6515) ) ;
    buf_clk cell_4673 ( .C (clk), .D (signal_6522), .Q (signal_6523) ) ;
    buf_clk cell_4681 ( .C (clk), .D (signal_6530), .Q (signal_6531) ) ;
    buf_clk cell_4689 ( .C (clk), .D (signal_6538), .Q (signal_6539) ) ;
    buf_clk cell_4697 ( .C (clk), .D (signal_6546), .Q (signal_6547) ) ;
    buf_clk cell_4705 ( .C (clk), .D (signal_6554), .Q (signal_6555) ) ;
    buf_clk cell_4713 ( .C (clk), .D (signal_6562), .Q (signal_6563) ) ;
    buf_clk cell_4721 ( .C (clk), .D (signal_6570), .Q (signal_6571) ) ;
    buf_clk cell_4729 ( .C (clk), .D (signal_6578), .Q (signal_6579) ) ;
    buf_clk cell_4737 ( .C (clk), .D (signal_6586), .Q (signal_6587) ) ;
    buf_clk cell_4745 ( .C (clk), .D (signal_6594), .Q (signal_6595) ) ;
    buf_clk cell_4753 ( .C (clk), .D (signal_6602), .Q (signal_6603) ) ;
    buf_clk cell_4761 ( .C (clk), .D (signal_6610), .Q (signal_6611) ) ;
    buf_clk cell_4769 ( .C (clk), .D (signal_6618), .Q (signal_6619) ) ;
    buf_clk cell_4777 ( .C (clk), .D (signal_6626), .Q (signal_6627) ) ;
    buf_clk cell_4785 ( .C (clk), .D (signal_6634), .Q (signal_6635) ) ;
    buf_clk cell_4793 ( .C (clk), .D (signal_6642), .Q (signal_6643) ) ;
    buf_clk cell_4801 ( .C (clk), .D (signal_6650), .Q (signal_6651) ) ;
    buf_clk cell_4809 ( .C (clk), .D (signal_6658), .Q (signal_6659) ) ;
    buf_clk cell_4817 ( .C (clk), .D (signal_6666), .Q (signal_6667) ) ;
    buf_clk cell_4825 ( .C (clk), .D (signal_6674), .Q (signal_6675) ) ;
    buf_clk cell_4833 ( .C (clk), .D (signal_6682), .Q (signal_6683) ) ;
    buf_clk cell_4841 ( .C (clk), .D (signal_6690), .Q (signal_6691) ) ;
    buf_clk cell_4849 ( .C (clk), .D (signal_6698), .Q (signal_6699) ) ;
    buf_clk cell_4857 ( .C (clk), .D (signal_6706), .Q (signal_6707) ) ;
    buf_clk cell_4865 ( .C (clk), .D (signal_6714), .Q (signal_6715) ) ;
    buf_clk cell_4873 ( .C (clk), .D (signal_6722), .Q (signal_6723) ) ;
    buf_clk cell_4881 ( .C (clk), .D (signal_6730), .Q (signal_6731) ) ;
    buf_clk cell_4889 ( .C (clk), .D (signal_6738), .Q (signal_6739) ) ;
    buf_clk cell_4897 ( .C (clk), .D (signal_6746), .Q (signal_6747) ) ;
    buf_clk cell_4905 ( .C (clk), .D (signal_6754), .Q (signal_6755) ) ;
    buf_clk cell_4913 ( .C (clk), .D (signal_6762), .Q (signal_6763) ) ;
    buf_clk cell_4921 ( .C (clk), .D (signal_6770), .Q (signal_6771) ) ;
    buf_clk cell_4929 ( .C (clk), .D (signal_6778), .Q (signal_6779) ) ;
    buf_clk cell_4937 ( .C (clk), .D (signal_6786), .Q (signal_6787) ) ;
    buf_clk cell_4945 ( .C (clk), .D (signal_6794), .Q (signal_6795) ) ;
    buf_clk cell_4953 ( .C (clk), .D (signal_6802), .Q (signal_6803) ) ;
    buf_clk cell_4961 ( .C (clk), .D (signal_6810), .Q (signal_6811) ) ;
    buf_clk cell_4969 ( .C (clk), .D (signal_6818), .Q (signal_6819) ) ;
    buf_clk cell_4977 ( .C (clk), .D (signal_6826), .Q (signal_6827) ) ;
    buf_clk cell_4985 ( .C (clk), .D (signal_6834), .Q (signal_6835) ) ;
    buf_clk cell_4993 ( .C (clk), .D (signal_6842), .Q (signal_6843) ) ;
    buf_clk cell_5001 ( .C (clk), .D (signal_6850), .Q (signal_6851) ) ;
    buf_clk cell_5009 ( .C (clk), .D (signal_6858), .Q (signal_6859) ) ;
    buf_clk cell_5017 ( .C (clk), .D (signal_6866), .Q (signal_6867) ) ;
    buf_clk cell_5025 ( .C (clk), .D (signal_6874), .Q (signal_6875) ) ;
    buf_clk cell_5033 ( .C (clk), .D (signal_6882), .Q (signal_6883) ) ;
    buf_clk cell_5041 ( .C (clk), .D (signal_6890), .Q (signal_6891) ) ;
    buf_clk cell_5049 ( .C (clk), .D (signal_6898), .Q (signal_6899) ) ;
    buf_clk cell_5057 ( .C (clk), .D (signal_6906), .Q (signal_6907) ) ;
    buf_clk cell_5065 ( .C (clk), .D (signal_6914), .Q (signal_6915) ) ;
    buf_clk cell_5073 ( .C (clk), .D (signal_6922), .Q (signal_6923) ) ;
    buf_clk cell_5081 ( .C (clk), .D (signal_6930), .Q (signal_6931) ) ;
    buf_clk cell_5089 ( .C (clk), .D (signal_6938), .Q (signal_6939) ) ;
    buf_clk cell_5097 ( .C (clk), .D (signal_6946), .Q (signal_6947) ) ;
    buf_clk cell_5105 ( .C (clk), .D (signal_6954), .Q (signal_6955) ) ;
    buf_clk cell_5113 ( .C (clk), .D (signal_6962), .Q (signal_6963) ) ;
    buf_clk cell_5121 ( .C (clk), .D (signal_6970), .Q (signal_6971) ) ;
    buf_clk cell_5129 ( .C (clk), .D (signal_6978), .Q (signal_6979) ) ;
    buf_clk cell_5137 ( .C (clk), .D (signal_6986), .Q (signal_6987) ) ;
    buf_clk cell_5145 ( .C (clk), .D (signal_6994), .Q (signal_6995) ) ;
    buf_clk cell_5153 ( .C (clk), .D (signal_7002), .Q (signal_7003) ) ;
    buf_clk cell_5161 ( .C (clk), .D (signal_7010), .Q (signal_7011) ) ;
    buf_clk cell_5169 ( .C (clk), .D (signal_7018), .Q (signal_7019) ) ;
    buf_clk cell_5177 ( .C (clk), .D (signal_7026), .Q (signal_7027) ) ;
    buf_clk cell_5185 ( .C (clk), .D (signal_7034), .Q (signal_7035) ) ;
    buf_clk cell_5193 ( .C (clk), .D (signal_7042), .Q (signal_7043) ) ;
    buf_clk cell_5201 ( .C (clk), .D (signal_7050), .Q (signal_7051) ) ;
    buf_clk cell_5209 ( .C (clk), .D (signal_7058), .Q (signal_7059) ) ;
    buf_clk cell_5217 ( .C (clk), .D (signal_7066), .Q (signal_7067) ) ;
    buf_clk cell_5225 ( .C (clk), .D (signal_7074), .Q (signal_7075) ) ;
    buf_clk cell_5233 ( .C (clk), .D (signal_7082), .Q (signal_7083) ) ;
    buf_clk cell_5241 ( .C (clk), .D (signal_7090), .Q (signal_7091) ) ;
    buf_clk cell_5249 ( .C (clk), .D (signal_7098), .Q (signal_7099) ) ;
    buf_clk cell_5257 ( .C (clk), .D (signal_7106), .Q (signal_7107) ) ;
    buf_clk cell_5265 ( .C (clk), .D (signal_7114), .Q (signal_7115) ) ;
    buf_clk cell_5273 ( .C (clk), .D (signal_7122), .Q (signal_7123) ) ;
    buf_clk cell_5281 ( .C (clk), .D (signal_7130), .Q (signal_7131) ) ;
    buf_clk cell_5289 ( .C (clk), .D (signal_7138), .Q (signal_7139) ) ;
    buf_clk cell_5297 ( .C (clk), .D (signal_7146), .Q (signal_7147) ) ;
    buf_clk cell_5305 ( .C (clk), .D (signal_7154), .Q (signal_7155) ) ;
    buf_clk cell_5313 ( .C (clk), .D (signal_7162), .Q (signal_7163) ) ;
    buf_clk cell_5321 ( .C (clk), .D (signal_7170), .Q (signal_7171) ) ;
    buf_clk cell_5329 ( .C (clk), .D (signal_7178), .Q (signal_7179) ) ;
    buf_clk cell_5337 ( .C (clk), .D (signal_7186), .Q (signal_7187) ) ;
    buf_clk cell_5345 ( .C (clk), .D (signal_7194), .Q (signal_7195) ) ;
    buf_clk cell_5353 ( .C (clk), .D (signal_7202), .Q (signal_7203) ) ;
    buf_clk cell_5361 ( .C (clk), .D (signal_7210), .Q (signal_7211) ) ;
    buf_clk cell_5369 ( .C (clk), .D (signal_7218), .Q (signal_7219) ) ;
    buf_clk cell_5377 ( .C (clk), .D (signal_7226), .Q (signal_7227) ) ;
    buf_clk cell_5385 ( .C (clk), .D (signal_7234), .Q (signal_7235) ) ;
    buf_clk cell_5393 ( .C (clk), .D (signal_7242), .Q (signal_7243) ) ;
    buf_clk cell_5401 ( .C (clk), .D (signal_7250), .Q (signal_7251) ) ;
    buf_clk cell_5409 ( .C (clk), .D (signal_7258), .Q (signal_7259) ) ;
    buf_clk cell_5417 ( .C (clk), .D (signal_7266), .Q (signal_7267) ) ;
    buf_clk cell_5425 ( .C (clk), .D (signal_7274), .Q (signal_7275) ) ;
    buf_clk cell_5433 ( .C (clk), .D (signal_7282), .Q (signal_7283) ) ;
    buf_clk cell_5441 ( .C (clk), .D (signal_7290), .Q (signal_7291) ) ;
    buf_clk cell_5449 ( .C (clk), .D (signal_7298), .Q (signal_7299) ) ;
    buf_clk cell_5457 ( .C (clk), .D (signal_7306), .Q (signal_7307) ) ;
    buf_clk cell_5465 ( .C (clk), .D (signal_7314), .Q (signal_7315) ) ;
    buf_clk cell_5473 ( .C (clk), .D (signal_7322), .Q (signal_7323) ) ;
    buf_clk cell_5481 ( .C (clk), .D (signal_7330), .Q (signal_7331) ) ;
    buf_clk cell_5489 ( .C (clk), .D (signal_7338), .Q (signal_7339) ) ;
    buf_clk cell_5497 ( .C (clk), .D (signal_7346), .Q (signal_7347) ) ;
    buf_clk cell_5505 ( .C (clk), .D (signal_7354), .Q (signal_7355) ) ;
    buf_clk cell_5513 ( .C (clk), .D (signal_7362), .Q (signal_7363) ) ;
    buf_clk cell_5521 ( .C (clk), .D (signal_7370), .Q (signal_7371) ) ;
    buf_clk cell_5529 ( .C (clk), .D (signal_7378), .Q (signal_7379) ) ;
    buf_clk cell_5537 ( .C (clk), .D (signal_7386), .Q (signal_7387) ) ;
    buf_clk cell_5545 ( .C (clk), .D (signal_7394), .Q (signal_7395) ) ;
    buf_clk cell_5553 ( .C (clk), .D (signal_7402), .Q (signal_7403) ) ;
    buf_clk cell_5561 ( .C (clk), .D (signal_7410), .Q (signal_7411) ) ;
    buf_clk cell_5569 ( .C (clk), .D (signal_7418), .Q (signal_7419) ) ;
    buf_clk cell_5577 ( .C (clk), .D (signal_7426), .Q (signal_7427) ) ;
    buf_clk cell_5585 ( .C (clk), .D (signal_7434), .Q (signal_7435) ) ;
    buf_clk cell_5593 ( .C (clk), .D (signal_7442), .Q (signal_7443) ) ;
    buf_clk cell_5601 ( .C (clk), .D (signal_7450), .Q (signal_7451) ) ;
    buf_clk cell_5609 ( .C (clk), .D (signal_7458), .Q (signal_7459) ) ;
    buf_clk cell_5617 ( .C (clk), .D (signal_7466), .Q (signal_7467) ) ;
    buf_clk cell_5625 ( .C (clk), .D (signal_7474), .Q (signal_7475) ) ;
    buf_clk cell_5633 ( .C (clk), .D (signal_7482), .Q (signal_7483) ) ;
    buf_clk cell_5641 ( .C (clk), .D (signal_7490), .Q (signal_7491) ) ;
    buf_clk cell_5649 ( .C (clk), .D (signal_7498), .Q (signal_7499) ) ;
    buf_clk cell_5657 ( .C (clk), .D (signal_7506), .Q (signal_7507) ) ;
    buf_clk cell_5665 ( .C (clk), .D (signal_7514), .Q (signal_7515) ) ;
    buf_clk cell_5673 ( .C (clk), .D (signal_7522), .Q (signal_7523) ) ;
    buf_clk cell_5681 ( .C (clk), .D (signal_7530), .Q (signal_7531) ) ;
    buf_clk cell_5689 ( .C (clk), .D (signal_7538), .Q (signal_7539) ) ;
    buf_clk cell_5697 ( .C (clk), .D (signal_7546), .Q (signal_7547) ) ;
    buf_clk cell_5705 ( .C (clk), .D (signal_7554), .Q (signal_7555) ) ;
    buf_clk cell_5713 ( .C (clk), .D (signal_7562), .Q (signal_7563) ) ;
    buf_clk cell_5721 ( .C (clk), .D (signal_7570), .Q (signal_7571) ) ;
    buf_clk cell_5729 ( .C (clk), .D (signal_7578), .Q (signal_7579) ) ;
    buf_clk cell_5737 ( .C (clk), .D (signal_7586), .Q (signal_7587) ) ;
    buf_clk cell_5745 ( .C (clk), .D (signal_7594), .Q (signal_7595) ) ;
    buf_clk cell_5753 ( .C (clk), .D (signal_7602), .Q (signal_7603) ) ;
    buf_clk cell_5761 ( .C (clk), .D (signal_7610), .Q (signal_7611) ) ;
    buf_clk cell_5769 ( .C (clk), .D (signal_7618), .Q (signal_7619) ) ;
    buf_clk cell_5777 ( .C (clk), .D (signal_7626), .Q (signal_7627) ) ;
    buf_clk cell_5785 ( .C (clk), .D (signal_7634), .Q (signal_7635) ) ;
    buf_clk cell_5793 ( .C (clk), .D (signal_7642), .Q (signal_7643) ) ;
    buf_clk cell_5801 ( .C (clk), .D (signal_7650), .Q (signal_7651) ) ;
    buf_clk cell_5809 ( .C (clk), .D (signal_7658), .Q (signal_7659) ) ;
    buf_clk cell_5817 ( .C (clk), .D (signal_7666), .Q (signal_7667) ) ;
    buf_clk cell_5825 ( .C (clk), .D (signal_7674), .Q (signal_7675) ) ;
    buf_clk cell_5833 ( .C (clk), .D (signal_7682), .Q (signal_7683) ) ;
    buf_clk cell_5841 ( .C (clk), .D (signal_7690), .Q (signal_7691) ) ;
    buf_clk cell_5849 ( .C (clk), .D (signal_7698), .Q (signal_7699) ) ;
    buf_clk cell_5857 ( .C (clk), .D (signal_7706), .Q (signal_7707) ) ;
    buf_clk cell_5865 ( .C (clk), .D (signal_7714), .Q (signal_7715) ) ;
    buf_clk cell_5873 ( .C (clk), .D (signal_7722), .Q (signal_7723) ) ;
    buf_clk cell_5881 ( .C (clk), .D (signal_7730), .Q (signal_7731) ) ;
    buf_clk cell_5889 ( .C (clk), .D (signal_7738), .Q (signal_7739) ) ;
    buf_clk cell_5897 ( .C (clk), .D (signal_7746), .Q (signal_7747) ) ;
    buf_clk cell_5905 ( .C (clk), .D (signal_7754), .Q (signal_7755) ) ;
    buf_clk cell_5913 ( .C (clk), .D (signal_7762), .Q (signal_7763) ) ;
    buf_clk cell_5921 ( .C (clk), .D (signal_7770), .Q (signal_7771) ) ;
    buf_clk cell_5929 ( .C (clk), .D (signal_7778), .Q (signal_7779) ) ;
    buf_clk cell_5937 ( .C (clk), .D (signal_7786), .Q (signal_7787) ) ;
    buf_clk cell_5945 ( .C (clk), .D (signal_7794), .Q (signal_7795) ) ;
    buf_clk cell_5953 ( .C (clk), .D (signal_7802), .Q (signal_7803) ) ;
    buf_clk cell_5961 ( .C (clk), .D (signal_7810), .Q (signal_7811) ) ;
    buf_clk cell_5969 ( .C (clk), .D (signal_7818), .Q (signal_7819) ) ;
    buf_clk cell_5977 ( .C (clk), .D (signal_7826), .Q (signal_7827) ) ;
    buf_clk cell_5985 ( .C (clk), .D (signal_7834), .Q (signal_7835) ) ;
    buf_clk cell_5993 ( .C (clk), .D (signal_7842), .Q (signal_7843) ) ;
    buf_clk cell_6001 ( .C (clk), .D (signal_7850), .Q (signal_7851) ) ;
    buf_clk cell_6009 ( .C (clk), .D (signal_7858), .Q (signal_7859) ) ;
    buf_clk cell_6017 ( .C (clk), .D (signal_7866), .Q (signal_7867) ) ;
    buf_clk cell_6025 ( .C (clk), .D (signal_7874), .Q (signal_7875) ) ;
    buf_clk cell_6033 ( .C (clk), .D (signal_7882), .Q (signal_7883) ) ;
    buf_clk cell_6041 ( .C (clk), .D (signal_7890), .Q (signal_7891) ) ;
    buf_clk cell_6049 ( .C (clk), .D (signal_7898), .Q (signal_7899) ) ;
    buf_clk cell_6057 ( .C (clk), .D (signal_7906), .Q (signal_7907) ) ;
    buf_clk cell_6065 ( .C (clk), .D (signal_7914), .Q (signal_7915) ) ;
    buf_clk cell_6073 ( .C (clk), .D (signal_7922), .Q (signal_7923) ) ;
    buf_clk cell_6081 ( .C (clk), .D (signal_7930), .Q (signal_7931) ) ;
    buf_clk cell_6089 ( .C (clk), .D (signal_7938), .Q (signal_7939) ) ;
    buf_clk cell_6097 ( .C (clk), .D (signal_7946), .Q (signal_7947) ) ;
    buf_clk cell_6105 ( .C (clk), .D (signal_7954), .Q (signal_7955) ) ;
    buf_clk cell_6113 ( .C (clk), .D (signal_7962), .Q (signal_7963) ) ;
    buf_clk cell_6121 ( .C (clk), .D (signal_7970), .Q (signal_7971) ) ;
    buf_clk cell_6129 ( .C (clk), .D (signal_7978), .Q (signal_7979) ) ;
    buf_clk cell_6137 ( .C (clk), .D (signal_7986), .Q (signal_7987) ) ;
    buf_clk cell_6145 ( .C (clk), .D (signal_7994), .Q (signal_7995) ) ;
    buf_clk cell_6153 ( .C (clk), .D (signal_8002), .Q (signal_8003) ) ;
    buf_clk cell_6161 ( .C (clk), .D (signal_8010), .Q (signal_8011) ) ;
    buf_clk cell_6169 ( .C (clk), .D (signal_8018), .Q (signal_8019) ) ;
    buf_clk cell_6177 ( .C (clk), .D (signal_8026), .Q (signal_8027) ) ;
    buf_clk cell_6185 ( .C (clk), .D (signal_8034), .Q (signal_8035) ) ;
    buf_clk cell_6193 ( .C (clk), .D (signal_8042), .Q (signal_8043) ) ;
    buf_clk cell_6201 ( .C (clk), .D (signal_8050), .Q (signal_8051) ) ;
    buf_clk cell_6209 ( .C (clk), .D (signal_8058), .Q (signal_8059) ) ;
    buf_clk cell_6217 ( .C (clk), .D (signal_8066), .Q (signal_8067) ) ;
    buf_clk cell_6225 ( .C (clk), .D (signal_8074), .Q (signal_8075) ) ;
    buf_clk cell_6233 ( .C (clk), .D (signal_8082), .Q (signal_8083) ) ;
    buf_clk cell_6241 ( .C (clk), .D (signal_8090), .Q (signal_8091) ) ;
    buf_clk cell_6249 ( .C (clk), .D (signal_8098), .Q (signal_8099) ) ;
    buf_clk cell_6257 ( .C (clk), .D (signal_8106), .Q (signal_8107) ) ;
    buf_clk cell_6265 ( .C (clk), .D (signal_8114), .Q (signal_8115) ) ;
    buf_clk cell_6273 ( .C (clk), .D (signal_8122), .Q (signal_8123) ) ;
    buf_clk cell_6281 ( .C (clk), .D (signal_8130), .Q (signal_8131) ) ;
    buf_clk cell_6289 ( .C (clk), .D (signal_8138), .Q (signal_8139) ) ;
    buf_clk cell_6297 ( .C (clk), .D (signal_8146), .Q (signal_8147) ) ;
    buf_clk cell_6305 ( .C (clk), .D (signal_8154), .Q (signal_8155) ) ;
    buf_clk cell_6313 ( .C (clk), .D (signal_8162), .Q (signal_8163) ) ;
    buf_clk cell_6321 ( .C (clk), .D (signal_8170), .Q (signal_8171) ) ;
    buf_clk cell_6329 ( .C (clk), .D (signal_8178), .Q (signal_8179) ) ;
    buf_clk cell_6337 ( .C (clk), .D (signal_8186), .Q (signal_8187) ) ;
    buf_clk cell_6345 ( .C (clk), .D (signal_8194), .Q (signal_8195) ) ;
    buf_clk cell_6353 ( .C (clk), .D (signal_8202), .Q (signal_8203) ) ;
    buf_clk cell_6361 ( .C (clk), .D (signal_8210), .Q (signal_8211) ) ;
    buf_clk cell_6369 ( .C (clk), .D (signal_8218), .Q (signal_8219) ) ;
    buf_clk cell_6377 ( .C (clk), .D (signal_8226), .Q (signal_8227) ) ;
    buf_clk cell_6385 ( .C (clk), .D (signal_8234), .Q (signal_8235) ) ;
    buf_clk cell_6393 ( .C (clk), .D (signal_8242), .Q (signal_8243) ) ;
    buf_clk cell_6401 ( .C (clk), .D (signal_8250), .Q (signal_8251) ) ;
    buf_clk cell_6409 ( .C (clk), .D (signal_8258), .Q (signal_8259) ) ;
    buf_clk cell_6417 ( .C (clk), .D (signal_8266), .Q (signal_8267) ) ;
    buf_clk cell_6425 ( .C (clk), .D (signal_8274), .Q (signal_8275) ) ;
    buf_clk cell_6433 ( .C (clk), .D (signal_8282), .Q (signal_8283) ) ;
    buf_clk cell_6441 ( .C (clk), .D (signal_8290), .Q (signal_8291) ) ;
    buf_clk cell_6449 ( .C (clk), .D (signal_8298), .Q (signal_8299) ) ;
    buf_clk cell_6457 ( .C (clk), .D (signal_8306), .Q (signal_8307) ) ;
    buf_clk cell_6465 ( .C (clk), .D (signal_8314), .Q (signal_8315) ) ;
    buf_clk cell_6473 ( .C (clk), .D (signal_8322), .Q (signal_8323) ) ;
    buf_clk cell_6481 ( .C (clk), .D (signal_8330), .Q (signal_8331) ) ;
    buf_clk cell_6489 ( .C (clk), .D (signal_8338), .Q (signal_8339) ) ;
    buf_clk cell_6497 ( .C (clk), .D (signal_8346), .Q (signal_8347) ) ;
    buf_clk cell_6505 ( .C (clk), .D (signal_8354), .Q (signal_8355) ) ;
    buf_clk cell_6513 ( .C (clk), .D (signal_8362), .Q (signal_8363) ) ;
    buf_clk cell_6521 ( .C (clk), .D (signal_8370), .Q (signal_8371) ) ;
    buf_clk cell_6529 ( .C (clk), .D (signal_8378), .Q (signal_8379) ) ;
    buf_clk cell_6537 ( .C (clk), .D (signal_8386), .Q (signal_8387) ) ;
    buf_clk cell_6545 ( .C (clk), .D (signal_8394), .Q (signal_8395) ) ;
    buf_clk cell_6553 ( .C (clk), .D (signal_8402), .Q (signal_8403) ) ;
    buf_clk cell_6561 ( .C (clk), .D (signal_8410), .Q (signal_8411) ) ;
    buf_clk cell_6569 ( .C (clk), .D (signal_8418), .Q (signal_8419) ) ;
    buf_clk cell_6577 ( .C (clk), .D (signal_8426), .Q (signal_8427) ) ;
    buf_clk cell_6585 ( .C (clk), .D (signal_8434), .Q (signal_8435) ) ;
    buf_clk cell_6593 ( .C (clk), .D (signal_8442), .Q (signal_8443) ) ;
    buf_clk cell_6601 ( .C (clk), .D (signal_8450), .Q (signal_8451) ) ;
    buf_clk cell_6609 ( .C (clk), .D (signal_8458), .Q (signal_8459) ) ;
    buf_clk cell_6617 ( .C (clk), .D (signal_8466), .Q (signal_8467) ) ;
    buf_clk cell_6625 ( .C (clk), .D (signal_8474), .Q (signal_8475) ) ;
    buf_clk cell_6633 ( .C (clk), .D (signal_8482), .Q (signal_8483) ) ;
    buf_clk cell_6641 ( .C (clk), .D (signal_8490), .Q (signal_8491) ) ;
    buf_clk cell_6649 ( .C (clk), .D (signal_8498), .Q (signal_8499) ) ;
    buf_clk cell_6657 ( .C (clk), .D (signal_8506), .Q (signal_8507) ) ;
    buf_clk cell_6665 ( .C (clk), .D (signal_8514), .Q (signal_8515) ) ;
    buf_clk cell_6673 ( .C (clk), .D (signal_8522), .Q (signal_8523) ) ;
    buf_clk cell_6681 ( .C (clk), .D (signal_8530), .Q (signal_8531) ) ;
    buf_clk cell_6689 ( .C (clk), .D (signal_8538), .Q (signal_8539) ) ;
    buf_clk cell_6697 ( .C (clk), .D (signal_8546), .Q (signal_8547) ) ;
    buf_clk cell_6705 ( .C (clk), .D (signal_8554), .Q (signal_8555) ) ;
    buf_clk cell_6713 ( .C (clk), .D (signal_8562), .Q (signal_8563) ) ;
    buf_clk cell_6721 ( .C (clk), .D (signal_8570), .Q (signal_8571) ) ;
    buf_clk cell_6729 ( .C (clk), .D (signal_8578), .Q (signal_8579) ) ;
    buf_clk cell_6737 ( .C (clk), .D (signal_8586), .Q (signal_8587) ) ;
    buf_clk cell_6745 ( .C (clk), .D (signal_8594), .Q (signal_8595) ) ;
    buf_clk cell_6753 ( .C (clk), .D (signal_8602), .Q (signal_8603) ) ;
    buf_clk cell_6761 ( .C (clk), .D (signal_8610), .Q (signal_8611) ) ;
    buf_clk cell_6769 ( .C (clk), .D (signal_8618), .Q (signal_8619) ) ;
    buf_clk cell_6777 ( .C (clk), .D (signal_8626), .Q (signal_8627) ) ;
    buf_clk cell_6785 ( .C (clk), .D (signal_8634), .Q (signal_8635) ) ;
    buf_clk cell_6793 ( .C (clk), .D (signal_8642), .Q (signal_8643) ) ;
    buf_clk cell_6801 ( .C (clk), .D (signal_8650), .Q (signal_8651) ) ;
    buf_clk cell_6809 ( .C (clk), .D (signal_8658), .Q (signal_8659) ) ;
    buf_clk cell_6817 ( .C (clk), .D (signal_8666), .Q (signal_8667) ) ;
    buf_clk cell_6825 ( .C (clk), .D (signal_8674), .Q (signal_8675) ) ;
    buf_clk cell_6833 ( .C (clk), .D (signal_8682), .Q (signal_8683) ) ;
    buf_clk cell_6841 ( .C (clk), .D (signal_8690), .Q (signal_8691) ) ;
    buf_clk cell_6849 ( .C (clk), .D (signal_8698), .Q (signal_8699) ) ;
    buf_clk cell_6857 ( .C (clk), .D (signal_8706), .Q (signal_8707) ) ;
    buf_clk cell_6865 ( .C (clk), .D (signal_8714), .Q (signal_8715) ) ;
    buf_clk cell_6873 ( .C (clk), .D (signal_8722), .Q (signal_8723) ) ;
    buf_clk cell_6881 ( .C (clk), .D (signal_8730), .Q (signal_8731) ) ;
    buf_clk cell_6889 ( .C (clk), .D (signal_8738), .Q (signal_8739) ) ;
    buf_clk cell_6897 ( .C (clk), .D (signal_8746), .Q (signal_8747) ) ;
    buf_clk cell_6905 ( .C (clk), .D (signal_8754), .Q (signal_8755) ) ;
    buf_clk cell_6913 ( .C (clk), .D (signal_8762), .Q (signal_8763) ) ;
    buf_clk cell_6921 ( .C (clk), .D (signal_8770), .Q (signal_8771) ) ;
    buf_clk cell_6929 ( .C (clk), .D (signal_8778), .Q (signal_8779) ) ;
    buf_clk cell_6937 ( .C (clk), .D (signal_8786), .Q (signal_8787) ) ;
    buf_clk cell_6945 ( .C (clk), .D (signal_8794), .Q (signal_8795) ) ;
    buf_clk cell_6953 ( .C (clk), .D (signal_8802), .Q (signal_8803) ) ;
    buf_clk cell_6961 ( .C (clk), .D (signal_8810), .Q (signal_8811) ) ;
    buf_clk cell_6969 ( .C (clk), .D (signal_8818), .Q (signal_8819) ) ;
    buf_clk cell_6977 ( .C (clk), .D (signal_8826), .Q (signal_8827) ) ;
    buf_clk cell_6985 ( .C (clk), .D (signal_8834), .Q (signal_8835) ) ;
    buf_clk cell_6993 ( .C (clk), .D (signal_8842), .Q (signal_8843) ) ;
    buf_clk cell_7001 ( .C (clk), .D (signal_8850), .Q (signal_8851) ) ;
    buf_clk cell_7009 ( .C (clk), .D (signal_8858), .Q (signal_8859) ) ;
    buf_clk cell_7017 ( .C (clk), .D (signal_8866), .Q (signal_8867) ) ;
    buf_clk cell_7025 ( .C (clk), .D (signal_8874), .Q (signal_8875) ) ;
    buf_clk cell_7033 ( .C (clk), .D (signal_8882), .Q (signal_8883) ) ;
    buf_clk cell_7041 ( .C (clk), .D (signal_8890), .Q (signal_8891) ) ;
    buf_clk cell_7049 ( .C (clk), .D (signal_8898), .Q (signal_8899) ) ;
    buf_clk cell_7057 ( .C (clk), .D (signal_8906), .Q (signal_8907) ) ;
    buf_clk cell_7065 ( .C (clk), .D (signal_8914), .Q (signal_8915) ) ;
    buf_clk cell_7073 ( .C (clk), .D (signal_8922), .Q (signal_8923) ) ;
    buf_clk cell_7081 ( .C (clk), .D (signal_8930), .Q (signal_8931) ) ;
    buf_clk cell_7089 ( .C (clk), .D (signal_8938), .Q (signal_8939) ) ;
    buf_clk cell_7097 ( .C (clk), .D (signal_8946), .Q (signal_8947) ) ;

    /* cells in depth 5 */
    buf_clk cell_1878 ( .C (clk), .D (signal_3713), .Q (signal_3728) ) ;
    buf_clk cell_1880 ( .C (clk), .D (signal_3715), .Q (signal_3730) ) ;
    buf_clk cell_1882 ( .C (clk), .D (signal_2039), .Q (signal_3732) ) ;
    buf_clk cell_1884 ( .C (clk), .D (signal_3515), .Q (signal_3734) ) ;
    buf_clk cell_1886 ( .C (clk), .D (signal_3717), .Q (signal_3736) ) ;
    buf_clk cell_1888 ( .C (clk), .D (signal_3719), .Q (signal_3738) ) ;
    buf_clk cell_1890 ( .C (clk), .D (signal_2044), .Q (signal_3740) ) ;
    buf_clk cell_1892 ( .C (clk), .D (signal_3520), .Q (signal_3742) ) ;
    buf_clk cell_1898 ( .C (clk), .D (signal_3747), .Q (signal_3748) ) ;
    buf_clk cell_1906 ( .C (clk), .D (signal_3755), .Q (signal_3756) ) ;
    buf_clk cell_1914 ( .C (clk), .D (signal_3763), .Q (signal_3764) ) ;
    buf_clk cell_1922 ( .C (clk), .D (signal_3771), .Q (signal_3772) ) ;
    buf_clk cell_1930 ( .C (clk), .D (signal_3779), .Q (signal_3780) ) ;
    buf_clk cell_1938 ( .C (clk), .D (signal_3787), .Q (signal_3788) ) ;
    buf_clk cell_1946 ( .C (clk), .D (signal_3795), .Q (signal_3796) ) ;
    buf_clk cell_1954 ( .C (clk), .D (signal_3803), .Q (signal_3804) ) ;
    buf_clk cell_1962 ( .C (clk), .D (signal_3811), .Q (signal_3812) ) ;
    buf_clk cell_1970 ( .C (clk), .D (signal_3819), .Q (signal_3820) ) ;
    buf_clk cell_1978 ( .C (clk), .D (signal_3827), .Q (signal_3828) ) ;
    buf_clk cell_1986 ( .C (clk), .D (signal_3835), .Q (signal_3836) ) ;
    buf_clk cell_1994 ( .C (clk), .D (signal_3843), .Q (signal_3844) ) ;
    buf_clk cell_2002 ( .C (clk), .D (signal_3851), .Q (signal_3852) ) ;
    buf_clk cell_2010 ( .C (clk), .D (signal_3859), .Q (signal_3860) ) ;
    buf_clk cell_2018 ( .C (clk), .D (signal_3867), .Q (signal_3868) ) ;
    buf_clk cell_2026 ( .C (clk), .D (signal_3875), .Q (signal_3876) ) ;
    buf_clk cell_2034 ( .C (clk), .D (signal_3883), .Q (signal_3884) ) ;
    buf_clk cell_2042 ( .C (clk), .D (signal_3891), .Q (signal_3892) ) ;
    buf_clk cell_2050 ( .C (clk), .D (signal_3899), .Q (signal_3900) ) ;
    buf_clk cell_2058 ( .C (clk), .D (signal_3907), .Q (signal_3908) ) ;
    buf_clk cell_2066 ( .C (clk), .D (signal_3915), .Q (signal_3916) ) ;
    buf_clk cell_2074 ( .C (clk), .D (signal_3923), .Q (signal_3924) ) ;
    buf_clk cell_2082 ( .C (clk), .D (signal_3931), .Q (signal_3932) ) ;
    buf_clk cell_2090 ( .C (clk), .D (signal_3939), .Q (signal_3940) ) ;
    buf_clk cell_2098 ( .C (clk), .D (signal_3947), .Q (signal_3948) ) ;
    buf_clk cell_2106 ( .C (clk), .D (signal_3955), .Q (signal_3956) ) ;
    buf_clk cell_2114 ( .C (clk), .D (signal_3963), .Q (signal_3964) ) ;
    buf_clk cell_2122 ( .C (clk), .D (signal_3971), .Q (signal_3972) ) ;
    buf_clk cell_2130 ( .C (clk), .D (signal_3979), .Q (signal_3980) ) ;
    buf_clk cell_2138 ( .C (clk), .D (signal_3987), .Q (signal_3988) ) ;
    buf_clk cell_2146 ( .C (clk), .D (signal_3995), .Q (signal_3996) ) ;
    buf_clk cell_2154 ( .C (clk), .D (signal_4003), .Q (signal_4004) ) ;
    buf_clk cell_2162 ( .C (clk), .D (signal_4011), .Q (signal_4012) ) ;
    buf_clk cell_2170 ( .C (clk), .D (signal_4019), .Q (signal_4020) ) ;
    buf_clk cell_2178 ( .C (clk), .D (signal_4027), .Q (signal_4028) ) ;
    buf_clk cell_2186 ( .C (clk), .D (signal_4035), .Q (signal_4036) ) ;
    buf_clk cell_2194 ( .C (clk), .D (signal_4043), .Q (signal_4044) ) ;
    buf_clk cell_2202 ( .C (clk), .D (signal_4051), .Q (signal_4052) ) ;
    buf_clk cell_2210 ( .C (clk), .D (signal_4059), .Q (signal_4060) ) ;
    buf_clk cell_2218 ( .C (clk), .D (signal_4067), .Q (signal_4068) ) ;
    buf_clk cell_2226 ( .C (clk), .D (signal_4075), .Q (signal_4076) ) ;
    buf_clk cell_2234 ( .C (clk), .D (signal_4083), .Q (signal_4084) ) ;
    buf_clk cell_2242 ( .C (clk), .D (signal_4091), .Q (signal_4092) ) ;
    buf_clk cell_2250 ( .C (clk), .D (signal_4099), .Q (signal_4100) ) ;
    buf_clk cell_2258 ( .C (clk), .D (signal_4107), .Q (signal_4108) ) ;
    buf_clk cell_2266 ( .C (clk), .D (signal_4115), .Q (signal_4116) ) ;
    buf_clk cell_2274 ( .C (clk), .D (signal_4123), .Q (signal_4124) ) ;
    buf_clk cell_2282 ( .C (clk), .D (signal_4131), .Q (signal_4132) ) ;
    buf_clk cell_2290 ( .C (clk), .D (signal_4139), .Q (signal_4140) ) ;
    buf_clk cell_2298 ( .C (clk), .D (signal_4147), .Q (signal_4148) ) ;
    buf_clk cell_2306 ( .C (clk), .D (signal_4155), .Q (signal_4156) ) ;
    buf_clk cell_2314 ( .C (clk), .D (signal_4163), .Q (signal_4164) ) ;
    buf_clk cell_2322 ( .C (clk), .D (signal_4171), .Q (signal_4172) ) ;
    buf_clk cell_2330 ( .C (clk), .D (signal_4179), .Q (signal_4180) ) ;
    buf_clk cell_2338 ( .C (clk), .D (signal_4187), .Q (signal_4188) ) ;
    buf_clk cell_2346 ( .C (clk), .D (signal_4195), .Q (signal_4196) ) ;
    buf_clk cell_2354 ( .C (clk), .D (signal_4203), .Q (signal_4204) ) ;
    buf_clk cell_2362 ( .C (clk), .D (signal_4211), .Q (signal_4212) ) ;
    buf_clk cell_2370 ( .C (clk), .D (signal_4219), .Q (signal_4220) ) ;
    buf_clk cell_2378 ( .C (clk), .D (signal_4227), .Q (signal_4228) ) ;
    buf_clk cell_2386 ( .C (clk), .D (signal_4235), .Q (signal_4236) ) ;
    buf_clk cell_2394 ( .C (clk), .D (signal_4243), .Q (signal_4244) ) ;
    buf_clk cell_2402 ( .C (clk), .D (signal_4251), .Q (signal_4252) ) ;
    buf_clk cell_2410 ( .C (clk), .D (signal_4259), .Q (signal_4260) ) ;
    buf_clk cell_2418 ( .C (clk), .D (signal_4267), .Q (signal_4268) ) ;
    buf_clk cell_2426 ( .C (clk), .D (signal_4275), .Q (signal_4276) ) ;
    buf_clk cell_2434 ( .C (clk), .D (signal_4283), .Q (signal_4284) ) ;
    buf_clk cell_2442 ( .C (clk), .D (signal_4291), .Q (signal_4292) ) ;
    buf_clk cell_2450 ( .C (clk), .D (signal_4299), .Q (signal_4300) ) ;
    buf_clk cell_2458 ( .C (clk), .D (signal_4307), .Q (signal_4308) ) ;
    buf_clk cell_2466 ( .C (clk), .D (signal_4315), .Q (signal_4316) ) ;
    buf_clk cell_2474 ( .C (clk), .D (signal_4323), .Q (signal_4324) ) ;
    buf_clk cell_2482 ( .C (clk), .D (signal_4331), .Q (signal_4332) ) ;
    buf_clk cell_2490 ( .C (clk), .D (signal_4339), .Q (signal_4340) ) ;
    buf_clk cell_2498 ( .C (clk), .D (signal_4347), .Q (signal_4348) ) ;
    buf_clk cell_2506 ( .C (clk), .D (signal_4355), .Q (signal_4356) ) ;
    buf_clk cell_2514 ( .C (clk), .D (signal_4363), .Q (signal_4364) ) ;
    buf_clk cell_2522 ( .C (clk), .D (signal_4371), .Q (signal_4372) ) ;
    buf_clk cell_2530 ( .C (clk), .D (signal_4379), .Q (signal_4380) ) ;
    buf_clk cell_2538 ( .C (clk), .D (signal_4387), .Q (signal_4388) ) ;
    buf_clk cell_2546 ( .C (clk), .D (signal_4395), .Q (signal_4396) ) ;
    buf_clk cell_2554 ( .C (clk), .D (signal_4403), .Q (signal_4404) ) ;
    buf_clk cell_2562 ( .C (clk), .D (signal_4411), .Q (signal_4412) ) ;
    buf_clk cell_2570 ( .C (clk), .D (signal_4419), .Q (signal_4420) ) ;
    buf_clk cell_2578 ( .C (clk), .D (signal_4427), .Q (signal_4428) ) ;
    buf_clk cell_2586 ( .C (clk), .D (signal_4435), .Q (signal_4436) ) ;
    buf_clk cell_2594 ( .C (clk), .D (signal_4443), .Q (signal_4444) ) ;
    buf_clk cell_2602 ( .C (clk), .D (signal_4451), .Q (signal_4452) ) ;
    buf_clk cell_2610 ( .C (clk), .D (signal_4459), .Q (signal_4460) ) ;
    buf_clk cell_2618 ( .C (clk), .D (signal_4467), .Q (signal_4468) ) ;
    buf_clk cell_2626 ( .C (clk), .D (signal_4475), .Q (signal_4476) ) ;
    buf_clk cell_2634 ( .C (clk), .D (signal_4483), .Q (signal_4484) ) ;
    buf_clk cell_2642 ( .C (clk), .D (signal_4491), .Q (signal_4492) ) ;
    buf_clk cell_2650 ( .C (clk), .D (signal_4499), .Q (signal_4500) ) ;
    buf_clk cell_2658 ( .C (clk), .D (signal_4507), .Q (signal_4508) ) ;
    buf_clk cell_2666 ( .C (clk), .D (signal_4515), .Q (signal_4516) ) ;
    buf_clk cell_2674 ( .C (clk), .D (signal_4523), .Q (signal_4524) ) ;
    buf_clk cell_2682 ( .C (clk), .D (signal_4531), .Q (signal_4532) ) ;
    buf_clk cell_2690 ( .C (clk), .D (signal_4539), .Q (signal_4540) ) ;
    buf_clk cell_2698 ( .C (clk), .D (signal_4547), .Q (signal_4548) ) ;
    buf_clk cell_2706 ( .C (clk), .D (signal_4555), .Q (signal_4556) ) ;
    buf_clk cell_2714 ( .C (clk), .D (signal_4563), .Q (signal_4564) ) ;
    buf_clk cell_2722 ( .C (clk), .D (signal_4571), .Q (signal_4572) ) ;
    buf_clk cell_2730 ( .C (clk), .D (signal_4579), .Q (signal_4580) ) ;
    buf_clk cell_2738 ( .C (clk), .D (signal_4587), .Q (signal_4588) ) ;
    buf_clk cell_2746 ( .C (clk), .D (signal_4595), .Q (signal_4596) ) ;
    buf_clk cell_2754 ( .C (clk), .D (signal_4603), .Q (signal_4604) ) ;
    buf_clk cell_2762 ( .C (clk), .D (signal_4611), .Q (signal_4612) ) ;
    buf_clk cell_2770 ( .C (clk), .D (signal_4619), .Q (signal_4620) ) ;
    buf_clk cell_2778 ( .C (clk), .D (signal_4627), .Q (signal_4628) ) ;
    buf_clk cell_2786 ( .C (clk), .D (signal_4635), .Q (signal_4636) ) ;
    buf_clk cell_2794 ( .C (clk), .D (signal_4643), .Q (signal_4644) ) ;
    buf_clk cell_2802 ( .C (clk), .D (signal_4651), .Q (signal_4652) ) ;
    buf_clk cell_2810 ( .C (clk), .D (signal_4659), .Q (signal_4660) ) ;
    buf_clk cell_2818 ( .C (clk), .D (signal_4667), .Q (signal_4668) ) ;
    buf_clk cell_2826 ( .C (clk), .D (signal_4675), .Q (signal_4676) ) ;
    buf_clk cell_2834 ( .C (clk), .D (signal_4683), .Q (signal_4684) ) ;
    buf_clk cell_2842 ( .C (clk), .D (signal_4691), .Q (signal_4692) ) ;
    buf_clk cell_2850 ( .C (clk), .D (signal_4699), .Q (signal_4700) ) ;
    buf_clk cell_2858 ( .C (clk), .D (signal_4707), .Q (signal_4708) ) ;
    buf_clk cell_2866 ( .C (clk), .D (signal_4715), .Q (signal_4716) ) ;
    buf_clk cell_2874 ( .C (clk), .D (signal_4723), .Q (signal_4724) ) ;
    buf_clk cell_2882 ( .C (clk), .D (signal_4731), .Q (signal_4732) ) ;
    buf_clk cell_2890 ( .C (clk), .D (signal_4739), .Q (signal_4740) ) ;
    buf_clk cell_2898 ( .C (clk), .D (signal_4747), .Q (signal_4748) ) ;
    buf_clk cell_2906 ( .C (clk), .D (signal_4755), .Q (signal_4756) ) ;
    buf_clk cell_2912 ( .C (clk), .D (signal_4761), .Q (signal_4762) ) ;
    buf_clk cell_2918 ( .C (clk), .D (signal_4767), .Q (signal_4768) ) ;
    buf_clk cell_2924 ( .C (clk), .D (signal_4773), .Q (signal_4774) ) ;
    buf_clk cell_2930 ( .C (clk), .D (signal_4779), .Q (signal_4780) ) ;
    buf_clk cell_2936 ( .C (clk), .D (signal_4785), .Q (signal_4786) ) ;
    buf_clk cell_2942 ( .C (clk), .D (signal_4791), .Q (signal_4792) ) ;
    buf_clk cell_2948 ( .C (clk), .D (signal_4797), .Q (signal_4798) ) ;
    buf_clk cell_2954 ( .C (clk), .D (signal_4803), .Q (signal_4804) ) ;
    buf_clk cell_2960 ( .C (clk), .D (signal_4809), .Q (signal_4810) ) ;
    buf_clk cell_2966 ( .C (clk), .D (signal_4815), .Q (signal_4816) ) ;
    buf_clk cell_2972 ( .C (clk), .D (signal_4821), .Q (signal_4822) ) ;
    buf_clk cell_2978 ( .C (clk), .D (signal_4827), .Q (signal_4828) ) ;
    buf_clk cell_2984 ( .C (clk), .D (signal_4833), .Q (signal_4834) ) ;
    buf_clk cell_2990 ( .C (clk), .D (signal_4839), .Q (signal_4840) ) ;
    buf_clk cell_2996 ( .C (clk), .D (signal_4845), .Q (signal_4846) ) ;
    buf_clk cell_3002 ( .C (clk), .D (signal_4851), .Q (signal_4852) ) ;
    buf_clk cell_3008 ( .C (clk), .D (signal_4857), .Q (signal_4858) ) ;
    buf_clk cell_3014 ( .C (clk), .D (signal_4863), .Q (signal_4864) ) ;
    buf_clk cell_3020 ( .C (clk), .D (signal_4869), .Q (signal_4870) ) ;
    buf_clk cell_3026 ( .C (clk), .D (signal_4875), .Q (signal_4876) ) ;
    buf_clk cell_3032 ( .C (clk), .D (signal_4881), .Q (signal_4882) ) ;
    buf_clk cell_3038 ( .C (clk), .D (signal_4887), .Q (signal_4888) ) ;
    buf_clk cell_3044 ( .C (clk), .D (signal_4893), .Q (signal_4894) ) ;
    buf_clk cell_3050 ( .C (clk), .D (signal_4899), .Q (signal_4900) ) ;
    buf_clk cell_3056 ( .C (clk), .D (signal_4905), .Q (signal_4906) ) ;
    buf_clk cell_3062 ( .C (clk), .D (signal_4911), .Q (signal_4912) ) ;
    buf_clk cell_3068 ( .C (clk), .D (signal_4917), .Q (signal_4918) ) ;
    buf_clk cell_3074 ( .C (clk), .D (signal_4923), .Q (signal_4924) ) ;
    buf_clk cell_3080 ( .C (clk), .D (signal_4929), .Q (signal_4930) ) ;
    buf_clk cell_3086 ( .C (clk), .D (signal_4935), .Q (signal_4936) ) ;
    buf_clk cell_3092 ( .C (clk), .D (signal_4941), .Q (signal_4942) ) ;
    buf_clk cell_3098 ( .C (clk), .D (signal_4947), .Q (signal_4948) ) ;
    buf_clk cell_3104 ( .C (clk), .D (signal_4953), .Q (signal_4954) ) ;
    buf_clk cell_3110 ( .C (clk), .D (signal_4959), .Q (signal_4960) ) ;
    buf_clk cell_3116 ( .C (clk), .D (signal_4965), .Q (signal_4966) ) ;
    buf_clk cell_3122 ( .C (clk), .D (signal_4971), .Q (signal_4972) ) ;
    buf_clk cell_3130 ( .C (clk), .D (signal_4979), .Q (signal_4980) ) ;
    buf_clk cell_3138 ( .C (clk), .D (signal_4987), .Q (signal_4988) ) ;
    buf_clk cell_3146 ( .C (clk), .D (signal_4995), .Q (signal_4996) ) ;
    buf_clk cell_3154 ( .C (clk), .D (signal_5003), .Q (signal_5004) ) ;
    buf_clk cell_3162 ( .C (clk), .D (signal_5011), .Q (signal_5012) ) ;
    buf_clk cell_3170 ( .C (clk), .D (signal_5019), .Q (signal_5020) ) ;
    buf_clk cell_3178 ( .C (clk), .D (signal_5027), .Q (signal_5028) ) ;
    buf_clk cell_3186 ( .C (clk), .D (signal_5035), .Q (signal_5036) ) ;
    buf_clk cell_3194 ( .C (clk), .D (signal_5043), .Q (signal_5044) ) ;
    buf_clk cell_3202 ( .C (clk), .D (signal_5051), .Q (signal_5052) ) ;
    buf_clk cell_3210 ( .C (clk), .D (signal_5059), .Q (signal_5060) ) ;
    buf_clk cell_3218 ( .C (clk), .D (signal_5067), .Q (signal_5068) ) ;
    buf_clk cell_3226 ( .C (clk), .D (signal_5075), .Q (signal_5076) ) ;
    buf_clk cell_3234 ( .C (clk), .D (signal_5083), .Q (signal_5084) ) ;
    buf_clk cell_3242 ( .C (clk), .D (signal_5091), .Q (signal_5092) ) ;
    buf_clk cell_3250 ( .C (clk), .D (signal_5099), .Q (signal_5100) ) ;
    buf_clk cell_3258 ( .C (clk), .D (signal_5107), .Q (signal_5108) ) ;
    buf_clk cell_3266 ( .C (clk), .D (signal_5115), .Q (signal_5116) ) ;
    buf_clk cell_3274 ( .C (clk), .D (signal_5123), .Q (signal_5124) ) ;
    buf_clk cell_3282 ( .C (clk), .D (signal_5131), .Q (signal_5132) ) ;
    buf_clk cell_3290 ( .C (clk), .D (signal_5139), .Q (signal_5140) ) ;
    buf_clk cell_3298 ( .C (clk), .D (signal_5147), .Q (signal_5148) ) ;
    buf_clk cell_3306 ( .C (clk), .D (signal_5155), .Q (signal_5156) ) ;
    buf_clk cell_3314 ( .C (clk), .D (signal_5163), .Q (signal_5164) ) ;
    buf_clk cell_3322 ( .C (clk), .D (signal_5171), .Q (signal_5172) ) ;
    buf_clk cell_3330 ( .C (clk), .D (signal_5179), .Q (signal_5180) ) ;
    buf_clk cell_3338 ( .C (clk), .D (signal_5187), .Q (signal_5188) ) ;
    buf_clk cell_3346 ( .C (clk), .D (signal_5195), .Q (signal_5196) ) ;
    buf_clk cell_3354 ( .C (clk), .D (signal_5203), .Q (signal_5204) ) ;
    buf_clk cell_3362 ( .C (clk), .D (signal_5211), .Q (signal_5212) ) ;
    buf_clk cell_3370 ( .C (clk), .D (signal_5219), .Q (signal_5220) ) ;
    buf_clk cell_3378 ( .C (clk), .D (signal_5227), .Q (signal_5228) ) ;
    buf_clk cell_3386 ( .C (clk), .D (signal_5235), .Q (signal_5236) ) ;
    buf_clk cell_3394 ( .C (clk), .D (signal_5243), .Q (signal_5244) ) ;
    buf_clk cell_3402 ( .C (clk), .D (signal_5251), .Q (signal_5252) ) ;
    buf_clk cell_3410 ( .C (clk), .D (signal_5259), .Q (signal_5260) ) ;
    buf_clk cell_3418 ( .C (clk), .D (signal_5267), .Q (signal_5268) ) ;
    buf_clk cell_3426 ( .C (clk), .D (signal_5275), .Q (signal_5276) ) ;
    buf_clk cell_3434 ( .C (clk), .D (signal_5283), .Q (signal_5284) ) ;
    buf_clk cell_3442 ( .C (clk), .D (signal_5291), .Q (signal_5292) ) ;
    buf_clk cell_3450 ( .C (clk), .D (signal_5299), .Q (signal_5300) ) ;
    buf_clk cell_3458 ( .C (clk), .D (signal_5307), .Q (signal_5308) ) ;
    buf_clk cell_3466 ( .C (clk), .D (signal_5315), .Q (signal_5316) ) ;
    buf_clk cell_3474 ( .C (clk), .D (signal_5323), .Q (signal_5324) ) ;
    buf_clk cell_3482 ( .C (clk), .D (signal_5331), .Q (signal_5332) ) ;
    buf_clk cell_3490 ( .C (clk), .D (signal_5339), .Q (signal_5340) ) ;
    buf_clk cell_3498 ( .C (clk), .D (signal_5347), .Q (signal_5348) ) ;
    buf_clk cell_3506 ( .C (clk), .D (signal_5355), .Q (signal_5356) ) ;
    buf_clk cell_3514 ( .C (clk), .D (signal_5363), .Q (signal_5364) ) ;
    buf_clk cell_3522 ( .C (clk), .D (signal_5371), .Q (signal_5372) ) ;
    buf_clk cell_3530 ( .C (clk), .D (signal_5379), .Q (signal_5380) ) ;
    buf_clk cell_3538 ( .C (clk), .D (signal_5387), .Q (signal_5388) ) ;
    buf_clk cell_3546 ( .C (clk), .D (signal_5395), .Q (signal_5396) ) ;
    buf_clk cell_3554 ( .C (clk), .D (signal_5403), .Q (signal_5404) ) ;
    buf_clk cell_3562 ( .C (clk), .D (signal_5411), .Q (signal_5412) ) ;
    buf_clk cell_3570 ( .C (clk), .D (signal_5419), .Q (signal_5420) ) ;
    buf_clk cell_3578 ( .C (clk), .D (signal_5427), .Q (signal_5428) ) ;
    buf_clk cell_3586 ( .C (clk), .D (signal_5435), .Q (signal_5436) ) ;
    buf_clk cell_3594 ( .C (clk), .D (signal_5443), .Q (signal_5444) ) ;
    buf_clk cell_3602 ( .C (clk), .D (signal_5451), .Q (signal_5452) ) ;
    buf_clk cell_3610 ( .C (clk), .D (signal_5459), .Q (signal_5460) ) ;
    buf_clk cell_3618 ( .C (clk), .D (signal_5467), .Q (signal_5468) ) ;
    buf_clk cell_3626 ( .C (clk), .D (signal_5475), .Q (signal_5476) ) ;
    buf_clk cell_3634 ( .C (clk), .D (signal_5483), .Q (signal_5484) ) ;
    buf_clk cell_3642 ( .C (clk), .D (signal_5491), .Q (signal_5492) ) ;
    buf_clk cell_3650 ( .C (clk), .D (signal_5499), .Q (signal_5500) ) ;
    buf_clk cell_3658 ( .C (clk), .D (signal_5507), .Q (signal_5508) ) ;
    buf_clk cell_3666 ( .C (clk), .D (signal_5515), .Q (signal_5516) ) ;
    buf_clk cell_3674 ( .C (clk), .D (signal_5523), .Q (signal_5524) ) ;
    buf_clk cell_3682 ( .C (clk), .D (signal_5531), .Q (signal_5532) ) ;
    buf_clk cell_3690 ( .C (clk), .D (signal_5539), .Q (signal_5540) ) ;
    buf_clk cell_3698 ( .C (clk), .D (signal_5547), .Q (signal_5548) ) ;
    buf_clk cell_3706 ( .C (clk), .D (signal_5555), .Q (signal_5556) ) ;
    buf_clk cell_3714 ( .C (clk), .D (signal_5563), .Q (signal_5564) ) ;
    buf_clk cell_3722 ( .C (clk), .D (signal_5571), .Q (signal_5572) ) ;
    buf_clk cell_3730 ( .C (clk), .D (signal_5579), .Q (signal_5580) ) ;
    buf_clk cell_3738 ( .C (clk), .D (signal_5587), .Q (signal_5588) ) ;
    buf_clk cell_3746 ( .C (clk), .D (signal_5595), .Q (signal_5596) ) ;
    buf_clk cell_3754 ( .C (clk), .D (signal_5603), .Q (signal_5604) ) ;
    buf_clk cell_3762 ( .C (clk), .D (signal_5611), .Q (signal_5612) ) ;
    buf_clk cell_3770 ( .C (clk), .D (signal_5619), .Q (signal_5620) ) ;
    buf_clk cell_3778 ( .C (clk), .D (signal_5627), .Q (signal_5628) ) ;
    buf_clk cell_3786 ( .C (clk), .D (signal_5635), .Q (signal_5636) ) ;
    buf_clk cell_3794 ( .C (clk), .D (signal_5643), .Q (signal_5644) ) ;
    buf_clk cell_3802 ( .C (clk), .D (signal_5651), .Q (signal_5652) ) ;
    buf_clk cell_3810 ( .C (clk), .D (signal_5659), .Q (signal_5660) ) ;
    buf_clk cell_3818 ( .C (clk), .D (signal_5667), .Q (signal_5668) ) ;
    buf_clk cell_3826 ( .C (clk), .D (signal_5675), .Q (signal_5676) ) ;
    buf_clk cell_3834 ( .C (clk), .D (signal_5683), .Q (signal_5684) ) ;
    buf_clk cell_3842 ( .C (clk), .D (signal_5691), .Q (signal_5692) ) ;
    buf_clk cell_3850 ( .C (clk), .D (signal_5699), .Q (signal_5700) ) ;
    buf_clk cell_3858 ( .C (clk), .D (signal_5707), .Q (signal_5708) ) ;
    buf_clk cell_3866 ( .C (clk), .D (signal_5715), .Q (signal_5716) ) ;
    buf_clk cell_3874 ( .C (clk), .D (signal_5723), .Q (signal_5724) ) ;
    buf_clk cell_3882 ( .C (clk), .D (signal_5731), .Q (signal_5732) ) ;
    buf_clk cell_3890 ( .C (clk), .D (signal_5739), .Q (signal_5740) ) ;
    buf_clk cell_3898 ( .C (clk), .D (signal_5747), .Q (signal_5748) ) ;
    buf_clk cell_3906 ( .C (clk), .D (signal_5755), .Q (signal_5756) ) ;
    buf_clk cell_3914 ( .C (clk), .D (signal_5763), .Q (signal_5764) ) ;
    buf_clk cell_3922 ( .C (clk), .D (signal_5771), .Q (signal_5772) ) ;
    buf_clk cell_3930 ( .C (clk), .D (signal_5779), .Q (signal_5780) ) ;
    buf_clk cell_3938 ( .C (clk), .D (signal_5787), .Q (signal_5788) ) ;
    buf_clk cell_3946 ( .C (clk), .D (signal_5795), .Q (signal_5796) ) ;
    buf_clk cell_3954 ( .C (clk), .D (signal_5803), .Q (signal_5804) ) ;
    buf_clk cell_3962 ( .C (clk), .D (signal_5811), .Q (signal_5812) ) ;
    buf_clk cell_3970 ( .C (clk), .D (signal_5819), .Q (signal_5820) ) ;
    buf_clk cell_3978 ( .C (clk), .D (signal_5827), .Q (signal_5828) ) ;
    buf_clk cell_3986 ( .C (clk), .D (signal_5835), .Q (signal_5836) ) ;
    buf_clk cell_3994 ( .C (clk), .D (signal_5843), .Q (signal_5844) ) ;
    buf_clk cell_4002 ( .C (clk), .D (signal_5851), .Q (signal_5852) ) ;
    buf_clk cell_4010 ( .C (clk), .D (signal_5859), .Q (signal_5860) ) ;
    buf_clk cell_4018 ( .C (clk), .D (signal_5867), .Q (signal_5868) ) ;
    buf_clk cell_4026 ( .C (clk), .D (signal_5875), .Q (signal_5876) ) ;
    buf_clk cell_4034 ( .C (clk), .D (signal_5883), .Q (signal_5884) ) ;
    buf_clk cell_4042 ( .C (clk), .D (signal_5891), .Q (signal_5892) ) ;
    buf_clk cell_4050 ( .C (clk), .D (signal_5899), .Q (signal_5900) ) ;
    buf_clk cell_4058 ( .C (clk), .D (signal_5907), .Q (signal_5908) ) ;
    buf_clk cell_4066 ( .C (clk), .D (signal_5915), .Q (signal_5916) ) ;
    buf_clk cell_4074 ( .C (clk), .D (signal_5923), .Q (signal_5924) ) ;
    buf_clk cell_4082 ( .C (clk), .D (signal_5931), .Q (signal_5932) ) ;
    buf_clk cell_4090 ( .C (clk), .D (signal_5939), .Q (signal_5940) ) ;
    buf_clk cell_4098 ( .C (clk), .D (signal_5947), .Q (signal_5948) ) ;
    buf_clk cell_4106 ( .C (clk), .D (signal_5955), .Q (signal_5956) ) ;
    buf_clk cell_4114 ( .C (clk), .D (signal_5963), .Q (signal_5964) ) ;
    buf_clk cell_4122 ( .C (clk), .D (signal_5971), .Q (signal_5972) ) ;
    buf_clk cell_4130 ( .C (clk), .D (signal_5979), .Q (signal_5980) ) ;
    buf_clk cell_4138 ( .C (clk), .D (signal_5987), .Q (signal_5988) ) ;
    buf_clk cell_4146 ( .C (clk), .D (signal_5995), .Q (signal_5996) ) ;
    buf_clk cell_4154 ( .C (clk), .D (signal_6003), .Q (signal_6004) ) ;
    buf_clk cell_4162 ( .C (clk), .D (signal_6011), .Q (signal_6012) ) ;
    buf_clk cell_4170 ( .C (clk), .D (signal_6019), .Q (signal_6020) ) ;
    buf_clk cell_4178 ( .C (clk), .D (signal_6027), .Q (signal_6028) ) ;
    buf_clk cell_4186 ( .C (clk), .D (signal_6035), .Q (signal_6036) ) ;
    buf_clk cell_4194 ( .C (clk), .D (signal_6043), .Q (signal_6044) ) ;
    buf_clk cell_4202 ( .C (clk), .D (signal_6051), .Q (signal_6052) ) ;
    buf_clk cell_4210 ( .C (clk), .D (signal_6059), .Q (signal_6060) ) ;
    buf_clk cell_4218 ( .C (clk), .D (signal_6067), .Q (signal_6068) ) ;
    buf_clk cell_4226 ( .C (clk), .D (signal_6075), .Q (signal_6076) ) ;
    buf_clk cell_4234 ( .C (clk), .D (signal_6083), .Q (signal_6084) ) ;
    buf_clk cell_4242 ( .C (clk), .D (signal_6091), .Q (signal_6092) ) ;
    buf_clk cell_4250 ( .C (clk), .D (signal_6099), .Q (signal_6100) ) ;
    buf_clk cell_4258 ( .C (clk), .D (signal_6107), .Q (signal_6108) ) ;
    buf_clk cell_4266 ( .C (clk), .D (signal_6115), .Q (signal_6116) ) ;
    buf_clk cell_4274 ( .C (clk), .D (signal_6123), .Q (signal_6124) ) ;
    buf_clk cell_4282 ( .C (clk), .D (signal_6131), .Q (signal_6132) ) ;
    buf_clk cell_4290 ( .C (clk), .D (signal_6139), .Q (signal_6140) ) ;
    buf_clk cell_4298 ( .C (clk), .D (signal_6147), .Q (signal_6148) ) ;
    buf_clk cell_4306 ( .C (clk), .D (signal_6155), .Q (signal_6156) ) ;
    buf_clk cell_4314 ( .C (clk), .D (signal_6163), .Q (signal_6164) ) ;
    buf_clk cell_4322 ( .C (clk), .D (signal_6171), .Q (signal_6172) ) ;
    buf_clk cell_4330 ( .C (clk), .D (signal_6179), .Q (signal_6180) ) ;
    buf_clk cell_4338 ( .C (clk), .D (signal_6187), .Q (signal_6188) ) ;
    buf_clk cell_4346 ( .C (clk), .D (signal_6195), .Q (signal_6196) ) ;
    buf_clk cell_4354 ( .C (clk), .D (signal_6203), .Q (signal_6204) ) ;
    buf_clk cell_4362 ( .C (clk), .D (signal_6211), .Q (signal_6212) ) ;
    buf_clk cell_4370 ( .C (clk), .D (signal_6219), .Q (signal_6220) ) ;
    buf_clk cell_4378 ( .C (clk), .D (signal_6227), .Q (signal_6228) ) ;
    buf_clk cell_4386 ( .C (clk), .D (signal_6235), .Q (signal_6236) ) ;
    buf_clk cell_4394 ( .C (clk), .D (signal_6243), .Q (signal_6244) ) ;
    buf_clk cell_4402 ( .C (clk), .D (signal_6251), .Q (signal_6252) ) ;
    buf_clk cell_4410 ( .C (clk), .D (signal_6259), .Q (signal_6260) ) ;
    buf_clk cell_4418 ( .C (clk), .D (signal_6267), .Q (signal_6268) ) ;
    buf_clk cell_4426 ( .C (clk), .D (signal_6275), .Q (signal_6276) ) ;
    buf_clk cell_4434 ( .C (clk), .D (signal_6283), .Q (signal_6284) ) ;
    buf_clk cell_4442 ( .C (clk), .D (signal_6291), .Q (signal_6292) ) ;
    buf_clk cell_4450 ( .C (clk), .D (signal_6299), .Q (signal_6300) ) ;
    buf_clk cell_4458 ( .C (clk), .D (signal_6307), .Q (signal_6308) ) ;
    buf_clk cell_4466 ( .C (clk), .D (signal_6315), .Q (signal_6316) ) ;
    buf_clk cell_4474 ( .C (clk), .D (signal_6323), .Q (signal_6324) ) ;
    buf_clk cell_4482 ( .C (clk), .D (signal_6331), .Q (signal_6332) ) ;
    buf_clk cell_4490 ( .C (clk), .D (signal_6339), .Q (signal_6340) ) ;
    buf_clk cell_4498 ( .C (clk), .D (signal_6347), .Q (signal_6348) ) ;
    buf_clk cell_4506 ( .C (clk), .D (signal_6355), .Q (signal_6356) ) ;
    buf_clk cell_4514 ( .C (clk), .D (signal_6363), .Q (signal_6364) ) ;
    buf_clk cell_4522 ( .C (clk), .D (signal_6371), .Q (signal_6372) ) ;
    buf_clk cell_4530 ( .C (clk), .D (signal_6379), .Q (signal_6380) ) ;
    buf_clk cell_4538 ( .C (clk), .D (signal_6387), .Q (signal_6388) ) ;
    buf_clk cell_4546 ( .C (clk), .D (signal_6395), .Q (signal_6396) ) ;
    buf_clk cell_4554 ( .C (clk), .D (signal_6403), .Q (signal_6404) ) ;
    buf_clk cell_4562 ( .C (clk), .D (signal_6411), .Q (signal_6412) ) ;
    buf_clk cell_4570 ( .C (clk), .D (signal_6419), .Q (signal_6420) ) ;
    buf_clk cell_4578 ( .C (clk), .D (signal_6427), .Q (signal_6428) ) ;
    buf_clk cell_4586 ( .C (clk), .D (signal_6435), .Q (signal_6436) ) ;
    buf_clk cell_4594 ( .C (clk), .D (signal_6443), .Q (signal_6444) ) ;
    buf_clk cell_4602 ( .C (clk), .D (signal_6451), .Q (signal_6452) ) ;
    buf_clk cell_4610 ( .C (clk), .D (signal_6459), .Q (signal_6460) ) ;
    buf_clk cell_4618 ( .C (clk), .D (signal_6467), .Q (signal_6468) ) ;
    buf_clk cell_4626 ( .C (clk), .D (signal_6475), .Q (signal_6476) ) ;
    buf_clk cell_4634 ( .C (clk), .D (signal_6483), .Q (signal_6484) ) ;
    buf_clk cell_4642 ( .C (clk), .D (signal_6491), .Q (signal_6492) ) ;
    buf_clk cell_4650 ( .C (clk), .D (signal_6499), .Q (signal_6500) ) ;
    buf_clk cell_4658 ( .C (clk), .D (signal_6507), .Q (signal_6508) ) ;
    buf_clk cell_4666 ( .C (clk), .D (signal_6515), .Q (signal_6516) ) ;
    buf_clk cell_4674 ( .C (clk), .D (signal_6523), .Q (signal_6524) ) ;
    buf_clk cell_4682 ( .C (clk), .D (signal_6531), .Q (signal_6532) ) ;
    buf_clk cell_4690 ( .C (clk), .D (signal_6539), .Q (signal_6540) ) ;
    buf_clk cell_4698 ( .C (clk), .D (signal_6547), .Q (signal_6548) ) ;
    buf_clk cell_4706 ( .C (clk), .D (signal_6555), .Q (signal_6556) ) ;
    buf_clk cell_4714 ( .C (clk), .D (signal_6563), .Q (signal_6564) ) ;
    buf_clk cell_4722 ( .C (clk), .D (signal_6571), .Q (signal_6572) ) ;
    buf_clk cell_4730 ( .C (clk), .D (signal_6579), .Q (signal_6580) ) ;
    buf_clk cell_4738 ( .C (clk), .D (signal_6587), .Q (signal_6588) ) ;
    buf_clk cell_4746 ( .C (clk), .D (signal_6595), .Q (signal_6596) ) ;
    buf_clk cell_4754 ( .C (clk), .D (signal_6603), .Q (signal_6604) ) ;
    buf_clk cell_4762 ( .C (clk), .D (signal_6611), .Q (signal_6612) ) ;
    buf_clk cell_4770 ( .C (clk), .D (signal_6619), .Q (signal_6620) ) ;
    buf_clk cell_4778 ( .C (clk), .D (signal_6627), .Q (signal_6628) ) ;
    buf_clk cell_4786 ( .C (clk), .D (signal_6635), .Q (signal_6636) ) ;
    buf_clk cell_4794 ( .C (clk), .D (signal_6643), .Q (signal_6644) ) ;
    buf_clk cell_4802 ( .C (clk), .D (signal_6651), .Q (signal_6652) ) ;
    buf_clk cell_4810 ( .C (clk), .D (signal_6659), .Q (signal_6660) ) ;
    buf_clk cell_4818 ( .C (clk), .D (signal_6667), .Q (signal_6668) ) ;
    buf_clk cell_4826 ( .C (clk), .D (signal_6675), .Q (signal_6676) ) ;
    buf_clk cell_4834 ( .C (clk), .D (signal_6683), .Q (signal_6684) ) ;
    buf_clk cell_4842 ( .C (clk), .D (signal_6691), .Q (signal_6692) ) ;
    buf_clk cell_4850 ( .C (clk), .D (signal_6699), .Q (signal_6700) ) ;
    buf_clk cell_4858 ( .C (clk), .D (signal_6707), .Q (signal_6708) ) ;
    buf_clk cell_4866 ( .C (clk), .D (signal_6715), .Q (signal_6716) ) ;
    buf_clk cell_4874 ( .C (clk), .D (signal_6723), .Q (signal_6724) ) ;
    buf_clk cell_4882 ( .C (clk), .D (signal_6731), .Q (signal_6732) ) ;
    buf_clk cell_4890 ( .C (clk), .D (signal_6739), .Q (signal_6740) ) ;
    buf_clk cell_4898 ( .C (clk), .D (signal_6747), .Q (signal_6748) ) ;
    buf_clk cell_4906 ( .C (clk), .D (signal_6755), .Q (signal_6756) ) ;
    buf_clk cell_4914 ( .C (clk), .D (signal_6763), .Q (signal_6764) ) ;
    buf_clk cell_4922 ( .C (clk), .D (signal_6771), .Q (signal_6772) ) ;
    buf_clk cell_4930 ( .C (clk), .D (signal_6779), .Q (signal_6780) ) ;
    buf_clk cell_4938 ( .C (clk), .D (signal_6787), .Q (signal_6788) ) ;
    buf_clk cell_4946 ( .C (clk), .D (signal_6795), .Q (signal_6796) ) ;
    buf_clk cell_4954 ( .C (clk), .D (signal_6803), .Q (signal_6804) ) ;
    buf_clk cell_4962 ( .C (clk), .D (signal_6811), .Q (signal_6812) ) ;
    buf_clk cell_4970 ( .C (clk), .D (signal_6819), .Q (signal_6820) ) ;
    buf_clk cell_4978 ( .C (clk), .D (signal_6827), .Q (signal_6828) ) ;
    buf_clk cell_4986 ( .C (clk), .D (signal_6835), .Q (signal_6836) ) ;
    buf_clk cell_4994 ( .C (clk), .D (signal_6843), .Q (signal_6844) ) ;
    buf_clk cell_5002 ( .C (clk), .D (signal_6851), .Q (signal_6852) ) ;
    buf_clk cell_5010 ( .C (clk), .D (signal_6859), .Q (signal_6860) ) ;
    buf_clk cell_5018 ( .C (clk), .D (signal_6867), .Q (signal_6868) ) ;
    buf_clk cell_5026 ( .C (clk), .D (signal_6875), .Q (signal_6876) ) ;
    buf_clk cell_5034 ( .C (clk), .D (signal_6883), .Q (signal_6884) ) ;
    buf_clk cell_5042 ( .C (clk), .D (signal_6891), .Q (signal_6892) ) ;
    buf_clk cell_5050 ( .C (clk), .D (signal_6899), .Q (signal_6900) ) ;
    buf_clk cell_5058 ( .C (clk), .D (signal_6907), .Q (signal_6908) ) ;
    buf_clk cell_5066 ( .C (clk), .D (signal_6915), .Q (signal_6916) ) ;
    buf_clk cell_5074 ( .C (clk), .D (signal_6923), .Q (signal_6924) ) ;
    buf_clk cell_5082 ( .C (clk), .D (signal_6931), .Q (signal_6932) ) ;
    buf_clk cell_5090 ( .C (clk), .D (signal_6939), .Q (signal_6940) ) ;
    buf_clk cell_5098 ( .C (clk), .D (signal_6947), .Q (signal_6948) ) ;
    buf_clk cell_5106 ( .C (clk), .D (signal_6955), .Q (signal_6956) ) ;
    buf_clk cell_5114 ( .C (clk), .D (signal_6963), .Q (signal_6964) ) ;
    buf_clk cell_5122 ( .C (clk), .D (signal_6971), .Q (signal_6972) ) ;
    buf_clk cell_5130 ( .C (clk), .D (signal_6979), .Q (signal_6980) ) ;
    buf_clk cell_5138 ( .C (clk), .D (signal_6987), .Q (signal_6988) ) ;
    buf_clk cell_5146 ( .C (clk), .D (signal_6995), .Q (signal_6996) ) ;
    buf_clk cell_5154 ( .C (clk), .D (signal_7003), .Q (signal_7004) ) ;
    buf_clk cell_5162 ( .C (clk), .D (signal_7011), .Q (signal_7012) ) ;
    buf_clk cell_5170 ( .C (clk), .D (signal_7019), .Q (signal_7020) ) ;
    buf_clk cell_5178 ( .C (clk), .D (signal_7027), .Q (signal_7028) ) ;
    buf_clk cell_5186 ( .C (clk), .D (signal_7035), .Q (signal_7036) ) ;
    buf_clk cell_5194 ( .C (clk), .D (signal_7043), .Q (signal_7044) ) ;
    buf_clk cell_5202 ( .C (clk), .D (signal_7051), .Q (signal_7052) ) ;
    buf_clk cell_5210 ( .C (clk), .D (signal_7059), .Q (signal_7060) ) ;
    buf_clk cell_5218 ( .C (clk), .D (signal_7067), .Q (signal_7068) ) ;
    buf_clk cell_5226 ( .C (clk), .D (signal_7075), .Q (signal_7076) ) ;
    buf_clk cell_5234 ( .C (clk), .D (signal_7083), .Q (signal_7084) ) ;
    buf_clk cell_5242 ( .C (clk), .D (signal_7091), .Q (signal_7092) ) ;
    buf_clk cell_5250 ( .C (clk), .D (signal_7099), .Q (signal_7100) ) ;
    buf_clk cell_5258 ( .C (clk), .D (signal_7107), .Q (signal_7108) ) ;
    buf_clk cell_5266 ( .C (clk), .D (signal_7115), .Q (signal_7116) ) ;
    buf_clk cell_5274 ( .C (clk), .D (signal_7123), .Q (signal_7124) ) ;
    buf_clk cell_5282 ( .C (clk), .D (signal_7131), .Q (signal_7132) ) ;
    buf_clk cell_5290 ( .C (clk), .D (signal_7139), .Q (signal_7140) ) ;
    buf_clk cell_5298 ( .C (clk), .D (signal_7147), .Q (signal_7148) ) ;
    buf_clk cell_5306 ( .C (clk), .D (signal_7155), .Q (signal_7156) ) ;
    buf_clk cell_5314 ( .C (clk), .D (signal_7163), .Q (signal_7164) ) ;
    buf_clk cell_5322 ( .C (clk), .D (signal_7171), .Q (signal_7172) ) ;
    buf_clk cell_5330 ( .C (clk), .D (signal_7179), .Q (signal_7180) ) ;
    buf_clk cell_5338 ( .C (clk), .D (signal_7187), .Q (signal_7188) ) ;
    buf_clk cell_5346 ( .C (clk), .D (signal_7195), .Q (signal_7196) ) ;
    buf_clk cell_5354 ( .C (clk), .D (signal_7203), .Q (signal_7204) ) ;
    buf_clk cell_5362 ( .C (clk), .D (signal_7211), .Q (signal_7212) ) ;
    buf_clk cell_5370 ( .C (clk), .D (signal_7219), .Q (signal_7220) ) ;
    buf_clk cell_5378 ( .C (clk), .D (signal_7227), .Q (signal_7228) ) ;
    buf_clk cell_5386 ( .C (clk), .D (signal_7235), .Q (signal_7236) ) ;
    buf_clk cell_5394 ( .C (clk), .D (signal_7243), .Q (signal_7244) ) ;
    buf_clk cell_5402 ( .C (clk), .D (signal_7251), .Q (signal_7252) ) ;
    buf_clk cell_5410 ( .C (clk), .D (signal_7259), .Q (signal_7260) ) ;
    buf_clk cell_5418 ( .C (clk), .D (signal_7267), .Q (signal_7268) ) ;
    buf_clk cell_5426 ( .C (clk), .D (signal_7275), .Q (signal_7276) ) ;
    buf_clk cell_5434 ( .C (clk), .D (signal_7283), .Q (signal_7284) ) ;
    buf_clk cell_5442 ( .C (clk), .D (signal_7291), .Q (signal_7292) ) ;
    buf_clk cell_5450 ( .C (clk), .D (signal_7299), .Q (signal_7300) ) ;
    buf_clk cell_5458 ( .C (clk), .D (signal_7307), .Q (signal_7308) ) ;
    buf_clk cell_5466 ( .C (clk), .D (signal_7315), .Q (signal_7316) ) ;
    buf_clk cell_5474 ( .C (clk), .D (signal_7323), .Q (signal_7324) ) ;
    buf_clk cell_5482 ( .C (clk), .D (signal_7331), .Q (signal_7332) ) ;
    buf_clk cell_5490 ( .C (clk), .D (signal_7339), .Q (signal_7340) ) ;
    buf_clk cell_5498 ( .C (clk), .D (signal_7347), .Q (signal_7348) ) ;
    buf_clk cell_5506 ( .C (clk), .D (signal_7355), .Q (signal_7356) ) ;
    buf_clk cell_5514 ( .C (clk), .D (signal_7363), .Q (signal_7364) ) ;
    buf_clk cell_5522 ( .C (clk), .D (signal_7371), .Q (signal_7372) ) ;
    buf_clk cell_5530 ( .C (clk), .D (signal_7379), .Q (signal_7380) ) ;
    buf_clk cell_5538 ( .C (clk), .D (signal_7387), .Q (signal_7388) ) ;
    buf_clk cell_5546 ( .C (clk), .D (signal_7395), .Q (signal_7396) ) ;
    buf_clk cell_5554 ( .C (clk), .D (signal_7403), .Q (signal_7404) ) ;
    buf_clk cell_5562 ( .C (clk), .D (signal_7411), .Q (signal_7412) ) ;
    buf_clk cell_5570 ( .C (clk), .D (signal_7419), .Q (signal_7420) ) ;
    buf_clk cell_5578 ( .C (clk), .D (signal_7427), .Q (signal_7428) ) ;
    buf_clk cell_5586 ( .C (clk), .D (signal_7435), .Q (signal_7436) ) ;
    buf_clk cell_5594 ( .C (clk), .D (signal_7443), .Q (signal_7444) ) ;
    buf_clk cell_5602 ( .C (clk), .D (signal_7451), .Q (signal_7452) ) ;
    buf_clk cell_5610 ( .C (clk), .D (signal_7459), .Q (signal_7460) ) ;
    buf_clk cell_5618 ( .C (clk), .D (signal_7467), .Q (signal_7468) ) ;
    buf_clk cell_5626 ( .C (clk), .D (signal_7475), .Q (signal_7476) ) ;
    buf_clk cell_5634 ( .C (clk), .D (signal_7483), .Q (signal_7484) ) ;
    buf_clk cell_5642 ( .C (clk), .D (signal_7491), .Q (signal_7492) ) ;
    buf_clk cell_5650 ( .C (clk), .D (signal_7499), .Q (signal_7500) ) ;
    buf_clk cell_5658 ( .C (clk), .D (signal_7507), .Q (signal_7508) ) ;
    buf_clk cell_5666 ( .C (clk), .D (signal_7515), .Q (signal_7516) ) ;
    buf_clk cell_5674 ( .C (clk), .D (signal_7523), .Q (signal_7524) ) ;
    buf_clk cell_5682 ( .C (clk), .D (signal_7531), .Q (signal_7532) ) ;
    buf_clk cell_5690 ( .C (clk), .D (signal_7539), .Q (signal_7540) ) ;
    buf_clk cell_5698 ( .C (clk), .D (signal_7547), .Q (signal_7548) ) ;
    buf_clk cell_5706 ( .C (clk), .D (signal_7555), .Q (signal_7556) ) ;
    buf_clk cell_5714 ( .C (clk), .D (signal_7563), .Q (signal_7564) ) ;
    buf_clk cell_5722 ( .C (clk), .D (signal_7571), .Q (signal_7572) ) ;
    buf_clk cell_5730 ( .C (clk), .D (signal_7579), .Q (signal_7580) ) ;
    buf_clk cell_5738 ( .C (clk), .D (signal_7587), .Q (signal_7588) ) ;
    buf_clk cell_5746 ( .C (clk), .D (signal_7595), .Q (signal_7596) ) ;
    buf_clk cell_5754 ( .C (clk), .D (signal_7603), .Q (signal_7604) ) ;
    buf_clk cell_5762 ( .C (clk), .D (signal_7611), .Q (signal_7612) ) ;
    buf_clk cell_5770 ( .C (clk), .D (signal_7619), .Q (signal_7620) ) ;
    buf_clk cell_5778 ( .C (clk), .D (signal_7627), .Q (signal_7628) ) ;
    buf_clk cell_5786 ( .C (clk), .D (signal_7635), .Q (signal_7636) ) ;
    buf_clk cell_5794 ( .C (clk), .D (signal_7643), .Q (signal_7644) ) ;
    buf_clk cell_5802 ( .C (clk), .D (signal_7651), .Q (signal_7652) ) ;
    buf_clk cell_5810 ( .C (clk), .D (signal_7659), .Q (signal_7660) ) ;
    buf_clk cell_5818 ( .C (clk), .D (signal_7667), .Q (signal_7668) ) ;
    buf_clk cell_5826 ( .C (clk), .D (signal_7675), .Q (signal_7676) ) ;
    buf_clk cell_5834 ( .C (clk), .D (signal_7683), .Q (signal_7684) ) ;
    buf_clk cell_5842 ( .C (clk), .D (signal_7691), .Q (signal_7692) ) ;
    buf_clk cell_5850 ( .C (clk), .D (signal_7699), .Q (signal_7700) ) ;
    buf_clk cell_5858 ( .C (clk), .D (signal_7707), .Q (signal_7708) ) ;
    buf_clk cell_5866 ( .C (clk), .D (signal_7715), .Q (signal_7716) ) ;
    buf_clk cell_5874 ( .C (clk), .D (signal_7723), .Q (signal_7724) ) ;
    buf_clk cell_5882 ( .C (clk), .D (signal_7731), .Q (signal_7732) ) ;
    buf_clk cell_5890 ( .C (clk), .D (signal_7739), .Q (signal_7740) ) ;
    buf_clk cell_5898 ( .C (clk), .D (signal_7747), .Q (signal_7748) ) ;
    buf_clk cell_5906 ( .C (clk), .D (signal_7755), .Q (signal_7756) ) ;
    buf_clk cell_5914 ( .C (clk), .D (signal_7763), .Q (signal_7764) ) ;
    buf_clk cell_5922 ( .C (clk), .D (signal_7771), .Q (signal_7772) ) ;
    buf_clk cell_5930 ( .C (clk), .D (signal_7779), .Q (signal_7780) ) ;
    buf_clk cell_5938 ( .C (clk), .D (signal_7787), .Q (signal_7788) ) ;
    buf_clk cell_5946 ( .C (clk), .D (signal_7795), .Q (signal_7796) ) ;
    buf_clk cell_5954 ( .C (clk), .D (signal_7803), .Q (signal_7804) ) ;
    buf_clk cell_5962 ( .C (clk), .D (signal_7811), .Q (signal_7812) ) ;
    buf_clk cell_5970 ( .C (clk), .D (signal_7819), .Q (signal_7820) ) ;
    buf_clk cell_5978 ( .C (clk), .D (signal_7827), .Q (signal_7828) ) ;
    buf_clk cell_5986 ( .C (clk), .D (signal_7835), .Q (signal_7836) ) ;
    buf_clk cell_5994 ( .C (clk), .D (signal_7843), .Q (signal_7844) ) ;
    buf_clk cell_6002 ( .C (clk), .D (signal_7851), .Q (signal_7852) ) ;
    buf_clk cell_6010 ( .C (clk), .D (signal_7859), .Q (signal_7860) ) ;
    buf_clk cell_6018 ( .C (clk), .D (signal_7867), .Q (signal_7868) ) ;
    buf_clk cell_6026 ( .C (clk), .D (signal_7875), .Q (signal_7876) ) ;
    buf_clk cell_6034 ( .C (clk), .D (signal_7883), .Q (signal_7884) ) ;
    buf_clk cell_6042 ( .C (clk), .D (signal_7891), .Q (signal_7892) ) ;
    buf_clk cell_6050 ( .C (clk), .D (signal_7899), .Q (signal_7900) ) ;
    buf_clk cell_6058 ( .C (clk), .D (signal_7907), .Q (signal_7908) ) ;
    buf_clk cell_6066 ( .C (clk), .D (signal_7915), .Q (signal_7916) ) ;
    buf_clk cell_6074 ( .C (clk), .D (signal_7923), .Q (signal_7924) ) ;
    buf_clk cell_6082 ( .C (clk), .D (signal_7931), .Q (signal_7932) ) ;
    buf_clk cell_6090 ( .C (clk), .D (signal_7939), .Q (signal_7940) ) ;
    buf_clk cell_6098 ( .C (clk), .D (signal_7947), .Q (signal_7948) ) ;
    buf_clk cell_6106 ( .C (clk), .D (signal_7955), .Q (signal_7956) ) ;
    buf_clk cell_6114 ( .C (clk), .D (signal_7963), .Q (signal_7964) ) ;
    buf_clk cell_6122 ( .C (clk), .D (signal_7971), .Q (signal_7972) ) ;
    buf_clk cell_6130 ( .C (clk), .D (signal_7979), .Q (signal_7980) ) ;
    buf_clk cell_6138 ( .C (clk), .D (signal_7987), .Q (signal_7988) ) ;
    buf_clk cell_6146 ( .C (clk), .D (signal_7995), .Q (signal_7996) ) ;
    buf_clk cell_6154 ( .C (clk), .D (signal_8003), .Q (signal_8004) ) ;
    buf_clk cell_6162 ( .C (clk), .D (signal_8011), .Q (signal_8012) ) ;
    buf_clk cell_6170 ( .C (clk), .D (signal_8019), .Q (signal_8020) ) ;
    buf_clk cell_6178 ( .C (clk), .D (signal_8027), .Q (signal_8028) ) ;
    buf_clk cell_6186 ( .C (clk), .D (signal_8035), .Q (signal_8036) ) ;
    buf_clk cell_6194 ( .C (clk), .D (signal_8043), .Q (signal_8044) ) ;
    buf_clk cell_6202 ( .C (clk), .D (signal_8051), .Q (signal_8052) ) ;
    buf_clk cell_6210 ( .C (clk), .D (signal_8059), .Q (signal_8060) ) ;
    buf_clk cell_6218 ( .C (clk), .D (signal_8067), .Q (signal_8068) ) ;
    buf_clk cell_6226 ( .C (clk), .D (signal_8075), .Q (signal_8076) ) ;
    buf_clk cell_6234 ( .C (clk), .D (signal_8083), .Q (signal_8084) ) ;
    buf_clk cell_6242 ( .C (clk), .D (signal_8091), .Q (signal_8092) ) ;
    buf_clk cell_6250 ( .C (clk), .D (signal_8099), .Q (signal_8100) ) ;
    buf_clk cell_6258 ( .C (clk), .D (signal_8107), .Q (signal_8108) ) ;
    buf_clk cell_6266 ( .C (clk), .D (signal_8115), .Q (signal_8116) ) ;
    buf_clk cell_6274 ( .C (clk), .D (signal_8123), .Q (signal_8124) ) ;
    buf_clk cell_6282 ( .C (clk), .D (signal_8131), .Q (signal_8132) ) ;
    buf_clk cell_6290 ( .C (clk), .D (signal_8139), .Q (signal_8140) ) ;
    buf_clk cell_6298 ( .C (clk), .D (signal_8147), .Q (signal_8148) ) ;
    buf_clk cell_6306 ( .C (clk), .D (signal_8155), .Q (signal_8156) ) ;
    buf_clk cell_6314 ( .C (clk), .D (signal_8163), .Q (signal_8164) ) ;
    buf_clk cell_6322 ( .C (clk), .D (signal_8171), .Q (signal_8172) ) ;
    buf_clk cell_6330 ( .C (clk), .D (signal_8179), .Q (signal_8180) ) ;
    buf_clk cell_6338 ( .C (clk), .D (signal_8187), .Q (signal_8188) ) ;
    buf_clk cell_6346 ( .C (clk), .D (signal_8195), .Q (signal_8196) ) ;
    buf_clk cell_6354 ( .C (clk), .D (signal_8203), .Q (signal_8204) ) ;
    buf_clk cell_6362 ( .C (clk), .D (signal_8211), .Q (signal_8212) ) ;
    buf_clk cell_6370 ( .C (clk), .D (signal_8219), .Q (signal_8220) ) ;
    buf_clk cell_6378 ( .C (clk), .D (signal_8227), .Q (signal_8228) ) ;
    buf_clk cell_6386 ( .C (clk), .D (signal_8235), .Q (signal_8236) ) ;
    buf_clk cell_6394 ( .C (clk), .D (signal_8243), .Q (signal_8244) ) ;
    buf_clk cell_6402 ( .C (clk), .D (signal_8251), .Q (signal_8252) ) ;
    buf_clk cell_6410 ( .C (clk), .D (signal_8259), .Q (signal_8260) ) ;
    buf_clk cell_6418 ( .C (clk), .D (signal_8267), .Q (signal_8268) ) ;
    buf_clk cell_6426 ( .C (clk), .D (signal_8275), .Q (signal_8276) ) ;
    buf_clk cell_6434 ( .C (clk), .D (signal_8283), .Q (signal_8284) ) ;
    buf_clk cell_6442 ( .C (clk), .D (signal_8291), .Q (signal_8292) ) ;
    buf_clk cell_6450 ( .C (clk), .D (signal_8299), .Q (signal_8300) ) ;
    buf_clk cell_6458 ( .C (clk), .D (signal_8307), .Q (signal_8308) ) ;
    buf_clk cell_6466 ( .C (clk), .D (signal_8315), .Q (signal_8316) ) ;
    buf_clk cell_6474 ( .C (clk), .D (signal_8323), .Q (signal_8324) ) ;
    buf_clk cell_6482 ( .C (clk), .D (signal_8331), .Q (signal_8332) ) ;
    buf_clk cell_6490 ( .C (clk), .D (signal_8339), .Q (signal_8340) ) ;
    buf_clk cell_6498 ( .C (clk), .D (signal_8347), .Q (signal_8348) ) ;
    buf_clk cell_6506 ( .C (clk), .D (signal_8355), .Q (signal_8356) ) ;
    buf_clk cell_6514 ( .C (clk), .D (signal_8363), .Q (signal_8364) ) ;
    buf_clk cell_6522 ( .C (clk), .D (signal_8371), .Q (signal_8372) ) ;
    buf_clk cell_6530 ( .C (clk), .D (signal_8379), .Q (signal_8380) ) ;
    buf_clk cell_6538 ( .C (clk), .D (signal_8387), .Q (signal_8388) ) ;
    buf_clk cell_6546 ( .C (clk), .D (signal_8395), .Q (signal_8396) ) ;
    buf_clk cell_6554 ( .C (clk), .D (signal_8403), .Q (signal_8404) ) ;
    buf_clk cell_6562 ( .C (clk), .D (signal_8411), .Q (signal_8412) ) ;
    buf_clk cell_6570 ( .C (clk), .D (signal_8419), .Q (signal_8420) ) ;
    buf_clk cell_6578 ( .C (clk), .D (signal_8427), .Q (signal_8428) ) ;
    buf_clk cell_6586 ( .C (clk), .D (signal_8435), .Q (signal_8436) ) ;
    buf_clk cell_6594 ( .C (clk), .D (signal_8443), .Q (signal_8444) ) ;
    buf_clk cell_6602 ( .C (clk), .D (signal_8451), .Q (signal_8452) ) ;
    buf_clk cell_6610 ( .C (clk), .D (signal_8459), .Q (signal_8460) ) ;
    buf_clk cell_6618 ( .C (clk), .D (signal_8467), .Q (signal_8468) ) ;
    buf_clk cell_6626 ( .C (clk), .D (signal_8475), .Q (signal_8476) ) ;
    buf_clk cell_6634 ( .C (clk), .D (signal_8483), .Q (signal_8484) ) ;
    buf_clk cell_6642 ( .C (clk), .D (signal_8491), .Q (signal_8492) ) ;
    buf_clk cell_6650 ( .C (clk), .D (signal_8499), .Q (signal_8500) ) ;
    buf_clk cell_6658 ( .C (clk), .D (signal_8507), .Q (signal_8508) ) ;
    buf_clk cell_6666 ( .C (clk), .D (signal_8515), .Q (signal_8516) ) ;
    buf_clk cell_6674 ( .C (clk), .D (signal_8523), .Q (signal_8524) ) ;
    buf_clk cell_6682 ( .C (clk), .D (signal_8531), .Q (signal_8532) ) ;
    buf_clk cell_6690 ( .C (clk), .D (signal_8539), .Q (signal_8540) ) ;
    buf_clk cell_6698 ( .C (clk), .D (signal_8547), .Q (signal_8548) ) ;
    buf_clk cell_6706 ( .C (clk), .D (signal_8555), .Q (signal_8556) ) ;
    buf_clk cell_6714 ( .C (clk), .D (signal_8563), .Q (signal_8564) ) ;
    buf_clk cell_6722 ( .C (clk), .D (signal_8571), .Q (signal_8572) ) ;
    buf_clk cell_6730 ( .C (clk), .D (signal_8579), .Q (signal_8580) ) ;
    buf_clk cell_6738 ( .C (clk), .D (signal_8587), .Q (signal_8588) ) ;
    buf_clk cell_6746 ( .C (clk), .D (signal_8595), .Q (signal_8596) ) ;
    buf_clk cell_6754 ( .C (clk), .D (signal_8603), .Q (signal_8604) ) ;
    buf_clk cell_6762 ( .C (clk), .D (signal_8611), .Q (signal_8612) ) ;
    buf_clk cell_6770 ( .C (clk), .D (signal_8619), .Q (signal_8620) ) ;
    buf_clk cell_6778 ( .C (clk), .D (signal_8627), .Q (signal_8628) ) ;
    buf_clk cell_6786 ( .C (clk), .D (signal_8635), .Q (signal_8636) ) ;
    buf_clk cell_6794 ( .C (clk), .D (signal_8643), .Q (signal_8644) ) ;
    buf_clk cell_6802 ( .C (clk), .D (signal_8651), .Q (signal_8652) ) ;
    buf_clk cell_6810 ( .C (clk), .D (signal_8659), .Q (signal_8660) ) ;
    buf_clk cell_6818 ( .C (clk), .D (signal_8667), .Q (signal_8668) ) ;
    buf_clk cell_6826 ( .C (clk), .D (signal_8675), .Q (signal_8676) ) ;
    buf_clk cell_6834 ( .C (clk), .D (signal_8683), .Q (signal_8684) ) ;
    buf_clk cell_6842 ( .C (clk), .D (signal_8691), .Q (signal_8692) ) ;
    buf_clk cell_6850 ( .C (clk), .D (signal_8699), .Q (signal_8700) ) ;
    buf_clk cell_6858 ( .C (clk), .D (signal_8707), .Q (signal_8708) ) ;
    buf_clk cell_6866 ( .C (clk), .D (signal_8715), .Q (signal_8716) ) ;
    buf_clk cell_6874 ( .C (clk), .D (signal_8723), .Q (signal_8724) ) ;
    buf_clk cell_6882 ( .C (clk), .D (signal_8731), .Q (signal_8732) ) ;
    buf_clk cell_6890 ( .C (clk), .D (signal_8739), .Q (signal_8740) ) ;
    buf_clk cell_6898 ( .C (clk), .D (signal_8747), .Q (signal_8748) ) ;
    buf_clk cell_6906 ( .C (clk), .D (signal_8755), .Q (signal_8756) ) ;
    buf_clk cell_6914 ( .C (clk), .D (signal_8763), .Q (signal_8764) ) ;
    buf_clk cell_6922 ( .C (clk), .D (signal_8771), .Q (signal_8772) ) ;
    buf_clk cell_6930 ( .C (clk), .D (signal_8779), .Q (signal_8780) ) ;
    buf_clk cell_6938 ( .C (clk), .D (signal_8787), .Q (signal_8788) ) ;
    buf_clk cell_6946 ( .C (clk), .D (signal_8795), .Q (signal_8796) ) ;
    buf_clk cell_6954 ( .C (clk), .D (signal_8803), .Q (signal_8804) ) ;
    buf_clk cell_6962 ( .C (clk), .D (signal_8811), .Q (signal_8812) ) ;
    buf_clk cell_6970 ( .C (clk), .D (signal_8819), .Q (signal_8820) ) ;
    buf_clk cell_6978 ( .C (clk), .D (signal_8827), .Q (signal_8828) ) ;
    buf_clk cell_6986 ( .C (clk), .D (signal_8835), .Q (signal_8836) ) ;
    buf_clk cell_6994 ( .C (clk), .D (signal_8843), .Q (signal_8844) ) ;
    buf_clk cell_7002 ( .C (clk), .D (signal_8851), .Q (signal_8852) ) ;
    buf_clk cell_7010 ( .C (clk), .D (signal_8859), .Q (signal_8860) ) ;
    buf_clk cell_7018 ( .C (clk), .D (signal_8867), .Q (signal_8868) ) ;
    buf_clk cell_7026 ( .C (clk), .D (signal_8875), .Q (signal_8876) ) ;
    buf_clk cell_7034 ( .C (clk), .D (signal_8883), .Q (signal_8884) ) ;
    buf_clk cell_7042 ( .C (clk), .D (signal_8891), .Q (signal_8892) ) ;
    buf_clk cell_7050 ( .C (clk), .D (signal_8899), .Q (signal_8900) ) ;
    buf_clk cell_7058 ( .C (clk), .D (signal_8907), .Q (signal_8908) ) ;
    buf_clk cell_7066 ( .C (clk), .D (signal_8915), .Q (signal_8916) ) ;
    buf_clk cell_7074 ( .C (clk), .D (signal_8923), .Q (signal_8924) ) ;
    buf_clk cell_7082 ( .C (clk), .D (signal_8931), .Q (signal_8932) ) ;
    buf_clk cell_7090 ( .C (clk), .D (signal_8939), .Q (signal_8940) ) ;
    buf_clk cell_7098 ( .C (clk), .D (signal_8947), .Q (signal_8948) ) ;

    /* cells in depth 6 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1772 ( .a ({signal_3723, signal_3721}), .b ({signal_3514, signal_2038}), .clk (clk), .r (Fresh[12]), .c ({signal_3516, signal_2040}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1773 ( .a ({signal_3727, signal_3725}), .b ({signal_3513, signal_2037}), .clk (clk), .r (Fresh[13]), .c ({signal_3517, signal_2041}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1774 ( .a ({signal_3723, signal_3721}), .b ({signal_3511, signal_2035}), .clk (clk), .r (Fresh[14]), .c ({signal_3518, signal_2042}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1775 ( .a ({signal_3508, signal_2032}), .b ({signal_3727, signal_3725}), .clk (clk), .r (Fresh[15]), .c ({signal_3519, signal_2043}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1777 ( .a ({signal_3731, signal_3729}), .b ({signal_3516, signal_2040}), .c ({signal_3521, signal_2045}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1778 ( .a ({signal_3735, signal_3733}), .b ({signal_3518, signal_2042}), .c ({signal_3522, signal_2046}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1779 ( .a ({signal_3739, signal_3737}), .b ({signal_3517, signal_2041}), .c ({signal_3523, signal_2047}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1780 ( .a ({signal_3519, signal_2043}), .b ({signal_3743, signal_3741}), .c ({signal_3524, signal_2048}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1789 ( .a ({signal_3522, signal_2046}), .b ({signal_3524, signal_2048}), .c ({signal_3533, signal_2057}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1790 ( .a ({signal_3521, signal_2045}), .b ({signal_3523, signal_2047}), .c ({signal_3534, signal_2058}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1791 ( .a ({signal_3521, signal_2045}), .b ({signal_3522, signal_2046}), .c ({signal_3535, signal_2059}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1792 ( .a ({signal_3523, signal_2047}), .b ({signal_3524, signal_2048}), .c ({signal_3536, signal_2060}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1801 ( .a ({signal_3533, signal_2057}), .b ({signal_3534, signal_2058}), .c ({signal_3545, signal_2069}) ) ;
    buf_clk cell_1879 ( .C (clk), .D (signal_3728), .Q (signal_3729) ) ;
    buf_clk cell_1881 ( .C (clk), .D (signal_3730), .Q (signal_3731) ) ;
    buf_clk cell_1883 ( .C (clk), .D (signal_3732), .Q (signal_3733) ) ;
    buf_clk cell_1885 ( .C (clk), .D (signal_3734), .Q (signal_3735) ) ;
    buf_clk cell_1887 ( .C (clk), .D (signal_3736), .Q (signal_3737) ) ;
    buf_clk cell_1889 ( .C (clk), .D (signal_3738), .Q (signal_3739) ) ;
    buf_clk cell_1891 ( .C (clk), .D (signal_3740), .Q (signal_3741) ) ;
    buf_clk cell_1893 ( .C (clk), .D (signal_3742), .Q (signal_3743) ) ;
    buf_clk cell_1899 ( .C (clk), .D (signal_3748), .Q (signal_3749) ) ;
    buf_clk cell_1907 ( .C (clk), .D (signal_3756), .Q (signal_3757) ) ;
    buf_clk cell_1915 ( .C (clk), .D (signal_3764), .Q (signal_3765) ) ;
    buf_clk cell_1923 ( .C (clk), .D (signal_3772), .Q (signal_3773) ) ;
    buf_clk cell_1931 ( .C (clk), .D (signal_3780), .Q (signal_3781) ) ;
    buf_clk cell_1939 ( .C (clk), .D (signal_3788), .Q (signal_3789) ) ;
    buf_clk cell_1947 ( .C (clk), .D (signal_3796), .Q (signal_3797) ) ;
    buf_clk cell_1955 ( .C (clk), .D (signal_3804), .Q (signal_3805) ) ;
    buf_clk cell_1963 ( .C (clk), .D (signal_3812), .Q (signal_3813) ) ;
    buf_clk cell_1971 ( .C (clk), .D (signal_3820), .Q (signal_3821) ) ;
    buf_clk cell_1979 ( .C (clk), .D (signal_3828), .Q (signal_3829) ) ;
    buf_clk cell_1987 ( .C (clk), .D (signal_3836), .Q (signal_3837) ) ;
    buf_clk cell_1995 ( .C (clk), .D (signal_3844), .Q (signal_3845) ) ;
    buf_clk cell_2003 ( .C (clk), .D (signal_3852), .Q (signal_3853) ) ;
    buf_clk cell_2011 ( .C (clk), .D (signal_3860), .Q (signal_3861) ) ;
    buf_clk cell_2019 ( .C (clk), .D (signal_3868), .Q (signal_3869) ) ;
    buf_clk cell_2027 ( .C (clk), .D (signal_3876), .Q (signal_3877) ) ;
    buf_clk cell_2035 ( .C (clk), .D (signal_3884), .Q (signal_3885) ) ;
    buf_clk cell_2043 ( .C (clk), .D (signal_3892), .Q (signal_3893) ) ;
    buf_clk cell_2051 ( .C (clk), .D (signal_3900), .Q (signal_3901) ) ;
    buf_clk cell_2059 ( .C (clk), .D (signal_3908), .Q (signal_3909) ) ;
    buf_clk cell_2067 ( .C (clk), .D (signal_3916), .Q (signal_3917) ) ;
    buf_clk cell_2075 ( .C (clk), .D (signal_3924), .Q (signal_3925) ) ;
    buf_clk cell_2083 ( .C (clk), .D (signal_3932), .Q (signal_3933) ) ;
    buf_clk cell_2091 ( .C (clk), .D (signal_3940), .Q (signal_3941) ) ;
    buf_clk cell_2099 ( .C (clk), .D (signal_3948), .Q (signal_3949) ) ;
    buf_clk cell_2107 ( .C (clk), .D (signal_3956), .Q (signal_3957) ) ;
    buf_clk cell_2115 ( .C (clk), .D (signal_3964), .Q (signal_3965) ) ;
    buf_clk cell_2123 ( .C (clk), .D (signal_3972), .Q (signal_3973) ) ;
    buf_clk cell_2131 ( .C (clk), .D (signal_3980), .Q (signal_3981) ) ;
    buf_clk cell_2139 ( .C (clk), .D (signal_3988), .Q (signal_3989) ) ;
    buf_clk cell_2147 ( .C (clk), .D (signal_3996), .Q (signal_3997) ) ;
    buf_clk cell_2155 ( .C (clk), .D (signal_4004), .Q (signal_4005) ) ;
    buf_clk cell_2163 ( .C (clk), .D (signal_4012), .Q (signal_4013) ) ;
    buf_clk cell_2171 ( .C (clk), .D (signal_4020), .Q (signal_4021) ) ;
    buf_clk cell_2179 ( .C (clk), .D (signal_4028), .Q (signal_4029) ) ;
    buf_clk cell_2187 ( .C (clk), .D (signal_4036), .Q (signal_4037) ) ;
    buf_clk cell_2195 ( .C (clk), .D (signal_4044), .Q (signal_4045) ) ;
    buf_clk cell_2203 ( .C (clk), .D (signal_4052), .Q (signal_4053) ) ;
    buf_clk cell_2211 ( .C (clk), .D (signal_4060), .Q (signal_4061) ) ;
    buf_clk cell_2219 ( .C (clk), .D (signal_4068), .Q (signal_4069) ) ;
    buf_clk cell_2227 ( .C (clk), .D (signal_4076), .Q (signal_4077) ) ;
    buf_clk cell_2235 ( .C (clk), .D (signal_4084), .Q (signal_4085) ) ;
    buf_clk cell_2243 ( .C (clk), .D (signal_4092), .Q (signal_4093) ) ;
    buf_clk cell_2251 ( .C (clk), .D (signal_4100), .Q (signal_4101) ) ;
    buf_clk cell_2259 ( .C (clk), .D (signal_4108), .Q (signal_4109) ) ;
    buf_clk cell_2267 ( .C (clk), .D (signal_4116), .Q (signal_4117) ) ;
    buf_clk cell_2275 ( .C (clk), .D (signal_4124), .Q (signal_4125) ) ;
    buf_clk cell_2283 ( .C (clk), .D (signal_4132), .Q (signal_4133) ) ;
    buf_clk cell_2291 ( .C (clk), .D (signal_4140), .Q (signal_4141) ) ;
    buf_clk cell_2299 ( .C (clk), .D (signal_4148), .Q (signal_4149) ) ;
    buf_clk cell_2307 ( .C (clk), .D (signal_4156), .Q (signal_4157) ) ;
    buf_clk cell_2315 ( .C (clk), .D (signal_4164), .Q (signal_4165) ) ;
    buf_clk cell_2323 ( .C (clk), .D (signal_4172), .Q (signal_4173) ) ;
    buf_clk cell_2331 ( .C (clk), .D (signal_4180), .Q (signal_4181) ) ;
    buf_clk cell_2339 ( .C (clk), .D (signal_4188), .Q (signal_4189) ) ;
    buf_clk cell_2347 ( .C (clk), .D (signal_4196), .Q (signal_4197) ) ;
    buf_clk cell_2355 ( .C (clk), .D (signal_4204), .Q (signal_4205) ) ;
    buf_clk cell_2363 ( .C (clk), .D (signal_4212), .Q (signal_4213) ) ;
    buf_clk cell_2371 ( .C (clk), .D (signal_4220), .Q (signal_4221) ) ;
    buf_clk cell_2379 ( .C (clk), .D (signal_4228), .Q (signal_4229) ) ;
    buf_clk cell_2387 ( .C (clk), .D (signal_4236), .Q (signal_4237) ) ;
    buf_clk cell_2395 ( .C (clk), .D (signal_4244), .Q (signal_4245) ) ;
    buf_clk cell_2403 ( .C (clk), .D (signal_4252), .Q (signal_4253) ) ;
    buf_clk cell_2411 ( .C (clk), .D (signal_4260), .Q (signal_4261) ) ;
    buf_clk cell_2419 ( .C (clk), .D (signal_4268), .Q (signal_4269) ) ;
    buf_clk cell_2427 ( .C (clk), .D (signal_4276), .Q (signal_4277) ) ;
    buf_clk cell_2435 ( .C (clk), .D (signal_4284), .Q (signal_4285) ) ;
    buf_clk cell_2443 ( .C (clk), .D (signal_4292), .Q (signal_4293) ) ;
    buf_clk cell_2451 ( .C (clk), .D (signal_4300), .Q (signal_4301) ) ;
    buf_clk cell_2459 ( .C (clk), .D (signal_4308), .Q (signal_4309) ) ;
    buf_clk cell_2467 ( .C (clk), .D (signal_4316), .Q (signal_4317) ) ;
    buf_clk cell_2475 ( .C (clk), .D (signal_4324), .Q (signal_4325) ) ;
    buf_clk cell_2483 ( .C (clk), .D (signal_4332), .Q (signal_4333) ) ;
    buf_clk cell_2491 ( .C (clk), .D (signal_4340), .Q (signal_4341) ) ;
    buf_clk cell_2499 ( .C (clk), .D (signal_4348), .Q (signal_4349) ) ;
    buf_clk cell_2507 ( .C (clk), .D (signal_4356), .Q (signal_4357) ) ;
    buf_clk cell_2515 ( .C (clk), .D (signal_4364), .Q (signal_4365) ) ;
    buf_clk cell_2523 ( .C (clk), .D (signal_4372), .Q (signal_4373) ) ;
    buf_clk cell_2531 ( .C (clk), .D (signal_4380), .Q (signal_4381) ) ;
    buf_clk cell_2539 ( .C (clk), .D (signal_4388), .Q (signal_4389) ) ;
    buf_clk cell_2547 ( .C (clk), .D (signal_4396), .Q (signal_4397) ) ;
    buf_clk cell_2555 ( .C (clk), .D (signal_4404), .Q (signal_4405) ) ;
    buf_clk cell_2563 ( .C (clk), .D (signal_4412), .Q (signal_4413) ) ;
    buf_clk cell_2571 ( .C (clk), .D (signal_4420), .Q (signal_4421) ) ;
    buf_clk cell_2579 ( .C (clk), .D (signal_4428), .Q (signal_4429) ) ;
    buf_clk cell_2587 ( .C (clk), .D (signal_4436), .Q (signal_4437) ) ;
    buf_clk cell_2595 ( .C (clk), .D (signal_4444), .Q (signal_4445) ) ;
    buf_clk cell_2603 ( .C (clk), .D (signal_4452), .Q (signal_4453) ) ;
    buf_clk cell_2611 ( .C (clk), .D (signal_4460), .Q (signal_4461) ) ;
    buf_clk cell_2619 ( .C (clk), .D (signal_4468), .Q (signal_4469) ) ;
    buf_clk cell_2627 ( .C (clk), .D (signal_4476), .Q (signal_4477) ) ;
    buf_clk cell_2635 ( .C (clk), .D (signal_4484), .Q (signal_4485) ) ;
    buf_clk cell_2643 ( .C (clk), .D (signal_4492), .Q (signal_4493) ) ;
    buf_clk cell_2651 ( .C (clk), .D (signal_4500), .Q (signal_4501) ) ;
    buf_clk cell_2659 ( .C (clk), .D (signal_4508), .Q (signal_4509) ) ;
    buf_clk cell_2667 ( .C (clk), .D (signal_4516), .Q (signal_4517) ) ;
    buf_clk cell_2675 ( .C (clk), .D (signal_4524), .Q (signal_4525) ) ;
    buf_clk cell_2683 ( .C (clk), .D (signal_4532), .Q (signal_4533) ) ;
    buf_clk cell_2691 ( .C (clk), .D (signal_4540), .Q (signal_4541) ) ;
    buf_clk cell_2699 ( .C (clk), .D (signal_4548), .Q (signal_4549) ) ;
    buf_clk cell_2707 ( .C (clk), .D (signal_4556), .Q (signal_4557) ) ;
    buf_clk cell_2715 ( .C (clk), .D (signal_4564), .Q (signal_4565) ) ;
    buf_clk cell_2723 ( .C (clk), .D (signal_4572), .Q (signal_4573) ) ;
    buf_clk cell_2731 ( .C (clk), .D (signal_4580), .Q (signal_4581) ) ;
    buf_clk cell_2739 ( .C (clk), .D (signal_4588), .Q (signal_4589) ) ;
    buf_clk cell_2747 ( .C (clk), .D (signal_4596), .Q (signal_4597) ) ;
    buf_clk cell_2755 ( .C (clk), .D (signal_4604), .Q (signal_4605) ) ;
    buf_clk cell_2763 ( .C (clk), .D (signal_4612), .Q (signal_4613) ) ;
    buf_clk cell_2771 ( .C (clk), .D (signal_4620), .Q (signal_4621) ) ;
    buf_clk cell_2779 ( .C (clk), .D (signal_4628), .Q (signal_4629) ) ;
    buf_clk cell_2787 ( .C (clk), .D (signal_4636), .Q (signal_4637) ) ;
    buf_clk cell_2795 ( .C (clk), .D (signal_4644), .Q (signal_4645) ) ;
    buf_clk cell_2803 ( .C (clk), .D (signal_4652), .Q (signal_4653) ) ;
    buf_clk cell_2811 ( .C (clk), .D (signal_4660), .Q (signal_4661) ) ;
    buf_clk cell_2819 ( .C (clk), .D (signal_4668), .Q (signal_4669) ) ;
    buf_clk cell_2827 ( .C (clk), .D (signal_4676), .Q (signal_4677) ) ;
    buf_clk cell_2835 ( .C (clk), .D (signal_4684), .Q (signal_4685) ) ;
    buf_clk cell_2843 ( .C (clk), .D (signal_4692), .Q (signal_4693) ) ;
    buf_clk cell_2851 ( .C (clk), .D (signal_4700), .Q (signal_4701) ) ;
    buf_clk cell_2859 ( .C (clk), .D (signal_4708), .Q (signal_4709) ) ;
    buf_clk cell_2867 ( .C (clk), .D (signal_4716), .Q (signal_4717) ) ;
    buf_clk cell_2875 ( .C (clk), .D (signal_4724), .Q (signal_4725) ) ;
    buf_clk cell_2883 ( .C (clk), .D (signal_4732), .Q (signal_4733) ) ;
    buf_clk cell_2891 ( .C (clk), .D (signal_4740), .Q (signal_4741) ) ;
    buf_clk cell_2899 ( .C (clk), .D (signal_4748), .Q (signal_4749) ) ;
    buf_clk cell_2907 ( .C (clk), .D (signal_4756), .Q (signal_4757) ) ;
    buf_clk cell_2913 ( .C (clk), .D (signal_4762), .Q (signal_4763) ) ;
    buf_clk cell_2919 ( .C (clk), .D (signal_4768), .Q (signal_4769) ) ;
    buf_clk cell_2925 ( .C (clk), .D (signal_4774), .Q (signal_4775) ) ;
    buf_clk cell_2931 ( .C (clk), .D (signal_4780), .Q (signal_4781) ) ;
    buf_clk cell_2937 ( .C (clk), .D (signal_4786), .Q (signal_4787) ) ;
    buf_clk cell_2943 ( .C (clk), .D (signal_4792), .Q (signal_4793) ) ;
    buf_clk cell_2949 ( .C (clk), .D (signal_4798), .Q (signal_4799) ) ;
    buf_clk cell_2955 ( .C (clk), .D (signal_4804), .Q (signal_4805) ) ;
    buf_clk cell_2961 ( .C (clk), .D (signal_4810), .Q (signal_4811) ) ;
    buf_clk cell_2967 ( .C (clk), .D (signal_4816), .Q (signal_4817) ) ;
    buf_clk cell_2973 ( .C (clk), .D (signal_4822), .Q (signal_4823) ) ;
    buf_clk cell_2979 ( .C (clk), .D (signal_4828), .Q (signal_4829) ) ;
    buf_clk cell_2985 ( .C (clk), .D (signal_4834), .Q (signal_4835) ) ;
    buf_clk cell_2991 ( .C (clk), .D (signal_4840), .Q (signal_4841) ) ;
    buf_clk cell_2997 ( .C (clk), .D (signal_4846), .Q (signal_4847) ) ;
    buf_clk cell_3003 ( .C (clk), .D (signal_4852), .Q (signal_4853) ) ;
    buf_clk cell_3009 ( .C (clk), .D (signal_4858), .Q (signal_4859) ) ;
    buf_clk cell_3015 ( .C (clk), .D (signal_4864), .Q (signal_4865) ) ;
    buf_clk cell_3021 ( .C (clk), .D (signal_4870), .Q (signal_4871) ) ;
    buf_clk cell_3027 ( .C (clk), .D (signal_4876), .Q (signal_4877) ) ;
    buf_clk cell_3033 ( .C (clk), .D (signal_4882), .Q (signal_4883) ) ;
    buf_clk cell_3039 ( .C (clk), .D (signal_4888), .Q (signal_4889) ) ;
    buf_clk cell_3045 ( .C (clk), .D (signal_4894), .Q (signal_4895) ) ;
    buf_clk cell_3051 ( .C (clk), .D (signal_4900), .Q (signal_4901) ) ;
    buf_clk cell_3057 ( .C (clk), .D (signal_4906), .Q (signal_4907) ) ;
    buf_clk cell_3063 ( .C (clk), .D (signal_4912), .Q (signal_4913) ) ;
    buf_clk cell_3069 ( .C (clk), .D (signal_4918), .Q (signal_4919) ) ;
    buf_clk cell_3075 ( .C (clk), .D (signal_4924), .Q (signal_4925) ) ;
    buf_clk cell_3081 ( .C (clk), .D (signal_4930), .Q (signal_4931) ) ;
    buf_clk cell_3087 ( .C (clk), .D (signal_4936), .Q (signal_4937) ) ;
    buf_clk cell_3093 ( .C (clk), .D (signal_4942), .Q (signal_4943) ) ;
    buf_clk cell_3099 ( .C (clk), .D (signal_4948), .Q (signal_4949) ) ;
    buf_clk cell_3105 ( .C (clk), .D (signal_4954), .Q (signal_4955) ) ;
    buf_clk cell_3111 ( .C (clk), .D (signal_4960), .Q (signal_4961) ) ;
    buf_clk cell_3117 ( .C (clk), .D (signal_4966), .Q (signal_4967) ) ;
    buf_clk cell_3123 ( .C (clk), .D (signal_4972), .Q (signal_4973) ) ;
    buf_clk cell_3131 ( .C (clk), .D (signal_4980), .Q (signal_4981) ) ;
    buf_clk cell_3139 ( .C (clk), .D (signal_4988), .Q (signal_4989) ) ;
    buf_clk cell_3147 ( .C (clk), .D (signal_4996), .Q (signal_4997) ) ;
    buf_clk cell_3155 ( .C (clk), .D (signal_5004), .Q (signal_5005) ) ;
    buf_clk cell_3163 ( .C (clk), .D (signal_5012), .Q (signal_5013) ) ;
    buf_clk cell_3171 ( .C (clk), .D (signal_5020), .Q (signal_5021) ) ;
    buf_clk cell_3179 ( .C (clk), .D (signal_5028), .Q (signal_5029) ) ;
    buf_clk cell_3187 ( .C (clk), .D (signal_5036), .Q (signal_5037) ) ;
    buf_clk cell_3195 ( .C (clk), .D (signal_5044), .Q (signal_5045) ) ;
    buf_clk cell_3203 ( .C (clk), .D (signal_5052), .Q (signal_5053) ) ;
    buf_clk cell_3211 ( .C (clk), .D (signal_5060), .Q (signal_5061) ) ;
    buf_clk cell_3219 ( .C (clk), .D (signal_5068), .Q (signal_5069) ) ;
    buf_clk cell_3227 ( .C (clk), .D (signal_5076), .Q (signal_5077) ) ;
    buf_clk cell_3235 ( .C (clk), .D (signal_5084), .Q (signal_5085) ) ;
    buf_clk cell_3243 ( .C (clk), .D (signal_5092), .Q (signal_5093) ) ;
    buf_clk cell_3251 ( .C (clk), .D (signal_5100), .Q (signal_5101) ) ;
    buf_clk cell_3259 ( .C (clk), .D (signal_5108), .Q (signal_5109) ) ;
    buf_clk cell_3267 ( .C (clk), .D (signal_5116), .Q (signal_5117) ) ;
    buf_clk cell_3275 ( .C (clk), .D (signal_5124), .Q (signal_5125) ) ;
    buf_clk cell_3283 ( .C (clk), .D (signal_5132), .Q (signal_5133) ) ;
    buf_clk cell_3291 ( .C (clk), .D (signal_5140), .Q (signal_5141) ) ;
    buf_clk cell_3299 ( .C (clk), .D (signal_5148), .Q (signal_5149) ) ;
    buf_clk cell_3307 ( .C (clk), .D (signal_5156), .Q (signal_5157) ) ;
    buf_clk cell_3315 ( .C (clk), .D (signal_5164), .Q (signal_5165) ) ;
    buf_clk cell_3323 ( .C (clk), .D (signal_5172), .Q (signal_5173) ) ;
    buf_clk cell_3331 ( .C (clk), .D (signal_5180), .Q (signal_5181) ) ;
    buf_clk cell_3339 ( .C (clk), .D (signal_5188), .Q (signal_5189) ) ;
    buf_clk cell_3347 ( .C (clk), .D (signal_5196), .Q (signal_5197) ) ;
    buf_clk cell_3355 ( .C (clk), .D (signal_5204), .Q (signal_5205) ) ;
    buf_clk cell_3363 ( .C (clk), .D (signal_5212), .Q (signal_5213) ) ;
    buf_clk cell_3371 ( .C (clk), .D (signal_5220), .Q (signal_5221) ) ;
    buf_clk cell_3379 ( .C (clk), .D (signal_5228), .Q (signal_5229) ) ;
    buf_clk cell_3387 ( .C (clk), .D (signal_5236), .Q (signal_5237) ) ;
    buf_clk cell_3395 ( .C (clk), .D (signal_5244), .Q (signal_5245) ) ;
    buf_clk cell_3403 ( .C (clk), .D (signal_5252), .Q (signal_5253) ) ;
    buf_clk cell_3411 ( .C (clk), .D (signal_5260), .Q (signal_5261) ) ;
    buf_clk cell_3419 ( .C (clk), .D (signal_5268), .Q (signal_5269) ) ;
    buf_clk cell_3427 ( .C (clk), .D (signal_5276), .Q (signal_5277) ) ;
    buf_clk cell_3435 ( .C (clk), .D (signal_5284), .Q (signal_5285) ) ;
    buf_clk cell_3443 ( .C (clk), .D (signal_5292), .Q (signal_5293) ) ;
    buf_clk cell_3451 ( .C (clk), .D (signal_5300), .Q (signal_5301) ) ;
    buf_clk cell_3459 ( .C (clk), .D (signal_5308), .Q (signal_5309) ) ;
    buf_clk cell_3467 ( .C (clk), .D (signal_5316), .Q (signal_5317) ) ;
    buf_clk cell_3475 ( .C (clk), .D (signal_5324), .Q (signal_5325) ) ;
    buf_clk cell_3483 ( .C (clk), .D (signal_5332), .Q (signal_5333) ) ;
    buf_clk cell_3491 ( .C (clk), .D (signal_5340), .Q (signal_5341) ) ;
    buf_clk cell_3499 ( .C (clk), .D (signal_5348), .Q (signal_5349) ) ;
    buf_clk cell_3507 ( .C (clk), .D (signal_5356), .Q (signal_5357) ) ;
    buf_clk cell_3515 ( .C (clk), .D (signal_5364), .Q (signal_5365) ) ;
    buf_clk cell_3523 ( .C (clk), .D (signal_5372), .Q (signal_5373) ) ;
    buf_clk cell_3531 ( .C (clk), .D (signal_5380), .Q (signal_5381) ) ;
    buf_clk cell_3539 ( .C (clk), .D (signal_5388), .Q (signal_5389) ) ;
    buf_clk cell_3547 ( .C (clk), .D (signal_5396), .Q (signal_5397) ) ;
    buf_clk cell_3555 ( .C (clk), .D (signal_5404), .Q (signal_5405) ) ;
    buf_clk cell_3563 ( .C (clk), .D (signal_5412), .Q (signal_5413) ) ;
    buf_clk cell_3571 ( .C (clk), .D (signal_5420), .Q (signal_5421) ) ;
    buf_clk cell_3579 ( .C (clk), .D (signal_5428), .Q (signal_5429) ) ;
    buf_clk cell_3587 ( .C (clk), .D (signal_5436), .Q (signal_5437) ) ;
    buf_clk cell_3595 ( .C (clk), .D (signal_5444), .Q (signal_5445) ) ;
    buf_clk cell_3603 ( .C (clk), .D (signal_5452), .Q (signal_5453) ) ;
    buf_clk cell_3611 ( .C (clk), .D (signal_5460), .Q (signal_5461) ) ;
    buf_clk cell_3619 ( .C (clk), .D (signal_5468), .Q (signal_5469) ) ;
    buf_clk cell_3627 ( .C (clk), .D (signal_5476), .Q (signal_5477) ) ;
    buf_clk cell_3635 ( .C (clk), .D (signal_5484), .Q (signal_5485) ) ;
    buf_clk cell_3643 ( .C (clk), .D (signal_5492), .Q (signal_5493) ) ;
    buf_clk cell_3651 ( .C (clk), .D (signal_5500), .Q (signal_5501) ) ;
    buf_clk cell_3659 ( .C (clk), .D (signal_5508), .Q (signal_5509) ) ;
    buf_clk cell_3667 ( .C (clk), .D (signal_5516), .Q (signal_5517) ) ;
    buf_clk cell_3675 ( .C (clk), .D (signal_5524), .Q (signal_5525) ) ;
    buf_clk cell_3683 ( .C (clk), .D (signal_5532), .Q (signal_5533) ) ;
    buf_clk cell_3691 ( .C (clk), .D (signal_5540), .Q (signal_5541) ) ;
    buf_clk cell_3699 ( .C (clk), .D (signal_5548), .Q (signal_5549) ) ;
    buf_clk cell_3707 ( .C (clk), .D (signal_5556), .Q (signal_5557) ) ;
    buf_clk cell_3715 ( .C (clk), .D (signal_5564), .Q (signal_5565) ) ;
    buf_clk cell_3723 ( .C (clk), .D (signal_5572), .Q (signal_5573) ) ;
    buf_clk cell_3731 ( .C (clk), .D (signal_5580), .Q (signal_5581) ) ;
    buf_clk cell_3739 ( .C (clk), .D (signal_5588), .Q (signal_5589) ) ;
    buf_clk cell_3747 ( .C (clk), .D (signal_5596), .Q (signal_5597) ) ;
    buf_clk cell_3755 ( .C (clk), .D (signal_5604), .Q (signal_5605) ) ;
    buf_clk cell_3763 ( .C (clk), .D (signal_5612), .Q (signal_5613) ) ;
    buf_clk cell_3771 ( .C (clk), .D (signal_5620), .Q (signal_5621) ) ;
    buf_clk cell_3779 ( .C (clk), .D (signal_5628), .Q (signal_5629) ) ;
    buf_clk cell_3787 ( .C (clk), .D (signal_5636), .Q (signal_5637) ) ;
    buf_clk cell_3795 ( .C (clk), .D (signal_5644), .Q (signal_5645) ) ;
    buf_clk cell_3803 ( .C (clk), .D (signal_5652), .Q (signal_5653) ) ;
    buf_clk cell_3811 ( .C (clk), .D (signal_5660), .Q (signal_5661) ) ;
    buf_clk cell_3819 ( .C (clk), .D (signal_5668), .Q (signal_5669) ) ;
    buf_clk cell_3827 ( .C (clk), .D (signal_5676), .Q (signal_5677) ) ;
    buf_clk cell_3835 ( .C (clk), .D (signal_5684), .Q (signal_5685) ) ;
    buf_clk cell_3843 ( .C (clk), .D (signal_5692), .Q (signal_5693) ) ;
    buf_clk cell_3851 ( .C (clk), .D (signal_5700), .Q (signal_5701) ) ;
    buf_clk cell_3859 ( .C (clk), .D (signal_5708), .Q (signal_5709) ) ;
    buf_clk cell_3867 ( .C (clk), .D (signal_5716), .Q (signal_5717) ) ;
    buf_clk cell_3875 ( .C (clk), .D (signal_5724), .Q (signal_5725) ) ;
    buf_clk cell_3883 ( .C (clk), .D (signal_5732), .Q (signal_5733) ) ;
    buf_clk cell_3891 ( .C (clk), .D (signal_5740), .Q (signal_5741) ) ;
    buf_clk cell_3899 ( .C (clk), .D (signal_5748), .Q (signal_5749) ) ;
    buf_clk cell_3907 ( .C (clk), .D (signal_5756), .Q (signal_5757) ) ;
    buf_clk cell_3915 ( .C (clk), .D (signal_5764), .Q (signal_5765) ) ;
    buf_clk cell_3923 ( .C (clk), .D (signal_5772), .Q (signal_5773) ) ;
    buf_clk cell_3931 ( .C (clk), .D (signal_5780), .Q (signal_5781) ) ;
    buf_clk cell_3939 ( .C (clk), .D (signal_5788), .Q (signal_5789) ) ;
    buf_clk cell_3947 ( .C (clk), .D (signal_5796), .Q (signal_5797) ) ;
    buf_clk cell_3955 ( .C (clk), .D (signal_5804), .Q (signal_5805) ) ;
    buf_clk cell_3963 ( .C (clk), .D (signal_5812), .Q (signal_5813) ) ;
    buf_clk cell_3971 ( .C (clk), .D (signal_5820), .Q (signal_5821) ) ;
    buf_clk cell_3979 ( .C (clk), .D (signal_5828), .Q (signal_5829) ) ;
    buf_clk cell_3987 ( .C (clk), .D (signal_5836), .Q (signal_5837) ) ;
    buf_clk cell_3995 ( .C (clk), .D (signal_5844), .Q (signal_5845) ) ;
    buf_clk cell_4003 ( .C (clk), .D (signal_5852), .Q (signal_5853) ) ;
    buf_clk cell_4011 ( .C (clk), .D (signal_5860), .Q (signal_5861) ) ;
    buf_clk cell_4019 ( .C (clk), .D (signal_5868), .Q (signal_5869) ) ;
    buf_clk cell_4027 ( .C (clk), .D (signal_5876), .Q (signal_5877) ) ;
    buf_clk cell_4035 ( .C (clk), .D (signal_5884), .Q (signal_5885) ) ;
    buf_clk cell_4043 ( .C (clk), .D (signal_5892), .Q (signal_5893) ) ;
    buf_clk cell_4051 ( .C (clk), .D (signal_5900), .Q (signal_5901) ) ;
    buf_clk cell_4059 ( .C (clk), .D (signal_5908), .Q (signal_5909) ) ;
    buf_clk cell_4067 ( .C (clk), .D (signal_5916), .Q (signal_5917) ) ;
    buf_clk cell_4075 ( .C (clk), .D (signal_5924), .Q (signal_5925) ) ;
    buf_clk cell_4083 ( .C (clk), .D (signal_5932), .Q (signal_5933) ) ;
    buf_clk cell_4091 ( .C (clk), .D (signal_5940), .Q (signal_5941) ) ;
    buf_clk cell_4099 ( .C (clk), .D (signal_5948), .Q (signal_5949) ) ;
    buf_clk cell_4107 ( .C (clk), .D (signal_5956), .Q (signal_5957) ) ;
    buf_clk cell_4115 ( .C (clk), .D (signal_5964), .Q (signal_5965) ) ;
    buf_clk cell_4123 ( .C (clk), .D (signal_5972), .Q (signal_5973) ) ;
    buf_clk cell_4131 ( .C (clk), .D (signal_5980), .Q (signal_5981) ) ;
    buf_clk cell_4139 ( .C (clk), .D (signal_5988), .Q (signal_5989) ) ;
    buf_clk cell_4147 ( .C (clk), .D (signal_5996), .Q (signal_5997) ) ;
    buf_clk cell_4155 ( .C (clk), .D (signal_6004), .Q (signal_6005) ) ;
    buf_clk cell_4163 ( .C (clk), .D (signal_6012), .Q (signal_6013) ) ;
    buf_clk cell_4171 ( .C (clk), .D (signal_6020), .Q (signal_6021) ) ;
    buf_clk cell_4179 ( .C (clk), .D (signal_6028), .Q (signal_6029) ) ;
    buf_clk cell_4187 ( .C (clk), .D (signal_6036), .Q (signal_6037) ) ;
    buf_clk cell_4195 ( .C (clk), .D (signal_6044), .Q (signal_6045) ) ;
    buf_clk cell_4203 ( .C (clk), .D (signal_6052), .Q (signal_6053) ) ;
    buf_clk cell_4211 ( .C (clk), .D (signal_6060), .Q (signal_6061) ) ;
    buf_clk cell_4219 ( .C (clk), .D (signal_6068), .Q (signal_6069) ) ;
    buf_clk cell_4227 ( .C (clk), .D (signal_6076), .Q (signal_6077) ) ;
    buf_clk cell_4235 ( .C (clk), .D (signal_6084), .Q (signal_6085) ) ;
    buf_clk cell_4243 ( .C (clk), .D (signal_6092), .Q (signal_6093) ) ;
    buf_clk cell_4251 ( .C (clk), .D (signal_6100), .Q (signal_6101) ) ;
    buf_clk cell_4259 ( .C (clk), .D (signal_6108), .Q (signal_6109) ) ;
    buf_clk cell_4267 ( .C (clk), .D (signal_6116), .Q (signal_6117) ) ;
    buf_clk cell_4275 ( .C (clk), .D (signal_6124), .Q (signal_6125) ) ;
    buf_clk cell_4283 ( .C (clk), .D (signal_6132), .Q (signal_6133) ) ;
    buf_clk cell_4291 ( .C (clk), .D (signal_6140), .Q (signal_6141) ) ;
    buf_clk cell_4299 ( .C (clk), .D (signal_6148), .Q (signal_6149) ) ;
    buf_clk cell_4307 ( .C (clk), .D (signal_6156), .Q (signal_6157) ) ;
    buf_clk cell_4315 ( .C (clk), .D (signal_6164), .Q (signal_6165) ) ;
    buf_clk cell_4323 ( .C (clk), .D (signal_6172), .Q (signal_6173) ) ;
    buf_clk cell_4331 ( .C (clk), .D (signal_6180), .Q (signal_6181) ) ;
    buf_clk cell_4339 ( .C (clk), .D (signal_6188), .Q (signal_6189) ) ;
    buf_clk cell_4347 ( .C (clk), .D (signal_6196), .Q (signal_6197) ) ;
    buf_clk cell_4355 ( .C (clk), .D (signal_6204), .Q (signal_6205) ) ;
    buf_clk cell_4363 ( .C (clk), .D (signal_6212), .Q (signal_6213) ) ;
    buf_clk cell_4371 ( .C (clk), .D (signal_6220), .Q (signal_6221) ) ;
    buf_clk cell_4379 ( .C (clk), .D (signal_6228), .Q (signal_6229) ) ;
    buf_clk cell_4387 ( .C (clk), .D (signal_6236), .Q (signal_6237) ) ;
    buf_clk cell_4395 ( .C (clk), .D (signal_6244), .Q (signal_6245) ) ;
    buf_clk cell_4403 ( .C (clk), .D (signal_6252), .Q (signal_6253) ) ;
    buf_clk cell_4411 ( .C (clk), .D (signal_6260), .Q (signal_6261) ) ;
    buf_clk cell_4419 ( .C (clk), .D (signal_6268), .Q (signal_6269) ) ;
    buf_clk cell_4427 ( .C (clk), .D (signal_6276), .Q (signal_6277) ) ;
    buf_clk cell_4435 ( .C (clk), .D (signal_6284), .Q (signal_6285) ) ;
    buf_clk cell_4443 ( .C (clk), .D (signal_6292), .Q (signal_6293) ) ;
    buf_clk cell_4451 ( .C (clk), .D (signal_6300), .Q (signal_6301) ) ;
    buf_clk cell_4459 ( .C (clk), .D (signal_6308), .Q (signal_6309) ) ;
    buf_clk cell_4467 ( .C (clk), .D (signal_6316), .Q (signal_6317) ) ;
    buf_clk cell_4475 ( .C (clk), .D (signal_6324), .Q (signal_6325) ) ;
    buf_clk cell_4483 ( .C (clk), .D (signal_6332), .Q (signal_6333) ) ;
    buf_clk cell_4491 ( .C (clk), .D (signal_6340), .Q (signal_6341) ) ;
    buf_clk cell_4499 ( .C (clk), .D (signal_6348), .Q (signal_6349) ) ;
    buf_clk cell_4507 ( .C (clk), .D (signal_6356), .Q (signal_6357) ) ;
    buf_clk cell_4515 ( .C (clk), .D (signal_6364), .Q (signal_6365) ) ;
    buf_clk cell_4523 ( .C (clk), .D (signal_6372), .Q (signal_6373) ) ;
    buf_clk cell_4531 ( .C (clk), .D (signal_6380), .Q (signal_6381) ) ;
    buf_clk cell_4539 ( .C (clk), .D (signal_6388), .Q (signal_6389) ) ;
    buf_clk cell_4547 ( .C (clk), .D (signal_6396), .Q (signal_6397) ) ;
    buf_clk cell_4555 ( .C (clk), .D (signal_6404), .Q (signal_6405) ) ;
    buf_clk cell_4563 ( .C (clk), .D (signal_6412), .Q (signal_6413) ) ;
    buf_clk cell_4571 ( .C (clk), .D (signal_6420), .Q (signal_6421) ) ;
    buf_clk cell_4579 ( .C (clk), .D (signal_6428), .Q (signal_6429) ) ;
    buf_clk cell_4587 ( .C (clk), .D (signal_6436), .Q (signal_6437) ) ;
    buf_clk cell_4595 ( .C (clk), .D (signal_6444), .Q (signal_6445) ) ;
    buf_clk cell_4603 ( .C (clk), .D (signal_6452), .Q (signal_6453) ) ;
    buf_clk cell_4611 ( .C (clk), .D (signal_6460), .Q (signal_6461) ) ;
    buf_clk cell_4619 ( .C (clk), .D (signal_6468), .Q (signal_6469) ) ;
    buf_clk cell_4627 ( .C (clk), .D (signal_6476), .Q (signal_6477) ) ;
    buf_clk cell_4635 ( .C (clk), .D (signal_6484), .Q (signal_6485) ) ;
    buf_clk cell_4643 ( .C (clk), .D (signal_6492), .Q (signal_6493) ) ;
    buf_clk cell_4651 ( .C (clk), .D (signal_6500), .Q (signal_6501) ) ;
    buf_clk cell_4659 ( .C (clk), .D (signal_6508), .Q (signal_6509) ) ;
    buf_clk cell_4667 ( .C (clk), .D (signal_6516), .Q (signal_6517) ) ;
    buf_clk cell_4675 ( .C (clk), .D (signal_6524), .Q (signal_6525) ) ;
    buf_clk cell_4683 ( .C (clk), .D (signal_6532), .Q (signal_6533) ) ;
    buf_clk cell_4691 ( .C (clk), .D (signal_6540), .Q (signal_6541) ) ;
    buf_clk cell_4699 ( .C (clk), .D (signal_6548), .Q (signal_6549) ) ;
    buf_clk cell_4707 ( .C (clk), .D (signal_6556), .Q (signal_6557) ) ;
    buf_clk cell_4715 ( .C (clk), .D (signal_6564), .Q (signal_6565) ) ;
    buf_clk cell_4723 ( .C (clk), .D (signal_6572), .Q (signal_6573) ) ;
    buf_clk cell_4731 ( .C (clk), .D (signal_6580), .Q (signal_6581) ) ;
    buf_clk cell_4739 ( .C (clk), .D (signal_6588), .Q (signal_6589) ) ;
    buf_clk cell_4747 ( .C (clk), .D (signal_6596), .Q (signal_6597) ) ;
    buf_clk cell_4755 ( .C (clk), .D (signal_6604), .Q (signal_6605) ) ;
    buf_clk cell_4763 ( .C (clk), .D (signal_6612), .Q (signal_6613) ) ;
    buf_clk cell_4771 ( .C (clk), .D (signal_6620), .Q (signal_6621) ) ;
    buf_clk cell_4779 ( .C (clk), .D (signal_6628), .Q (signal_6629) ) ;
    buf_clk cell_4787 ( .C (clk), .D (signal_6636), .Q (signal_6637) ) ;
    buf_clk cell_4795 ( .C (clk), .D (signal_6644), .Q (signal_6645) ) ;
    buf_clk cell_4803 ( .C (clk), .D (signal_6652), .Q (signal_6653) ) ;
    buf_clk cell_4811 ( .C (clk), .D (signal_6660), .Q (signal_6661) ) ;
    buf_clk cell_4819 ( .C (clk), .D (signal_6668), .Q (signal_6669) ) ;
    buf_clk cell_4827 ( .C (clk), .D (signal_6676), .Q (signal_6677) ) ;
    buf_clk cell_4835 ( .C (clk), .D (signal_6684), .Q (signal_6685) ) ;
    buf_clk cell_4843 ( .C (clk), .D (signal_6692), .Q (signal_6693) ) ;
    buf_clk cell_4851 ( .C (clk), .D (signal_6700), .Q (signal_6701) ) ;
    buf_clk cell_4859 ( .C (clk), .D (signal_6708), .Q (signal_6709) ) ;
    buf_clk cell_4867 ( .C (clk), .D (signal_6716), .Q (signal_6717) ) ;
    buf_clk cell_4875 ( .C (clk), .D (signal_6724), .Q (signal_6725) ) ;
    buf_clk cell_4883 ( .C (clk), .D (signal_6732), .Q (signal_6733) ) ;
    buf_clk cell_4891 ( .C (clk), .D (signal_6740), .Q (signal_6741) ) ;
    buf_clk cell_4899 ( .C (clk), .D (signal_6748), .Q (signal_6749) ) ;
    buf_clk cell_4907 ( .C (clk), .D (signal_6756), .Q (signal_6757) ) ;
    buf_clk cell_4915 ( .C (clk), .D (signal_6764), .Q (signal_6765) ) ;
    buf_clk cell_4923 ( .C (clk), .D (signal_6772), .Q (signal_6773) ) ;
    buf_clk cell_4931 ( .C (clk), .D (signal_6780), .Q (signal_6781) ) ;
    buf_clk cell_4939 ( .C (clk), .D (signal_6788), .Q (signal_6789) ) ;
    buf_clk cell_4947 ( .C (clk), .D (signal_6796), .Q (signal_6797) ) ;
    buf_clk cell_4955 ( .C (clk), .D (signal_6804), .Q (signal_6805) ) ;
    buf_clk cell_4963 ( .C (clk), .D (signal_6812), .Q (signal_6813) ) ;
    buf_clk cell_4971 ( .C (clk), .D (signal_6820), .Q (signal_6821) ) ;
    buf_clk cell_4979 ( .C (clk), .D (signal_6828), .Q (signal_6829) ) ;
    buf_clk cell_4987 ( .C (clk), .D (signal_6836), .Q (signal_6837) ) ;
    buf_clk cell_4995 ( .C (clk), .D (signal_6844), .Q (signal_6845) ) ;
    buf_clk cell_5003 ( .C (clk), .D (signal_6852), .Q (signal_6853) ) ;
    buf_clk cell_5011 ( .C (clk), .D (signal_6860), .Q (signal_6861) ) ;
    buf_clk cell_5019 ( .C (clk), .D (signal_6868), .Q (signal_6869) ) ;
    buf_clk cell_5027 ( .C (clk), .D (signal_6876), .Q (signal_6877) ) ;
    buf_clk cell_5035 ( .C (clk), .D (signal_6884), .Q (signal_6885) ) ;
    buf_clk cell_5043 ( .C (clk), .D (signal_6892), .Q (signal_6893) ) ;
    buf_clk cell_5051 ( .C (clk), .D (signal_6900), .Q (signal_6901) ) ;
    buf_clk cell_5059 ( .C (clk), .D (signal_6908), .Q (signal_6909) ) ;
    buf_clk cell_5067 ( .C (clk), .D (signal_6916), .Q (signal_6917) ) ;
    buf_clk cell_5075 ( .C (clk), .D (signal_6924), .Q (signal_6925) ) ;
    buf_clk cell_5083 ( .C (clk), .D (signal_6932), .Q (signal_6933) ) ;
    buf_clk cell_5091 ( .C (clk), .D (signal_6940), .Q (signal_6941) ) ;
    buf_clk cell_5099 ( .C (clk), .D (signal_6948), .Q (signal_6949) ) ;
    buf_clk cell_5107 ( .C (clk), .D (signal_6956), .Q (signal_6957) ) ;
    buf_clk cell_5115 ( .C (clk), .D (signal_6964), .Q (signal_6965) ) ;
    buf_clk cell_5123 ( .C (clk), .D (signal_6972), .Q (signal_6973) ) ;
    buf_clk cell_5131 ( .C (clk), .D (signal_6980), .Q (signal_6981) ) ;
    buf_clk cell_5139 ( .C (clk), .D (signal_6988), .Q (signal_6989) ) ;
    buf_clk cell_5147 ( .C (clk), .D (signal_6996), .Q (signal_6997) ) ;
    buf_clk cell_5155 ( .C (clk), .D (signal_7004), .Q (signal_7005) ) ;
    buf_clk cell_5163 ( .C (clk), .D (signal_7012), .Q (signal_7013) ) ;
    buf_clk cell_5171 ( .C (clk), .D (signal_7020), .Q (signal_7021) ) ;
    buf_clk cell_5179 ( .C (clk), .D (signal_7028), .Q (signal_7029) ) ;
    buf_clk cell_5187 ( .C (clk), .D (signal_7036), .Q (signal_7037) ) ;
    buf_clk cell_5195 ( .C (clk), .D (signal_7044), .Q (signal_7045) ) ;
    buf_clk cell_5203 ( .C (clk), .D (signal_7052), .Q (signal_7053) ) ;
    buf_clk cell_5211 ( .C (clk), .D (signal_7060), .Q (signal_7061) ) ;
    buf_clk cell_5219 ( .C (clk), .D (signal_7068), .Q (signal_7069) ) ;
    buf_clk cell_5227 ( .C (clk), .D (signal_7076), .Q (signal_7077) ) ;
    buf_clk cell_5235 ( .C (clk), .D (signal_7084), .Q (signal_7085) ) ;
    buf_clk cell_5243 ( .C (clk), .D (signal_7092), .Q (signal_7093) ) ;
    buf_clk cell_5251 ( .C (clk), .D (signal_7100), .Q (signal_7101) ) ;
    buf_clk cell_5259 ( .C (clk), .D (signal_7108), .Q (signal_7109) ) ;
    buf_clk cell_5267 ( .C (clk), .D (signal_7116), .Q (signal_7117) ) ;
    buf_clk cell_5275 ( .C (clk), .D (signal_7124), .Q (signal_7125) ) ;
    buf_clk cell_5283 ( .C (clk), .D (signal_7132), .Q (signal_7133) ) ;
    buf_clk cell_5291 ( .C (clk), .D (signal_7140), .Q (signal_7141) ) ;
    buf_clk cell_5299 ( .C (clk), .D (signal_7148), .Q (signal_7149) ) ;
    buf_clk cell_5307 ( .C (clk), .D (signal_7156), .Q (signal_7157) ) ;
    buf_clk cell_5315 ( .C (clk), .D (signal_7164), .Q (signal_7165) ) ;
    buf_clk cell_5323 ( .C (clk), .D (signal_7172), .Q (signal_7173) ) ;
    buf_clk cell_5331 ( .C (clk), .D (signal_7180), .Q (signal_7181) ) ;
    buf_clk cell_5339 ( .C (clk), .D (signal_7188), .Q (signal_7189) ) ;
    buf_clk cell_5347 ( .C (clk), .D (signal_7196), .Q (signal_7197) ) ;
    buf_clk cell_5355 ( .C (clk), .D (signal_7204), .Q (signal_7205) ) ;
    buf_clk cell_5363 ( .C (clk), .D (signal_7212), .Q (signal_7213) ) ;
    buf_clk cell_5371 ( .C (clk), .D (signal_7220), .Q (signal_7221) ) ;
    buf_clk cell_5379 ( .C (clk), .D (signal_7228), .Q (signal_7229) ) ;
    buf_clk cell_5387 ( .C (clk), .D (signal_7236), .Q (signal_7237) ) ;
    buf_clk cell_5395 ( .C (clk), .D (signal_7244), .Q (signal_7245) ) ;
    buf_clk cell_5403 ( .C (clk), .D (signal_7252), .Q (signal_7253) ) ;
    buf_clk cell_5411 ( .C (clk), .D (signal_7260), .Q (signal_7261) ) ;
    buf_clk cell_5419 ( .C (clk), .D (signal_7268), .Q (signal_7269) ) ;
    buf_clk cell_5427 ( .C (clk), .D (signal_7276), .Q (signal_7277) ) ;
    buf_clk cell_5435 ( .C (clk), .D (signal_7284), .Q (signal_7285) ) ;
    buf_clk cell_5443 ( .C (clk), .D (signal_7292), .Q (signal_7293) ) ;
    buf_clk cell_5451 ( .C (clk), .D (signal_7300), .Q (signal_7301) ) ;
    buf_clk cell_5459 ( .C (clk), .D (signal_7308), .Q (signal_7309) ) ;
    buf_clk cell_5467 ( .C (clk), .D (signal_7316), .Q (signal_7317) ) ;
    buf_clk cell_5475 ( .C (clk), .D (signal_7324), .Q (signal_7325) ) ;
    buf_clk cell_5483 ( .C (clk), .D (signal_7332), .Q (signal_7333) ) ;
    buf_clk cell_5491 ( .C (clk), .D (signal_7340), .Q (signal_7341) ) ;
    buf_clk cell_5499 ( .C (clk), .D (signal_7348), .Q (signal_7349) ) ;
    buf_clk cell_5507 ( .C (clk), .D (signal_7356), .Q (signal_7357) ) ;
    buf_clk cell_5515 ( .C (clk), .D (signal_7364), .Q (signal_7365) ) ;
    buf_clk cell_5523 ( .C (clk), .D (signal_7372), .Q (signal_7373) ) ;
    buf_clk cell_5531 ( .C (clk), .D (signal_7380), .Q (signal_7381) ) ;
    buf_clk cell_5539 ( .C (clk), .D (signal_7388), .Q (signal_7389) ) ;
    buf_clk cell_5547 ( .C (clk), .D (signal_7396), .Q (signal_7397) ) ;
    buf_clk cell_5555 ( .C (clk), .D (signal_7404), .Q (signal_7405) ) ;
    buf_clk cell_5563 ( .C (clk), .D (signal_7412), .Q (signal_7413) ) ;
    buf_clk cell_5571 ( .C (clk), .D (signal_7420), .Q (signal_7421) ) ;
    buf_clk cell_5579 ( .C (clk), .D (signal_7428), .Q (signal_7429) ) ;
    buf_clk cell_5587 ( .C (clk), .D (signal_7436), .Q (signal_7437) ) ;
    buf_clk cell_5595 ( .C (clk), .D (signal_7444), .Q (signal_7445) ) ;
    buf_clk cell_5603 ( .C (clk), .D (signal_7452), .Q (signal_7453) ) ;
    buf_clk cell_5611 ( .C (clk), .D (signal_7460), .Q (signal_7461) ) ;
    buf_clk cell_5619 ( .C (clk), .D (signal_7468), .Q (signal_7469) ) ;
    buf_clk cell_5627 ( .C (clk), .D (signal_7476), .Q (signal_7477) ) ;
    buf_clk cell_5635 ( .C (clk), .D (signal_7484), .Q (signal_7485) ) ;
    buf_clk cell_5643 ( .C (clk), .D (signal_7492), .Q (signal_7493) ) ;
    buf_clk cell_5651 ( .C (clk), .D (signal_7500), .Q (signal_7501) ) ;
    buf_clk cell_5659 ( .C (clk), .D (signal_7508), .Q (signal_7509) ) ;
    buf_clk cell_5667 ( .C (clk), .D (signal_7516), .Q (signal_7517) ) ;
    buf_clk cell_5675 ( .C (clk), .D (signal_7524), .Q (signal_7525) ) ;
    buf_clk cell_5683 ( .C (clk), .D (signal_7532), .Q (signal_7533) ) ;
    buf_clk cell_5691 ( .C (clk), .D (signal_7540), .Q (signal_7541) ) ;
    buf_clk cell_5699 ( .C (clk), .D (signal_7548), .Q (signal_7549) ) ;
    buf_clk cell_5707 ( .C (clk), .D (signal_7556), .Q (signal_7557) ) ;
    buf_clk cell_5715 ( .C (clk), .D (signal_7564), .Q (signal_7565) ) ;
    buf_clk cell_5723 ( .C (clk), .D (signal_7572), .Q (signal_7573) ) ;
    buf_clk cell_5731 ( .C (clk), .D (signal_7580), .Q (signal_7581) ) ;
    buf_clk cell_5739 ( .C (clk), .D (signal_7588), .Q (signal_7589) ) ;
    buf_clk cell_5747 ( .C (clk), .D (signal_7596), .Q (signal_7597) ) ;
    buf_clk cell_5755 ( .C (clk), .D (signal_7604), .Q (signal_7605) ) ;
    buf_clk cell_5763 ( .C (clk), .D (signal_7612), .Q (signal_7613) ) ;
    buf_clk cell_5771 ( .C (clk), .D (signal_7620), .Q (signal_7621) ) ;
    buf_clk cell_5779 ( .C (clk), .D (signal_7628), .Q (signal_7629) ) ;
    buf_clk cell_5787 ( .C (clk), .D (signal_7636), .Q (signal_7637) ) ;
    buf_clk cell_5795 ( .C (clk), .D (signal_7644), .Q (signal_7645) ) ;
    buf_clk cell_5803 ( .C (clk), .D (signal_7652), .Q (signal_7653) ) ;
    buf_clk cell_5811 ( .C (clk), .D (signal_7660), .Q (signal_7661) ) ;
    buf_clk cell_5819 ( .C (clk), .D (signal_7668), .Q (signal_7669) ) ;
    buf_clk cell_5827 ( .C (clk), .D (signal_7676), .Q (signal_7677) ) ;
    buf_clk cell_5835 ( .C (clk), .D (signal_7684), .Q (signal_7685) ) ;
    buf_clk cell_5843 ( .C (clk), .D (signal_7692), .Q (signal_7693) ) ;
    buf_clk cell_5851 ( .C (clk), .D (signal_7700), .Q (signal_7701) ) ;
    buf_clk cell_5859 ( .C (clk), .D (signal_7708), .Q (signal_7709) ) ;
    buf_clk cell_5867 ( .C (clk), .D (signal_7716), .Q (signal_7717) ) ;
    buf_clk cell_5875 ( .C (clk), .D (signal_7724), .Q (signal_7725) ) ;
    buf_clk cell_5883 ( .C (clk), .D (signal_7732), .Q (signal_7733) ) ;
    buf_clk cell_5891 ( .C (clk), .D (signal_7740), .Q (signal_7741) ) ;
    buf_clk cell_5899 ( .C (clk), .D (signal_7748), .Q (signal_7749) ) ;
    buf_clk cell_5907 ( .C (clk), .D (signal_7756), .Q (signal_7757) ) ;
    buf_clk cell_5915 ( .C (clk), .D (signal_7764), .Q (signal_7765) ) ;
    buf_clk cell_5923 ( .C (clk), .D (signal_7772), .Q (signal_7773) ) ;
    buf_clk cell_5931 ( .C (clk), .D (signal_7780), .Q (signal_7781) ) ;
    buf_clk cell_5939 ( .C (clk), .D (signal_7788), .Q (signal_7789) ) ;
    buf_clk cell_5947 ( .C (clk), .D (signal_7796), .Q (signal_7797) ) ;
    buf_clk cell_5955 ( .C (clk), .D (signal_7804), .Q (signal_7805) ) ;
    buf_clk cell_5963 ( .C (clk), .D (signal_7812), .Q (signal_7813) ) ;
    buf_clk cell_5971 ( .C (clk), .D (signal_7820), .Q (signal_7821) ) ;
    buf_clk cell_5979 ( .C (clk), .D (signal_7828), .Q (signal_7829) ) ;
    buf_clk cell_5987 ( .C (clk), .D (signal_7836), .Q (signal_7837) ) ;
    buf_clk cell_5995 ( .C (clk), .D (signal_7844), .Q (signal_7845) ) ;
    buf_clk cell_6003 ( .C (clk), .D (signal_7852), .Q (signal_7853) ) ;
    buf_clk cell_6011 ( .C (clk), .D (signal_7860), .Q (signal_7861) ) ;
    buf_clk cell_6019 ( .C (clk), .D (signal_7868), .Q (signal_7869) ) ;
    buf_clk cell_6027 ( .C (clk), .D (signal_7876), .Q (signal_7877) ) ;
    buf_clk cell_6035 ( .C (clk), .D (signal_7884), .Q (signal_7885) ) ;
    buf_clk cell_6043 ( .C (clk), .D (signal_7892), .Q (signal_7893) ) ;
    buf_clk cell_6051 ( .C (clk), .D (signal_7900), .Q (signal_7901) ) ;
    buf_clk cell_6059 ( .C (clk), .D (signal_7908), .Q (signal_7909) ) ;
    buf_clk cell_6067 ( .C (clk), .D (signal_7916), .Q (signal_7917) ) ;
    buf_clk cell_6075 ( .C (clk), .D (signal_7924), .Q (signal_7925) ) ;
    buf_clk cell_6083 ( .C (clk), .D (signal_7932), .Q (signal_7933) ) ;
    buf_clk cell_6091 ( .C (clk), .D (signal_7940), .Q (signal_7941) ) ;
    buf_clk cell_6099 ( .C (clk), .D (signal_7948), .Q (signal_7949) ) ;
    buf_clk cell_6107 ( .C (clk), .D (signal_7956), .Q (signal_7957) ) ;
    buf_clk cell_6115 ( .C (clk), .D (signal_7964), .Q (signal_7965) ) ;
    buf_clk cell_6123 ( .C (clk), .D (signal_7972), .Q (signal_7973) ) ;
    buf_clk cell_6131 ( .C (clk), .D (signal_7980), .Q (signal_7981) ) ;
    buf_clk cell_6139 ( .C (clk), .D (signal_7988), .Q (signal_7989) ) ;
    buf_clk cell_6147 ( .C (clk), .D (signal_7996), .Q (signal_7997) ) ;
    buf_clk cell_6155 ( .C (clk), .D (signal_8004), .Q (signal_8005) ) ;
    buf_clk cell_6163 ( .C (clk), .D (signal_8012), .Q (signal_8013) ) ;
    buf_clk cell_6171 ( .C (clk), .D (signal_8020), .Q (signal_8021) ) ;
    buf_clk cell_6179 ( .C (clk), .D (signal_8028), .Q (signal_8029) ) ;
    buf_clk cell_6187 ( .C (clk), .D (signal_8036), .Q (signal_8037) ) ;
    buf_clk cell_6195 ( .C (clk), .D (signal_8044), .Q (signal_8045) ) ;
    buf_clk cell_6203 ( .C (clk), .D (signal_8052), .Q (signal_8053) ) ;
    buf_clk cell_6211 ( .C (clk), .D (signal_8060), .Q (signal_8061) ) ;
    buf_clk cell_6219 ( .C (clk), .D (signal_8068), .Q (signal_8069) ) ;
    buf_clk cell_6227 ( .C (clk), .D (signal_8076), .Q (signal_8077) ) ;
    buf_clk cell_6235 ( .C (clk), .D (signal_8084), .Q (signal_8085) ) ;
    buf_clk cell_6243 ( .C (clk), .D (signal_8092), .Q (signal_8093) ) ;
    buf_clk cell_6251 ( .C (clk), .D (signal_8100), .Q (signal_8101) ) ;
    buf_clk cell_6259 ( .C (clk), .D (signal_8108), .Q (signal_8109) ) ;
    buf_clk cell_6267 ( .C (clk), .D (signal_8116), .Q (signal_8117) ) ;
    buf_clk cell_6275 ( .C (clk), .D (signal_8124), .Q (signal_8125) ) ;
    buf_clk cell_6283 ( .C (clk), .D (signal_8132), .Q (signal_8133) ) ;
    buf_clk cell_6291 ( .C (clk), .D (signal_8140), .Q (signal_8141) ) ;
    buf_clk cell_6299 ( .C (clk), .D (signal_8148), .Q (signal_8149) ) ;
    buf_clk cell_6307 ( .C (clk), .D (signal_8156), .Q (signal_8157) ) ;
    buf_clk cell_6315 ( .C (clk), .D (signal_8164), .Q (signal_8165) ) ;
    buf_clk cell_6323 ( .C (clk), .D (signal_8172), .Q (signal_8173) ) ;
    buf_clk cell_6331 ( .C (clk), .D (signal_8180), .Q (signal_8181) ) ;
    buf_clk cell_6339 ( .C (clk), .D (signal_8188), .Q (signal_8189) ) ;
    buf_clk cell_6347 ( .C (clk), .D (signal_8196), .Q (signal_8197) ) ;
    buf_clk cell_6355 ( .C (clk), .D (signal_8204), .Q (signal_8205) ) ;
    buf_clk cell_6363 ( .C (clk), .D (signal_8212), .Q (signal_8213) ) ;
    buf_clk cell_6371 ( .C (clk), .D (signal_8220), .Q (signal_8221) ) ;
    buf_clk cell_6379 ( .C (clk), .D (signal_8228), .Q (signal_8229) ) ;
    buf_clk cell_6387 ( .C (clk), .D (signal_8236), .Q (signal_8237) ) ;
    buf_clk cell_6395 ( .C (clk), .D (signal_8244), .Q (signal_8245) ) ;
    buf_clk cell_6403 ( .C (clk), .D (signal_8252), .Q (signal_8253) ) ;
    buf_clk cell_6411 ( .C (clk), .D (signal_8260), .Q (signal_8261) ) ;
    buf_clk cell_6419 ( .C (clk), .D (signal_8268), .Q (signal_8269) ) ;
    buf_clk cell_6427 ( .C (clk), .D (signal_8276), .Q (signal_8277) ) ;
    buf_clk cell_6435 ( .C (clk), .D (signal_8284), .Q (signal_8285) ) ;
    buf_clk cell_6443 ( .C (clk), .D (signal_8292), .Q (signal_8293) ) ;
    buf_clk cell_6451 ( .C (clk), .D (signal_8300), .Q (signal_8301) ) ;
    buf_clk cell_6459 ( .C (clk), .D (signal_8308), .Q (signal_8309) ) ;
    buf_clk cell_6467 ( .C (clk), .D (signal_8316), .Q (signal_8317) ) ;
    buf_clk cell_6475 ( .C (clk), .D (signal_8324), .Q (signal_8325) ) ;
    buf_clk cell_6483 ( .C (clk), .D (signal_8332), .Q (signal_8333) ) ;
    buf_clk cell_6491 ( .C (clk), .D (signal_8340), .Q (signal_8341) ) ;
    buf_clk cell_6499 ( .C (clk), .D (signal_8348), .Q (signal_8349) ) ;
    buf_clk cell_6507 ( .C (clk), .D (signal_8356), .Q (signal_8357) ) ;
    buf_clk cell_6515 ( .C (clk), .D (signal_8364), .Q (signal_8365) ) ;
    buf_clk cell_6523 ( .C (clk), .D (signal_8372), .Q (signal_8373) ) ;
    buf_clk cell_6531 ( .C (clk), .D (signal_8380), .Q (signal_8381) ) ;
    buf_clk cell_6539 ( .C (clk), .D (signal_8388), .Q (signal_8389) ) ;
    buf_clk cell_6547 ( .C (clk), .D (signal_8396), .Q (signal_8397) ) ;
    buf_clk cell_6555 ( .C (clk), .D (signal_8404), .Q (signal_8405) ) ;
    buf_clk cell_6563 ( .C (clk), .D (signal_8412), .Q (signal_8413) ) ;
    buf_clk cell_6571 ( .C (clk), .D (signal_8420), .Q (signal_8421) ) ;
    buf_clk cell_6579 ( .C (clk), .D (signal_8428), .Q (signal_8429) ) ;
    buf_clk cell_6587 ( .C (clk), .D (signal_8436), .Q (signal_8437) ) ;
    buf_clk cell_6595 ( .C (clk), .D (signal_8444), .Q (signal_8445) ) ;
    buf_clk cell_6603 ( .C (clk), .D (signal_8452), .Q (signal_8453) ) ;
    buf_clk cell_6611 ( .C (clk), .D (signal_8460), .Q (signal_8461) ) ;
    buf_clk cell_6619 ( .C (clk), .D (signal_8468), .Q (signal_8469) ) ;
    buf_clk cell_6627 ( .C (clk), .D (signal_8476), .Q (signal_8477) ) ;
    buf_clk cell_6635 ( .C (clk), .D (signal_8484), .Q (signal_8485) ) ;
    buf_clk cell_6643 ( .C (clk), .D (signal_8492), .Q (signal_8493) ) ;
    buf_clk cell_6651 ( .C (clk), .D (signal_8500), .Q (signal_8501) ) ;
    buf_clk cell_6659 ( .C (clk), .D (signal_8508), .Q (signal_8509) ) ;
    buf_clk cell_6667 ( .C (clk), .D (signal_8516), .Q (signal_8517) ) ;
    buf_clk cell_6675 ( .C (clk), .D (signal_8524), .Q (signal_8525) ) ;
    buf_clk cell_6683 ( .C (clk), .D (signal_8532), .Q (signal_8533) ) ;
    buf_clk cell_6691 ( .C (clk), .D (signal_8540), .Q (signal_8541) ) ;
    buf_clk cell_6699 ( .C (clk), .D (signal_8548), .Q (signal_8549) ) ;
    buf_clk cell_6707 ( .C (clk), .D (signal_8556), .Q (signal_8557) ) ;
    buf_clk cell_6715 ( .C (clk), .D (signal_8564), .Q (signal_8565) ) ;
    buf_clk cell_6723 ( .C (clk), .D (signal_8572), .Q (signal_8573) ) ;
    buf_clk cell_6731 ( .C (clk), .D (signal_8580), .Q (signal_8581) ) ;
    buf_clk cell_6739 ( .C (clk), .D (signal_8588), .Q (signal_8589) ) ;
    buf_clk cell_6747 ( .C (clk), .D (signal_8596), .Q (signal_8597) ) ;
    buf_clk cell_6755 ( .C (clk), .D (signal_8604), .Q (signal_8605) ) ;
    buf_clk cell_6763 ( .C (clk), .D (signal_8612), .Q (signal_8613) ) ;
    buf_clk cell_6771 ( .C (clk), .D (signal_8620), .Q (signal_8621) ) ;
    buf_clk cell_6779 ( .C (clk), .D (signal_8628), .Q (signal_8629) ) ;
    buf_clk cell_6787 ( .C (clk), .D (signal_8636), .Q (signal_8637) ) ;
    buf_clk cell_6795 ( .C (clk), .D (signal_8644), .Q (signal_8645) ) ;
    buf_clk cell_6803 ( .C (clk), .D (signal_8652), .Q (signal_8653) ) ;
    buf_clk cell_6811 ( .C (clk), .D (signal_8660), .Q (signal_8661) ) ;
    buf_clk cell_6819 ( .C (clk), .D (signal_8668), .Q (signal_8669) ) ;
    buf_clk cell_6827 ( .C (clk), .D (signal_8676), .Q (signal_8677) ) ;
    buf_clk cell_6835 ( .C (clk), .D (signal_8684), .Q (signal_8685) ) ;
    buf_clk cell_6843 ( .C (clk), .D (signal_8692), .Q (signal_8693) ) ;
    buf_clk cell_6851 ( .C (clk), .D (signal_8700), .Q (signal_8701) ) ;
    buf_clk cell_6859 ( .C (clk), .D (signal_8708), .Q (signal_8709) ) ;
    buf_clk cell_6867 ( .C (clk), .D (signal_8716), .Q (signal_8717) ) ;
    buf_clk cell_6875 ( .C (clk), .D (signal_8724), .Q (signal_8725) ) ;
    buf_clk cell_6883 ( .C (clk), .D (signal_8732), .Q (signal_8733) ) ;
    buf_clk cell_6891 ( .C (clk), .D (signal_8740), .Q (signal_8741) ) ;
    buf_clk cell_6899 ( .C (clk), .D (signal_8748), .Q (signal_8749) ) ;
    buf_clk cell_6907 ( .C (clk), .D (signal_8756), .Q (signal_8757) ) ;
    buf_clk cell_6915 ( .C (clk), .D (signal_8764), .Q (signal_8765) ) ;
    buf_clk cell_6923 ( .C (clk), .D (signal_8772), .Q (signal_8773) ) ;
    buf_clk cell_6931 ( .C (clk), .D (signal_8780), .Q (signal_8781) ) ;
    buf_clk cell_6939 ( .C (clk), .D (signal_8788), .Q (signal_8789) ) ;
    buf_clk cell_6947 ( .C (clk), .D (signal_8796), .Q (signal_8797) ) ;
    buf_clk cell_6955 ( .C (clk), .D (signal_8804), .Q (signal_8805) ) ;
    buf_clk cell_6963 ( .C (clk), .D (signal_8812), .Q (signal_8813) ) ;
    buf_clk cell_6971 ( .C (clk), .D (signal_8820), .Q (signal_8821) ) ;
    buf_clk cell_6979 ( .C (clk), .D (signal_8828), .Q (signal_8829) ) ;
    buf_clk cell_6987 ( .C (clk), .D (signal_8836), .Q (signal_8837) ) ;
    buf_clk cell_6995 ( .C (clk), .D (signal_8844), .Q (signal_8845) ) ;
    buf_clk cell_7003 ( .C (clk), .D (signal_8852), .Q (signal_8853) ) ;
    buf_clk cell_7011 ( .C (clk), .D (signal_8860), .Q (signal_8861) ) ;
    buf_clk cell_7019 ( .C (clk), .D (signal_8868), .Q (signal_8869) ) ;
    buf_clk cell_7027 ( .C (clk), .D (signal_8876), .Q (signal_8877) ) ;
    buf_clk cell_7035 ( .C (clk), .D (signal_8884), .Q (signal_8885) ) ;
    buf_clk cell_7043 ( .C (clk), .D (signal_8892), .Q (signal_8893) ) ;
    buf_clk cell_7051 ( .C (clk), .D (signal_8900), .Q (signal_8901) ) ;
    buf_clk cell_7059 ( .C (clk), .D (signal_8908), .Q (signal_8909) ) ;
    buf_clk cell_7067 ( .C (clk), .D (signal_8916), .Q (signal_8917) ) ;
    buf_clk cell_7075 ( .C (clk), .D (signal_8924), .Q (signal_8925) ) ;
    buf_clk cell_7083 ( .C (clk), .D (signal_8932), .Q (signal_8933) ) ;
    buf_clk cell_7091 ( .C (clk), .D (signal_8940), .Q (signal_8941) ) ;
    buf_clk cell_7099 ( .C (clk), .D (signal_8948), .Q (signal_8949) ) ;

    /* cells in depth 7 */
    buf_clk cell_1900 ( .C (clk), .D (signal_3749), .Q (signal_3750) ) ;
    buf_clk cell_1908 ( .C (clk), .D (signal_3757), .Q (signal_3758) ) ;
    buf_clk cell_1916 ( .C (clk), .D (signal_3765), .Q (signal_3766) ) ;
    buf_clk cell_1924 ( .C (clk), .D (signal_3773), .Q (signal_3774) ) ;
    buf_clk cell_1932 ( .C (clk), .D (signal_3781), .Q (signal_3782) ) ;
    buf_clk cell_1940 ( .C (clk), .D (signal_3789), .Q (signal_3790) ) ;
    buf_clk cell_1948 ( .C (clk), .D (signal_3797), .Q (signal_3798) ) ;
    buf_clk cell_1956 ( .C (clk), .D (signal_3805), .Q (signal_3806) ) ;
    buf_clk cell_1964 ( .C (clk), .D (signal_3813), .Q (signal_3814) ) ;
    buf_clk cell_1972 ( .C (clk), .D (signal_3821), .Q (signal_3822) ) ;
    buf_clk cell_1980 ( .C (clk), .D (signal_3829), .Q (signal_3830) ) ;
    buf_clk cell_1988 ( .C (clk), .D (signal_3837), .Q (signal_3838) ) ;
    buf_clk cell_1996 ( .C (clk), .D (signal_3845), .Q (signal_3846) ) ;
    buf_clk cell_2004 ( .C (clk), .D (signal_3853), .Q (signal_3854) ) ;
    buf_clk cell_2012 ( .C (clk), .D (signal_3861), .Q (signal_3862) ) ;
    buf_clk cell_2020 ( .C (clk), .D (signal_3869), .Q (signal_3870) ) ;
    buf_clk cell_2028 ( .C (clk), .D (signal_3877), .Q (signal_3878) ) ;
    buf_clk cell_2036 ( .C (clk), .D (signal_3885), .Q (signal_3886) ) ;
    buf_clk cell_2044 ( .C (clk), .D (signal_3893), .Q (signal_3894) ) ;
    buf_clk cell_2052 ( .C (clk), .D (signal_3901), .Q (signal_3902) ) ;
    buf_clk cell_2060 ( .C (clk), .D (signal_3909), .Q (signal_3910) ) ;
    buf_clk cell_2068 ( .C (clk), .D (signal_3917), .Q (signal_3918) ) ;
    buf_clk cell_2076 ( .C (clk), .D (signal_3925), .Q (signal_3926) ) ;
    buf_clk cell_2084 ( .C (clk), .D (signal_3933), .Q (signal_3934) ) ;
    buf_clk cell_2092 ( .C (clk), .D (signal_3941), .Q (signal_3942) ) ;
    buf_clk cell_2100 ( .C (clk), .D (signal_3949), .Q (signal_3950) ) ;
    buf_clk cell_2108 ( .C (clk), .D (signal_3957), .Q (signal_3958) ) ;
    buf_clk cell_2116 ( .C (clk), .D (signal_3965), .Q (signal_3966) ) ;
    buf_clk cell_2124 ( .C (clk), .D (signal_3973), .Q (signal_3974) ) ;
    buf_clk cell_2132 ( .C (clk), .D (signal_3981), .Q (signal_3982) ) ;
    buf_clk cell_2140 ( .C (clk), .D (signal_3989), .Q (signal_3990) ) ;
    buf_clk cell_2148 ( .C (clk), .D (signal_3997), .Q (signal_3998) ) ;
    buf_clk cell_2156 ( .C (clk), .D (signal_4005), .Q (signal_4006) ) ;
    buf_clk cell_2164 ( .C (clk), .D (signal_4013), .Q (signal_4014) ) ;
    buf_clk cell_2172 ( .C (clk), .D (signal_4021), .Q (signal_4022) ) ;
    buf_clk cell_2180 ( .C (clk), .D (signal_4029), .Q (signal_4030) ) ;
    buf_clk cell_2188 ( .C (clk), .D (signal_4037), .Q (signal_4038) ) ;
    buf_clk cell_2196 ( .C (clk), .D (signal_4045), .Q (signal_4046) ) ;
    buf_clk cell_2204 ( .C (clk), .D (signal_4053), .Q (signal_4054) ) ;
    buf_clk cell_2212 ( .C (clk), .D (signal_4061), .Q (signal_4062) ) ;
    buf_clk cell_2220 ( .C (clk), .D (signal_4069), .Q (signal_4070) ) ;
    buf_clk cell_2228 ( .C (clk), .D (signal_4077), .Q (signal_4078) ) ;
    buf_clk cell_2236 ( .C (clk), .D (signal_4085), .Q (signal_4086) ) ;
    buf_clk cell_2244 ( .C (clk), .D (signal_4093), .Q (signal_4094) ) ;
    buf_clk cell_2252 ( .C (clk), .D (signal_4101), .Q (signal_4102) ) ;
    buf_clk cell_2260 ( .C (clk), .D (signal_4109), .Q (signal_4110) ) ;
    buf_clk cell_2268 ( .C (clk), .D (signal_4117), .Q (signal_4118) ) ;
    buf_clk cell_2276 ( .C (clk), .D (signal_4125), .Q (signal_4126) ) ;
    buf_clk cell_2284 ( .C (clk), .D (signal_4133), .Q (signal_4134) ) ;
    buf_clk cell_2292 ( .C (clk), .D (signal_4141), .Q (signal_4142) ) ;
    buf_clk cell_2300 ( .C (clk), .D (signal_4149), .Q (signal_4150) ) ;
    buf_clk cell_2308 ( .C (clk), .D (signal_4157), .Q (signal_4158) ) ;
    buf_clk cell_2316 ( .C (clk), .D (signal_4165), .Q (signal_4166) ) ;
    buf_clk cell_2324 ( .C (clk), .D (signal_4173), .Q (signal_4174) ) ;
    buf_clk cell_2332 ( .C (clk), .D (signal_4181), .Q (signal_4182) ) ;
    buf_clk cell_2340 ( .C (clk), .D (signal_4189), .Q (signal_4190) ) ;
    buf_clk cell_2348 ( .C (clk), .D (signal_4197), .Q (signal_4198) ) ;
    buf_clk cell_2356 ( .C (clk), .D (signal_4205), .Q (signal_4206) ) ;
    buf_clk cell_2364 ( .C (clk), .D (signal_4213), .Q (signal_4214) ) ;
    buf_clk cell_2372 ( .C (clk), .D (signal_4221), .Q (signal_4222) ) ;
    buf_clk cell_2380 ( .C (clk), .D (signal_4229), .Q (signal_4230) ) ;
    buf_clk cell_2388 ( .C (clk), .D (signal_4237), .Q (signal_4238) ) ;
    buf_clk cell_2396 ( .C (clk), .D (signal_4245), .Q (signal_4246) ) ;
    buf_clk cell_2404 ( .C (clk), .D (signal_4253), .Q (signal_4254) ) ;
    buf_clk cell_2412 ( .C (clk), .D (signal_4261), .Q (signal_4262) ) ;
    buf_clk cell_2420 ( .C (clk), .D (signal_4269), .Q (signal_4270) ) ;
    buf_clk cell_2428 ( .C (clk), .D (signal_4277), .Q (signal_4278) ) ;
    buf_clk cell_2436 ( .C (clk), .D (signal_4285), .Q (signal_4286) ) ;
    buf_clk cell_2444 ( .C (clk), .D (signal_4293), .Q (signal_4294) ) ;
    buf_clk cell_2452 ( .C (clk), .D (signal_4301), .Q (signal_4302) ) ;
    buf_clk cell_2460 ( .C (clk), .D (signal_4309), .Q (signal_4310) ) ;
    buf_clk cell_2468 ( .C (clk), .D (signal_4317), .Q (signal_4318) ) ;
    buf_clk cell_2476 ( .C (clk), .D (signal_4325), .Q (signal_4326) ) ;
    buf_clk cell_2484 ( .C (clk), .D (signal_4333), .Q (signal_4334) ) ;
    buf_clk cell_2492 ( .C (clk), .D (signal_4341), .Q (signal_4342) ) ;
    buf_clk cell_2500 ( .C (clk), .D (signal_4349), .Q (signal_4350) ) ;
    buf_clk cell_2508 ( .C (clk), .D (signal_4357), .Q (signal_4358) ) ;
    buf_clk cell_2516 ( .C (clk), .D (signal_4365), .Q (signal_4366) ) ;
    buf_clk cell_2524 ( .C (clk), .D (signal_4373), .Q (signal_4374) ) ;
    buf_clk cell_2532 ( .C (clk), .D (signal_4381), .Q (signal_4382) ) ;
    buf_clk cell_2540 ( .C (clk), .D (signal_4389), .Q (signal_4390) ) ;
    buf_clk cell_2548 ( .C (clk), .D (signal_4397), .Q (signal_4398) ) ;
    buf_clk cell_2556 ( .C (clk), .D (signal_4405), .Q (signal_4406) ) ;
    buf_clk cell_2564 ( .C (clk), .D (signal_4413), .Q (signal_4414) ) ;
    buf_clk cell_2572 ( .C (clk), .D (signal_4421), .Q (signal_4422) ) ;
    buf_clk cell_2580 ( .C (clk), .D (signal_4429), .Q (signal_4430) ) ;
    buf_clk cell_2588 ( .C (clk), .D (signal_4437), .Q (signal_4438) ) ;
    buf_clk cell_2596 ( .C (clk), .D (signal_4445), .Q (signal_4446) ) ;
    buf_clk cell_2604 ( .C (clk), .D (signal_4453), .Q (signal_4454) ) ;
    buf_clk cell_2612 ( .C (clk), .D (signal_4461), .Q (signal_4462) ) ;
    buf_clk cell_2620 ( .C (clk), .D (signal_4469), .Q (signal_4470) ) ;
    buf_clk cell_2628 ( .C (clk), .D (signal_4477), .Q (signal_4478) ) ;
    buf_clk cell_2636 ( .C (clk), .D (signal_4485), .Q (signal_4486) ) ;
    buf_clk cell_2644 ( .C (clk), .D (signal_4493), .Q (signal_4494) ) ;
    buf_clk cell_2652 ( .C (clk), .D (signal_4501), .Q (signal_4502) ) ;
    buf_clk cell_2660 ( .C (clk), .D (signal_4509), .Q (signal_4510) ) ;
    buf_clk cell_2668 ( .C (clk), .D (signal_4517), .Q (signal_4518) ) ;
    buf_clk cell_2676 ( .C (clk), .D (signal_4525), .Q (signal_4526) ) ;
    buf_clk cell_2684 ( .C (clk), .D (signal_4533), .Q (signal_4534) ) ;
    buf_clk cell_2692 ( .C (clk), .D (signal_4541), .Q (signal_4542) ) ;
    buf_clk cell_2700 ( .C (clk), .D (signal_4549), .Q (signal_4550) ) ;
    buf_clk cell_2708 ( .C (clk), .D (signal_4557), .Q (signal_4558) ) ;
    buf_clk cell_2716 ( .C (clk), .D (signal_4565), .Q (signal_4566) ) ;
    buf_clk cell_2724 ( .C (clk), .D (signal_4573), .Q (signal_4574) ) ;
    buf_clk cell_2732 ( .C (clk), .D (signal_4581), .Q (signal_4582) ) ;
    buf_clk cell_2740 ( .C (clk), .D (signal_4589), .Q (signal_4590) ) ;
    buf_clk cell_2748 ( .C (clk), .D (signal_4597), .Q (signal_4598) ) ;
    buf_clk cell_2756 ( .C (clk), .D (signal_4605), .Q (signal_4606) ) ;
    buf_clk cell_2764 ( .C (clk), .D (signal_4613), .Q (signal_4614) ) ;
    buf_clk cell_2772 ( .C (clk), .D (signal_4621), .Q (signal_4622) ) ;
    buf_clk cell_2780 ( .C (clk), .D (signal_4629), .Q (signal_4630) ) ;
    buf_clk cell_2788 ( .C (clk), .D (signal_4637), .Q (signal_4638) ) ;
    buf_clk cell_2796 ( .C (clk), .D (signal_4645), .Q (signal_4646) ) ;
    buf_clk cell_2804 ( .C (clk), .D (signal_4653), .Q (signal_4654) ) ;
    buf_clk cell_2812 ( .C (clk), .D (signal_4661), .Q (signal_4662) ) ;
    buf_clk cell_2820 ( .C (clk), .D (signal_4669), .Q (signal_4670) ) ;
    buf_clk cell_2828 ( .C (clk), .D (signal_4677), .Q (signal_4678) ) ;
    buf_clk cell_2836 ( .C (clk), .D (signal_4685), .Q (signal_4686) ) ;
    buf_clk cell_2844 ( .C (clk), .D (signal_4693), .Q (signal_4694) ) ;
    buf_clk cell_2852 ( .C (clk), .D (signal_4701), .Q (signal_4702) ) ;
    buf_clk cell_2860 ( .C (clk), .D (signal_4709), .Q (signal_4710) ) ;
    buf_clk cell_2868 ( .C (clk), .D (signal_4717), .Q (signal_4718) ) ;
    buf_clk cell_2876 ( .C (clk), .D (signal_4725), .Q (signal_4726) ) ;
    buf_clk cell_2884 ( .C (clk), .D (signal_4733), .Q (signal_4734) ) ;
    buf_clk cell_2892 ( .C (clk), .D (signal_4741), .Q (signal_4742) ) ;
    buf_clk cell_2900 ( .C (clk), .D (signal_4749), .Q (signal_4750) ) ;
    buf_clk cell_3124 ( .C (clk), .D (signal_4973), .Q (signal_4974) ) ;
    buf_clk cell_3132 ( .C (clk), .D (signal_4981), .Q (signal_4982) ) ;
    buf_clk cell_3140 ( .C (clk), .D (signal_4989), .Q (signal_4990) ) ;
    buf_clk cell_3148 ( .C (clk), .D (signal_4997), .Q (signal_4998) ) ;
    buf_clk cell_3156 ( .C (clk), .D (signal_5005), .Q (signal_5006) ) ;
    buf_clk cell_3164 ( .C (clk), .D (signal_5013), .Q (signal_5014) ) ;
    buf_clk cell_3172 ( .C (clk), .D (signal_5021), .Q (signal_5022) ) ;
    buf_clk cell_3180 ( .C (clk), .D (signal_5029), .Q (signal_5030) ) ;
    buf_clk cell_3188 ( .C (clk), .D (signal_5037), .Q (signal_5038) ) ;
    buf_clk cell_3196 ( .C (clk), .D (signal_5045), .Q (signal_5046) ) ;
    buf_clk cell_3204 ( .C (clk), .D (signal_5053), .Q (signal_5054) ) ;
    buf_clk cell_3212 ( .C (clk), .D (signal_5061), .Q (signal_5062) ) ;
    buf_clk cell_3220 ( .C (clk), .D (signal_5069), .Q (signal_5070) ) ;
    buf_clk cell_3228 ( .C (clk), .D (signal_5077), .Q (signal_5078) ) ;
    buf_clk cell_3236 ( .C (clk), .D (signal_5085), .Q (signal_5086) ) ;
    buf_clk cell_3244 ( .C (clk), .D (signal_5093), .Q (signal_5094) ) ;
    buf_clk cell_3252 ( .C (clk), .D (signal_5101), .Q (signal_5102) ) ;
    buf_clk cell_3260 ( .C (clk), .D (signal_5109), .Q (signal_5110) ) ;
    buf_clk cell_3268 ( .C (clk), .D (signal_5117), .Q (signal_5118) ) ;
    buf_clk cell_3276 ( .C (clk), .D (signal_5125), .Q (signal_5126) ) ;
    buf_clk cell_3284 ( .C (clk), .D (signal_5133), .Q (signal_5134) ) ;
    buf_clk cell_3292 ( .C (clk), .D (signal_5141), .Q (signal_5142) ) ;
    buf_clk cell_3300 ( .C (clk), .D (signal_5149), .Q (signal_5150) ) ;
    buf_clk cell_3308 ( .C (clk), .D (signal_5157), .Q (signal_5158) ) ;
    buf_clk cell_3316 ( .C (clk), .D (signal_5165), .Q (signal_5166) ) ;
    buf_clk cell_3324 ( .C (clk), .D (signal_5173), .Q (signal_5174) ) ;
    buf_clk cell_3332 ( .C (clk), .D (signal_5181), .Q (signal_5182) ) ;
    buf_clk cell_3340 ( .C (clk), .D (signal_5189), .Q (signal_5190) ) ;
    buf_clk cell_3348 ( .C (clk), .D (signal_5197), .Q (signal_5198) ) ;
    buf_clk cell_3356 ( .C (clk), .D (signal_5205), .Q (signal_5206) ) ;
    buf_clk cell_3364 ( .C (clk), .D (signal_5213), .Q (signal_5214) ) ;
    buf_clk cell_3372 ( .C (clk), .D (signal_5221), .Q (signal_5222) ) ;
    buf_clk cell_3380 ( .C (clk), .D (signal_5229), .Q (signal_5230) ) ;
    buf_clk cell_3388 ( .C (clk), .D (signal_5237), .Q (signal_5238) ) ;
    buf_clk cell_3396 ( .C (clk), .D (signal_5245), .Q (signal_5246) ) ;
    buf_clk cell_3404 ( .C (clk), .D (signal_5253), .Q (signal_5254) ) ;
    buf_clk cell_3412 ( .C (clk), .D (signal_5261), .Q (signal_5262) ) ;
    buf_clk cell_3420 ( .C (clk), .D (signal_5269), .Q (signal_5270) ) ;
    buf_clk cell_3428 ( .C (clk), .D (signal_5277), .Q (signal_5278) ) ;
    buf_clk cell_3436 ( .C (clk), .D (signal_5285), .Q (signal_5286) ) ;
    buf_clk cell_3444 ( .C (clk), .D (signal_5293), .Q (signal_5294) ) ;
    buf_clk cell_3452 ( .C (clk), .D (signal_5301), .Q (signal_5302) ) ;
    buf_clk cell_3460 ( .C (clk), .D (signal_5309), .Q (signal_5310) ) ;
    buf_clk cell_3468 ( .C (clk), .D (signal_5317), .Q (signal_5318) ) ;
    buf_clk cell_3476 ( .C (clk), .D (signal_5325), .Q (signal_5326) ) ;
    buf_clk cell_3484 ( .C (clk), .D (signal_5333), .Q (signal_5334) ) ;
    buf_clk cell_3492 ( .C (clk), .D (signal_5341), .Q (signal_5342) ) ;
    buf_clk cell_3500 ( .C (clk), .D (signal_5349), .Q (signal_5350) ) ;
    buf_clk cell_3508 ( .C (clk), .D (signal_5357), .Q (signal_5358) ) ;
    buf_clk cell_3516 ( .C (clk), .D (signal_5365), .Q (signal_5366) ) ;
    buf_clk cell_3524 ( .C (clk), .D (signal_5373), .Q (signal_5374) ) ;
    buf_clk cell_3532 ( .C (clk), .D (signal_5381), .Q (signal_5382) ) ;
    buf_clk cell_3540 ( .C (clk), .D (signal_5389), .Q (signal_5390) ) ;
    buf_clk cell_3548 ( .C (clk), .D (signal_5397), .Q (signal_5398) ) ;
    buf_clk cell_3556 ( .C (clk), .D (signal_5405), .Q (signal_5406) ) ;
    buf_clk cell_3564 ( .C (clk), .D (signal_5413), .Q (signal_5414) ) ;
    buf_clk cell_3572 ( .C (clk), .D (signal_5421), .Q (signal_5422) ) ;
    buf_clk cell_3580 ( .C (clk), .D (signal_5429), .Q (signal_5430) ) ;
    buf_clk cell_3588 ( .C (clk), .D (signal_5437), .Q (signal_5438) ) ;
    buf_clk cell_3596 ( .C (clk), .D (signal_5445), .Q (signal_5446) ) ;
    buf_clk cell_3604 ( .C (clk), .D (signal_5453), .Q (signal_5454) ) ;
    buf_clk cell_3612 ( .C (clk), .D (signal_5461), .Q (signal_5462) ) ;
    buf_clk cell_3620 ( .C (clk), .D (signal_5469), .Q (signal_5470) ) ;
    buf_clk cell_3628 ( .C (clk), .D (signal_5477), .Q (signal_5478) ) ;
    buf_clk cell_3636 ( .C (clk), .D (signal_5485), .Q (signal_5486) ) ;
    buf_clk cell_3644 ( .C (clk), .D (signal_5493), .Q (signal_5494) ) ;
    buf_clk cell_3652 ( .C (clk), .D (signal_5501), .Q (signal_5502) ) ;
    buf_clk cell_3660 ( .C (clk), .D (signal_5509), .Q (signal_5510) ) ;
    buf_clk cell_3668 ( .C (clk), .D (signal_5517), .Q (signal_5518) ) ;
    buf_clk cell_3676 ( .C (clk), .D (signal_5525), .Q (signal_5526) ) ;
    buf_clk cell_3684 ( .C (clk), .D (signal_5533), .Q (signal_5534) ) ;
    buf_clk cell_3692 ( .C (clk), .D (signal_5541), .Q (signal_5542) ) ;
    buf_clk cell_3700 ( .C (clk), .D (signal_5549), .Q (signal_5550) ) ;
    buf_clk cell_3708 ( .C (clk), .D (signal_5557), .Q (signal_5558) ) ;
    buf_clk cell_3716 ( .C (clk), .D (signal_5565), .Q (signal_5566) ) ;
    buf_clk cell_3724 ( .C (clk), .D (signal_5573), .Q (signal_5574) ) ;
    buf_clk cell_3732 ( .C (clk), .D (signal_5581), .Q (signal_5582) ) ;
    buf_clk cell_3740 ( .C (clk), .D (signal_5589), .Q (signal_5590) ) ;
    buf_clk cell_3748 ( .C (clk), .D (signal_5597), .Q (signal_5598) ) ;
    buf_clk cell_3756 ( .C (clk), .D (signal_5605), .Q (signal_5606) ) ;
    buf_clk cell_3764 ( .C (clk), .D (signal_5613), .Q (signal_5614) ) ;
    buf_clk cell_3772 ( .C (clk), .D (signal_5621), .Q (signal_5622) ) ;
    buf_clk cell_3780 ( .C (clk), .D (signal_5629), .Q (signal_5630) ) ;
    buf_clk cell_3788 ( .C (clk), .D (signal_5637), .Q (signal_5638) ) ;
    buf_clk cell_3796 ( .C (clk), .D (signal_5645), .Q (signal_5646) ) ;
    buf_clk cell_3804 ( .C (clk), .D (signal_5653), .Q (signal_5654) ) ;
    buf_clk cell_3812 ( .C (clk), .D (signal_5661), .Q (signal_5662) ) ;
    buf_clk cell_3820 ( .C (clk), .D (signal_5669), .Q (signal_5670) ) ;
    buf_clk cell_3828 ( .C (clk), .D (signal_5677), .Q (signal_5678) ) ;
    buf_clk cell_3836 ( .C (clk), .D (signal_5685), .Q (signal_5686) ) ;
    buf_clk cell_3844 ( .C (clk), .D (signal_5693), .Q (signal_5694) ) ;
    buf_clk cell_3852 ( .C (clk), .D (signal_5701), .Q (signal_5702) ) ;
    buf_clk cell_3860 ( .C (clk), .D (signal_5709), .Q (signal_5710) ) ;
    buf_clk cell_3868 ( .C (clk), .D (signal_5717), .Q (signal_5718) ) ;
    buf_clk cell_3876 ( .C (clk), .D (signal_5725), .Q (signal_5726) ) ;
    buf_clk cell_3884 ( .C (clk), .D (signal_5733), .Q (signal_5734) ) ;
    buf_clk cell_3892 ( .C (clk), .D (signal_5741), .Q (signal_5742) ) ;
    buf_clk cell_3900 ( .C (clk), .D (signal_5749), .Q (signal_5750) ) ;
    buf_clk cell_3908 ( .C (clk), .D (signal_5757), .Q (signal_5758) ) ;
    buf_clk cell_3916 ( .C (clk), .D (signal_5765), .Q (signal_5766) ) ;
    buf_clk cell_3924 ( .C (clk), .D (signal_5773), .Q (signal_5774) ) ;
    buf_clk cell_3932 ( .C (clk), .D (signal_5781), .Q (signal_5782) ) ;
    buf_clk cell_3940 ( .C (clk), .D (signal_5789), .Q (signal_5790) ) ;
    buf_clk cell_3948 ( .C (clk), .D (signal_5797), .Q (signal_5798) ) ;
    buf_clk cell_3956 ( .C (clk), .D (signal_5805), .Q (signal_5806) ) ;
    buf_clk cell_3964 ( .C (clk), .D (signal_5813), .Q (signal_5814) ) ;
    buf_clk cell_3972 ( .C (clk), .D (signal_5821), .Q (signal_5822) ) ;
    buf_clk cell_3980 ( .C (clk), .D (signal_5829), .Q (signal_5830) ) ;
    buf_clk cell_3988 ( .C (clk), .D (signal_5837), .Q (signal_5838) ) ;
    buf_clk cell_3996 ( .C (clk), .D (signal_5845), .Q (signal_5846) ) ;
    buf_clk cell_4004 ( .C (clk), .D (signal_5853), .Q (signal_5854) ) ;
    buf_clk cell_4012 ( .C (clk), .D (signal_5861), .Q (signal_5862) ) ;
    buf_clk cell_4020 ( .C (clk), .D (signal_5869), .Q (signal_5870) ) ;
    buf_clk cell_4028 ( .C (clk), .D (signal_5877), .Q (signal_5878) ) ;
    buf_clk cell_4036 ( .C (clk), .D (signal_5885), .Q (signal_5886) ) ;
    buf_clk cell_4044 ( .C (clk), .D (signal_5893), .Q (signal_5894) ) ;
    buf_clk cell_4052 ( .C (clk), .D (signal_5901), .Q (signal_5902) ) ;
    buf_clk cell_4060 ( .C (clk), .D (signal_5909), .Q (signal_5910) ) ;
    buf_clk cell_4068 ( .C (clk), .D (signal_5917), .Q (signal_5918) ) ;
    buf_clk cell_4076 ( .C (clk), .D (signal_5925), .Q (signal_5926) ) ;
    buf_clk cell_4084 ( .C (clk), .D (signal_5933), .Q (signal_5934) ) ;
    buf_clk cell_4092 ( .C (clk), .D (signal_5941), .Q (signal_5942) ) ;
    buf_clk cell_4100 ( .C (clk), .D (signal_5949), .Q (signal_5950) ) ;
    buf_clk cell_4108 ( .C (clk), .D (signal_5957), .Q (signal_5958) ) ;
    buf_clk cell_4116 ( .C (clk), .D (signal_5965), .Q (signal_5966) ) ;
    buf_clk cell_4124 ( .C (clk), .D (signal_5973), .Q (signal_5974) ) ;
    buf_clk cell_4132 ( .C (clk), .D (signal_5981), .Q (signal_5982) ) ;
    buf_clk cell_4140 ( .C (clk), .D (signal_5989), .Q (signal_5990) ) ;
    buf_clk cell_4148 ( .C (clk), .D (signal_5997), .Q (signal_5998) ) ;
    buf_clk cell_4156 ( .C (clk), .D (signal_6005), .Q (signal_6006) ) ;
    buf_clk cell_4164 ( .C (clk), .D (signal_6013), .Q (signal_6014) ) ;
    buf_clk cell_4172 ( .C (clk), .D (signal_6021), .Q (signal_6022) ) ;
    buf_clk cell_4180 ( .C (clk), .D (signal_6029), .Q (signal_6030) ) ;
    buf_clk cell_4188 ( .C (clk), .D (signal_6037), .Q (signal_6038) ) ;
    buf_clk cell_4196 ( .C (clk), .D (signal_6045), .Q (signal_6046) ) ;
    buf_clk cell_4204 ( .C (clk), .D (signal_6053), .Q (signal_6054) ) ;
    buf_clk cell_4212 ( .C (clk), .D (signal_6061), .Q (signal_6062) ) ;
    buf_clk cell_4220 ( .C (clk), .D (signal_6069), .Q (signal_6070) ) ;
    buf_clk cell_4228 ( .C (clk), .D (signal_6077), .Q (signal_6078) ) ;
    buf_clk cell_4236 ( .C (clk), .D (signal_6085), .Q (signal_6086) ) ;
    buf_clk cell_4244 ( .C (clk), .D (signal_6093), .Q (signal_6094) ) ;
    buf_clk cell_4252 ( .C (clk), .D (signal_6101), .Q (signal_6102) ) ;
    buf_clk cell_4260 ( .C (clk), .D (signal_6109), .Q (signal_6110) ) ;
    buf_clk cell_4268 ( .C (clk), .D (signal_6117), .Q (signal_6118) ) ;
    buf_clk cell_4276 ( .C (clk), .D (signal_6125), .Q (signal_6126) ) ;
    buf_clk cell_4284 ( .C (clk), .D (signal_6133), .Q (signal_6134) ) ;
    buf_clk cell_4292 ( .C (clk), .D (signal_6141), .Q (signal_6142) ) ;
    buf_clk cell_4300 ( .C (clk), .D (signal_6149), .Q (signal_6150) ) ;
    buf_clk cell_4308 ( .C (clk), .D (signal_6157), .Q (signal_6158) ) ;
    buf_clk cell_4316 ( .C (clk), .D (signal_6165), .Q (signal_6166) ) ;
    buf_clk cell_4324 ( .C (clk), .D (signal_6173), .Q (signal_6174) ) ;
    buf_clk cell_4332 ( .C (clk), .D (signal_6181), .Q (signal_6182) ) ;
    buf_clk cell_4340 ( .C (clk), .D (signal_6189), .Q (signal_6190) ) ;
    buf_clk cell_4348 ( .C (clk), .D (signal_6197), .Q (signal_6198) ) ;
    buf_clk cell_4356 ( .C (clk), .D (signal_6205), .Q (signal_6206) ) ;
    buf_clk cell_4364 ( .C (clk), .D (signal_6213), .Q (signal_6214) ) ;
    buf_clk cell_4372 ( .C (clk), .D (signal_6221), .Q (signal_6222) ) ;
    buf_clk cell_4380 ( .C (clk), .D (signal_6229), .Q (signal_6230) ) ;
    buf_clk cell_4388 ( .C (clk), .D (signal_6237), .Q (signal_6238) ) ;
    buf_clk cell_4396 ( .C (clk), .D (signal_6245), .Q (signal_6246) ) ;
    buf_clk cell_4404 ( .C (clk), .D (signal_6253), .Q (signal_6254) ) ;
    buf_clk cell_4412 ( .C (clk), .D (signal_6261), .Q (signal_6262) ) ;
    buf_clk cell_4420 ( .C (clk), .D (signal_6269), .Q (signal_6270) ) ;
    buf_clk cell_4428 ( .C (clk), .D (signal_6277), .Q (signal_6278) ) ;
    buf_clk cell_4436 ( .C (clk), .D (signal_6285), .Q (signal_6286) ) ;
    buf_clk cell_4444 ( .C (clk), .D (signal_6293), .Q (signal_6294) ) ;
    buf_clk cell_4452 ( .C (clk), .D (signal_6301), .Q (signal_6302) ) ;
    buf_clk cell_4460 ( .C (clk), .D (signal_6309), .Q (signal_6310) ) ;
    buf_clk cell_4468 ( .C (clk), .D (signal_6317), .Q (signal_6318) ) ;
    buf_clk cell_4476 ( .C (clk), .D (signal_6325), .Q (signal_6326) ) ;
    buf_clk cell_4484 ( .C (clk), .D (signal_6333), .Q (signal_6334) ) ;
    buf_clk cell_4492 ( .C (clk), .D (signal_6341), .Q (signal_6342) ) ;
    buf_clk cell_4500 ( .C (clk), .D (signal_6349), .Q (signal_6350) ) ;
    buf_clk cell_4508 ( .C (clk), .D (signal_6357), .Q (signal_6358) ) ;
    buf_clk cell_4516 ( .C (clk), .D (signal_6365), .Q (signal_6366) ) ;
    buf_clk cell_4524 ( .C (clk), .D (signal_6373), .Q (signal_6374) ) ;
    buf_clk cell_4532 ( .C (clk), .D (signal_6381), .Q (signal_6382) ) ;
    buf_clk cell_4540 ( .C (clk), .D (signal_6389), .Q (signal_6390) ) ;
    buf_clk cell_4548 ( .C (clk), .D (signal_6397), .Q (signal_6398) ) ;
    buf_clk cell_4556 ( .C (clk), .D (signal_6405), .Q (signal_6406) ) ;
    buf_clk cell_4564 ( .C (clk), .D (signal_6413), .Q (signal_6414) ) ;
    buf_clk cell_4572 ( .C (clk), .D (signal_6421), .Q (signal_6422) ) ;
    buf_clk cell_4580 ( .C (clk), .D (signal_6429), .Q (signal_6430) ) ;
    buf_clk cell_4588 ( .C (clk), .D (signal_6437), .Q (signal_6438) ) ;
    buf_clk cell_4596 ( .C (clk), .D (signal_6445), .Q (signal_6446) ) ;
    buf_clk cell_4604 ( .C (clk), .D (signal_6453), .Q (signal_6454) ) ;
    buf_clk cell_4612 ( .C (clk), .D (signal_6461), .Q (signal_6462) ) ;
    buf_clk cell_4620 ( .C (clk), .D (signal_6469), .Q (signal_6470) ) ;
    buf_clk cell_4628 ( .C (clk), .D (signal_6477), .Q (signal_6478) ) ;
    buf_clk cell_4636 ( .C (clk), .D (signal_6485), .Q (signal_6486) ) ;
    buf_clk cell_4644 ( .C (clk), .D (signal_6493), .Q (signal_6494) ) ;
    buf_clk cell_4652 ( .C (clk), .D (signal_6501), .Q (signal_6502) ) ;
    buf_clk cell_4660 ( .C (clk), .D (signal_6509), .Q (signal_6510) ) ;
    buf_clk cell_4668 ( .C (clk), .D (signal_6517), .Q (signal_6518) ) ;
    buf_clk cell_4676 ( .C (clk), .D (signal_6525), .Q (signal_6526) ) ;
    buf_clk cell_4684 ( .C (clk), .D (signal_6533), .Q (signal_6534) ) ;
    buf_clk cell_4692 ( .C (clk), .D (signal_6541), .Q (signal_6542) ) ;
    buf_clk cell_4700 ( .C (clk), .D (signal_6549), .Q (signal_6550) ) ;
    buf_clk cell_4708 ( .C (clk), .D (signal_6557), .Q (signal_6558) ) ;
    buf_clk cell_4716 ( .C (clk), .D (signal_6565), .Q (signal_6566) ) ;
    buf_clk cell_4724 ( .C (clk), .D (signal_6573), .Q (signal_6574) ) ;
    buf_clk cell_4732 ( .C (clk), .D (signal_6581), .Q (signal_6582) ) ;
    buf_clk cell_4740 ( .C (clk), .D (signal_6589), .Q (signal_6590) ) ;
    buf_clk cell_4748 ( .C (clk), .D (signal_6597), .Q (signal_6598) ) ;
    buf_clk cell_4756 ( .C (clk), .D (signal_6605), .Q (signal_6606) ) ;
    buf_clk cell_4764 ( .C (clk), .D (signal_6613), .Q (signal_6614) ) ;
    buf_clk cell_4772 ( .C (clk), .D (signal_6621), .Q (signal_6622) ) ;
    buf_clk cell_4780 ( .C (clk), .D (signal_6629), .Q (signal_6630) ) ;
    buf_clk cell_4788 ( .C (clk), .D (signal_6637), .Q (signal_6638) ) ;
    buf_clk cell_4796 ( .C (clk), .D (signal_6645), .Q (signal_6646) ) ;
    buf_clk cell_4804 ( .C (clk), .D (signal_6653), .Q (signal_6654) ) ;
    buf_clk cell_4812 ( .C (clk), .D (signal_6661), .Q (signal_6662) ) ;
    buf_clk cell_4820 ( .C (clk), .D (signal_6669), .Q (signal_6670) ) ;
    buf_clk cell_4828 ( .C (clk), .D (signal_6677), .Q (signal_6678) ) ;
    buf_clk cell_4836 ( .C (clk), .D (signal_6685), .Q (signal_6686) ) ;
    buf_clk cell_4844 ( .C (clk), .D (signal_6693), .Q (signal_6694) ) ;
    buf_clk cell_4852 ( .C (clk), .D (signal_6701), .Q (signal_6702) ) ;
    buf_clk cell_4860 ( .C (clk), .D (signal_6709), .Q (signal_6710) ) ;
    buf_clk cell_4868 ( .C (clk), .D (signal_6717), .Q (signal_6718) ) ;
    buf_clk cell_4876 ( .C (clk), .D (signal_6725), .Q (signal_6726) ) ;
    buf_clk cell_4884 ( .C (clk), .D (signal_6733), .Q (signal_6734) ) ;
    buf_clk cell_4892 ( .C (clk), .D (signal_6741), .Q (signal_6742) ) ;
    buf_clk cell_4900 ( .C (clk), .D (signal_6749), .Q (signal_6750) ) ;
    buf_clk cell_4908 ( .C (clk), .D (signal_6757), .Q (signal_6758) ) ;
    buf_clk cell_4916 ( .C (clk), .D (signal_6765), .Q (signal_6766) ) ;
    buf_clk cell_4924 ( .C (clk), .D (signal_6773), .Q (signal_6774) ) ;
    buf_clk cell_4932 ( .C (clk), .D (signal_6781), .Q (signal_6782) ) ;
    buf_clk cell_4940 ( .C (clk), .D (signal_6789), .Q (signal_6790) ) ;
    buf_clk cell_4948 ( .C (clk), .D (signal_6797), .Q (signal_6798) ) ;
    buf_clk cell_4956 ( .C (clk), .D (signal_6805), .Q (signal_6806) ) ;
    buf_clk cell_4964 ( .C (clk), .D (signal_6813), .Q (signal_6814) ) ;
    buf_clk cell_4972 ( .C (clk), .D (signal_6821), .Q (signal_6822) ) ;
    buf_clk cell_4980 ( .C (clk), .D (signal_6829), .Q (signal_6830) ) ;
    buf_clk cell_4988 ( .C (clk), .D (signal_6837), .Q (signal_6838) ) ;
    buf_clk cell_4996 ( .C (clk), .D (signal_6845), .Q (signal_6846) ) ;
    buf_clk cell_5004 ( .C (clk), .D (signal_6853), .Q (signal_6854) ) ;
    buf_clk cell_5012 ( .C (clk), .D (signal_6861), .Q (signal_6862) ) ;
    buf_clk cell_5020 ( .C (clk), .D (signal_6869), .Q (signal_6870) ) ;
    buf_clk cell_5028 ( .C (clk), .D (signal_6877), .Q (signal_6878) ) ;
    buf_clk cell_5036 ( .C (clk), .D (signal_6885), .Q (signal_6886) ) ;
    buf_clk cell_5044 ( .C (clk), .D (signal_6893), .Q (signal_6894) ) ;
    buf_clk cell_5052 ( .C (clk), .D (signal_6901), .Q (signal_6902) ) ;
    buf_clk cell_5060 ( .C (clk), .D (signal_6909), .Q (signal_6910) ) ;
    buf_clk cell_5068 ( .C (clk), .D (signal_6917), .Q (signal_6918) ) ;
    buf_clk cell_5076 ( .C (clk), .D (signal_6925), .Q (signal_6926) ) ;
    buf_clk cell_5084 ( .C (clk), .D (signal_6933), .Q (signal_6934) ) ;
    buf_clk cell_5092 ( .C (clk), .D (signal_6941), .Q (signal_6942) ) ;
    buf_clk cell_5100 ( .C (clk), .D (signal_6949), .Q (signal_6950) ) ;
    buf_clk cell_5108 ( .C (clk), .D (signal_6957), .Q (signal_6958) ) ;
    buf_clk cell_5116 ( .C (clk), .D (signal_6965), .Q (signal_6966) ) ;
    buf_clk cell_5124 ( .C (clk), .D (signal_6973), .Q (signal_6974) ) ;
    buf_clk cell_5132 ( .C (clk), .D (signal_6981), .Q (signal_6982) ) ;
    buf_clk cell_5140 ( .C (clk), .D (signal_6989), .Q (signal_6990) ) ;
    buf_clk cell_5148 ( .C (clk), .D (signal_6997), .Q (signal_6998) ) ;
    buf_clk cell_5156 ( .C (clk), .D (signal_7005), .Q (signal_7006) ) ;
    buf_clk cell_5164 ( .C (clk), .D (signal_7013), .Q (signal_7014) ) ;
    buf_clk cell_5172 ( .C (clk), .D (signal_7021), .Q (signal_7022) ) ;
    buf_clk cell_5180 ( .C (clk), .D (signal_7029), .Q (signal_7030) ) ;
    buf_clk cell_5188 ( .C (clk), .D (signal_7037), .Q (signal_7038) ) ;
    buf_clk cell_5196 ( .C (clk), .D (signal_7045), .Q (signal_7046) ) ;
    buf_clk cell_5204 ( .C (clk), .D (signal_7053), .Q (signal_7054) ) ;
    buf_clk cell_5212 ( .C (clk), .D (signal_7061), .Q (signal_7062) ) ;
    buf_clk cell_5220 ( .C (clk), .D (signal_7069), .Q (signal_7070) ) ;
    buf_clk cell_5228 ( .C (clk), .D (signal_7077), .Q (signal_7078) ) ;
    buf_clk cell_5236 ( .C (clk), .D (signal_7085), .Q (signal_7086) ) ;
    buf_clk cell_5244 ( .C (clk), .D (signal_7093), .Q (signal_7094) ) ;
    buf_clk cell_5252 ( .C (clk), .D (signal_7101), .Q (signal_7102) ) ;
    buf_clk cell_5260 ( .C (clk), .D (signal_7109), .Q (signal_7110) ) ;
    buf_clk cell_5268 ( .C (clk), .D (signal_7117), .Q (signal_7118) ) ;
    buf_clk cell_5276 ( .C (clk), .D (signal_7125), .Q (signal_7126) ) ;
    buf_clk cell_5284 ( .C (clk), .D (signal_7133), .Q (signal_7134) ) ;
    buf_clk cell_5292 ( .C (clk), .D (signal_7141), .Q (signal_7142) ) ;
    buf_clk cell_5300 ( .C (clk), .D (signal_7149), .Q (signal_7150) ) ;
    buf_clk cell_5308 ( .C (clk), .D (signal_7157), .Q (signal_7158) ) ;
    buf_clk cell_5316 ( .C (clk), .D (signal_7165), .Q (signal_7166) ) ;
    buf_clk cell_5324 ( .C (clk), .D (signal_7173), .Q (signal_7174) ) ;
    buf_clk cell_5332 ( .C (clk), .D (signal_7181), .Q (signal_7182) ) ;
    buf_clk cell_5340 ( .C (clk), .D (signal_7189), .Q (signal_7190) ) ;
    buf_clk cell_5348 ( .C (clk), .D (signal_7197), .Q (signal_7198) ) ;
    buf_clk cell_5356 ( .C (clk), .D (signal_7205), .Q (signal_7206) ) ;
    buf_clk cell_5364 ( .C (clk), .D (signal_7213), .Q (signal_7214) ) ;
    buf_clk cell_5372 ( .C (clk), .D (signal_7221), .Q (signal_7222) ) ;
    buf_clk cell_5380 ( .C (clk), .D (signal_7229), .Q (signal_7230) ) ;
    buf_clk cell_5388 ( .C (clk), .D (signal_7237), .Q (signal_7238) ) ;
    buf_clk cell_5396 ( .C (clk), .D (signal_7245), .Q (signal_7246) ) ;
    buf_clk cell_5404 ( .C (clk), .D (signal_7253), .Q (signal_7254) ) ;
    buf_clk cell_5412 ( .C (clk), .D (signal_7261), .Q (signal_7262) ) ;
    buf_clk cell_5420 ( .C (clk), .D (signal_7269), .Q (signal_7270) ) ;
    buf_clk cell_5428 ( .C (clk), .D (signal_7277), .Q (signal_7278) ) ;
    buf_clk cell_5436 ( .C (clk), .D (signal_7285), .Q (signal_7286) ) ;
    buf_clk cell_5444 ( .C (clk), .D (signal_7293), .Q (signal_7294) ) ;
    buf_clk cell_5452 ( .C (clk), .D (signal_7301), .Q (signal_7302) ) ;
    buf_clk cell_5460 ( .C (clk), .D (signal_7309), .Q (signal_7310) ) ;
    buf_clk cell_5468 ( .C (clk), .D (signal_7317), .Q (signal_7318) ) ;
    buf_clk cell_5476 ( .C (clk), .D (signal_7325), .Q (signal_7326) ) ;
    buf_clk cell_5484 ( .C (clk), .D (signal_7333), .Q (signal_7334) ) ;
    buf_clk cell_5492 ( .C (clk), .D (signal_7341), .Q (signal_7342) ) ;
    buf_clk cell_5500 ( .C (clk), .D (signal_7349), .Q (signal_7350) ) ;
    buf_clk cell_5508 ( .C (clk), .D (signal_7357), .Q (signal_7358) ) ;
    buf_clk cell_5516 ( .C (clk), .D (signal_7365), .Q (signal_7366) ) ;
    buf_clk cell_5524 ( .C (clk), .D (signal_7373), .Q (signal_7374) ) ;
    buf_clk cell_5532 ( .C (clk), .D (signal_7381), .Q (signal_7382) ) ;
    buf_clk cell_5540 ( .C (clk), .D (signal_7389), .Q (signal_7390) ) ;
    buf_clk cell_5548 ( .C (clk), .D (signal_7397), .Q (signal_7398) ) ;
    buf_clk cell_5556 ( .C (clk), .D (signal_7405), .Q (signal_7406) ) ;
    buf_clk cell_5564 ( .C (clk), .D (signal_7413), .Q (signal_7414) ) ;
    buf_clk cell_5572 ( .C (clk), .D (signal_7421), .Q (signal_7422) ) ;
    buf_clk cell_5580 ( .C (clk), .D (signal_7429), .Q (signal_7430) ) ;
    buf_clk cell_5588 ( .C (clk), .D (signal_7437), .Q (signal_7438) ) ;
    buf_clk cell_5596 ( .C (clk), .D (signal_7445), .Q (signal_7446) ) ;
    buf_clk cell_5604 ( .C (clk), .D (signal_7453), .Q (signal_7454) ) ;
    buf_clk cell_5612 ( .C (clk), .D (signal_7461), .Q (signal_7462) ) ;
    buf_clk cell_5620 ( .C (clk), .D (signal_7469), .Q (signal_7470) ) ;
    buf_clk cell_5628 ( .C (clk), .D (signal_7477), .Q (signal_7478) ) ;
    buf_clk cell_5636 ( .C (clk), .D (signal_7485), .Q (signal_7486) ) ;
    buf_clk cell_5644 ( .C (clk), .D (signal_7493), .Q (signal_7494) ) ;
    buf_clk cell_5652 ( .C (clk), .D (signal_7501), .Q (signal_7502) ) ;
    buf_clk cell_5660 ( .C (clk), .D (signal_7509), .Q (signal_7510) ) ;
    buf_clk cell_5668 ( .C (clk), .D (signal_7517), .Q (signal_7518) ) ;
    buf_clk cell_5676 ( .C (clk), .D (signal_7525), .Q (signal_7526) ) ;
    buf_clk cell_5684 ( .C (clk), .D (signal_7533), .Q (signal_7534) ) ;
    buf_clk cell_5692 ( .C (clk), .D (signal_7541), .Q (signal_7542) ) ;
    buf_clk cell_5700 ( .C (clk), .D (signal_7549), .Q (signal_7550) ) ;
    buf_clk cell_5708 ( .C (clk), .D (signal_7557), .Q (signal_7558) ) ;
    buf_clk cell_5716 ( .C (clk), .D (signal_7565), .Q (signal_7566) ) ;
    buf_clk cell_5724 ( .C (clk), .D (signal_7573), .Q (signal_7574) ) ;
    buf_clk cell_5732 ( .C (clk), .D (signal_7581), .Q (signal_7582) ) ;
    buf_clk cell_5740 ( .C (clk), .D (signal_7589), .Q (signal_7590) ) ;
    buf_clk cell_5748 ( .C (clk), .D (signal_7597), .Q (signal_7598) ) ;
    buf_clk cell_5756 ( .C (clk), .D (signal_7605), .Q (signal_7606) ) ;
    buf_clk cell_5764 ( .C (clk), .D (signal_7613), .Q (signal_7614) ) ;
    buf_clk cell_5772 ( .C (clk), .D (signal_7621), .Q (signal_7622) ) ;
    buf_clk cell_5780 ( .C (clk), .D (signal_7629), .Q (signal_7630) ) ;
    buf_clk cell_5788 ( .C (clk), .D (signal_7637), .Q (signal_7638) ) ;
    buf_clk cell_5796 ( .C (clk), .D (signal_7645), .Q (signal_7646) ) ;
    buf_clk cell_5804 ( .C (clk), .D (signal_7653), .Q (signal_7654) ) ;
    buf_clk cell_5812 ( .C (clk), .D (signal_7661), .Q (signal_7662) ) ;
    buf_clk cell_5820 ( .C (clk), .D (signal_7669), .Q (signal_7670) ) ;
    buf_clk cell_5828 ( .C (clk), .D (signal_7677), .Q (signal_7678) ) ;
    buf_clk cell_5836 ( .C (clk), .D (signal_7685), .Q (signal_7686) ) ;
    buf_clk cell_5844 ( .C (clk), .D (signal_7693), .Q (signal_7694) ) ;
    buf_clk cell_5852 ( .C (clk), .D (signal_7701), .Q (signal_7702) ) ;
    buf_clk cell_5860 ( .C (clk), .D (signal_7709), .Q (signal_7710) ) ;
    buf_clk cell_5868 ( .C (clk), .D (signal_7717), .Q (signal_7718) ) ;
    buf_clk cell_5876 ( .C (clk), .D (signal_7725), .Q (signal_7726) ) ;
    buf_clk cell_5884 ( .C (clk), .D (signal_7733), .Q (signal_7734) ) ;
    buf_clk cell_5892 ( .C (clk), .D (signal_7741), .Q (signal_7742) ) ;
    buf_clk cell_5900 ( .C (clk), .D (signal_7749), .Q (signal_7750) ) ;
    buf_clk cell_5908 ( .C (clk), .D (signal_7757), .Q (signal_7758) ) ;
    buf_clk cell_5916 ( .C (clk), .D (signal_7765), .Q (signal_7766) ) ;
    buf_clk cell_5924 ( .C (clk), .D (signal_7773), .Q (signal_7774) ) ;
    buf_clk cell_5932 ( .C (clk), .D (signal_7781), .Q (signal_7782) ) ;
    buf_clk cell_5940 ( .C (clk), .D (signal_7789), .Q (signal_7790) ) ;
    buf_clk cell_5948 ( .C (clk), .D (signal_7797), .Q (signal_7798) ) ;
    buf_clk cell_5956 ( .C (clk), .D (signal_7805), .Q (signal_7806) ) ;
    buf_clk cell_5964 ( .C (clk), .D (signal_7813), .Q (signal_7814) ) ;
    buf_clk cell_5972 ( .C (clk), .D (signal_7821), .Q (signal_7822) ) ;
    buf_clk cell_5980 ( .C (clk), .D (signal_7829), .Q (signal_7830) ) ;
    buf_clk cell_5988 ( .C (clk), .D (signal_7837), .Q (signal_7838) ) ;
    buf_clk cell_5996 ( .C (clk), .D (signal_7845), .Q (signal_7846) ) ;
    buf_clk cell_6004 ( .C (clk), .D (signal_7853), .Q (signal_7854) ) ;
    buf_clk cell_6012 ( .C (clk), .D (signal_7861), .Q (signal_7862) ) ;
    buf_clk cell_6020 ( .C (clk), .D (signal_7869), .Q (signal_7870) ) ;
    buf_clk cell_6028 ( .C (clk), .D (signal_7877), .Q (signal_7878) ) ;
    buf_clk cell_6036 ( .C (clk), .D (signal_7885), .Q (signal_7886) ) ;
    buf_clk cell_6044 ( .C (clk), .D (signal_7893), .Q (signal_7894) ) ;
    buf_clk cell_6052 ( .C (clk), .D (signal_7901), .Q (signal_7902) ) ;
    buf_clk cell_6060 ( .C (clk), .D (signal_7909), .Q (signal_7910) ) ;
    buf_clk cell_6068 ( .C (clk), .D (signal_7917), .Q (signal_7918) ) ;
    buf_clk cell_6076 ( .C (clk), .D (signal_7925), .Q (signal_7926) ) ;
    buf_clk cell_6084 ( .C (clk), .D (signal_7933), .Q (signal_7934) ) ;
    buf_clk cell_6092 ( .C (clk), .D (signal_7941), .Q (signal_7942) ) ;
    buf_clk cell_6100 ( .C (clk), .D (signal_7949), .Q (signal_7950) ) ;
    buf_clk cell_6108 ( .C (clk), .D (signal_7957), .Q (signal_7958) ) ;
    buf_clk cell_6116 ( .C (clk), .D (signal_7965), .Q (signal_7966) ) ;
    buf_clk cell_6124 ( .C (clk), .D (signal_7973), .Q (signal_7974) ) ;
    buf_clk cell_6132 ( .C (clk), .D (signal_7981), .Q (signal_7982) ) ;
    buf_clk cell_6140 ( .C (clk), .D (signal_7989), .Q (signal_7990) ) ;
    buf_clk cell_6148 ( .C (clk), .D (signal_7997), .Q (signal_7998) ) ;
    buf_clk cell_6156 ( .C (clk), .D (signal_8005), .Q (signal_8006) ) ;
    buf_clk cell_6164 ( .C (clk), .D (signal_8013), .Q (signal_8014) ) ;
    buf_clk cell_6172 ( .C (clk), .D (signal_8021), .Q (signal_8022) ) ;
    buf_clk cell_6180 ( .C (clk), .D (signal_8029), .Q (signal_8030) ) ;
    buf_clk cell_6188 ( .C (clk), .D (signal_8037), .Q (signal_8038) ) ;
    buf_clk cell_6196 ( .C (clk), .D (signal_8045), .Q (signal_8046) ) ;
    buf_clk cell_6204 ( .C (clk), .D (signal_8053), .Q (signal_8054) ) ;
    buf_clk cell_6212 ( .C (clk), .D (signal_8061), .Q (signal_8062) ) ;
    buf_clk cell_6220 ( .C (clk), .D (signal_8069), .Q (signal_8070) ) ;
    buf_clk cell_6228 ( .C (clk), .D (signal_8077), .Q (signal_8078) ) ;
    buf_clk cell_6236 ( .C (clk), .D (signal_8085), .Q (signal_8086) ) ;
    buf_clk cell_6244 ( .C (clk), .D (signal_8093), .Q (signal_8094) ) ;
    buf_clk cell_6252 ( .C (clk), .D (signal_8101), .Q (signal_8102) ) ;
    buf_clk cell_6260 ( .C (clk), .D (signal_8109), .Q (signal_8110) ) ;
    buf_clk cell_6268 ( .C (clk), .D (signal_8117), .Q (signal_8118) ) ;
    buf_clk cell_6276 ( .C (clk), .D (signal_8125), .Q (signal_8126) ) ;
    buf_clk cell_6284 ( .C (clk), .D (signal_8133), .Q (signal_8134) ) ;
    buf_clk cell_6292 ( .C (clk), .D (signal_8141), .Q (signal_8142) ) ;
    buf_clk cell_6300 ( .C (clk), .D (signal_8149), .Q (signal_8150) ) ;
    buf_clk cell_6308 ( .C (clk), .D (signal_8157), .Q (signal_8158) ) ;
    buf_clk cell_6316 ( .C (clk), .D (signal_8165), .Q (signal_8166) ) ;
    buf_clk cell_6324 ( .C (clk), .D (signal_8173), .Q (signal_8174) ) ;
    buf_clk cell_6332 ( .C (clk), .D (signal_8181), .Q (signal_8182) ) ;
    buf_clk cell_6340 ( .C (clk), .D (signal_8189), .Q (signal_8190) ) ;
    buf_clk cell_6348 ( .C (clk), .D (signal_8197), .Q (signal_8198) ) ;
    buf_clk cell_6356 ( .C (clk), .D (signal_8205), .Q (signal_8206) ) ;
    buf_clk cell_6364 ( .C (clk), .D (signal_8213), .Q (signal_8214) ) ;
    buf_clk cell_6372 ( .C (clk), .D (signal_8221), .Q (signal_8222) ) ;
    buf_clk cell_6380 ( .C (clk), .D (signal_8229), .Q (signal_8230) ) ;
    buf_clk cell_6388 ( .C (clk), .D (signal_8237), .Q (signal_8238) ) ;
    buf_clk cell_6396 ( .C (clk), .D (signal_8245), .Q (signal_8246) ) ;
    buf_clk cell_6404 ( .C (clk), .D (signal_8253), .Q (signal_8254) ) ;
    buf_clk cell_6412 ( .C (clk), .D (signal_8261), .Q (signal_8262) ) ;
    buf_clk cell_6420 ( .C (clk), .D (signal_8269), .Q (signal_8270) ) ;
    buf_clk cell_6428 ( .C (clk), .D (signal_8277), .Q (signal_8278) ) ;
    buf_clk cell_6436 ( .C (clk), .D (signal_8285), .Q (signal_8286) ) ;
    buf_clk cell_6444 ( .C (clk), .D (signal_8293), .Q (signal_8294) ) ;
    buf_clk cell_6452 ( .C (clk), .D (signal_8301), .Q (signal_8302) ) ;
    buf_clk cell_6460 ( .C (clk), .D (signal_8309), .Q (signal_8310) ) ;
    buf_clk cell_6468 ( .C (clk), .D (signal_8317), .Q (signal_8318) ) ;
    buf_clk cell_6476 ( .C (clk), .D (signal_8325), .Q (signal_8326) ) ;
    buf_clk cell_6484 ( .C (clk), .D (signal_8333), .Q (signal_8334) ) ;
    buf_clk cell_6492 ( .C (clk), .D (signal_8341), .Q (signal_8342) ) ;
    buf_clk cell_6500 ( .C (clk), .D (signal_8349), .Q (signal_8350) ) ;
    buf_clk cell_6508 ( .C (clk), .D (signal_8357), .Q (signal_8358) ) ;
    buf_clk cell_6516 ( .C (clk), .D (signal_8365), .Q (signal_8366) ) ;
    buf_clk cell_6524 ( .C (clk), .D (signal_8373), .Q (signal_8374) ) ;
    buf_clk cell_6532 ( .C (clk), .D (signal_8381), .Q (signal_8382) ) ;
    buf_clk cell_6540 ( .C (clk), .D (signal_8389), .Q (signal_8390) ) ;
    buf_clk cell_6548 ( .C (clk), .D (signal_8397), .Q (signal_8398) ) ;
    buf_clk cell_6556 ( .C (clk), .D (signal_8405), .Q (signal_8406) ) ;
    buf_clk cell_6564 ( .C (clk), .D (signal_8413), .Q (signal_8414) ) ;
    buf_clk cell_6572 ( .C (clk), .D (signal_8421), .Q (signal_8422) ) ;
    buf_clk cell_6580 ( .C (clk), .D (signal_8429), .Q (signal_8430) ) ;
    buf_clk cell_6588 ( .C (clk), .D (signal_8437), .Q (signal_8438) ) ;
    buf_clk cell_6596 ( .C (clk), .D (signal_8445), .Q (signal_8446) ) ;
    buf_clk cell_6604 ( .C (clk), .D (signal_8453), .Q (signal_8454) ) ;
    buf_clk cell_6612 ( .C (clk), .D (signal_8461), .Q (signal_8462) ) ;
    buf_clk cell_6620 ( .C (clk), .D (signal_8469), .Q (signal_8470) ) ;
    buf_clk cell_6628 ( .C (clk), .D (signal_8477), .Q (signal_8478) ) ;
    buf_clk cell_6636 ( .C (clk), .D (signal_8485), .Q (signal_8486) ) ;
    buf_clk cell_6644 ( .C (clk), .D (signal_8493), .Q (signal_8494) ) ;
    buf_clk cell_6652 ( .C (clk), .D (signal_8501), .Q (signal_8502) ) ;
    buf_clk cell_6660 ( .C (clk), .D (signal_8509), .Q (signal_8510) ) ;
    buf_clk cell_6668 ( .C (clk), .D (signal_8517), .Q (signal_8518) ) ;
    buf_clk cell_6676 ( .C (clk), .D (signal_8525), .Q (signal_8526) ) ;
    buf_clk cell_6684 ( .C (clk), .D (signal_8533), .Q (signal_8534) ) ;
    buf_clk cell_6692 ( .C (clk), .D (signal_8541), .Q (signal_8542) ) ;
    buf_clk cell_6700 ( .C (clk), .D (signal_8549), .Q (signal_8550) ) ;
    buf_clk cell_6708 ( .C (clk), .D (signal_8557), .Q (signal_8558) ) ;
    buf_clk cell_6716 ( .C (clk), .D (signal_8565), .Q (signal_8566) ) ;
    buf_clk cell_6724 ( .C (clk), .D (signal_8573), .Q (signal_8574) ) ;
    buf_clk cell_6732 ( .C (clk), .D (signal_8581), .Q (signal_8582) ) ;
    buf_clk cell_6740 ( .C (clk), .D (signal_8589), .Q (signal_8590) ) ;
    buf_clk cell_6748 ( .C (clk), .D (signal_8597), .Q (signal_8598) ) ;
    buf_clk cell_6756 ( .C (clk), .D (signal_8605), .Q (signal_8606) ) ;
    buf_clk cell_6764 ( .C (clk), .D (signal_8613), .Q (signal_8614) ) ;
    buf_clk cell_6772 ( .C (clk), .D (signal_8621), .Q (signal_8622) ) ;
    buf_clk cell_6780 ( .C (clk), .D (signal_8629), .Q (signal_8630) ) ;
    buf_clk cell_6788 ( .C (clk), .D (signal_8637), .Q (signal_8638) ) ;
    buf_clk cell_6796 ( .C (clk), .D (signal_8645), .Q (signal_8646) ) ;
    buf_clk cell_6804 ( .C (clk), .D (signal_8653), .Q (signal_8654) ) ;
    buf_clk cell_6812 ( .C (clk), .D (signal_8661), .Q (signal_8662) ) ;
    buf_clk cell_6820 ( .C (clk), .D (signal_8669), .Q (signal_8670) ) ;
    buf_clk cell_6828 ( .C (clk), .D (signal_8677), .Q (signal_8678) ) ;
    buf_clk cell_6836 ( .C (clk), .D (signal_8685), .Q (signal_8686) ) ;
    buf_clk cell_6844 ( .C (clk), .D (signal_8693), .Q (signal_8694) ) ;
    buf_clk cell_6852 ( .C (clk), .D (signal_8701), .Q (signal_8702) ) ;
    buf_clk cell_6860 ( .C (clk), .D (signal_8709), .Q (signal_8710) ) ;
    buf_clk cell_6868 ( .C (clk), .D (signal_8717), .Q (signal_8718) ) ;
    buf_clk cell_6876 ( .C (clk), .D (signal_8725), .Q (signal_8726) ) ;
    buf_clk cell_6884 ( .C (clk), .D (signal_8733), .Q (signal_8734) ) ;
    buf_clk cell_6892 ( .C (clk), .D (signal_8741), .Q (signal_8742) ) ;
    buf_clk cell_6900 ( .C (clk), .D (signal_8749), .Q (signal_8750) ) ;
    buf_clk cell_6908 ( .C (clk), .D (signal_8757), .Q (signal_8758) ) ;
    buf_clk cell_6916 ( .C (clk), .D (signal_8765), .Q (signal_8766) ) ;
    buf_clk cell_6924 ( .C (clk), .D (signal_8773), .Q (signal_8774) ) ;
    buf_clk cell_6932 ( .C (clk), .D (signal_8781), .Q (signal_8782) ) ;
    buf_clk cell_6940 ( .C (clk), .D (signal_8789), .Q (signal_8790) ) ;
    buf_clk cell_6948 ( .C (clk), .D (signal_8797), .Q (signal_8798) ) ;
    buf_clk cell_6956 ( .C (clk), .D (signal_8805), .Q (signal_8806) ) ;
    buf_clk cell_6964 ( .C (clk), .D (signal_8813), .Q (signal_8814) ) ;
    buf_clk cell_6972 ( .C (clk), .D (signal_8821), .Q (signal_8822) ) ;
    buf_clk cell_6980 ( .C (clk), .D (signal_8829), .Q (signal_8830) ) ;
    buf_clk cell_6988 ( .C (clk), .D (signal_8837), .Q (signal_8838) ) ;
    buf_clk cell_6996 ( .C (clk), .D (signal_8845), .Q (signal_8846) ) ;
    buf_clk cell_7004 ( .C (clk), .D (signal_8853), .Q (signal_8854) ) ;
    buf_clk cell_7012 ( .C (clk), .D (signal_8861), .Q (signal_8862) ) ;
    buf_clk cell_7020 ( .C (clk), .D (signal_8869), .Q (signal_8870) ) ;
    buf_clk cell_7028 ( .C (clk), .D (signal_8877), .Q (signal_8878) ) ;
    buf_clk cell_7036 ( .C (clk), .D (signal_8885), .Q (signal_8886) ) ;
    buf_clk cell_7044 ( .C (clk), .D (signal_8893), .Q (signal_8894) ) ;
    buf_clk cell_7052 ( .C (clk), .D (signal_8901), .Q (signal_8902) ) ;
    buf_clk cell_7060 ( .C (clk), .D (signal_8909), .Q (signal_8910) ) ;
    buf_clk cell_7068 ( .C (clk), .D (signal_8917), .Q (signal_8918) ) ;
    buf_clk cell_7076 ( .C (clk), .D (signal_8925), .Q (signal_8926) ) ;
    buf_clk cell_7084 ( .C (clk), .D (signal_8933), .Q (signal_8934) ) ;
    buf_clk cell_7092 ( .C (clk), .D (signal_8941), .Q (signal_8942) ) ;
    buf_clk cell_7100 ( .C (clk), .D (signal_8949), .Q (signal_8950) ) ;

    /* cells in depth 8 */
    mux2_masked #(.security_order(1), .pipeline(1)) cell_56 ( .s (signal_3751), .b ({signal_3579, signal_1405}), .a ({signal_3767, signal_3759}), .c ({signal_3587, signal_1421}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_57 ( .s (signal_3751), .b ({signal_3599, signal_1404}), .a ({signal_3783, signal_3775}), .c ({signal_3600, signal_1420}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_58 ( .s (signal_3751), .b ({signal_3585, signal_1403}), .a ({signal_3799, signal_3791}), .c ({signal_3588, signal_1419}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_59 ( .s (signal_3751), .b ({signal_3584, signal_1402}), .a ({signal_3815, signal_3807}), .c ({signal_3589, signal_1418}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_60 ( .s (signal_3751), .b ({signal_3583, signal_1401}), .a ({signal_3831, signal_3823}), .c ({signal_3590, signal_1417}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_61 ( .s (signal_3751), .b ({signal_3598, signal_1400}), .a ({signal_3847, signal_3839}), .c ({signal_3601, signal_1416}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_62 ( .s (signal_3751), .b ({signal_3597, signal_1399}), .a ({signal_3863, signal_3855}), .c ({signal_3602, signal_1415}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_63 ( .s (signal_3751), .b ({signal_3580, signal_1398}), .a ({signal_3879, signal_3871}), .c ({signal_3591, signal_1414}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_445 ( .s (signal_3887), .b ({signal_3620, signal_1557}), .a ({signal_3903, signal_3895}), .c ({signal_3637, signal_705}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_448 ( .s (signal_3887), .b ({signal_3643, signal_1556}), .a ({signal_3919, signal_3911}), .c ({signal_3656, signal_707}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_451 ( .s (signal_3887), .b ({signal_3622, signal_1555}), .a ({signal_3935, signal_3927}), .c ({signal_3638, signal_709}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_454 ( .s (signal_3887), .b ({signal_3624, signal_1554}), .a ({signal_3951, signal_3943}), .c ({signal_3639, signal_711}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_457 ( .s (signal_3887), .b ({signal_3626, signal_1553}), .a ({signal_3967, signal_3959}), .c ({signal_3640, signal_713}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_460 ( .s (signal_3887), .b ({signal_3645, signal_1552}), .a ({signal_3983, signal_3975}), .c ({signal_3657, signal_715}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_463 ( .s (signal_3887), .b ({signal_3647, signal_1551}), .a ({signal_3999, signal_3991}), .c ({signal_3658, signal_717}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_466 ( .s (signal_3887), .b ({signal_3628, signal_1550}), .a ({signal_4015, signal_4007}), .c ({signal_3641, signal_719}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_613 ( .s (signal_4023), .b ({signal_3587, signal_1421}), .a ({signal_4039, signal_4031}), .c ({signal_3603, signal_1525}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_614 ( .s (signal_4023), .b ({signal_3600, signal_1420}), .a ({signal_4055, signal_4047}), .c ({signal_3616, signal_1524}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_615 ( .s (signal_4023), .b ({signal_3588, signal_1419}), .a ({signal_4071, signal_4063}), .c ({signal_3604, signal_1523}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_616 ( .s (signal_4023), .b ({signal_3589, signal_1418}), .a ({signal_4087, signal_4079}), .c ({signal_3605, signal_1522}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_617 ( .s (signal_4023), .b ({signal_3590, signal_1417}), .a ({signal_4103, signal_4095}), .c ({signal_3606, signal_1521}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_618 ( .s (signal_4023), .b ({signal_3601, signal_1416}), .a ({signal_4119, signal_4111}), .c ({signal_3617, signal_1520}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_619 ( .s (signal_4023), .b ({signal_3602, signal_1415}), .a ({signal_4135, signal_4127}), .c ({signal_3618, signal_1519}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_620 ( .s (signal_4023), .b ({signal_3591, signal_1414}), .a ({signal_4151, signal_4143}), .c ({signal_3607, signal_1518}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_621 ( .s (signal_4159), .b ({signal_4175, signal_4167}), .a ({signal_3603, signal_1525}), .c ({signal_3620, signal_1557}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_622 ( .s (signal_4159), .b ({signal_4191, signal_4183}), .a ({signal_3616, signal_1524}), .c ({signal_3643, signal_1556}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_623 ( .s (signal_4159), .b ({signal_4207, signal_4199}), .a ({signal_3604, signal_1523}), .c ({signal_3622, signal_1555}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_624 ( .s (signal_4159), .b ({signal_4223, signal_4215}), .a ({signal_3605, signal_1522}), .c ({signal_3624, signal_1554}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_625 ( .s (signal_4159), .b ({signal_4239, signal_4231}), .a ({signal_3606, signal_1521}), .c ({signal_3626, signal_1553}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_626 ( .s (signal_4159), .b ({signal_4255, signal_4247}), .a ({signal_3617, signal_1520}), .c ({signal_3645, signal_1552}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_627 ( .s (signal_4159), .b ({signal_4271, signal_4263}), .a ({signal_3618, signal_1519}), .c ({signal_3647, signal_1551}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_628 ( .s (signal_4159), .b ({signal_4287, signal_4279}), .a ({signal_3607, signal_1518}), .c ({signal_3628, signal_1550}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_672 ( .a ({signal_3592, signal_724}), .b ({signal_4303, signal_4295}), .c ({signal_3608, signal_1750}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_673 ( .a ({1'b0, signal_4311}), .b ({signal_3580, signal_1398}), .c ({signal_3592, signal_724}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_674 ( .a ({signal_3609, signal_725}), .b ({signal_4327, signal_4319}), .c ({signal_3629, signal_1751}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_675 ( .a ({1'b0, signal_4335}), .b ({signal_3597, signal_1399}), .c ({signal_3609, signal_725}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_676 ( .a ({signal_3610, signal_726}), .b ({signal_4351, signal_4343}), .c ({signal_3630, signal_1752}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_677 ( .a ({1'b0, signal_4359}), .b ({signal_3598, signal_1400}), .c ({signal_3610, signal_726}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_678 ( .a ({signal_3593, signal_727}), .b ({signal_4375, signal_4367}), .c ({signal_3611, signal_1753}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_679 ( .a ({1'b0, signal_4383}), .b ({signal_3583, signal_1401}), .c ({signal_3593, signal_727}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_680 ( .a ({signal_3594, signal_728}), .b ({signal_4399, signal_4391}), .c ({signal_3612, signal_1754}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_681 ( .a ({1'b0, signal_4407}), .b ({signal_3584, signal_1402}), .c ({signal_3594, signal_728}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_682 ( .a ({signal_3595, signal_729}), .b ({signal_4423, signal_4415}), .c ({signal_3613, signal_1755}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_683 ( .a ({1'b0, signal_4431}), .b ({signal_3585, signal_1403}), .c ({signal_3595, signal_729}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_684 ( .a ({signal_3614, signal_730}), .b ({signal_4447, signal_4439}), .c ({signal_3631, signal_1756}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_685 ( .a ({1'b0, signal_4455}), .b ({signal_3599, signal_1404}), .c ({signal_3614, signal_730}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_686 ( .a ({signal_3596, signal_731}), .b ({signal_4471, signal_4463}), .c ({signal_3615, signal_1757}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_687 ( .a ({1'b0, signal_4479}), .b ({signal_3579, signal_1405}), .c ({signal_3596, signal_731}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1098 ( .s (signal_4487), .b ({signal_4503, signal_4495}), .a ({signal_3632, signal_1055}), .c ({signal_3648, signal_1054}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1099 ( .s (signal_4511), .b ({signal_4527, signal_4519}), .a ({signal_3615, signal_1757}), .c ({signal_3632, signal_1055}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1102 ( .s (signal_4487), .b ({signal_4543, signal_4535}), .a ({signal_3649, signal_1058}), .c ({signal_3659, signal_1057}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1103 ( .s (signal_4511), .b ({signal_4559, signal_4551}), .a ({signal_3631, signal_1756}), .c ({signal_3649, signal_1058}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1106 ( .s (signal_4487), .b ({signal_4575, signal_4567}), .a ({signal_3633, signal_1061}), .c ({signal_3650, signal_1060}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1107 ( .s (signal_4511), .b ({signal_4591, signal_4583}), .a ({signal_3613, signal_1755}), .c ({signal_3633, signal_1061}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1110 ( .s (signal_4487), .b ({signal_4607, signal_4599}), .a ({signal_3634, signal_1064}), .c ({signal_3651, signal_1063}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1111 ( .s (signal_4511), .b ({signal_4623, signal_4615}), .a ({signal_3612, signal_1754}), .c ({signal_3634, signal_1064}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1114 ( .s (signal_4487), .b ({signal_4639, signal_4631}), .a ({signal_3635, signal_1067}), .c ({signal_3652, signal_1066}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1115 ( .s (signal_4511), .b ({signal_4655, signal_4647}), .a ({signal_3611, signal_1753}), .c ({signal_3635, signal_1067}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1118 ( .s (signal_4487), .b ({signal_4671, signal_4663}), .a ({signal_3653, signal_1070}), .c ({signal_3660, signal_1069}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1119 ( .s (signal_4511), .b ({signal_4687, signal_4679}), .a ({signal_3630, signal_1752}), .c ({signal_3653, signal_1070}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1122 ( .s (signal_4487), .b ({signal_4703, signal_4695}), .a ({signal_3654, signal_1073}), .c ({signal_3661, signal_1072}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1123 ( .s (signal_4511), .b ({signal_4719, signal_4711}), .a ({signal_3629, signal_1751}), .c ({signal_3654, signal_1073}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1126 ( .s (signal_4487), .b ({signal_4735, signal_4727}), .a ({signal_3636, signal_1076}), .c ({signal_3655, signal_1075}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1127 ( .s (signal_4511), .b ({signal_4751, signal_4743}), .a ({signal_3608, signal_1750}), .c ({signal_3636, signal_1076}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1781 ( .a ({signal_4763, signal_4757}), .b ({signal_3524, signal_2048}), .clk (clk), .r (Fresh[16]), .c ({signal_3525, signal_2049}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1782 ( .a ({signal_4775, signal_4769}), .b ({signal_3523, signal_2047}), .clk (clk), .r (Fresh[17]), .c ({signal_3526, signal_2050}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1783 ( .a ({signal_4787, signal_4781}), .b ({signal_3522, signal_2046}), .clk (clk), .r (Fresh[18]), .c ({signal_3527, signal_2051}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1784 ( .a ({signal_4799, signal_4793}), .b ({signal_3521, signal_2045}), .clk (clk), .r (Fresh[19]), .c ({signal_3528, signal_2052}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1785 ( .a ({signal_4811, signal_4805}), .b ({signal_3524, signal_2048}), .clk (clk), .r (Fresh[20]), .c ({signal_3529, signal_2053}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1786 ( .a ({signal_4823, signal_4817}), .b ({signal_3523, signal_2047}), .clk (clk), .r (Fresh[21]), .c ({signal_3530, signal_2054}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1787 ( .a ({signal_4835, signal_4829}), .b ({signal_3522, signal_2046}), .clk (clk), .r (Fresh[22]), .c ({signal_3531, signal_2055}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1788 ( .a ({signal_4847, signal_4841}), .b ({signal_3521, signal_2045}), .clk (clk), .r (Fresh[23]), .c ({signal_3532, signal_2056}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1793 ( .a ({signal_4859, signal_4853}), .b ({signal_3536, signal_2060}), .clk (clk), .r (Fresh[24]), .c ({signal_3537, signal_2061}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1794 ( .a ({signal_4871, signal_4865}), .b ({signal_3535, signal_2059}), .clk (clk), .r (Fresh[25]), .c ({signal_3538, signal_2062}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1795 ( .a ({signal_4883, signal_4877}), .b ({signal_3534, signal_2058}), .clk (clk), .r (Fresh[26]), .c ({signal_3539, signal_2063}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1796 ( .a ({signal_4895, signal_4889}), .b ({signal_3533, signal_2057}), .clk (clk), .r (Fresh[27]), .c ({signal_3540, signal_2064}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1797 ( .a ({signal_4907, signal_4901}), .b ({signal_3536, signal_2060}), .clk (clk), .r (Fresh[28]), .c ({signal_3541, signal_2065}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1798 ( .a ({signal_4919, signal_4913}), .b ({signal_3535, signal_2059}), .clk (clk), .r (Fresh[29]), .c ({signal_3542, signal_2066}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1799 ( .a ({signal_4931, signal_4925}), .b ({signal_3534, signal_2058}), .clk (clk), .r (Fresh[30]), .c ({signal_3543, signal_2067}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1800 ( .a ({signal_4943, signal_4937}), .b ({signal_3533, signal_2057}), .clk (clk), .r (Fresh[31]), .c ({signal_3544, signal_2068}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1802 ( .a ({signal_3527, signal_2051}), .b ({signal_3529, signal_2053}), .c ({signal_3546, signal_2070}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1803 ( .a ({signal_3528, signal_2052}), .b ({signal_3531, signal_2055}), .c ({signal_3547, signal_2071}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1804 ( .a ({signal_3526, signal_2050}), .b ({signal_3528, signal_2052}), .c ({signal_3548, signal_2072}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1805 ( .a ({signal_4955, signal_4949}), .b ({signal_3545, signal_2069}), .clk (clk), .r (Fresh[32]), .c ({signal_3549, signal_2073}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1806 ( .a ({signal_4967, signal_4961}), .b ({signal_3545, signal_2069}), .clk (clk), .r (Fresh[33]), .c ({signal_3550, signal_2074}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1807 ( .a ({signal_3526, signal_2050}), .b ({signal_3537, signal_2061}), .c ({signal_3551, signal_2075}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1808 ( .a ({signal_3525, signal_2049}), .b ({signal_3541, signal_2065}), .c ({signal_3552, signal_2076}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1809 ( .a ({signal_3540, signal_2064}), .b ({signal_3542, signal_2066}), .c ({signal_3553, signal_2077}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1810 ( .a ({signal_3538, signal_2062}), .b ({signal_3543, signal_2067}), .c ({signal_3554, signal_2078}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1811 ( .a ({signal_3539, signal_2063}), .b ({signal_3543, signal_2067}), .c ({signal_3555, signal_2079}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1812 ( .a ({signal_3541, signal_2065}), .b ({signal_3546, signal_2070}), .c ({signal_3556, signal_2080}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1813 ( .a ({signal_3530, signal_2054}), .b ({signal_3546, signal_2070}), .c ({signal_3557, signal_2081}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1814 ( .a ({signal_3542, signal_2066}), .b ({signal_3547, signal_2071}), .c ({signal_3558, signal_2082}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1815 ( .a ({signal_3543, signal_2067}), .b ({signal_3550, signal_2074}), .c ({signal_3559, signal_2083}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1816 ( .a ({signal_3550, signal_2074}), .b ({signal_3554, signal_2078}), .c ({signal_3560, signal_2084}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1817 ( .a ({signal_3537, signal_2061}), .b ({signal_3552, signal_2076}), .c ({signal_3561, signal_2085}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1818 ( .a ({signal_3539, signal_2063}), .b ({signal_3549, signal_2073}), .c ({signal_3562, signal_2086}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1819 ( .a ({signal_3549, signal_2073}), .b ({signal_3553, signal_2077}), .c ({signal_3563, signal_2087}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1820 ( .a ({signal_3532, signal_2056}), .b ({signal_3551, signal_2075}), .c ({signal_3564, signal_2088}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1821 ( .a ({signal_3544, signal_2068}), .b ({signal_3553, signal_2077}), .c ({signal_3565, signal_2089}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1822 ( .a ({signal_3548, signal_2072}), .b ({signal_3552, signal_2076}), .c ({signal_3566, signal_2090}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1823 ( .a ({signal_3551, signal_2075}), .b ({signal_3558, signal_2082}), .c ({signal_3567, signal_2091}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1824 ( .a ({signal_3527, signal_2051}), .b ({signal_3559, signal_2083}), .c ({signal_3568, signal_2092}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1825 ( .a ({signal_3529, signal_2053}), .b ({signal_3559, signal_2083}), .c ({signal_3569, signal_2093}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1826 ( .a ({signal_3546, signal_2070}), .b ({signal_3559, signal_2083}), .c ({signal_3570, signal_2094}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1827 ( .a ({signal_3546, signal_2070}), .b ({signal_3561, signal_2085}), .c ({signal_3571, signal_2095}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1828 ( .a ({signal_3556, signal_2080}), .b ({signal_3562, signal_2086}), .c ({signal_3572, signal_2096}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1829 ( .a ({signal_3560, signal_2084}), .b ({signal_3563, signal_2087}), .c ({signal_3573, signal_2097}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1830 ( .a ({signal_3561, signal_2085}), .b ({signal_3562, signal_2086}), .c ({signal_3574, signal_2098}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1831 ( .a ({signal_3547, signal_2071}), .b ({signal_3563, signal_2087}), .c ({signal_3575, signal_2099}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1832 ( .a ({signal_3555, signal_2079}), .b ({signal_3564, signal_2088}), .c ({signal_3576, signal_2100}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1833 ( .a ({signal_3557, signal_2081}), .b ({signal_3564, signal_2088}), .c ({signal_3577, signal_2101}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1834 ( .a ({signal_3560, signal_2084}), .b ({signal_3567, signal_2091}), .c ({signal_3578, signal_2102}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1835 ( .a ({signal_3578, signal_2102}), .b ({signal_3579, signal_1405}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1836 ( .a ({signal_3560, signal_2084}), .b ({signal_3572, signal_2096}), .c ({signal_3580, signal_1398}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1837 ( .a ({signal_3569, signal_2093}), .b ({signal_3574, signal_2098}), .c ({signal_3581, signal_2103}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1838 ( .a ({signal_3565, signal_2089}), .b ({signal_3576, signal_2100}), .c ({signal_3582, signal_2104}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1839 ( .a ({signal_3560, signal_2084}), .b ({signal_3571, signal_2095}), .c ({signal_3583, signal_1401}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1840 ( .a ({signal_3566, signal_2090}), .b ({signal_3570, signal_2094}), .c ({signal_3584, signal_1402}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1841 ( .a ({signal_3573, signal_2097}), .b ({signal_3577, signal_2101}), .c ({signal_3585, signal_1403}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1842 ( .a ({signal_3568, signal_2092}), .b ({signal_3575, signal_2099}), .c ({signal_3586, signal_2105}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1843 ( .a ({signal_3581, signal_2103}), .b ({signal_3597, signal_1399}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1844 ( .a ({signal_3582, signal_2104}), .b ({signal_3598, signal_1400}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1845 ( .a ({signal_3586, signal_2105}), .b ({signal_3599, signal_1404}) ) ;
    buf_clk cell_1901 ( .C (clk), .D (signal_3750), .Q (signal_3751) ) ;
    buf_clk cell_1909 ( .C (clk), .D (signal_3758), .Q (signal_3759) ) ;
    buf_clk cell_1917 ( .C (clk), .D (signal_3766), .Q (signal_3767) ) ;
    buf_clk cell_1925 ( .C (clk), .D (signal_3774), .Q (signal_3775) ) ;
    buf_clk cell_1933 ( .C (clk), .D (signal_3782), .Q (signal_3783) ) ;
    buf_clk cell_1941 ( .C (clk), .D (signal_3790), .Q (signal_3791) ) ;
    buf_clk cell_1949 ( .C (clk), .D (signal_3798), .Q (signal_3799) ) ;
    buf_clk cell_1957 ( .C (clk), .D (signal_3806), .Q (signal_3807) ) ;
    buf_clk cell_1965 ( .C (clk), .D (signal_3814), .Q (signal_3815) ) ;
    buf_clk cell_1973 ( .C (clk), .D (signal_3822), .Q (signal_3823) ) ;
    buf_clk cell_1981 ( .C (clk), .D (signal_3830), .Q (signal_3831) ) ;
    buf_clk cell_1989 ( .C (clk), .D (signal_3838), .Q (signal_3839) ) ;
    buf_clk cell_1997 ( .C (clk), .D (signal_3846), .Q (signal_3847) ) ;
    buf_clk cell_2005 ( .C (clk), .D (signal_3854), .Q (signal_3855) ) ;
    buf_clk cell_2013 ( .C (clk), .D (signal_3862), .Q (signal_3863) ) ;
    buf_clk cell_2021 ( .C (clk), .D (signal_3870), .Q (signal_3871) ) ;
    buf_clk cell_2029 ( .C (clk), .D (signal_3878), .Q (signal_3879) ) ;
    buf_clk cell_2037 ( .C (clk), .D (signal_3886), .Q (signal_3887) ) ;
    buf_clk cell_2045 ( .C (clk), .D (signal_3894), .Q (signal_3895) ) ;
    buf_clk cell_2053 ( .C (clk), .D (signal_3902), .Q (signal_3903) ) ;
    buf_clk cell_2061 ( .C (clk), .D (signal_3910), .Q (signal_3911) ) ;
    buf_clk cell_2069 ( .C (clk), .D (signal_3918), .Q (signal_3919) ) ;
    buf_clk cell_2077 ( .C (clk), .D (signal_3926), .Q (signal_3927) ) ;
    buf_clk cell_2085 ( .C (clk), .D (signal_3934), .Q (signal_3935) ) ;
    buf_clk cell_2093 ( .C (clk), .D (signal_3942), .Q (signal_3943) ) ;
    buf_clk cell_2101 ( .C (clk), .D (signal_3950), .Q (signal_3951) ) ;
    buf_clk cell_2109 ( .C (clk), .D (signal_3958), .Q (signal_3959) ) ;
    buf_clk cell_2117 ( .C (clk), .D (signal_3966), .Q (signal_3967) ) ;
    buf_clk cell_2125 ( .C (clk), .D (signal_3974), .Q (signal_3975) ) ;
    buf_clk cell_2133 ( .C (clk), .D (signal_3982), .Q (signal_3983) ) ;
    buf_clk cell_2141 ( .C (clk), .D (signal_3990), .Q (signal_3991) ) ;
    buf_clk cell_2149 ( .C (clk), .D (signal_3998), .Q (signal_3999) ) ;
    buf_clk cell_2157 ( .C (clk), .D (signal_4006), .Q (signal_4007) ) ;
    buf_clk cell_2165 ( .C (clk), .D (signal_4014), .Q (signal_4015) ) ;
    buf_clk cell_2173 ( .C (clk), .D (signal_4022), .Q (signal_4023) ) ;
    buf_clk cell_2181 ( .C (clk), .D (signal_4030), .Q (signal_4031) ) ;
    buf_clk cell_2189 ( .C (clk), .D (signal_4038), .Q (signal_4039) ) ;
    buf_clk cell_2197 ( .C (clk), .D (signal_4046), .Q (signal_4047) ) ;
    buf_clk cell_2205 ( .C (clk), .D (signal_4054), .Q (signal_4055) ) ;
    buf_clk cell_2213 ( .C (clk), .D (signal_4062), .Q (signal_4063) ) ;
    buf_clk cell_2221 ( .C (clk), .D (signal_4070), .Q (signal_4071) ) ;
    buf_clk cell_2229 ( .C (clk), .D (signal_4078), .Q (signal_4079) ) ;
    buf_clk cell_2237 ( .C (clk), .D (signal_4086), .Q (signal_4087) ) ;
    buf_clk cell_2245 ( .C (clk), .D (signal_4094), .Q (signal_4095) ) ;
    buf_clk cell_2253 ( .C (clk), .D (signal_4102), .Q (signal_4103) ) ;
    buf_clk cell_2261 ( .C (clk), .D (signal_4110), .Q (signal_4111) ) ;
    buf_clk cell_2269 ( .C (clk), .D (signal_4118), .Q (signal_4119) ) ;
    buf_clk cell_2277 ( .C (clk), .D (signal_4126), .Q (signal_4127) ) ;
    buf_clk cell_2285 ( .C (clk), .D (signal_4134), .Q (signal_4135) ) ;
    buf_clk cell_2293 ( .C (clk), .D (signal_4142), .Q (signal_4143) ) ;
    buf_clk cell_2301 ( .C (clk), .D (signal_4150), .Q (signal_4151) ) ;
    buf_clk cell_2309 ( .C (clk), .D (signal_4158), .Q (signal_4159) ) ;
    buf_clk cell_2317 ( .C (clk), .D (signal_4166), .Q (signal_4167) ) ;
    buf_clk cell_2325 ( .C (clk), .D (signal_4174), .Q (signal_4175) ) ;
    buf_clk cell_2333 ( .C (clk), .D (signal_4182), .Q (signal_4183) ) ;
    buf_clk cell_2341 ( .C (clk), .D (signal_4190), .Q (signal_4191) ) ;
    buf_clk cell_2349 ( .C (clk), .D (signal_4198), .Q (signal_4199) ) ;
    buf_clk cell_2357 ( .C (clk), .D (signal_4206), .Q (signal_4207) ) ;
    buf_clk cell_2365 ( .C (clk), .D (signal_4214), .Q (signal_4215) ) ;
    buf_clk cell_2373 ( .C (clk), .D (signal_4222), .Q (signal_4223) ) ;
    buf_clk cell_2381 ( .C (clk), .D (signal_4230), .Q (signal_4231) ) ;
    buf_clk cell_2389 ( .C (clk), .D (signal_4238), .Q (signal_4239) ) ;
    buf_clk cell_2397 ( .C (clk), .D (signal_4246), .Q (signal_4247) ) ;
    buf_clk cell_2405 ( .C (clk), .D (signal_4254), .Q (signal_4255) ) ;
    buf_clk cell_2413 ( .C (clk), .D (signal_4262), .Q (signal_4263) ) ;
    buf_clk cell_2421 ( .C (clk), .D (signal_4270), .Q (signal_4271) ) ;
    buf_clk cell_2429 ( .C (clk), .D (signal_4278), .Q (signal_4279) ) ;
    buf_clk cell_2437 ( .C (clk), .D (signal_4286), .Q (signal_4287) ) ;
    buf_clk cell_2445 ( .C (clk), .D (signal_4294), .Q (signal_4295) ) ;
    buf_clk cell_2453 ( .C (clk), .D (signal_4302), .Q (signal_4303) ) ;
    buf_clk cell_2461 ( .C (clk), .D (signal_4310), .Q (signal_4311) ) ;
    buf_clk cell_2469 ( .C (clk), .D (signal_4318), .Q (signal_4319) ) ;
    buf_clk cell_2477 ( .C (clk), .D (signal_4326), .Q (signal_4327) ) ;
    buf_clk cell_2485 ( .C (clk), .D (signal_4334), .Q (signal_4335) ) ;
    buf_clk cell_2493 ( .C (clk), .D (signal_4342), .Q (signal_4343) ) ;
    buf_clk cell_2501 ( .C (clk), .D (signal_4350), .Q (signal_4351) ) ;
    buf_clk cell_2509 ( .C (clk), .D (signal_4358), .Q (signal_4359) ) ;
    buf_clk cell_2517 ( .C (clk), .D (signal_4366), .Q (signal_4367) ) ;
    buf_clk cell_2525 ( .C (clk), .D (signal_4374), .Q (signal_4375) ) ;
    buf_clk cell_2533 ( .C (clk), .D (signal_4382), .Q (signal_4383) ) ;
    buf_clk cell_2541 ( .C (clk), .D (signal_4390), .Q (signal_4391) ) ;
    buf_clk cell_2549 ( .C (clk), .D (signal_4398), .Q (signal_4399) ) ;
    buf_clk cell_2557 ( .C (clk), .D (signal_4406), .Q (signal_4407) ) ;
    buf_clk cell_2565 ( .C (clk), .D (signal_4414), .Q (signal_4415) ) ;
    buf_clk cell_2573 ( .C (clk), .D (signal_4422), .Q (signal_4423) ) ;
    buf_clk cell_2581 ( .C (clk), .D (signal_4430), .Q (signal_4431) ) ;
    buf_clk cell_2589 ( .C (clk), .D (signal_4438), .Q (signal_4439) ) ;
    buf_clk cell_2597 ( .C (clk), .D (signal_4446), .Q (signal_4447) ) ;
    buf_clk cell_2605 ( .C (clk), .D (signal_4454), .Q (signal_4455) ) ;
    buf_clk cell_2613 ( .C (clk), .D (signal_4462), .Q (signal_4463) ) ;
    buf_clk cell_2621 ( .C (clk), .D (signal_4470), .Q (signal_4471) ) ;
    buf_clk cell_2629 ( .C (clk), .D (signal_4478), .Q (signal_4479) ) ;
    buf_clk cell_2637 ( .C (clk), .D (signal_4486), .Q (signal_4487) ) ;
    buf_clk cell_2645 ( .C (clk), .D (signal_4494), .Q (signal_4495) ) ;
    buf_clk cell_2653 ( .C (clk), .D (signal_4502), .Q (signal_4503) ) ;
    buf_clk cell_2661 ( .C (clk), .D (signal_4510), .Q (signal_4511) ) ;
    buf_clk cell_2669 ( .C (clk), .D (signal_4518), .Q (signal_4519) ) ;
    buf_clk cell_2677 ( .C (clk), .D (signal_4526), .Q (signal_4527) ) ;
    buf_clk cell_2685 ( .C (clk), .D (signal_4534), .Q (signal_4535) ) ;
    buf_clk cell_2693 ( .C (clk), .D (signal_4542), .Q (signal_4543) ) ;
    buf_clk cell_2701 ( .C (clk), .D (signal_4550), .Q (signal_4551) ) ;
    buf_clk cell_2709 ( .C (clk), .D (signal_4558), .Q (signal_4559) ) ;
    buf_clk cell_2717 ( .C (clk), .D (signal_4566), .Q (signal_4567) ) ;
    buf_clk cell_2725 ( .C (clk), .D (signal_4574), .Q (signal_4575) ) ;
    buf_clk cell_2733 ( .C (clk), .D (signal_4582), .Q (signal_4583) ) ;
    buf_clk cell_2741 ( .C (clk), .D (signal_4590), .Q (signal_4591) ) ;
    buf_clk cell_2749 ( .C (clk), .D (signal_4598), .Q (signal_4599) ) ;
    buf_clk cell_2757 ( .C (clk), .D (signal_4606), .Q (signal_4607) ) ;
    buf_clk cell_2765 ( .C (clk), .D (signal_4614), .Q (signal_4615) ) ;
    buf_clk cell_2773 ( .C (clk), .D (signal_4622), .Q (signal_4623) ) ;
    buf_clk cell_2781 ( .C (clk), .D (signal_4630), .Q (signal_4631) ) ;
    buf_clk cell_2789 ( .C (clk), .D (signal_4638), .Q (signal_4639) ) ;
    buf_clk cell_2797 ( .C (clk), .D (signal_4646), .Q (signal_4647) ) ;
    buf_clk cell_2805 ( .C (clk), .D (signal_4654), .Q (signal_4655) ) ;
    buf_clk cell_2813 ( .C (clk), .D (signal_4662), .Q (signal_4663) ) ;
    buf_clk cell_2821 ( .C (clk), .D (signal_4670), .Q (signal_4671) ) ;
    buf_clk cell_2829 ( .C (clk), .D (signal_4678), .Q (signal_4679) ) ;
    buf_clk cell_2837 ( .C (clk), .D (signal_4686), .Q (signal_4687) ) ;
    buf_clk cell_2845 ( .C (clk), .D (signal_4694), .Q (signal_4695) ) ;
    buf_clk cell_2853 ( .C (clk), .D (signal_4702), .Q (signal_4703) ) ;
    buf_clk cell_2861 ( .C (clk), .D (signal_4710), .Q (signal_4711) ) ;
    buf_clk cell_2869 ( .C (clk), .D (signal_4718), .Q (signal_4719) ) ;
    buf_clk cell_2877 ( .C (clk), .D (signal_4726), .Q (signal_4727) ) ;
    buf_clk cell_2885 ( .C (clk), .D (signal_4734), .Q (signal_4735) ) ;
    buf_clk cell_2893 ( .C (clk), .D (signal_4742), .Q (signal_4743) ) ;
    buf_clk cell_2901 ( .C (clk), .D (signal_4750), .Q (signal_4751) ) ;
    buf_clk cell_3125 ( .C (clk), .D (signal_4974), .Q (signal_4975) ) ;
    buf_clk cell_3133 ( .C (clk), .D (signal_4982), .Q (signal_4983) ) ;
    buf_clk cell_3141 ( .C (clk), .D (signal_4990), .Q (signal_4991) ) ;
    buf_clk cell_3149 ( .C (clk), .D (signal_4998), .Q (signal_4999) ) ;
    buf_clk cell_3157 ( .C (clk), .D (signal_5006), .Q (signal_5007) ) ;
    buf_clk cell_3165 ( .C (clk), .D (signal_5014), .Q (signal_5015) ) ;
    buf_clk cell_3173 ( .C (clk), .D (signal_5022), .Q (signal_5023) ) ;
    buf_clk cell_3181 ( .C (clk), .D (signal_5030), .Q (signal_5031) ) ;
    buf_clk cell_3189 ( .C (clk), .D (signal_5038), .Q (signal_5039) ) ;
    buf_clk cell_3197 ( .C (clk), .D (signal_5046), .Q (signal_5047) ) ;
    buf_clk cell_3205 ( .C (clk), .D (signal_5054), .Q (signal_5055) ) ;
    buf_clk cell_3213 ( .C (clk), .D (signal_5062), .Q (signal_5063) ) ;
    buf_clk cell_3221 ( .C (clk), .D (signal_5070), .Q (signal_5071) ) ;
    buf_clk cell_3229 ( .C (clk), .D (signal_5078), .Q (signal_5079) ) ;
    buf_clk cell_3237 ( .C (clk), .D (signal_5086), .Q (signal_5087) ) ;
    buf_clk cell_3245 ( .C (clk), .D (signal_5094), .Q (signal_5095) ) ;
    buf_clk cell_3253 ( .C (clk), .D (signal_5102), .Q (signal_5103) ) ;
    buf_clk cell_3261 ( .C (clk), .D (signal_5110), .Q (signal_5111) ) ;
    buf_clk cell_3269 ( .C (clk), .D (signal_5118), .Q (signal_5119) ) ;
    buf_clk cell_3277 ( .C (clk), .D (signal_5126), .Q (signal_5127) ) ;
    buf_clk cell_3285 ( .C (clk), .D (signal_5134), .Q (signal_5135) ) ;
    buf_clk cell_3293 ( .C (clk), .D (signal_5142), .Q (signal_5143) ) ;
    buf_clk cell_3301 ( .C (clk), .D (signal_5150), .Q (signal_5151) ) ;
    buf_clk cell_3309 ( .C (clk), .D (signal_5158), .Q (signal_5159) ) ;
    buf_clk cell_3317 ( .C (clk), .D (signal_5166), .Q (signal_5167) ) ;
    buf_clk cell_3325 ( .C (clk), .D (signal_5174), .Q (signal_5175) ) ;
    buf_clk cell_3333 ( .C (clk), .D (signal_5182), .Q (signal_5183) ) ;
    buf_clk cell_3341 ( .C (clk), .D (signal_5190), .Q (signal_5191) ) ;
    buf_clk cell_3349 ( .C (clk), .D (signal_5198), .Q (signal_5199) ) ;
    buf_clk cell_3357 ( .C (clk), .D (signal_5206), .Q (signal_5207) ) ;
    buf_clk cell_3365 ( .C (clk), .D (signal_5214), .Q (signal_5215) ) ;
    buf_clk cell_3373 ( .C (clk), .D (signal_5222), .Q (signal_5223) ) ;
    buf_clk cell_3381 ( .C (clk), .D (signal_5230), .Q (signal_5231) ) ;
    buf_clk cell_3389 ( .C (clk), .D (signal_5238), .Q (signal_5239) ) ;
    buf_clk cell_3397 ( .C (clk), .D (signal_5246), .Q (signal_5247) ) ;
    buf_clk cell_3405 ( .C (clk), .D (signal_5254), .Q (signal_5255) ) ;
    buf_clk cell_3413 ( .C (clk), .D (signal_5262), .Q (signal_5263) ) ;
    buf_clk cell_3421 ( .C (clk), .D (signal_5270), .Q (signal_5271) ) ;
    buf_clk cell_3429 ( .C (clk), .D (signal_5278), .Q (signal_5279) ) ;
    buf_clk cell_3437 ( .C (clk), .D (signal_5286), .Q (signal_5287) ) ;
    buf_clk cell_3445 ( .C (clk), .D (signal_5294), .Q (signal_5295) ) ;
    buf_clk cell_3453 ( .C (clk), .D (signal_5302), .Q (signal_5303) ) ;
    buf_clk cell_3461 ( .C (clk), .D (signal_5310), .Q (signal_5311) ) ;
    buf_clk cell_3469 ( .C (clk), .D (signal_5318), .Q (signal_5319) ) ;
    buf_clk cell_3477 ( .C (clk), .D (signal_5326), .Q (signal_5327) ) ;
    buf_clk cell_3485 ( .C (clk), .D (signal_5334), .Q (signal_5335) ) ;
    buf_clk cell_3493 ( .C (clk), .D (signal_5342), .Q (signal_5343) ) ;
    buf_clk cell_3501 ( .C (clk), .D (signal_5350), .Q (signal_5351) ) ;
    buf_clk cell_3509 ( .C (clk), .D (signal_5358), .Q (signal_5359) ) ;
    buf_clk cell_3517 ( .C (clk), .D (signal_5366), .Q (signal_5367) ) ;
    buf_clk cell_3525 ( .C (clk), .D (signal_5374), .Q (signal_5375) ) ;
    buf_clk cell_3533 ( .C (clk), .D (signal_5382), .Q (signal_5383) ) ;
    buf_clk cell_3541 ( .C (clk), .D (signal_5390), .Q (signal_5391) ) ;
    buf_clk cell_3549 ( .C (clk), .D (signal_5398), .Q (signal_5399) ) ;
    buf_clk cell_3557 ( .C (clk), .D (signal_5406), .Q (signal_5407) ) ;
    buf_clk cell_3565 ( .C (clk), .D (signal_5414), .Q (signal_5415) ) ;
    buf_clk cell_3573 ( .C (clk), .D (signal_5422), .Q (signal_5423) ) ;
    buf_clk cell_3581 ( .C (clk), .D (signal_5430), .Q (signal_5431) ) ;
    buf_clk cell_3589 ( .C (clk), .D (signal_5438), .Q (signal_5439) ) ;
    buf_clk cell_3597 ( .C (clk), .D (signal_5446), .Q (signal_5447) ) ;
    buf_clk cell_3605 ( .C (clk), .D (signal_5454), .Q (signal_5455) ) ;
    buf_clk cell_3613 ( .C (clk), .D (signal_5462), .Q (signal_5463) ) ;
    buf_clk cell_3621 ( .C (clk), .D (signal_5470), .Q (signal_5471) ) ;
    buf_clk cell_3629 ( .C (clk), .D (signal_5478), .Q (signal_5479) ) ;
    buf_clk cell_3637 ( .C (clk), .D (signal_5486), .Q (signal_5487) ) ;
    buf_clk cell_3645 ( .C (clk), .D (signal_5494), .Q (signal_5495) ) ;
    buf_clk cell_3653 ( .C (clk), .D (signal_5502), .Q (signal_5503) ) ;
    buf_clk cell_3661 ( .C (clk), .D (signal_5510), .Q (signal_5511) ) ;
    buf_clk cell_3669 ( .C (clk), .D (signal_5518), .Q (signal_5519) ) ;
    buf_clk cell_3677 ( .C (clk), .D (signal_5526), .Q (signal_5527) ) ;
    buf_clk cell_3685 ( .C (clk), .D (signal_5534), .Q (signal_5535) ) ;
    buf_clk cell_3693 ( .C (clk), .D (signal_5542), .Q (signal_5543) ) ;
    buf_clk cell_3701 ( .C (clk), .D (signal_5550), .Q (signal_5551) ) ;
    buf_clk cell_3709 ( .C (clk), .D (signal_5558), .Q (signal_5559) ) ;
    buf_clk cell_3717 ( .C (clk), .D (signal_5566), .Q (signal_5567) ) ;
    buf_clk cell_3725 ( .C (clk), .D (signal_5574), .Q (signal_5575) ) ;
    buf_clk cell_3733 ( .C (clk), .D (signal_5582), .Q (signal_5583) ) ;
    buf_clk cell_3741 ( .C (clk), .D (signal_5590), .Q (signal_5591) ) ;
    buf_clk cell_3749 ( .C (clk), .D (signal_5598), .Q (signal_5599) ) ;
    buf_clk cell_3757 ( .C (clk), .D (signal_5606), .Q (signal_5607) ) ;
    buf_clk cell_3765 ( .C (clk), .D (signal_5614), .Q (signal_5615) ) ;
    buf_clk cell_3773 ( .C (clk), .D (signal_5622), .Q (signal_5623) ) ;
    buf_clk cell_3781 ( .C (clk), .D (signal_5630), .Q (signal_5631) ) ;
    buf_clk cell_3789 ( .C (clk), .D (signal_5638), .Q (signal_5639) ) ;
    buf_clk cell_3797 ( .C (clk), .D (signal_5646), .Q (signal_5647) ) ;
    buf_clk cell_3805 ( .C (clk), .D (signal_5654), .Q (signal_5655) ) ;
    buf_clk cell_3813 ( .C (clk), .D (signal_5662), .Q (signal_5663) ) ;
    buf_clk cell_3821 ( .C (clk), .D (signal_5670), .Q (signal_5671) ) ;
    buf_clk cell_3829 ( .C (clk), .D (signal_5678), .Q (signal_5679) ) ;
    buf_clk cell_3837 ( .C (clk), .D (signal_5686), .Q (signal_5687) ) ;
    buf_clk cell_3845 ( .C (clk), .D (signal_5694), .Q (signal_5695) ) ;
    buf_clk cell_3853 ( .C (clk), .D (signal_5702), .Q (signal_5703) ) ;
    buf_clk cell_3861 ( .C (clk), .D (signal_5710), .Q (signal_5711) ) ;
    buf_clk cell_3869 ( .C (clk), .D (signal_5718), .Q (signal_5719) ) ;
    buf_clk cell_3877 ( .C (clk), .D (signal_5726), .Q (signal_5727) ) ;
    buf_clk cell_3885 ( .C (clk), .D (signal_5734), .Q (signal_5735) ) ;
    buf_clk cell_3893 ( .C (clk), .D (signal_5742), .Q (signal_5743) ) ;
    buf_clk cell_3901 ( .C (clk), .D (signal_5750), .Q (signal_5751) ) ;
    buf_clk cell_3909 ( .C (clk), .D (signal_5758), .Q (signal_5759) ) ;
    buf_clk cell_3917 ( .C (clk), .D (signal_5766), .Q (signal_5767) ) ;
    buf_clk cell_3925 ( .C (clk), .D (signal_5774), .Q (signal_5775) ) ;
    buf_clk cell_3933 ( .C (clk), .D (signal_5782), .Q (signal_5783) ) ;
    buf_clk cell_3941 ( .C (clk), .D (signal_5790), .Q (signal_5791) ) ;
    buf_clk cell_3949 ( .C (clk), .D (signal_5798), .Q (signal_5799) ) ;
    buf_clk cell_3957 ( .C (clk), .D (signal_5806), .Q (signal_5807) ) ;
    buf_clk cell_3965 ( .C (clk), .D (signal_5814), .Q (signal_5815) ) ;
    buf_clk cell_3973 ( .C (clk), .D (signal_5822), .Q (signal_5823) ) ;
    buf_clk cell_3981 ( .C (clk), .D (signal_5830), .Q (signal_5831) ) ;
    buf_clk cell_3989 ( .C (clk), .D (signal_5838), .Q (signal_5839) ) ;
    buf_clk cell_3997 ( .C (clk), .D (signal_5846), .Q (signal_5847) ) ;
    buf_clk cell_4005 ( .C (clk), .D (signal_5854), .Q (signal_5855) ) ;
    buf_clk cell_4013 ( .C (clk), .D (signal_5862), .Q (signal_5863) ) ;
    buf_clk cell_4021 ( .C (clk), .D (signal_5870), .Q (signal_5871) ) ;
    buf_clk cell_4029 ( .C (clk), .D (signal_5878), .Q (signal_5879) ) ;
    buf_clk cell_4037 ( .C (clk), .D (signal_5886), .Q (signal_5887) ) ;
    buf_clk cell_4045 ( .C (clk), .D (signal_5894), .Q (signal_5895) ) ;
    buf_clk cell_4053 ( .C (clk), .D (signal_5902), .Q (signal_5903) ) ;
    buf_clk cell_4061 ( .C (clk), .D (signal_5910), .Q (signal_5911) ) ;
    buf_clk cell_4069 ( .C (clk), .D (signal_5918), .Q (signal_5919) ) ;
    buf_clk cell_4077 ( .C (clk), .D (signal_5926), .Q (signal_5927) ) ;
    buf_clk cell_4085 ( .C (clk), .D (signal_5934), .Q (signal_5935) ) ;
    buf_clk cell_4093 ( .C (clk), .D (signal_5942), .Q (signal_5943) ) ;
    buf_clk cell_4101 ( .C (clk), .D (signal_5950), .Q (signal_5951) ) ;
    buf_clk cell_4109 ( .C (clk), .D (signal_5958), .Q (signal_5959) ) ;
    buf_clk cell_4117 ( .C (clk), .D (signal_5966), .Q (signal_5967) ) ;
    buf_clk cell_4125 ( .C (clk), .D (signal_5974), .Q (signal_5975) ) ;
    buf_clk cell_4133 ( .C (clk), .D (signal_5982), .Q (signal_5983) ) ;
    buf_clk cell_4141 ( .C (clk), .D (signal_5990), .Q (signal_5991) ) ;
    buf_clk cell_4149 ( .C (clk), .D (signal_5998), .Q (signal_5999) ) ;
    buf_clk cell_4157 ( .C (clk), .D (signal_6006), .Q (signal_6007) ) ;
    buf_clk cell_4165 ( .C (clk), .D (signal_6014), .Q (signal_6015) ) ;
    buf_clk cell_4173 ( .C (clk), .D (signal_6022), .Q (signal_6023) ) ;
    buf_clk cell_4181 ( .C (clk), .D (signal_6030), .Q (signal_6031) ) ;
    buf_clk cell_4189 ( .C (clk), .D (signal_6038), .Q (signal_6039) ) ;
    buf_clk cell_4197 ( .C (clk), .D (signal_6046), .Q (signal_6047) ) ;
    buf_clk cell_4205 ( .C (clk), .D (signal_6054), .Q (signal_6055) ) ;
    buf_clk cell_4213 ( .C (clk), .D (signal_6062), .Q (signal_6063) ) ;
    buf_clk cell_4221 ( .C (clk), .D (signal_6070), .Q (signal_6071) ) ;
    buf_clk cell_4229 ( .C (clk), .D (signal_6078), .Q (signal_6079) ) ;
    buf_clk cell_4237 ( .C (clk), .D (signal_6086), .Q (signal_6087) ) ;
    buf_clk cell_4245 ( .C (clk), .D (signal_6094), .Q (signal_6095) ) ;
    buf_clk cell_4253 ( .C (clk), .D (signal_6102), .Q (signal_6103) ) ;
    buf_clk cell_4261 ( .C (clk), .D (signal_6110), .Q (signal_6111) ) ;
    buf_clk cell_4269 ( .C (clk), .D (signal_6118), .Q (signal_6119) ) ;
    buf_clk cell_4277 ( .C (clk), .D (signal_6126), .Q (signal_6127) ) ;
    buf_clk cell_4285 ( .C (clk), .D (signal_6134), .Q (signal_6135) ) ;
    buf_clk cell_4293 ( .C (clk), .D (signal_6142), .Q (signal_6143) ) ;
    buf_clk cell_4301 ( .C (clk), .D (signal_6150), .Q (signal_6151) ) ;
    buf_clk cell_4309 ( .C (clk), .D (signal_6158), .Q (signal_6159) ) ;
    buf_clk cell_4317 ( .C (clk), .D (signal_6166), .Q (signal_6167) ) ;
    buf_clk cell_4325 ( .C (clk), .D (signal_6174), .Q (signal_6175) ) ;
    buf_clk cell_4333 ( .C (clk), .D (signal_6182), .Q (signal_6183) ) ;
    buf_clk cell_4341 ( .C (clk), .D (signal_6190), .Q (signal_6191) ) ;
    buf_clk cell_4349 ( .C (clk), .D (signal_6198), .Q (signal_6199) ) ;
    buf_clk cell_4357 ( .C (clk), .D (signal_6206), .Q (signal_6207) ) ;
    buf_clk cell_4365 ( .C (clk), .D (signal_6214), .Q (signal_6215) ) ;
    buf_clk cell_4373 ( .C (clk), .D (signal_6222), .Q (signal_6223) ) ;
    buf_clk cell_4381 ( .C (clk), .D (signal_6230), .Q (signal_6231) ) ;
    buf_clk cell_4389 ( .C (clk), .D (signal_6238), .Q (signal_6239) ) ;
    buf_clk cell_4397 ( .C (clk), .D (signal_6246), .Q (signal_6247) ) ;
    buf_clk cell_4405 ( .C (clk), .D (signal_6254), .Q (signal_6255) ) ;
    buf_clk cell_4413 ( .C (clk), .D (signal_6262), .Q (signal_6263) ) ;
    buf_clk cell_4421 ( .C (clk), .D (signal_6270), .Q (signal_6271) ) ;
    buf_clk cell_4429 ( .C (clk), .D (signal_6278), .Q (signal_6279) ) ;
    buf_clk cell_4437 ( .C (clk), .D (signal_6286), .Q (signal_6287) ) ;
    buf_clk cell_4445 ( .C (clk), .D (signal_6294), .Q (signal_6295) ) ;
    buf_clk cell_4453 ( .C (clk), .D (signal_6302), .Q (signal_6303) ) ;
    buf_clk cell_4461 ( .C (clk), .D (signal_6310), .Q (signal_6311) ) ;
    buf_clk cell_4469 ( .C (clk), .D (signal_6318), .Q (signal_6319) ) ;
    buf_clk cell_4477 ( .C (clk), .D (signal_6326), .Q (signal_6327) ) ;
    buf_clk cell_4485 ( .C (clk), .D (signal_6334), .Q (signal_6335) ) ;
    buf_clk cell_4493 ( .C (clk), .D (signal_6342), .Q (signal_6343) ) ;
    buf_clk cell_4501 ( .C (clk), .D (signal_6350), .Q (signal_6351) ) ;
    buf_clk cell_4509 ( .C (clk), .D (signal_6358), .Q (signal_6359) ) ;
    buf_clk cell_4517 ( .C (clk), .D (signal_6366), .Q (signal_6367) ) ;
    buf_clk cell_4525 ( .C (clk), .D (signal_6374), .Q (signal_6375) ) ;
    buf_clk cell_4533 ( .C (clk), .D (signal_6382), .Q (signal_6383) ) ;
    buf_clk cell_4541 ( .C (clk), .D (signal_6390), .Q (signal_6391) ) ;
    buf_clk cell_4549 ( .C (clk), .D (signal_6398), .Q (signal_6399) ) ;
    buf_clk cell_4557 ( .C (clk), .D (signal_6406), .Q (signal_6407) ) ;
    buf_clk cell_4565 ( .C (clk), .D (signal_6414), .Q (signal_6415) ) ;
    buf_clk cell_4573 ( .C (clk), .D (signal_6422), .Q (signal_6423) ) ;
    buf_clk cell_4581 ( .C (clk), .D (signal_6430), .Q (signal_6431) ) ;
    buf_clk cell_4589 ( .C (clk), .D (signal_6438), .Q (signal_6439) ) ;
    buf_clk cell_4597 ( .C (clk), .D (signal_6446), .Q (signal_6447) ) ;
    buf_clk cell_4605 ( .C (clk), .D (signal_6454), .Q (signal_6455) ) ;
    buf_clk cell_4613 ( .C (clk), .D (signal_6462), .Q (signal_6463) ) ;
    buf_clk cell_4621 ( .C (clk), .D (signal_6470), .Q (signal_6471) ) ;
    buf_clk cell_4629 ( .C (clk), .D (signal_6478), .Q (signal_6479) ) ;
    buf_clk cell_4637 ( .C (clk), .D (signal_6486), .Q (signal_6487) ) ;
    buf_clk cell_4645 ( .C (clk), .D (signal_6494), .Q (signal_6495) ) ;
    buf_clk cell_4653 ( .C (clk), .D (signal_6502), .Q (signal_6503) ) ;
    buf_clk cell_4661 ( .C (clk), .D (signal_6510), .Q (signal_6511) ) ;
    buf_clk cell_4669 ( .C (clk), .D (signal_6518), .Q (signal_6519) ) ;
    buf_clk cell_4677 ( .C (clk), .D (signal_6526), .Q (signal_6527) ) ;
    buf_clk cell_4685 ( .C (clk), .D (signal_6534), .Q (signal_6535) ) ;
    buf_clk cell_4693 ( .C (clk), .D (signal_6542), .Q (signal_6543) ) ;
    buf_clk cell_4701 ( .C (clk), .D (signal_6550), .Q (signal_6551) ) ;
    buf_clk cell_4709 ( .C (clk), .D (signal_6558), .Q (signal_6559) ) ;
    buf_clk cell_4717 ( .C (clk), .D (signal_6566), .Q (signal_6567) ) ;
    buf_clk cell_4725 ( .C (clk), .D (signal_6574), .Q (signal_6575) ) ;
    buf_clk cell_4733 ( .C (clk), .D (signal_6582), .Q (signal_6583) ) ;
    buf_clk cell_4741 ( .C (clk), .D (signal_6590), .Q (signal_6591) ) ;
    buf_clk cell_4749 ( .C (clk), .D (signal_6598), .Q (signal_6599) ) ;
    buf_clk cell_4757 ( .C (clk), .D (signal_6606), .Q (signal_6607) ) ;
    buf_clk cell_4765 ( .C (clk), .D (signal_6614), .Q (signal_6615) ) ;
    buf_clk cell_4773 ( .C (clk), .D (signal_6622), .Q (signal_6623) ) ;
    buf_clk cell_4781 ( .C (clk), .D (signal_6630), .Q (signal_6631) ) ;
    buf_clk cell_4789 ( .C (clk), .D (signal_6638), .Q (signal_6639) ) ;
    buf_clk cell_4797 ( .C (clk), .D (signal_6646), .Q (signal_6647) ) ;
    buf_clk cell_4805 ( .C (clk), .D (signal_6654), .Q (signal_6655) ) ;
    buf_clk cell_4813 ( .C (clk), .D (signal_6662), .Q (signal_6663) ) ;
    buf_clk cell_4821 ( .C (clk), .D (signal_6670), .Q (signal_6671) ) ;
    buf_clk cell_4829 ( .C (clk), .D (signal_6678), .Q (signal_6679) ) ;
    buf_clk cell_4837 ( .C (clk), .D (signal_6686), .Q (signal_6687) ) ;
    buf_clk cell_4845 ( .C (clk), .D (signal_6694), .Q (signal_6695) ) ;
    buf_clk cell_4853 ( .C (clk), .D (signal_6702), .Q (signal_6703) ) ;
    buf_clk cell_4861 ( .C (clk), .D (signal_6710), .Q (signal_6711) ) ;
    buf_clk cell_4869 ( .C (clk), .D (signal_6718), .Q (signal_6719) ) ;
    buf_clk cell_4877 ( .C (clk), .D (signal_6726), .Q (signal_6727) ) ;
    buf_clk cell_4885 ( .C (clk), .D (signal_6734), .Q (signal_6735) ) ;
    buf_clk cell_4893 ( .C (clk), .D (signal_6742), .Q (signal_6743) ) ;
    buf_clk cell_4901 ( .C (clk), .D (signal_6750), .Q (signal_6751) ) ;
    buf_clk cell_4909 ( .C (clk), .D (signal_6758), .Q (signal_6759) ) ;
    buf_clk cell_4917 ( .C (clk), .D (signal_6766), .Q (signal_6767) ) ;
    buf_clk cell_4925 ( .C (clk), .D (signal_6774), .Q (signal_6775) ) ;
    buf_clk cell_4933 ( .C (clk), .D (signal_6782), .Q (signal_6783) ) ;
    buf_clk cell_4941 ( .C (clk), .D (signal_6790), .Q (signal_6791) ) ;
    buf_clk cell_4949 ( .C (clk), .D (signal_6798), .Q (signal_6799) ) ;
    buf_clk cell_4957 ( .C (clk), .D (signal_6806), .Q (signal_6807) ) ;
    buf_clk cell_4965 ( .C (clk), .D (signal_6814), .Q (signal_6815) ) ;
    buf_clk cell_4973 ( .C (clk), .D (signal_6822), .Q (signal_6823) ) ;
    buf_clk cell_4981 ( .C (clk), .D (signal_6830), .Q (signal_6831) ) ;
    buf_clk cell_4989 ( .C (clk), .D (signal_6838), .Q (signal_6839) ) ;
    buf_clk cell_4997 ( .C (clk), .D (signal_6846), .Q (signal_6847) ) ;
    buf_clk cell_5005 ( .C (clk), .D (signal_6854), .Q (signal_6855) ) ;
    buf_clk cell_5013 ( .C (clk), .D (signal_6862), .Q (signal_6863) ) ;
    buf_clk cell_5021 ( .C (clk), .D (signal_6870), .Q (signal_6871) ) ;
    buf_clk cell_5029 ( .C (clk), .D (signal_6878), .Q (signal_6879) ) ;
    buf_clk cell_5037 ( .C (clk), .D (signal_6886), .Q (signal_6887) ) ;
    buf_clk cell_5045 ( .C (clk), .D (signal_6894), .Q (signal_6895) ) ;
    buf_clk cell_5053 ( .C (clk), .D (signal_6902), .Q (signal_6903) ) ;
    buf_clk cell_5061 ( .C (clk), .D (signal_6910), .Q (signal_6911) ) ;
    buf_clk cell_5069 ( .C (clk), .D (signal_6918), .Q (signal_6919) ) ;
    buf_clk cell_5077 ( .C (clk), .D (signal_6926), .Q (signal_6927) ) ;
    buf_clk cell_5085 ( .C (clk), .D (signal_6934), .Q (signal_6935) ) ;
    buf_clk cell_5093 ( .C (clk), .D (signal_6942), .Q (signal_6943) ) ;
    buf_clk cell_5101 ( .C (clk), .D (signal_6950), .Q (signal_6951) ) ;
    buf_clk cell_5109 ( .C (clk), .D (signal_6958), .Q (signal_6959) ) ;
    buf_clk cell_5117 ( .C (clk), .D (signal_6966), .Q (signal_6967) ) ;
    buf_clk cell_5125 ( .C (clk), .D (signal_6974), .Q (signal_6975) ) ;
    buf_clk cell_5133 ( .C (clk), .D (signal_6982), .Q (signal_6983) ) ;
    buf_clk cell_5141 ( .C (clk), .D (signal_6990), .Q (signal_6991) ) ;
    buf_clk cell_5149 ( .C (clk), .D (signal_6998), .Q (signal_6999) ) ;
    buf_clk cell_5157 ( .C (clk), .D (signal_7006), .Q (signal_7007) ) ;
    buf_clk cell_5165 ( .C (clk), .D (signal_7014), .Q (signal_7015) ) ;
    buf_clk cell_5173 ( .C (clk), .D (signal_7022), .Q (signal_7023) ) ;
    buf_clk cell_5181 ( .C (clk), .D (signal_7030), .Q (signal_7031) ) ;
    buf_clk cell_5189 ( .C (clk), .D (signal_7038), .Q (signal_7039) ) ;
    buf_clk cell_5197 ( .C (clk), .D (signal_7046), .Q (signal_7047) ) ;
    buf_clk cell_5205 ( .C (clk), .D (signal_7054), .Q (signal_7055) ) ;
    buf_clk cell_5213 ( .C (clk), .D (signal_7062), .Q (signal_7063) ) ;
    buf_clk cell_5221 ( .C (clk), .D (signal_7070), .Q (signal_7071) ) ;
    buf_clk cell_5229 ( .C (clk), .D (signal_7078), .Q (signal_7079) ) ;
    buf_clk cell_5237 ( .C (clk), .D (signal_7086), .Q (signal_7087) ) ;
    buf_clk cell_5245 ( .C (clk), .D (signal_7094), .Q (signal_7095) ) ;
    buf_clk cell_5253 ( .C (clk), .D (signal_7102), .Q (signal_7103) ) ;
    buf_clk cell_5261 ( .C (clk), .D (signal_7110), .Q (signal_7111) ) ;
    buf_clk cell_5269 ( .C (clk), .D (signal_7118), .Q (signal_7119) ) ;
    buf_clk cell_5277 ( .C (clk), .D (signal_7126), .Q (signal_7127) ) ;
    buf_clk cell_5285 ( .C (clk), .D (signal_7134), .Q (signal_7135) ) ;
    buf_clk cell_5293 ( .C (clk), .D (signal_7142), .Q (signal_7143) ) ;
    buf_clk cell_5301 ( .C (clk), .D (signal_7150), .Q (signal_7151) ) ;
    buf_clk cell_5309 ( .C (clk), .D (signal_7158), .Q (signal_7159) ) ;
    buf_clk cell_5317 ( .C (clk), .D (signal_7166), .Q (signal_7167) ) ;
    buf_clk cell_5325 ( .C (clk), .D (signal_7174), .Q (signal_7175) ) ;
    buf_clk cell_5333 ( .C (clk), .D (signal_7182), .Q (signal_7183) ) ;
    buf_clk cell_5341 ( .C (clk), .D (signal_7190), .Q (signal_7191) ) ;
    buf_clk cell_5349 ( .C (clk), .D (signal_7198), .Q (signal_7199) ) ;
    buf_clk cell_5357 ( .C (clk), .D (signal_7206), .Q (signal_7207) ) ;
    buf_clk cell_5365 ( .C (clk), .D (signal_7214), .Q (signal_7215) ) ;
    buf_clk cell_5373 ( .C (clk), .D (signal_7222), .Q (signal_7223) ) ;
    buf_clk cell_5381 ( .C (clk), .D (signal_7230), .Q (signal_7231) ) ;
    buf_clk cell_5389 ( .C (clk), .D (signal_7238), .Q (signal_7239) ) ;
    buf_clk cell_5397 ( .C (clk), .D (signal_7246), .Q (signal_7247) ) ;
    buf_clk cell_5405 ( .C (clk), .D (signal_7254), .Q (signal_7255) ) ;
    buf_clk cell_5413 ( .C (clk), .D (signal_7262), .Q (signal_7263) ) ;
    buf_clk cell_5421 ( .C (clk), .D (signal_7270), .Q (signal_7271) ) ;
    buf_clk cell_5429 ( .C (clk), .D (signal_7278), .Q (signal_7279) ) ;
    buf_clk cell_5437 ( .C (clk), .D (signal_7286), .Q (signal_7287) ) ;
    buf_clk cell_5445 ( .C (clk), .D (signal_7294), .Q (signal_7295) ) ;
    buf_clk cell_5453 ( .C (clk), .D (signal_7302), .Q (signal_7303) ) ;
    buf_clk cell_5461 ( .C (clk), .D (signal_7310), .Q (signal_7311) ) ;
    buf_clk cell_5469 ( .C (clk), .D (signal_7318), .Q (signal_7319) ) ;
    buf_clk cell_5477 ( .C (clk), .D (signal_7326), .Q (signal_7327) ) ;
    buf_clk cell_5485 ( .C (clk), .D (signal_7334), .Q (signal_7335) ) ;
    buf_clk cell_5493 ( .C (clk), .D (signal_7342), .Q (signal_7343) ) ;
    buf_clk cell_5501 ( .C (clk), .D (signal_7350), .Q (signal_7351) ) ;
    buf_clk cell_5509 ( .C (clk), .D (signal_7358), .Q (signal_7359) ) ;
    buf_clk cell_5517 ( .C (clk), .D (signal_7366), .Q (signal_7367) ) ;
    buf_clk cell_5525 ( .C (clk), .D (signal_7374), .Q (signal_7375) ) ;
    buf_clk cell_5533 ( .C (clk), .D (signal_7382), .Q (signal_7383) ) ;
    buf_clk cell_5541 ( .C (clk), .D (signal_7390), .Q (signal_7391) ) ;
    buf_clk cell_5549 ( .C (clk), .D (signal_7398), .Q (signal_7399) ) ;
    buf_clk cell_5557 ( .C (clk), .D (signal_7406), .Q (signal_7407) ) ;
    buf_clk cell_5565 ( .C (clk), .D (signal_7414), .Q (signal_7415) ) ;
    buf_clk cell_5573 ( .C (clk), .D (signal_7422), .Q (signal_7423) ) ;
    buf_clk cell_5581 ( .C (clk), .D (signal_7430), .Q (signal_7431) ) ;
    buf_clk cell_5589 ( .C (clk), .D (signal_7438), .Q (signal_7439) ) ;
    buf_clk cell_5597 ( .C (clk), .D (signal_7446), .Q (signal_7447) ) ;
    buf_clk cell_5605 ( .C (clk), .D (signal_7454), .Q (signal_7455) ) ;
    buf_clk cell_5613 ( .C (clk), .D (signal_7462), .Q (signal_7463) ) ;
    buf_clk cell_5621 ( .C (clk), .D (signal_7470), .Q (signal_7471) ) ;
    buf_clk cell_5629 ( .C (clk), .D (signal_7478), .Q (signal_7479) ) ;
    buf_clk cell_5637 ( .C (clk), .D (signal_7486), .Q (signal_7487) ) ;
    buf_clk cell_5645 ( .C (clk), .D (signal_7494), .Q (signal_7495) ) ;
    buf_clk cell_5653 ( .C (clk), .D (signal_7502), .Q (signal_7503) ) ;
    buf_clk cell_5661 ( .C (clk), .D (signal_7510), .Q (signal_7511) ) ;
    buf_clk cell_5669 ( .C (clk), .D (signal_7518), .Q (signal_7519) ) ;
    buf_clk cell_5677 ( .C (clk), .D (signal_7526), .Q (signal_7527) ) ;
    buf_clk cell_5685 ( .C (clk), .D (signal_7534), .Q (signal_7535) ) ;
    buf_clk cell_5693 ( .C (clk), .D (signal_7542), .Q (signal_7543) ) ;
    buf_clk cell_5701 ( .C (clk), .D (signal_7550), .Q (signal_7551) ) ;
    buf_clk cell_5709 ( .C (clk), .D (signal_7558), .Q (signal_7559) ) ;
    buf_clk cell_5717 ( .C (clk), .D (signal_7566), .Q (signal_7567) ) ;
    buf_clk cell_5725 ( .C (clk), .D (signal_7574), .Q (signal_7575) ) ;
    buf_clk cell_5733 ( .C (clk), .D (signal_7582), .Q (signal_7583) ) ;
    buf_clk cell_5741 ( .C (clk), .D (signal_7590), .Q (signal_7591) ) ;
    buf_clk cell_5749 ( .C (clk), .D (signal_7598), .Q (signal_7599) ) ;
    buf_clk cell_5757 ( .C (clk), .D (signal_7606), .Q (signal_7607) ) ;
    buf_clk cell_5765 ( .C (clk), .D (signal_7614), .Q (signal_7615) ) ;
    buf_clk cell_5773 ( .C (clk), .D (signal_7622), .Q (signal_7623) ) ;
    buf_clk cell_5781 ( .C (clk), .D (signal_7630), .Q (signal_7631) ) ;
    buf_clk cell_5789 ( .C (clk), .D (signal_7638), .Q (signal_7639) ) ;
    buf_clk cell_5797 ( .C (clk), .D (signal_7646), .Q (signal_7647) ) ;
    buf_clk cell_5805 ( .C (clk), .D (signal_7654), .Q (signal_7655) ) ;
    buf_clk cell_5813 ( .C (clk), .D (signal_7662), .Q (signal_7663) ) ;
    buf_clk cell_5821 ( .C (clk), .D (signal_7670), .Q (signal_7671) ) ;
    buf_clk cell_5829 ( .C (clk), .D (signal_7678), .Q (signal_7679) ) ;
    buf_clk cell_5837 ( .C (clk), .D (signal_7686), .Q (signal_7687) ) ;
    buf_clk cell_5845 ( .C (clk), .D (signal_7694), .Q (signal_7695) ) ;
    buf_clk cell_5853 ( .C (clk), .D (signal_7702), .Q (signal_7703) ) ;
    buf_clk cell_5861 ( .C (clk), .D (signal_7710), .Q (signal_7711) ) ;
    buf_clk cell_5869 ( .C (clk), .D (signal_7718), .Q (signal_7719) ) ;
    buf_clk cell_5877 ( .C (clk), .D (signal_7726), .Q (signal_7727) ) ;
    buf_clk cell_5885 ( .C (clk), .D (signal_7734), .Q (signal_7735) ) ;
    buf_clk cell_5893 ( .C (clk), .D (signal_7742), .Q (signal_7743) ) ;
    buf_clk cell_5901 ( .C (clk), .D (signal_7750), .Q (signal_7751) ) ;
    buf_clk cell_5909 ( .C (clk), .D (signal_7758), .Q (signal_7759) ) ;
    buf_clk cell_5917 ( .C (clk), .D (signal_7766), .Q (signal_7767) ) ;
    buf_clk cell_5925 ( .C (clk), .D (signal_7774), .Q (signal_7775) ) ;
    buf_clk cell_5933 ( .C (clk), .D (signal_7782), .Q (signal_7783) ) ;
    buf_clk cell_5941 ( .C (clk), .D (signal_7790), .Q (signal_7791) ) ;
    buf_clk cell_5949 ( .C (clk), .D (signal_7798), .Q (signal_7799) ) ;
    buf_clk cell_5957 ( .C (clk), .D (signal_7806), .Q (signal_7807) ) ;
    buf_clk cell_5965 ( .C (clk), .D (signal_7814), .Q (signal_7815) ) ;
    buf_clk cell_5973 ( .C (clk), .D (signal_7822), .Q (signal_7823) ) ;
    buf_clk cell_5981 ( .C (clk), .D (signal_7830), .Q (signal_7831) ) ;
    buf_clk cell_5989 ( .C (clk), .D (signal_7838), .Q (signal_7839) ) ;
    buf_clk cell_5997 ( .C (clk), .D (signal_7846), .Q (signal_7847) ) ;
    buf_clk cell_6005 ( .C (clk), .D (signal_7854), .Q (signal_7855) ) ;
    buf_clk cell_6013 ( .C (clk), .D (signal_7862), .Q (signal_7863) ) ;
    buf_clk cell_6021 ( .C (clk), .D (signal_7870), .Q (signal_7871) ) ;
    buf_clk cell_6029 ( .C (clk), .D (signal_7878), .Q (signal_7879) ) ;
    buf_clk cell_6037 ( .C (clk), .D (signal_7886), .Q (signal_7887) ) ;
    buf_clk cell_6045 ( .C (clk), .D (signal_7894), .Q (signal_7895) ) ;
    buf_clk cell_6053 ( .C (clk), .D (signal_7902), .Q (signal_7903) ) ;
    buf_clk cell_6061 ( .C (clk), .D (signal_7910), .Q (signal_7911) ) ;
    buf_clk cell_6069 ( .C (clk), .D (signal_7918), .Q (signal_7919) ) ;
    buf_clk cell_6077 ( .C (clk), .D (signal_7926), .Q (signal_7927) ) ;
    buf_clk cell_6085 ( .C (clk), .D (signal_7934), .Q (signal_7935) ) ;
    buf_clk cell_6093 ( .C (clk), .D (signal_7942), .Q (signal_7943) ) ;
    buf_clk cell_6101 ( .C (clk), .D (signal_7950), .Q (signal_7951) ) ;
    buf_clk cell_6109 ( .C (clk), .D (signal_7958), .Q (signal_7959) ) ;
    buf_clk cell_6117 ( .C (clk), .D (signal_7966), .Q (signal_7967) ) ;
    buf_clk cell_6125 ( .C (clk), .D (signal_7974), .Q (signal_7975) ) ;
    buf_clk cell_6133 ( .C (clk), .D (signal_7982), .Q (signal_7983) ) ;
    buf_clk cell_6141 ( .C (clk), .D (signal_7990), .Q (signal_7991) ) ;
    buf_clk cell_6149 ( .C (clk), .D (signal_7998), .Q (signal_7999) ) ;
    buf_clk cell_6157 ( .C (clk), .D (signal_8006), .Q (signal_8007) ) ;
    buf_clk cell_6165 ( .C (clk), .D (signal_8014), .Q (signal_8015) ) ;
    buf_clk cell_6173 ( .C (clk), .D (signal_8022), .Q (signal_8023) ) ;
    buf_clk cell_6181 ( .C (clk), .D (signal_8030), .Q (signal_8031) ) ;
    buf_clk cell_6189 ( .C (clk), .D (signal_8038), .Q (signal_8039) ) ;
    buf_clk cell_6197 ( .C (clk), .D (signal_8046), .Q (signal_8047) ) ;
    buf_clk cell_6205 ( .C (clk), .D (signal_8054), .Q (signal_8055) ) ;
    buf_clk cell_6213 ( .C (clk), .D (signal_8062), .Q (signal_8063) ) ;
    buf_clk cell_6221 ( .C (clk), .D (signal_8070), .Q (signal_8071) ) ;
    buf_clk cell_6229 ( .C (clk), .D (signal_8078), .Q (signal_8079) ) ;
    buf_clk cell_6237 ( .C (clk), .D (signal_8086), .Q (signal_8087) ) ;
    buf_clk cell_6245 ( .C (clk), .D (signal_8094), .Q (signal_8095) ) ;
    buf_clk cell_6253 ( .C (clk), .D (signal_8102), .Q (signal_8103) ) ;
    buf_clk cell_6261 ( .C (clk), .D (signal_8110), .Q (signal_8111) ) ;
    buf_clk cell_6269 ( .C (clk), .D (signal_8118), .Q (signal_8119) ) ;
    buf_clk cell_6277 ( .C (clk), .D (signal_8126), .Q (signal_8127) ) ;
    buf_clk cell_6285 ( .C (clk), .D (signal_8134), .Q (signal_8135) ) ;
    buf_clk cell_6293 ( .C (clk), .D (signal_8142), .Q (signal_8143) ) ;
    buf_clk cell_6301 ( .C (clk), .D (signal_8150), .Q (signal_8151) ) ;
    buf_clk cell_6309 ( .C (clk), .D (signal_8158), .Q (signal_8159) ) ;
    buf_clk cell_6317 ( .C (clk), .D (signal_8166), .Q (signal_8167) ) ;
    buf_clk cell_6325 ( .C (clk), .D (signal_8174), .Q (signal_8175) ) ;
    buf_clk cell_6333 ( .C (clk), .D (signal_8182), .Q (signal_8183) ) ;
    buf_clk cell_6341 ( .C (clk), .D (signal_8190), .Q (signal_8191) ) ;
    buf_clk cell_6349 ( .C (clk), .D (signal_8198), .Q (signal_8199) ) ;
    buf_clk cell_6357 ( .C (clk), .D (signal_8206), .Q (signal_8207) ) ;
    buf_clk cell_6365 ( .C (clk), .D (signal_8214), .Q (signal_8215) ) ;
    buf_clk cell_6373 ( .C (clk), .D (signal_8222), .Q (signal_8223) ) ;
    buf_clk cell_6381 ( .C (clk), .D (signal_8230), .Q (signal_8231) ) ;
    buf_clk cell_6389 ( .C (clk), .D (signal_8238), .Q (signal_8239) ) ;
    buf_clk cell_6397 ( .C (clk), .D (signal_8246), .Q (signal_8247) ) ;
    buf_clk cell_6405 ( .C (clk), .D (signal_8254), .Q (signal_8255) ) ;
    buf_clk cell_6413 ( .C (clk), .D (signal_8262), .Q (signal_8263) ) ;
    buf_clk cell_6421 ( .C (clk), .D (signal_8270), .Q (signal_8271) ) ;
    buf_clk cell_6429 ( .C (clk), .D (signal_8278), .Q (signal_8279) ) ;
    buf_clk cell_6437 ( .C (clk), .D (signal_8286), .Q (signal_8287) ) ;
    buf_clk cell_6445 ( .C (clk), .D (signal_8294), .Q (signal_8295) ) ;
    buf_clk cell_6453 ( .C (clk), .D (signal_8302), .Q (signal_8303) ) ;
    buf_clk cell_6461 ( .C (clk), .D (signal_8310), .Q (signal_8311) ) ;
    buf_clk cell_6469 ( .C (clk), .D (signal_8318), .Q (signal_8319) ) ;
    buf_clk cell_6477 ( .C (clk), .D (signal_8326), .Q (signal_8327) ) ;
    buf_clk cell_6485 ( .C (clk), .D (signal_8334), .Q (signal_8335) ) ;
    buf_clk cell_6493 ( .C (clk), .D (signal_8342), .Q (signal_8343) ) ;
    buf_clk cell_6501 ( .C (clk), .D (signal_8350), .Q (signal_8351) ) ;
    buf_clk cell_6509 ( .C (clk), .D (signal_8358), .Q (signal_8359) ) ;
    buf_clk cell_6517 ( .C (clk), .D (signal_8366), .Q (signal_8367) ) ;
    buf_clk cell_6525 ( .C (clk), .D (signal_8374), .Q (signal_8375) ) ;
    buf_clk cell_6533 ( .C (clk), .D (signal_8382), .Q (signal_8383) ) ;
    buf_clk cell_6541 ( .C (clk), .D (signal_8390), .Q (signal_8391) ) ;
    buf_clk cell_6549 ( .C (clk), .D (signal_8398), .Q (signal_8399) ) ;
    buf_clk cell_6557 ( .C (clk), .D (signal_8406), .Q (signal_8407) ) ;
    buf_clk cell_6565 ( .C (clk), .D (signal_8414), .Q (signal_8415) ) ;
    buf_clk cell_6573 ( .C (clk), .D (signal_8422), .Q (signal_8423) ) ;
    buf_clk cell_6581 ( .C (clk), .D (signal_8430), .Q (signal_8431) ) ;
    buf_clk cell_6589 ( .C (clk), .D (signal_8438), .Q (signal_8439) ) ;
    buf_clk cell_6597 ( .C (clk), .D (signal_8446), .Q (signal_8447) ) ;
    buf_clk cell_6605 ( .C (clk), .D (signal_8454), .Q (signal_8455) ) ;
    buf_clk cell_6613 ( .C (clk), .D (signal_8462), .Q (signal_8463) ) ;
    buf_clk cell_6621 ( .C (clk), .D (signal_8470), .Q (signal_8471) ) ;
    buf_clk cell_6629 ( .C (clk), .D (signal_8478), .Q (signal_8479) ) ;
    buf_clk cell_6637 ( .C (clk), .D (signal_8486), .Q (signal_8487) ) ;
    buf_clk cell_6645 ( .C (clk), .D (signal_8494), .Q (signal_8495) ) ;
    buf_clk cell_6653 ( .C (clk), .D (signal_8502), .Q (signal_8503) ) ;
    buf_clk cell_6661 ( .C (clk), .D (signal_8510), .Q (signal_8511) ) ;
    buf_clk cell_6669 ( .C (clk), .D (signal_8518), .Q (signal_8519) ) ;
    buf_clk cell_6677 ( .C (clk), .D (signal_8526), .Q (signal_8527) ) ;
    buf_clk cell_6685 ( .C (clk), .D (signal_8534), .Q (signal_8535) ) ;
    buf_clk cell_6693 ( .C (clk), .D (signal_8542), .Q (signal_8543) ) ;
    buf_clk cell_6701 ( .C (clk), .D (signal_8550), .Q (signal_8551) ) ;
    buf_clk cell_6709 ( .C (clk), .D (signal_8558), .Q (signal_8559) ) ;
    buf_clk cell_6717 ( .C (clk), .D (signal_8566), .Q (signal_8567) ) ;
    buf_clk cell_6725 ( .C (clk), .D (signal_8574), .Q (signal_8575) ) ;
    buf_clk cell_6733 ( .C (clk), .D (signal_8582), .Q (signal_8583) ) ;
    buf_clk cell_6741 ( .C (clk), .D (signal_8590), .Q (signal_8591) ) ;
    buf_clk cell_6749 ( .C (clk), .D (signal_8598), .Q (signal_8599) ) ;
    buf_clk cell_6757 ( .C (clk), .D (signal_8606), .Q (signal_8607) ) ;
    buf_clk cell_6765 ( .C (clk), .D (signal_8614), .Q (signal_8615) ) ;
    buf_clk cell_6773 ( .C (clk), .D (signal_8622), .Q (signal_8623) ) ;
    buf_clk cell_6781 ( .C (clk), .D (signal_8630), .Q (signal_8631) ) ;
    buf_clk cell_6789 ( .C (clk), .D (signal_8638), .Q (signal_8639) ) ;
    buf_clk cell_6797 ( .C (clk), .D (signal_8646), .Q (signal_8647) ) ;
    buf_clk cell_6805 ( .C (clk), .D (signal_8654), .Q (signal_8655) ) ;
    buf_clk cell_6813 ( .C (clk), .D (signal_8662), .Q (signal_8663) ) ;
    buf_clk cell_6821 ( .C (clk), .D (signal_8670), .Q (signal_8671) ) ;
    buf_clk cell_6829 ( .C (clk), .D (signal_8678), .Q (signal_8679) ) ;
    buf_clk cell_6837 ( .C (clk), .D (signal_8686), .Q (signal_8687) ) ;
    buf_clk cell_6845 ( .C (clk), .D (signal_8694), .Q (signal_8695) ) ;
    buf_clk cell_6853 ( .C (clk), .D (signal_8702), .Q (signal_8703) ) ;
    buf_clk cell_6861 ( .C (clk), .D (signal_8710), .Q (signal_8711) ) ;
    buf_clk cell_6869 ( .C (clk), .D (signal_8718), .Q (signal_8719) ) ;
    buf_clk cell_6877 ( .C (clk), .D (signal_8726), .Q (signal_8727) ) ;
    buf_clk cell_6885 ( .C (clk), .D (signal_8734), .Q (signal_8735) ) ;
    buf_clk cell_6893 ( .C (clk), .D (signal_8742), .Q (signal_8743) ) ;
    buf_clk cell_6901 ( .C (clk), .D (signal_8750), .Q (signal_8751) ) ;
    buf_clk cell_6909 ( .C (clk), .D (signal_8758), .Q (signal_8759) ) ;
    buf_clk cell_6917 ( .C (clk), .D (signal_8766), .Q (signal_8767) ) ;
    buf_clk cell_6925 ( .C (clk), .D (signal_8774), .Q (signal_8775) ) ;
    buf_clk cell_6933 ( .C (clk), .D (signal_8782), .Q (signal_8783) ) ;
    buf_clk cell_6941 ( .C (clk), .D (signal_8790), .Q (signal_8791) ) ;
    buf_clk cell_6949 ( .C (clk), .D (signal_8798), .Q (signal_8799) ) ;
    buf_clk cell_6957 ( .C (clk), .D (signal_8806), .Q (signal_8807) ) ;
    buf_clk cell_6965 ( .C (clk), .D (signal_8814), .Q (signal_8815) ) ;
    buf_clk cell_6973 ( .C (clk), .D (signal_8822), .Q (signal_8823) ) ;
    buf_clk cell_6981 ( .C (clk), .D (signal_8830), .Q (signal_8831) ) ;
    buf_clk cell_6989 ( .C (clk), .D (signal_8838), .Q (signal_8839) ) ;
    buf_clk cell_6997 ( .C (clk), .D (signal_8846), .Q (signal_8847) ) ;
    buf_clk cell_7005 ( .C (clk), .D (signal_8854), .Q (signal_8855) ) ;
    buf_clk cell_7013 ( .C (clk), .D (signal_8862), .Q (signal_8863) ) ;
    buf_clk cell_7021 ( .C (clk), .D (signal_8870), .Q (signal_8871) ) ;
    buf_clk cell_7029 ( .C (clk), .D (signal_8878), .Q (signal_8879) ) ;
    buf_clk cell_7037 ( .C (clk), .D (signal_8886), .Q (signal_8887) ) ;
    buf_clk cell_7045 ( .C (clk), .D (signal_8894), .Q (signal_8895) ) ;
    buf_clk cell_7053 ( .C (clk), .D (signal_8902), .Q (signal_8903) ) ;
    buf_clk cell_7061 ( .C (clk), .D (signal_8910), .Q (signal_8911) ) ;
    buf_clk cell_7069 ( .C (clk), .D (signal_8918), .Q (signal_8919) ) ;
    buf_clk cell_7077 ( .C (clk), .D (signal_8926), .Q (signal_8927) ) ;
    buf_clk cell_7085 ( .C (clk), .D (signal_8934), .Q (signal_8935) ) ;
    buf_clk cell_7093 ( .C (clk), .D (signal_8942), .Q (signal_8943) ) ;
    buf_clk cell_7101 ( .C (clk), .D (signal_8950), .Q (signal_8951) ) ;

    /* register cells */
    DFF_X1 cell_33 ( .CK (clk), .D (signal_4975), .Q (signal_425), .QN () ) ;
    DFF_X1 cell_36 ( .CK (clk), .D (signal_4983), .Q (signal_426), .QN () ) ;
    DFF_X1 cell_39 ( .CK (clk), .D (signal_4991), .Q (signal_427), .QN () ) ;
    DFF_X1 cell_42 ( .CK (clk), .D (signal_4999), .Q (signal_428), .QN () ) ;
    DFF_X1 cell_45 ( .CK (clk), .D (signal_5007), .Q (signal_424), .QN () ) ;
    DFF_X1 cell_48 ( .CK (clk), .D (signal_5015), .Q (signal_421), .QN () ) ;
    DFF_X1 cell_51 ( .CK (clk), .D (signal_5023), .Q (signal_420), .QN () ) ;
    DFF_X1 cell_53 ( .CK (clk), .D (signal_5031), .Q (signal_418), .QN () ) ;
    DFF_X1 cell_55 ( .CK (clk), .D (signal_5039), .Q (signal_397), .QN () ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_87 ( .clk (clk), .D ({signal_5055, signal_5047}), .Q ({ciphertext_s1[120], ciphertext_s0[120]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_90 ( .clk (clk), .D ({signal_5071, signal_5063}), .Q ({ciphertext_s1[121], ciphertext_s0[121]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_93 ( .clk (clk), .D ({signal_5087, signal_5079}), .Q ({ciphertext_s1[122], ciphertext_s0[122]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_96 ( .clk (clk), .D ({signal_5103, signal_5095}), .Q ({ciphertext_s1[123], ciphertext_s0[123]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_99 ( .clk (clk), .D ({signal_5119, signal_5111}), .Q ({ciphertext_s1[124], ciphertext_s0[124]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_102 ( .clk (clk), .D ({signal_5135, signal_5127}), .Q ({ciphertext_s1[125], ciphertext_s0[125]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_105 ( .clk (clk), .D ({signal_5151, signal_5143}), .Q ({ciphertext_s1[126], ciphertext_s0[126]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_108 ( .clk (clk), .D ({signal_5167, signal_5159}), .Q ({ciphertext_s1[127], ciphertext_s0[127]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_111 ( .clk (clk), .D ({signal_5183, signal_5175}), .Q ({ciphertext_s1[112], ciphertext_s0[112]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_114 ( .clk (clk), .D ({signal_5199, signal_5191}), .Q ({ciphertext_s1[113], ciphertext_s0[113]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_117 ( .clk (clk), .D ({signal_5215, signal_5207}), .Q ({ciphertext_s1[114], ciphertext_s0[114]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_120 ( .clk (clk), .D ({signal_5231, signal_5223}), .Q ({ciphertext_s1[115], ciphertext_s0[115]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_123 ( .clk (clk), .D ({signal_5247, signal_5239}), .Q ({ciphertext_s1[116], ciphertext_s0[116]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_126 ( .clk (clk), .D ({signal_5263, signal_5255}), .Q ({ciphertext_s1[117], ciphertext_s0[117]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_129 ( .clk (clk), .D ({signal_5279, signal_5271}), .Q ({ciphertext_s1[118], ciphertext_s0[118]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_132 ( .clk (clk), .D ({signal_5295, signal_5287}), .Q ({ciphertext_s1[119], ciphertext_s0[119]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_135 ( .clk (clk), .D ({signal_5311, signal_5303}), .Q ({ciphertext_s1[104], ciphertext_s0[104]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_138 ( .clk (clk), .D ({signal_5327, signal_5319}), .Q ({ciphertext_s1[105], ciphertext_s0[105]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_141 ( .clk (clk), .D ({signal_5343, signal_5335}), .Q ({ciphertext_s1[106], ciphertext_s0[106]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_144 ( .clk (clk), .D ({signal_5359, signal_5351}), .Q ({ciphertext_s1[107], ciphertext_s0[107]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_147 ( .clk (clk), .D ({signal_5375, signal_5367}), .Q ({ciphertext_s1[108], ciphertext_s0[108]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_150 ( .clk (clk), .D ({signal_5391, signal_5383}), .Q ({ciphertext_s1[109], ciphertext_s0[109]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_153 ( .clk (clk), .D ({signal_5407, signal_5399}), .Q ({ciphertext_s1[110], ciphertext_s0[110]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_156 ( .clk (clk), .D ({signal_5423, signal_5415}), .Q ({ciphertext_s1[111], ciphertext_s0[111]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_159 ( .clk (clk), .D ({signal_5439, signal_5431}), .Q ({ciphertext_s1[96], ciphertext_s0[96]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_162 ( .clk (clk), .D ({signal_5455, signal_5447}), .Q ({ciphertext_s1[97], ciphertext_s0[97]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_165 ( .clk (clk), .D ({signal_5471, signal_5463}), .Q ({ciphertext_s1[98], ciphertext_s0[98]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_168 ( .clk (clk), .D ({signal_5487, signal_5479}), .Q ({ciphertext_s1[99], ciphertext_s0[99]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_171 ( .clk (clk), .D ({signal_5503, signal_5495}), .Q ({ciphertext_s1[100], ciphertext_s0[100]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_174 ( .clk (clk), .D ({signal_5519, signal_5511}), .Q ({ciphertext_s1[101], ciphertext_s0[101]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_177 ( .clk (clk), .D ({signal_5535, signal_5527}), .Q ({ciphertext_s1[102], ciphertext_s0[102]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_180 ( .clk (clk), .D ({signal_5551, signal_5543}), .Q ({ciphertext_s1[103], ciphertext_s0[103]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_183 ( .clk (clk), .D ({signal_5567, signal_5559}), .Q ({ciphertext_s1[88], ciphertext_s0[88]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_186 ( .clk (clk), .D ({signal_5583, signal_5575}), .Q ({ciphertext_s1[89], ciphertext_s0[89]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_189 ( .clk (clk), .D ({signal_5599, signal_5591}), .Q ({ciphertext_s1[90], ciphertext_s0[90]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_192 ( .clk (clk), .D ({signal_5615, signal_5607}), .Q ({ciphertext_s1[91], ciphertext_s0[91]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_195 ( .clk (clk), .D ({signal_5631, signal_5623}), .Q ({ciphertext_s1[92], ciphertext_s0[92]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_198 ( .clk (clk), .D ({signal_5647, signal_5639}), .Q ({ciphertext_s1[93], ciphertext_s0[93]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_201 ( .clk (clk), .D ({signal_5663, signal_5655}), .Q ({ciphertext_s1[94], ciphertext_s0[94]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_204 ( .clk (clk), .D ({signal_5679, signal_5671}), .Q ({ciphertext_s1[95], ciphertext_s0[95]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_207 ( .clk (clk), .D ({signal_5695, signal_5687}), .Q ({ciphertext_s1[80], ciphertext_s0[80]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_210 ( .clk (clk), .D ({signal_5711, signal_5703}), .Q ({ciphertext_s1[81], ciphertext_s0[81]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_213 ( .clk (clk), .D ({signal_5727, signal_5719}), .Q ({ciphertext_s1[82], ciphertext_s0[82]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_216 ( .clk (clk), .D ({signal_5743, signal_5735}), .Q ({ciphertext_s1[83], ciphertext_s0[83]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_219 ( .clk (clk), .D ({signal_5759, signal_5751}), .Q ({ciphertext_s1[84], ciphertext_s0[84]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_222 ( .clk (clk), .D ({signal_5775, signal_5767}), .Q ({ciphertext_s1[85], ciphertext_s0[85]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_225 ( .clk (clk), .D ({signal_5791, signal_5783}), .Q ({ciphertext_s1[86], ciphertext_s0[86]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_228 ( .clk (clk), .D ({signal_5807, signal_5799}), .Q ({ciphertext_s1[87], ciphertext_s0[87]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_231 ( .clk (clk), .D ({signal_5823, signal_5815}), .Q ({ciphertext_s1[72], ciphertext_s0[72]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_234 ( .clk (clk), .D ({signal_5839, signal_5831}), .Q ({ciphertext_s1[73], ciphertext_s0[73]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_237 ( .clk (clk), .D ({signal_5855, signal_5847}), .Q ({ciphertext_s1[74], ciphertext_s0[74]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_240 ( .clk (clk), .D ({signal_5871, signal_5863}), .Q ({ciphertext_s1[75], ciphertext_s0[75]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_243 ( .clk (clk), .D ({signal_5887, signal_5879}), .Q ({ciphertext_s1[76], ciphertext_s0[76]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_246 ( .clk (clk), .D ({signal_5903, signal_5895}), .Q ({ciphertext_s1[77], ciphertext_s0[77]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_249 ( .clk (clk), .D ({signal_5919, signal_5911}), .Q ({ciphertext_s1[78], ciphertext_s0[78]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_252 ( .clk (clk), .D ({signal_5935, signal_5927}), .Q ({ciphertext_s1[79], ciphertext_s0[79]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_255 ( .clk (clk), .D ({signal_5951, signal_5943}), .Q ({ciphertext_s1[64], ciphertext_s0[64]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_258 ( .clk (clk), .D ({signal_5967, signal_5959}), .Q ({ciphertext_s1[65], ciphertext_s0[65]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_261 ( .clk (clk), .D ({signal_5983, signal_5975}), .Q ({ciphertext_s1[66], ciphertext_s0[66]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_264 ( .clk (clk), .D ({signal_5999, signal_5991}), .Q ({ciphertext_s1[67], ciphertext_s0[67]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_267 ( .clk (clk), .D ({signal_6015, signal_6007}), .Q ({ciphertext_s1[68], ciphertext_s0[68]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_270 ( .clk (clk), .D ({signal_6031, signal_6023}), .Q ({ciphertext_s1[69], ciphertext_s0[69]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_273 ( .clk (clk), .D ({signal_6047, signal_6039}), .Q ({ciphertext_s1[70], ciphertext_s0[70]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_276 ( .clk (clk), .D ({signal_6063, signal_6055}), .Q ({ciphertext_s1[71], ciphertext_s0[71]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_279 ( .clk (clk), .D ({signal_6079, signal_6071}), .Q ({ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_282 ( .clk (clk), .D ({signal_6095, signal_6087}), .Q ({ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_285 ( .clk (clk), .D ({signal_6111, signal_6103}), .Q ({ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_288 ( .clk (clk), .D ({signal_6127, signal_6119}), .Q ({ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_291 ( .clk (clk), .D ({signal_6143, signal_6135}), .Q ({ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_294 ( .clk (clk), .D ({signal_6159, signal_6151}), .Q ({ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_297 ( .clk (clk), .D ({signal_6175, signal_6167}), .Q ({ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_300 ( .clk (clk), .D ({signal_6191, signal_6183}), .Q ({ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_303 ( .clk (clk), .D ({signal_6207, signal_6199}), .Q ({ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_306 ( .clk (clk), .D ({signal_6223, signal_6215}), .Q ({ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_309 ( .clk (clk), .D ({signal_6239, signal_6231}), .Q ({ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_312 ( .clk (clk), .D ({signal_6255, signal_6247}), .Q ({ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_315 ( .clk (clk), .D ({signal_6271, signal_6263}), .Q ({ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_318 ( .clk (clk), .D ({signal_6287, signal_6279}), .Q ({ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_321 ( .clk (clk), .D ({signal_6303, signal_6295}), .Q ({ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_324 ( .clk (clk), .D ({signal_6319, signal_6311}), .Q ({ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_327 ( .clk (clk), .D ({signal_6335, signal_6327}), .Q ({ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_330 ( .clk (clk), .D ({signal_6351, signal_6343}), .Q ({ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_333 ( .clk (clk), .D ({signal_6367, signal_6359}), .Q ({ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_336 ( .clk (clk), .D ({signal_6383, signal_6375}), .Q ({ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_339 ( .clk (clk), .D ({signal_6399, signal_6391}), .Q ({ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_342 ( .clk (clk), .D ({signal_6415, signal_6407}), .Q ({ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_345 ( .clk (clk), .D ({signal_6431, signal_6423}), .Q ({ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_348 ( .clk (clk), .D ({signal_6447, signal_6439}), .Q ({ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_351 ( .clk (clk), .D ({signal_6463, signal_6455}), .Q ({ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_354 ( .clk (clk), .D ({signal_6479, signal_6471}), .Q ({ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_357 ( .clk (clk), .D ({signal_6495, signal_6487}), .Q ({ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_360 ( .clk (clk), .D ({signal_6511, signal_6503}), .Q ({ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_363 ( .clk (clk), .D ({signal_6527, signal_6519}), .Q ({ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_366 ( .clk (clk), .D ({signal_6543, signal_6535}), .Q ({ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_369 ( .clk (clk), .D ({signal_6559, signal_6551}), .Q ({ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_372 ( .clk (clk), .D ({signal_6575, signal_6567}), .Q ({ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_375 ( .clk (clk), .D ({signal_6591, signal_6583}), .Q ({ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_378 ( .clk (clk), .D ({signal_6607, signal_6599}), .Q ({ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_381 ( .clk (clk), .D ({signal_6623, signal_6615}), .Q ({ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_384 ( .clk (clk), .D ({signal_6639, signal_6631}), .Q ({ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_387 ( .clk (clk), .D ({signal_6655, signal_6647}), .Q ({ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_390 ( .clk (clk), .D ({signal_6671, signal_6663}), .Q ({ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_393 ( .clk (clk), .D ({signal_6687, signal_6679}), .Q ({ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_396 ( .clk (clk), .D ({signal_6703, signal_6695}), .Q ({ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_399 ( .clk (clk), .D ({signal_6719, signal_6711}), .Q ({ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_402 ( .clk (clk), .D ({signal_6735, signal_6727}), .Q ({ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_405 ( .clk (clk), .D ({signal_6751, signal_6743}), .Q ({ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_408 ( .clk (clk), .D ({signal_6767, signal_6759}), .Q ({ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_411 ( .clk (clk), .D ({signal_6783, signal_6775}), .Q ({ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_414 ( .clk (clk), .D ({signal_6799, signal_6791}), .Q ({ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_417 ( .clk (clk), .D ({signal_6815, signal_6807}), .Q ({ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_420 ( .clk (clk), .D ({signal_6831, signal_6823}), .Q ({ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_423 ( .clk (clk), .D ({signal_6847, signal_6839}), .Q ({ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_426 ( .clk (clk), .D ({signal_6863, signal_6855}), .Q ({ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_429 ( .clk (clk), .D ({signal_6879, signal_6871}), .Q ({ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_432 ( .clk (clk), .D ({signal_6895, signal_6887}), .Q ({ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_435 ( .clk (clk), .D ({signal_6911, signal_6903}), .Q ({ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_438 ( .clk (clk), .D ({signal_6927, signal_6919}), .Q ({ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_441 ( .clk (clk), .D ({signal_6943, signal_6935}), .Q ({ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_444 ( .clk (clk), .D ({signal_6959, signal_6951}), .Q ({ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_447 ( .clk (clk), .D ({signal_3637, signal_705}), .Q ({ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_450 ( .clk (clk), .D ({signal_3656, signal_707}), .Q ({ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_453 ( .clk (clk), .D ({signal_3638, signal_709}), .Q ({ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_456 ( .clk (clk), .D ({signal_3639, signal_711}), .Q ({ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_459 ( .clk (clk), .D ({signal_3640, signal_713}), .Q ({ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_462 ( .clk (clk), .D ({signal_3657, signal_715}), .Q ({ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_465 ( .clk (clk), .D ({signal_3658, signal_717}), .Q ({ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_468 ( .clk (clk), .D ({signal_3641, signal_719}), .Q ({ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_717 ( .clk (clk), .D ({signal_6975, signal_6967}), .Q ({signal_2107, signal_1493}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_721 ( .clk (clk), .D ({signal_6991, signal_6983}), .Q ({signal_2110, signal_1492}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_725 ( .clk (clk), .D ({signal_7007, signal_6999}), .Q ({signal_2113, signal_1491}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_729 ( .clk (clk), .D ({signal_7023, signal_7015}), .Q ({signal_2116, signal_1490}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_733 ( .clk (clk), .D ({signal_7039, signal_7031}), .Q ({signal_2119, signal_1489}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_737 ( .clk (clk), .D ({signal_7055, signal_7047}), .Q ({signal_2122, signal_1488}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_741 ( .clk (clk), .D ({signal_7071, signal_7063}), .Q ({signal_2125, signal_1487}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_745 ( .clk (clk), .D ({signal_7087, signal_7079}), .Q ({signal_2128, signal_1486}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_749 ( .clk (clk), .D ({signal_7103, signal_7095}), .Q ({signal_2144, signal_758}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_753 ( .clk (clk), .D ({signal_7119, signal_7111}), .Q ({signal_2142, signal_759}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_757 ( .clk (clk), .D ({signal_7135, signal_7127}), .Q ({signal_2140, signal_760}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_761 ( .clk (clk), .D ({signal_7151, signal_7143}), .Q ({signal_2138, signal_761}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_765 ( .clk (clk), .D ({signal_7167, signal_7159}), .Q ({signal_2136, signal_762}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_769 ( .clk (clk), .D ({signal_7183, signal_7175}), .Q ({signal_2134, signal_763}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_773 ( .clk (clk), .D ({signal_7199, signal_7191}), .Q ({signal_2132, signal_764}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_777 ( .clk (clk), .D ({signal_7215, signal_7207}), .Q ({signal_2130, signal_765}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_781 ( .clk (clk), .D ({signal_7231, signal_7223}), .Q ({signal_2567, signal_1909}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_785 ( .clk (clk), .D ({signal_7247, signal_7239}), .Q ({signal_2570, signal_1908}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_789 ( .clk (clk), .D ({signal_7263, signal_7255}), .Q ({signal_2573, signal_1907}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_793 ( .clk (clk), .D ({signal_7279, signal_7271}), .Q ({signal_2576, signal_1906}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_797 ( .clk (clk), .D ({signal_7295, signal_7287}), .Q ({signal_2579, signal_1905}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_801 ( .clk (clk), .D ({signal_7311, signal_7303}), .Q ({signal_2582, signal_1904}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_805 ( .clk (clk), .D ({signal_7327, signal_7319}), .Q ({signal_2585, signal_1903}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_809 ( .clk (clk), .D ({signal_7343, signal_7335}), .Q ({signal_2588, signal_1902}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_813 ( .clk (clk), .D ({signal_7359, signal_7351}), .Q ({signal_2591, signal_1893}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_817 ( .clk (clk), .D ({signal_7375, signal_7367}), .Q ({signal_2594, signal_1892}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_821 ( .clk (clk), .D ({signal_7391, signal_7383}), .Q ({signal_2597, signal_1891}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_825 ( .clk (clk), .D ({signal_7407, signal_7399}), .Q ({signal_2600, signal_1890}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_829 ( .clk (clk), .D ({signal_7423, signal_7415}), .Q ({signal_2603, signal_1889}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_833 ( .clk (clk), .D ({signal_7439, signal_7431}), .Q ({signal_2606, signal_1888}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_837 ( .clk (clk), .D ({signal_7455, signal_7447}), .Q ({signal_2609, signal_1887}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_841 ( .clk (clk), .D ({signal_7471, signal_7463}), .Q ({signal_2612, signal_1886}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_845 ( .clk (clk), .D ({signal_7487, signal_7479}), .Q ({signal_2615, signal_1877}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_849 ( .clk (clk), .D ({signal_7503, signal_7495}), .Q ({signal_2618, signal_1876}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_853 ( .clk (clk), .D ({signal_7519, signal_7511}), .Q ({signal_2621, signal_1875}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_857 ( .clk (clk), .D ({signal_7535, signal_7527}), .Q ({signal_2624, signal_1874}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_861 ( .clk (clk), .D ({signal_7551, signal_7543}), .Q ({signal_2627, signal_1873}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_865 ( .clk (clk), .D ({signal_7567, signal_7559}), .Q ({signal_2630, signal_1872}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_869 ( .clk (clk), .D ({signal_7583, signal_7575}), .Q ({signal_2633, signal_1871}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_873 ( .clk (clk), .D ({signal_7599, signal_7591}), .Q ({signal_2636, signal_1870}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_877 ( .clk (clk), .D ({signal_7615, signal_7607}), .Q ({signal_2639, signal_1861}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_881 ( .clk (clk), .D ({signal_7631, signal_7623}), .Q ({signal_2642, signal_1860}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_885 ( .clk (clk), .D ({signal_7647, signal_7639}), .Q ({signal_2645, signal_1859}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_889 ( .clk (clk), .D ({signal_7663, signal_7655}), .Q ({signal_2648, signal_1858}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_893 ( .clk (clk), .D ({signal_7679, signal_7671}), .Q ({signal_2651, signal_1857}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_897 ( .clk (clk), .D ({signal_7695, signal_7687}), .Q ({signal_2654, signal_1856}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_901 ( .clk (clk), .D ({signal_7711, signal_7703}), .Q ({signal_2657, signal_1855}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_905 ( .clk (clk), .D ({signal_7727, signal_7719}), .Q ({signal_2660, signal_1854}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_909 ( .clk (clk), .D ({signal_7743, signal_7735}), .Q ({signal_2663, signal_1845}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_913 ( .clk (clk), .D ({signal_7759, signal_7751}), .Q ({signal_2666, signal_1844}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_917 ( .clk (clk), .D ({signal_7775, signal_7767}), .Q ({signal_2669, signal_1843}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_921 ( .clk (clk), .D ({signal_7791, signal_7783}), .Q ({signal_2672, signal_1842}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_925 ( .clk (clk), .D ({signal_7807, signal_7799}), .Q ({signal_2675, signal_1841}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_929 ( .clk (clk), .D ({signal_7823, signal_7815}), .Q ({signal_2678, signal_1840}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_933 ( .clk (clk), .D ({signal_7839, signal_7831}), .Q ({signal_2681, signal_1839}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_937 ( .clk (clk), .D ({signal_7855, signal_7847}), .Q ({signal_2684, signal_1838}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_941 ( .clk (clk), .D ({signal_7871, signal_7863}), .Q ({signal_2687, signal_1509}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_945 ( .clk (clk), .D ({signal_7887, signal_7879}), .Q ({signal_2690, signal_1508}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_949 ( .clk (clk), .D ({signal_7903, signal_7895}), .Q ({signal_2693, signal_1507}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_953 ( .clk (clk), .D ({signal_7919, signal_7911}), .Q ({signal_2696, signal_1506}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_957 ( .clk (clk), .D ({signal_7935, signal_7927}), .Q ({signal_2699, signal_1505}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_961 ( .clk (clk), .D ({signal_7951, signal_7943}), .Q ({signal_2702, signal_1504}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_965 ( .clk (clk), .D ({signal_7967, signal_7959}), .Q ({signal_2705, signal_1503}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_969 ( .clk (clk), .D ({signal_7983, signal_7975}), .Q ({signal_2708, signal_1502}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_973 ( .clk (clk), .D ({signal_7999, signal_7991}), .Q ({signal_2711, signal_1821}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_977 ( .clk (clk), .D ({signal_8015, signal_8007}), .Q ({signal_2714, signal_1820}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_981 ( .clk (clk), .D ({signal_8031, signal_8023}), .Q ({signal_2717, signal_1819}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_985 ( .clk (clk), .D ({signal_8047, signal_8039}), .Q ({signal_2720, signal_1818}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_989 ( .clk (clk), .D ({signal_8063, signal_8055}), .Q ({signal_2723, signal_1817}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_993 ( .clk (clk), .D ({signal_8079, signal_8071}), .Q ({signal_2726, signal_1816}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_997 ( .clk (clk), .D ({signal_8095, signal_8087}), .Q ({signal_2729, signal_1815}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1001 ( .clk (clk), .D ({signal_8111, signal_8103}), .Q ({signal_2732, signal_1814}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1005 ( .clk (clk), .D ({signal_8127, signal_8119}), .Q ({signal_2735, signal_1805}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1009 ( .clk (clk), .D ({signal_8143, signal_8135}), .Q ({signal_2738, signal_1804}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1013 ( .clk (clk), .D ({signal_8159, signal_8151}), .Q ({signal_2741, signal_1803}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1017 ( .clk (clk), .D ({signal_8175, signal_8167}), .Q ({signal_2744, signal_1802}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1021 ( .clk (clk), .D ({signal_8191, signal_8183}), .Q ({signal_2747, signal_1801}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1025 ( .clk (clk), .D ({signal_8207, signal_8199}), .Q ({signal_2750, signal_1800}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1029 ( .clk (clk), .D ({signal_8223, signal_8215}), .Q ({signal_2753, signal_1799}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1033 ( .clk (clk), .D ({signal_8239, signal_8231}), .Q ({signal_2756, signal_1798}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1037 ( .clk (clk), .D ({signal_8255, signal_8247}), .Q ({signal_2759, signal_1789}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1041 ( .clk (clk), .D ({signal_8271, signal_8263}), .Q ({signal_2762, signal_1788}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1045 ( .clk (clk), .D ({signal_8287, signal_8279}), .Q ({signal_2765, signal_1787}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1049 ( .clk (clk), .D ({signal_8303, signal_8295}), .Q ({signal_2768, signal_1786}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1053 ( .clk (clk), .D ({signal_8319, signal_8311}), .Q ({signal_2771, signal_1785}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1057 ( .clk (clk), .D ({signal_8335, signal_8327}), .Q ({signal_2774, signal_1784}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1061 ( .clk (clk), .D ({signal_8351, signal_8343}), .Q ({signal_2777, signal_1783}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1065 ( .clk (clk), .D ({signal_8367, signal_8359}), .Q ({signal_2780, signal_1782}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1069 ( .clk (clk), .D ({signal_8383, signal_8375}), .Q ({signal_2783, signal_1773}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1073 ( .clk (clk), .D ({signal_8399, signal_8391}), .Q ({signal_2786, signal_1772}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1077 ( .clk (clk), .D ({signal_8415, signal_8407}), .Q ({signal_2789, signal_1771}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1081 ( .clk (clk), .D ({signal_8431, signal_8423}), .Q ({signal_2792, signal_1770}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1085 ( .clk (clk), .D ({signal_8447, signal_8439}), .Q ({signal_2795, signal_1769}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1089 ( .clk (clk), .D ({signal_8463, signal_8455}), .Q ({signal_2798, signal_1768}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1093 ( .clk (clk), .D ({signal_8479, signal_8471}), .Q ({signal_2801, signal_1767}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1097 ( .clk (clk), .D ({signal_8495, signal_8487}), .Q ({signal_2804, signal_1766}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1101 ( .clk (clk), .D ({signal_3648, signal_1054}), .Q ({signal_2807, signal_1749}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1105 ( .clk (clk), .D ({signal_3659, signal_1057}), .Q ({signal_2810, signal_1748}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1109 ( .clk (clk), .D ({signal_3650, signal_1060}), .Q ({signal_2813, signal_1747}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1113 ( .clk (clk), .D ({signal_3651, signal_1063}), .Q ({signal_2816, signal_1746}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1117 ( .clk (clk), .D ({signal_3652, signal_1066}), .Q ({signal_2819, signal_1745}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1121 ( .clk (clk), .D ({signal_3660, signal_1069}), .Q ({signal_2822, signal_1744}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1125 ( .clk (clk), .D ({signal_3661, signal_1072}), .Q ({signal_2825, signal_1743}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1129 ( .clk (clk), .D ({signal_3655, signal_1075}), .Q ({signal_2828, signal_1742}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1133 ( .clk (clk), .D ({signal_8511, signal_8503}), .Q ({signal_2831, signal_1733}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1137 ( .clk (clk), .D ({signal_8527, signal_8519}), .Q ({signal_2834, signal_1732}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1141 ( .clk (clk), .D ({signal_8543, signal_8535}), .Q ({signal_2837, signal_1731}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1145 ( .clk (clk), .D ({signal_8559, signal_8551}), .Q ({signal_2840, signal_1730}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1149 ( .clk (clk), .D ({signal_8575, signal_8567}), .Q ({signal_2843, signal_1729}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1153 ( .clk (clk), .D ({signal_8591, signal_8583}), .Q ({signal_2846, signal_1728}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1157 ( .clk (clk), .D ({signal_8607, signal_8599}), .Q ({signal_2849, signal_1727}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1161 ( .clk (clk), .D ({signal_8623, signal_8615}), .Q ({signal_2852, signal_1726}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1165 ( .clk (clk), .D ({signal_8639, signal_8631}), .Q ({signal_2855, signal_1717}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1169 ( .clk (clk), .D ({signal_8655, signal_8647}), .Q ({signal_2858, signal_1716}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1173 ( .clk (clk), .D ({signal_8671, signal_8663}), .Q ({signal_2861, signal_1715}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1177 ( .clk (clk), .D ({signal_8687, signal_8679}), .Q ({signal_2864, signal_1714}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1181 ( .clk (clk), .D ({signal_8703, signal_8695}), .Q ({signal_2867, signal_1713}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1185 ( .clk (clk), .D ({signal_8719, signal_8711}), .Q ({signal_2870, signal_1712}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1189 ( .clk (clk), .D ({signal_8735, signal_8727}), .Q ({signal_2873, signal_1711}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1193 ( .clk (clk), .D ({signal_8751, signal_8743}), .Q ({signal_2876, signal_1710}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1197 ( .clk (clk), .D ({signal_8767, signal_8759}), .Q ({signal_2879, signal_1701}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1201 ( .clk (clk), .D ({signal_8783, signal_8775}), .Q ({signal_2882, signal_1700}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1205 ( .clk (clk), .D ({signal_8799, signal_8791}), .Q ({signal_2885, signal_1699}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1209 ( .clk (clk), .D ({signal_8815, signal_8807}), .Q ({signal_2888, signal_1698}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1213 ( .clk (clk), .D ({signal_8831, signal_8823}), .Q ({signal_2891, signal_1697}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1217 ( .clk (clk), .D ({signal_8847, signal_8839}), .Q ({signal_2894, signal_1696}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1221 ( .clk (clk), .D ({signal_8863, signal_8855}), .Q ({signal_2897, signal_1695}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1225 ( .clk (clk), .D ({signal_8879, signal_8871}), .Q ({signal_2900, signal_1694}) ) ;
    DFF_X1 cell_1561 ( .CK (clk), .D (signal_8887), .Q (signal_1268), .QN () ) ;
    DFF_X1 cell_1563 ( .CK (clk), .D (signal_8895), .Q (signal_1269), .QN () ) ;
    DFF_X1 cell_1565 ( .CK (clk), .D (signal_8903), .Q (signal_1270), .QN () ) ;
    DFF_X1 cell_1567 ( .CK (clk), .D (signal_8911), .Q (signal_1271), .QN () ) ;
    DFF_X1 cell_1569 ( .CK (clk), .D (signal_8919), .Q (signal_1272), .QN () ) ;
    DFF_X1 cell_1571 ( .CK (clk), .D (signal_8927), .Q (signal_1273), .QN () ) ;
    DFF_X1 cell_1573 ( .CK (clk), .D (signal_8935), .Q (signal_1274), .QN () ) ;
    DFF_X1 cell_1575 ( .CK (clk), .D (signal_8943), .Q (signal_1254), .QN () ) ;
    DFF_X1 cell_1713 ( .CK (clk), .D (signal_8951), .Q (signal_393), .QN () ) ;
endmodule
