/* modified netlist. Source: module Midori64 in file /Midori_round_based/AGEMA/Midori64.v */
/* clock gating is added to the circuit, the latency increased 8 time(s)  */

module Midori64_HPC2_ClockGating_d2 (DataIn_s0, key_s0, clk, reset, enc_dec, key_s1, key_s2, DataIn_s1, DataIn_s2, Fresh, DataOut_s0, done, DataOut_s1, DataOut_s2, Synch);
    input [63:0] DataIn_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input reset ;
    input enc_dec ;
    input [127:0] key_s1 ;
    input [127:0] key_s2 ;
    input [63:0] DataIn_s1 ;
    input [63:0] DataIn_s2 ;
    input [767:0] Fresh ;
    output [63:0] DataOut_s0 ;
    output done ;
    output [63:0] DataOut_s1 ;
    output [63:0] DataOut_s2 ;
    output Synch ;
    wire controller_n2 ;
    wire controller_n1 ;
    wire controller_roundCounter_n13 ;
    wire controller_roundCounter_n12 ;
    wire controller_roundCounter_n11 ;
    wire controller_roundCounter_n10 ;
    wire controller_roundCounter_n9 ;
    wire controller_roundCounter_n8 ;
    wire controller_roundCounter_n7 ;
    wire controller_roundCounter_n5 ;
    wire controller_roundCounter_n4 ;
    wire controller_roundCounter_n3 ;
    wire controller_roundCounter_n2 ;
    wire controller_roundCounter_n1 ;
    wire controller_roundCounter_N10 ;
    wire controller_roundCounter_n6 ;
    wire controller_roundCounter_N8 ;
    wire controller_roundCounter_N7 ;
    wire Midori_rounds_n16 ;
    wire Midori_rounds_n15 ;
    wire Midori_rounds_n14 ;
    wire Midori_rounds_n13 ;
    wire Midori_rounds_n12 ;
    wire Midori_rounds_n11 ;
    wire Midori_rounds_n10 ;
    wire Midori_rounds_n9 ;
    wire Midori_rounds_n8 ;
    wire Midori_rounds_n7 ;
    wire Midori_rounds_n6 ;
    wire Midori_rounds_n5 ;
    wire Midori_rounds_n4 ;
    wire Midori_rounds_n3 ;
    wire Midori_rounds_n2 ;
    wire Midori_rounds_n1 ;
    wire Midori_rounds_SelectedKey_0_ ;
    wire Midori_rounds_SelectedKey_1_ ;
    wire Midori_rounds_SelectedKey_2_ ;
    wire Midori_rounds_SelectedKey_3_ ;
    wire Midori_rounds_SelectedKey_4_ ;
    wire Midori_rounds_SelectedKey_5_ ;
    wire Midori_rounds_SelectedKey_6_ ;
    wire Midori_rounds_SelectedKey_7_ ;
    wire Midori_rounds_SelectedKey_8_ ;
    wire Midori_rounds_SelectedKey_9_ ;
    wire Midori_rounds_SelectedKey_10_ ;
    wire Midori_rounds_SelectedKey_11_ ;
    wire Midori_rounds_SelectedKey_12_ ;
    wire Midori_rounds_SelectedKey_13_ ;
    wire Midori_rounds_SelectedKey_14_ ;
    wire Midori_rounds_SelectedKey_15_ ;
    wire Midori_rounds_SelectedKey_16_ ;
    wire Midori_rounds_SelectedKey_17_ ;
    wire Midori_rounds_SelectedKey_18_ ;
    wire Midori_rounds_SelectedKey_19_ ;
    wire Midori_rounds_SelectedKey_20_ ;
    wire Midori_rounds_SelectedKey_21_ ;
    wire Midori_rounds_SelectedKey_22_ ;
    wire Midori_rounds_SelectedKey_23_ ;
    wire Midori_rounds_SelectedKey_24_ ;
    wire Midori_rounds_SelectedKey_25_ ;
    wire Midori_rounds_SelectedKey_26_ ;
    wire Midori_rounds_SelectedKey_27_ ;
    wire Midori_rounds_SelectedKey_28_ ;
    wire Midori_rounds_SelectedKey_29_ ;
    wire Midori_rounds_SelectedKey_30_ ;
    wire Midori_rounds_SelectedKey_31_ ;
    wire Midori_rounds_SelectedKey_32_ ;
    wire Midori_rounds_SelectedKey_33_ ;
    wire Midori_rounds_SelectedKey_34_ ;
    wire Midori_rounds_SelectedKey_35_ ;
    wire Midori_rounds_SelectedKey_36_ ;
    wire Midori_rounds_SelectedKey_37_ ;
    wire Midori_rounds_SelectedKey_38_ ;
    wire Midori_rounds_SelectedKey_39_ ;
    wire Midori_rounds_SelectedKey_40_ ;
    wire Midori_rounds_SelectedKey_41_ ;
    wire Midori_rounds_SelectedKey_42_ ;
    wire Midori_rounds_SelectedKey_43_ ;
    wire Midori_rounds_SelectedKey_44_ ;
    wire Midori_rounds_SelectedKey_45_ ;
    wire Midori_rounds_SelectedKey_46_ ;
    wire Midori_rounds_SelectedKey_47_ ;
    wire Midori_rounds_SelectedKey_48_ ;
    wire Midori_rounds_SelectedKey_49_ ;
    wire Midori_rounds_SelectedKey_50_ ;
    wire Midori_rounds_SelectedKey_51_ ;
    wire Midori_rounds_SelectedKey_52_ ;
    wire Midori_rounds_SelectedKey_53_ ;
    wire Midori_rounds_SelectedKey_54_ ;
    wire Midori_rounds_SelectedKey_55_ ;
    wire Midori_rounds_SelectedKey_56_ ;
    wire Midori_rounds_SelectedKey_57_ ;
    wire Midori_rounds_SelectedKey_58_ ;
    wire Midori_rounds_SelectedKey_59_ ;
    wire Midori_rounds_SelectedKey_60_ ;
    wire Midori_rounds_SelectedKey_61_ ;
    wire Midori_rounds_SelectedKey_62_ ;
    wire Midori_rounds_SelectedKey_63_ ;
    wire Midori_rounds_constant_MUX_n217 ;
    wire Midori_rounds_constant_MUX_n216 ;
    wire Midori_rounds_constant_MUX_n215 ;
    wire Midori_rounds_constant_MUX_n214 ;
    wire Midori_rounds_constant_MUX_n213 ;
    wire Midori_rounds_constant_MUX_n212 ;
    wire Midori_rounds_constant_MUX_n211 ;
    wire Midori_rounds_constant_MUX_n210 ;
    wire Midori_rounds_constant_MUX_n209 ;
    wire Midori_rounds_constant_MUX_n208 ;
    wire Midori_rounds_constant_MUX_n207 ;
    wire Midori_rounds_constant_MUX_n206 ;
    wire Midori_rounds_constant_MUX_n205 ;
    wire Midori_rounds_constant_MUX_n204 ;
    wire Midori_rounds_constant_MUX_n203 ;
    wire Midori_rounds_constant_MUX_n202 ;
    wire Midori_rounds_constant_MUX_n201 ;
    wire Midori_rounds_constant_MUX_n200 ;
    wire Midori_rounds_constant_MUX_n199 ;
    wire Midori_rounds_constant_MUX_n198 ;
    wire Midori_rounds_constant_MUX_n197 ;
    wire Midori_rounds_constant_MUX_n196 ;
    wire Midori_rounds_constant_MUX_n195 ;
    wire Midori_rounds_constant_MUX_n194 ;
    wire Midori_rounds_constant_MUX_n193 ;
    wire Midori_rounds_constant_MUX_n192 ;
    wire Midori_rounds_constant_MUX_n191 ;
    wire Midori_rounds_constant_MUX_n190 ;
    wire Midori_rounds_constant_MUX_n189 ;
    wire Midori_rounds_constant_MUX_n188 ;
    wire Midori_rounds_constant_MUX_n187 ;
    wire Midori_rounds_constant_MUX_n186 ;
    wire Midori_rounds_constant_MUX_n185 ;
    wire Midori_rounds_constant_MUX_n184 ;
    wire Midori_rounds_constant_MUX_n183 ;
    wire Midori_rounds_constant_MUX_n182 ;
    wire Midori_rounds_constant_MUX_n181 ;
    wire Midori_rounds_constant_MUX_n180 ;
    wire Midori_rounds_constant_MUX_n179 ;
    wire Midori_rounds_constant_MUX_n178 ;
    wire Midori_rounds_constant_MUX_n177 ;
    wire Midori_rounds_constant_MUX_n176 ;
    wire Midori_rounds_constant_MUX_n175 ;
    wire Midori_rounds_constant_MUX_n174 ;
    wire Midori_rounds_constant_MUX_n173 ;
    wire Midori_rounds_constant_MUX_n172 ;
    wire Midori_rounds_constant_MUX_n171 ;
    wire Midori_rounds_constant_MUX_n170 ;
    wire Midori_rounds_constant_MUX_n169 ;
    wire Midori_rounds_constant_MUX_n168 ;
    wire Midori_rounds_constant_MUX_n167 ;
    wire Midori_rounds_constant_MUX_n166 ;
    wire Midori_rounds_constant_MUX_n165 ;
    wire Midori_rounds_constant_MUX_n164 ;
    wire Midori_rounds_constant_MUX_n163 ;
    wire Midori_rounds_constant_MUX_n162 ;
    wire Midori_rounds_constant_MUX_n161 ;
    wire Midori_rounds_constant_MUX_n160 ;
    wire Midori_rounds_constant_MUX_n159 ;
    wire Midori_rounds_constant_MUX_n158 ;
    wire Midori_rounds_constant_MUX_n157 ;
    wire Midori_rounds_constant_MUX_n156 ;
    wire Midori_rounds_constant_MUX_n155 ;
    wire Midori_rounds_constant_MUX_n154 ;
    wire Midori_rounds_constant_MUX_n153 ;
    wire Midori_rounds_constant_MUX_n152 ;
    wire Midori_rounds_constant_MUX_n151 ;
    wire Midori_rounds_constant_MUX_n150 ;
    wire Midori_rounds_constant_MUX_n149 ;
    wire Midori_rounds_constant_MUX_n148 ;
    wire Midori_rounds_constant_MUX_n147 ;
    wire Midori_rounds_constant_MUX_n146 ;
    wire Midori_rounds_constant_MUX_n145 ;
    wire Midori_rounds_constant_MUX_n144 ;
    wire Midori_rounds_constant_MUX_n143 ;
    wire Midori_rounds_constant_MUX_n142 ;
    wire Midori_rounds_constant_MUX_n141 ;
    wire Midori_rounds_constant_MUX_n140 ;
    wire Midori_rounds_constant_MUX_n139 ;
    wire Midori_rounds_constant_MUX_n138 ;
    wire Midori_rounds_constant_MUX_n137 ;
    wire Midori_rounds_constant_MUX_n136 ;
    wire Midori_rounds_constant_MUX_n135 ;
    wire Midori_rounds_constant_MUX_n134 ;
    wire Midori_rounds_constant_MUX_n133 ;
    wire Midori_rounds_constant_MUX_n132 ;
    wire Midori_rounds_constant_MUX_n131 ;
    wire Midori_rounds_constant_MUX_n130 ;
    wire Midori_rounds_constant_MUX_n129 ;
    wire Midori_rounds_constant_MUX_n128 ;
    wire Midori_rounds_MUXInst_n11 ;
    wire Midori_rounds_MUXInst_n10 ;
    wire Midori_rounds_MUXInst_n9 ;
    wire Midori_rounds_MUXInst_n8 ;
    wire Midori_rounds_roundResult_Reg_SFF_0_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_1_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_2_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_3_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_4_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_5_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_6_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_7_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_8_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_9_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_10_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_11_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_12_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_13_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_14_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_15_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_16_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_17_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_18_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_19_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_20_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_21_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_22_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_23_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_24_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_25_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_26_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_27_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_28_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_29_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_30_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_31_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_32_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_33_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_34_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_35_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_36_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_37_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_38_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_39_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_40_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_41_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_42_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_43_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_44_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_45_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_46_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_47_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_48_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_49_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_50_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_51_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_52_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_53_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_54_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_55_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_56_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_57_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_58_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_59_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_60_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_61_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_62_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_63_DQ ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n1 ;
    wire Midori_rounds_mul_MC1_n8 ;
    wire Midori_rounds_mul_MC1_n7 ;
    wire Midori_rounds_mul_MC1_n6 ;
    wire Midori_rounds_mul_MC1_n5 ;
    wire Midori_rounds_mul_MC1_n4 ;
    wire Midori_rounds_mul_MC1_n3 ;
    wire Midori_rounds_mul_MC1_n2 ;
    wire Midori_rounds_mul_MC1_n1 ;
    wire Midori_rounds_mul_MC2_n8 ;
    wire Midori_rounds_mul_MC2_n7 ;
    wire Midori_rounds_mul_MC2_n6 ;
    wire Midori_rounds_mul_MC2_n5 ;
    wire Midori_rounds_mul_MC2_n4 ;
    wire Midori_rounds_mul_MC2_n3 ;
    wire Midori_rounds_mul_MC2_n2 ;
    wire Midori_rounds_mul_MC2_n1 ;
    wire Midori_rounds_mul_MC3_n8 ;
    wire Midori_rounds_mul_MC3_n7 ;
    wire Midori_rounds_mul_MC3_n6 ;
    wire Midori_rounds_mul_MC3_n5 ;
    wire Midori_rounds_mul_MC3_n4 ;
    wire Midori_rounds_mul_MC3_n3 ;
    wire Midori_rounds_mul_MC3_n2 ;
    wire Midori_rounds_mul_MC3_n1 ;
    wire Midori_rounds_mul_MC4_n8 ;
    wire Midori_rounds_mul_MC4_n7 ;
    wire Midori_rounds_mul_MC4_n6 ;
    wire Midori_rounds_mul_MC4_n5 ;
    wire Midori_rounds_mul_MC4_n4 ;
    wire Midori_rounds_mul_MC4_n3 ;
    wire Midori_rounds_mul_MC4_n2 ;
    wire Midori_rounds_mul_MC4_n1 ;
    wire [63:0] wk ;
    wire [3:0] round_Signal ;
    wire [63:0] Midori_add_Result_Start ;
    wire [63:0] Midori_rounds_mul_ResultXORkey ;
    wire [63:0] Midori_rounds_SR_Inv_Result ;
    wire [63:0] Midori_rounds_mul_input ;
    wire [63:0] Midori_rounds_sub_ResultXORkey ;
    wire [63:0] Midori_rounds_SR_Result ;
    wire [63:0] Midori_rounds_roundReg_out ;
    wire [63:0] Midori_rounds_round_Result ;
    wire [15:0] Midori_rounds_round_Constant ;
    wire new_AGEMA_signal_1460 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1502 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1520 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1563 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1581 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1593 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1599 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1653 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1701 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1870 ;
    wire new_AGEMA_signal_1871 ;
    wire new_AGEMA_signal_1872 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1880 ;
    wire new_AGEMA_signal_1881 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1888 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1896 ;
    wire new_AGEMA_signal_1897 ;
    wire new_AGEMA_signal_1898 ;
    wire new_AGEMA_signal_1899 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1906 ;
    wire new_AGEMA_signal_1907 ;
    wire new_AGEMA_signal_1908 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1914 ;
    wire new_AGEMA_signal_1915 ;
    wire new_AGEMA_signal_1916 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1923 ;
    wire new_AGEMA_signal_1924 ;
    wire new_AGEMA_signal_1925 ;
    wire new_AGEMA_signal_1926 ;
    wire new_AGEMA_signal_1927 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1931 ;
    wire new_AGEMA_signal_1932 ;
    wire new_AGEMA_signal_1933 ;
    wire new_AGEMA_signal_1934 ;
    wire new_AGEMA_signal_1935 ;
    wire new_AGEMA_signal_1936 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1938 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1940 ;
    wire new_AGEMA_signal_1941 ;
    wire new_AGEMA_signal_1942 ;
    wire new_AGEMA_signal_1943 ;
    wire new_AGEMA_signal_1944 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1947 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1949 ;
    wire new_AGEMA_signal_1950 ;
    wire new_AGEMA_signal_1951 ;
    wire new_AGEMA_signal_1952 ;
    wire new_AGEMA_signal_1953 ;
    wire new_AGEMA_signal_1954 ;
    wire new_AGEMA_signal_1955 ;
    wire new_AGEMA_signal_1956 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1958 ;
    wire new_AGEMA_signal_1959 ;
    wire new_AGEMA_signal_1960 ;
    wire new_AGEMA_signal_1961 ;
    wire new_AGEMA_signal_1962 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1967 ;
    wire new_AGEMA_signal_1968 ;
    wire new_AGEMA_signal_1969 ;
    wire new_AGEMA_signal_1970 ;
    wire new_AGEMA_signal_1971 ;
    wire new_AGEMA_signal_1972 ;
    wire new_AGEMA_signal_1973 ;
    wire new_AGEMA_signal_1974 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1976 ;
    wire new_AGEMA_signal_1977 ;
    wire new_AGEMA_signal_1978 ;
    wire new_AGEMA_signal_1979 ;
    wire new_AGEMA_signal_1980 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1985 ;
    wire new_AGEMA_signal_1986 ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1988 ;
    wire new_AGEMA_signal_1989 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1995 ;
    wire new_AGEMA_signal_1996 ;
    wire new_AGEMA_signal_1997 ;
    wire new_AGEMA_signal_1998 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2003 ;
    wire new_AGEMA_signal_2004 ;
    wire new_AGEMA_signal_2005 ;
    wire new_AGEMA_signal_2006 ;
    wire new_AGEMA_signal_2007 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2014 ;
    wire new_AGEMA_signal_2015 ;
    wire new_AGEMA_signal_2016 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2022 ;
    wire new_AGEMA_signal_2023 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2025 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2032 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2034 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2041 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2043 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2050 ;
    wire new_AGEMA_signal_2051 ;
    wire new_AGEMA_signal_2052 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2059 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2061 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2086 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2097 ;
    wire new_AGEMA_signal_2098 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2102 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2104 ;
    wire new_AGEMA_signal_2105 ;
    wire new_AGEMA_signal_2106 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2114 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2116 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2120 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2124 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2133 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2140 ;
    wire new_AGEMA_signal_2141 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2156 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2160 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2168 ;
    wire new_AGEMA_signal_2169 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2176 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2188 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2205 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2209 ;
    wire new_AGEMA_signal_2212 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2221 ;
    wire new_AGEMA_signal_2224 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2228 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2232 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2236 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2240 ;
    wire new_AGEMA_signal_2241 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2248 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2260 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2264 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2268 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2272 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2276 ;
    wire new_AGEMA_signal_2277 ;
    wire new_AGEMA_signal_2280 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2284 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2296 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2300 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2304 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2308 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2312 ;
    wire new_AGEMA_signal_2313 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2320 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2324 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2332 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2392 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2826 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2914 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2926 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2934 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2942 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2950 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3132 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3139 ;
    wire new_AGEMA_signal_3140 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3248 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3256 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3374 ;
    wire new_AGEMA_signal_3375 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3391 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3411 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3418 ;
    wire new_AGEMA_signal_3419 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3423 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3427 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3447 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3483 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3502 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3561 ;
    wire new_AGEMA_signal_3562 ;
    wire new_AGEMA_signal_3563 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3567 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3569 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3571 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3579 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3583 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3587 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3590 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3615 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3617 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3623 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3634 ;
    wire new_AGEMA_signal_3635 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3659 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_3723 ;
    wire new_AGEMA_signal_3724 ;
    wire new_AGEMA_signal_3725 ;
    wire new_AGEMA_signal_3726 ;
    wire new_AGEMA_signal_3727 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3730 ;
    wire new_AGEMA_signal_3731 ;
    wire new_AGEMA_signal_3732 ;
    wire new_AGEMA_signal_3733 ;
    wire new_AGEMA_signal_3734 ;
    wire new_AGEMA_signal_3735 ;
    wire new_AGEMA_signal_3736 ;
    wire new_AGEMA_signal_3737 ;
    wire new_AGEMA_signal_3738 ;
    wire new_AGEMA_signal_3739 ;
    wire new_AGEMA_signal_3740 ;
    wire new_AGEMA_signal_3741 ;
    wire new_AGEMA_signal_3742 ;
    wire new_AGEMA_signal_3743 ;
    wire new_AGEMA_signal_3744 ;
    wire new_AGEMA_signal_3745 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3747 ;
    wire new_AGEMA_signal_3748 ;
    wire new_AGEMA_signal_3749 ;
    wire new_AGEMA_signal_3750 ;
    wire new_AGEMA_signal_3751 ;
    wire new_AGEMA_signal_3752 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3754 ;
    wire new_AGEMA_signal_3755 ;
    wire new_AGEMA_signal_3756 ;
    wire new_AGEMA_signal_3757 ;
    wire new_AGEMA_signal_3758 ;
    wire new_AGEMA_signal_3759 ;
    wire new_AGEMA_signal_3760 ;
    wire new_AGEMA_signal_3761 ;
    wire new_AGEMA_signal_3762 ;
    wire new_AGEMA_signal_3763 ;
    wire new_AGEMA_signal_3764 ;
    wire new_AGEMA_signal_3765 ;
    wire new_AGEMA_signal_3766 ;
    wire new_AGEMA_signal_3767 ;
    wire new_AGEMA_signal_3768 ;
    wire new_AGEMA_signal_3769 ;
    wire new_AGEMA_signal_3770 ;
    wire new_AGEMA_signal_3771 ;
    wire new_AGEMA_signal_3772 ;
    wire new_AGEMA_signal_3773 ;
    wire new_AGEMA_signal_3774 ;
    wire new_AGEMA_signal_3775 ;
    wire new_AGEMA_signal_3776 ;
    wire new_AGEMA_signal_3777 ;
    wire new_AGEMA_signal_3778 ;
    wire new_AGEMA_signal_3779 ;
    wire new_AGEMA_signal_3780 ;
    wire new_AGEMA_signal_3781 ;
    wire new_AGEMA_signal_3782 ;
    wire new_AGEMA_signal_3783 ;
    wire new_AGEMA_signal_3784 ;
    wire new_AGEMA_signal_3785 ;
    wire new_AGEMA_signal_3786 ;
    wire new_AGEMA_signal_3787 ;
    wire new_AGEMA_signal_3788 ;
    wire new_AGEMA_signal_3789 ;
    wire new_AGEMA_signal_3790 ;
    wire new_AGEMA_signal_3791 ;
    wire new_AGEMA_signal_3792 ;
    wire new_AGEMA_signal_3793 ;
    wire new_AGEMA_signal_3794 ;
    wire new_AGEMA_signal_3795 ;
    wire new_AGEMA_signal_3796 ;
    wire new_AGEMA_signal_3797 ;
    wire new_AGEMA_signal_3798 ;
    wire new_AGEMA_signal_3799 ;
    wire new_AGEMA_signal_3800 ;
    wire new_AGEMA_signal_3801 ;
    wire new_AGEMA_signal_3802 ;
    wire new_AGEMA_signal_3803 ;
    wire new_AGEMA_signal_3804 ;
    wire new_AGEMA_signal_3805 ;
    wire new_AGEMA_signal_3806 ;
    wire new_AGEMA_signal_3807 ;
    wire new_AGEMA_signal_3808 ;
    wire new_AGEMA_signal_3809 ;
    wire new_AGEMA_signal_3810 ;
    wire new_AGEMA_signal_3811 ;
    wire new_AGEMA_signal_3812 ;
    wire new_AGEMA_signal_3813 ;
    wire new_AGEMA_signal_3814 ;
    wire new_AGEMA_signal_3815 ;
    wire new_AGEMA_signal_3816 ;
    wire new_AGEMA_signal_3817 ;
    wire new_AGEMA_signal_3818 ;
    wire new_AGEMA_signal_3819 ;
    wire new_AGEMA_signal_3820 ;
    wire new_AGEMA_signal_3821 ;
    wire new_AGEMA_signal_3822 ;
    wire new_AGEMA_signal_3823 ;
    wire new_AGEMA_signal_3824 ;
    wire new_AGEMA_signal_3825 ;
    wire new_AGEMA_signal_3826 ;
    wire new_AGEMA_signal_3827 ;
    wire new_AGEMA_signal_3828 ;
    wire new_AGEMA_signal_3829 ;
    wire new_AGEMA_signal_3830 ;
    wire new_AGEMA_signal_3831 ;
    wire new_AGEMA_signal_3832 ;
    wire new_AGEMA_signal_3833 ;
    wire new_AGEMA_signal_3834 ;
    wire new_AGEMA_signal_3835 ;
    wire new_AGEMA_signal_3836 ;
    wire new_AGEMA_signal_3837 ;
    wire new_AGEMA_signal_3838 ;
    wire new_AGEMA_signal_3839 ;
    wire new_AGEMA_signal_3840 ;
    wire new_AGEMA_signal_3841 ;
    wire new_AGEMA_signal_3842 ;
    wire new_AGEMA_signal_3843 ;
    wire new_AGEMA_signal_3844 ;
    wire new_AGEMA_signal_3845 ;
    wire new_AGEMA_signal_3846 ;
    wire new_AGEMA_signal_3847 ;
    wire new_AGEMA_signal_3848 ;
    wire new_AGEMA_signal_3849 ;
    wire new_AGEMA_signal_3850 ;
    wire new_AGEMA_signal_3851 ;
    wire new_AGEMA_signal_3852 ;
    wire new_AGEMA_signal_3853 ;
    wire new_AGEMA_signal_3854 ;
    wire new_AGEMA_signal_3855 ;
    wire new_AGEMA_signal_3856 ;
    wire new_AGEMA_signal_3857 ;
    wire new_AGEMA_signal_3858 ;
    wire new_AGEMA_signal_3859 ;
    wire new_AGEMA_signal_3860 ;
    wire new_AGEMA_signal_3861 ;
    wire new_AGEMA_signal_3862 ;
    wire new_AGEMA_signal_3863 ;
    wire new_AGEMA_signal_3864 ;
    wire new_AGEMA_signal_3865 ;
    wire new_AGEMA_signal_3866 ;
    wire new_AGEMA_signal_3867 ;
    wire new_AGEMA_signal_3868 ;
    wire new_AGEMA_signal_3869 ;
    wire new_AGEMA_signal_3870 ;
    wire new_AGEMA_signal_3871 ;
    wire new_AGEMA_signal_3872 ;
    wire new_AGEMA_signal_3873 ;
    wire new_AGEMA_signal_3874 ;
    wire new_AGEMA_signal_3875 ;
    wire new_AGEMA_signal_3876 ;
    wire new_AGEMA_signal_3877 ;
    wire new_AGEMA_signal_3878 ;
    wire new_AGEMA_signal_3879 ;
    wire new_AGEMA_signal_3880 ;
    wire new_AGEMA_signal_3881 ;
    wire new_AGEMA_signal_3882 ;
    wire new_AGEMA_signal_3883 ;
    wire new_AGEMA_signal_3884 ;
    wire new_AGEMA_signal_3885 ;
    wire new_AGEMA_signal_3886 ;
    wire new_AGEMA_signal_3887 ;
    wire new_AGEMA_signal_3888 ;
    wire new_AGEMA_signal_3889 ;
    wire new_AGEMA_signal_3890 ;
    wire new_AGEMA_signal_3891 ;
    wire new_AGEMA_signal_3892 ;
    wire new_AGEMA_signal_3893 ;
    wire new_AGEMA_signal_3894 ;
    wire new_AGEMA_signal_3895 ;
    wire new_AGEMA_signal_3896 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3898 ;
    wire new_AGEMA_signal_3899 ;
    wire new_AGEMA_signal_3900 ;
    wire new_AGEMA_signal_3901 ;
    wire new_AGEMA_signal_3902 ;
    wire new_AGEMA_signal_3903 ;
    wire new_AGEMA_signal_3904 ;
    wire new_AGEMA_signal_3905 ;
    wire new_AGEMA_signal_3906 ;
    wire new_AGEMA_signal_3907 ;
    wire new_AGEMA_signal_3908 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3910 ;
    wire new_AGEMA_signal_3911 ;
    wire new_AGEMA_signal_3912 ;
    wire new_AGEMA_signal_3913 ;
    wire new_AGEMA_signal_3914 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3916 ;
    wire new_AGEMA_signal_3917 ;
    wire new_AGEMA_signal_3918 ;
    wire new_AGEMA_signal_3919 ;
    wire new_AGEMA_signal_3920 ;
    wire new_AGEMA_signal_3921 ;
    wire new_AGEMA_signal_3922 ;
    wire new_AGEMA_signal_3923 ;
    wire new_AGEMA_signal_3924 ;
    wire new_AGEMA_signal_3925 ;
    wire new_AGEMA_signal_3926 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3928 ;
    wire new_AGEMA_signal_3929 ;
    wire new_AGEMA_signal_3930 ;
    wire new_AGEMA_signal_3931 ;
    wire new_AGEMA_signal_3932 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3934 ;
    wire new_AGEMA_signal_3935 ;
    wire new_AGEMA_signal_3936 ;
    wire new_AGEMA_signal_3937 ;
    wire new_AGEMA_signal_3938 ;
    wire new_AGEMA_signal_3939 ;
    wire new_AGEMA_signal_3940 ;
    wire new_AGEMA_signal_3941 ;
    wire new_AGEMA_signal_3942 ;
    wire new_AGEMA_signal_3943 ;
    wire new_AGEMA_signal_3944 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3946 ;
    wire new_AGEMA_signal_3947 ;
    wire new_AGEMA_signal_3948 ;
    wire new_AGEMA_signal_3949 ;
    wire new_AGEMA_signal_3950 ;
    wire new_AGEMA_signal_3951 ;
    wire clk_gated ;

    /* cells in depth 0 */
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U64 ( .a ({key_s2[73], key_s1[73], key_s0[73]}), .b ({key_s2[9], key_s1[9], key_s0[9]}), .c ({new_AGEMA_signal_1461, new_AGEMA_signal_1460, wk[9]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U63 ( .a ({key_s2[72], key_s1[72], key_s0[72]}), .b ({key_s2[8], key_s1[8], key_s0[8]}), .c ({new_AGEMA_signal_1467, new_AGEMA_signal_1466, wk[8]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U62 ( .a ({key_s2[71], key_s1[71], key_s0[71]}), .b ({key_s2[7], key_s1[7], key_s0[7]}), .c ({new_AGEMA_signal_1473, new_AGEMA_signal_1472, wk[7]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U61 ( .a ({key_s2[6], key_s1[6], key_s0[6]}), .b ({key_s2[70], key_s1[70], key_s0[70]}), .c ({new_AGEMA_signal_1479, new_AGEMA_signal_1478, wk[6]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U60 ( .a ({key_s2[127], key_s1[127], key_s0[127]}), .b ({key_s2[63], key_s1[63], key_s0[63]}), .c ({new_AGEMA_signal_1485, new_AGEMA_signal_1484, wk[63]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U59 ( .a ({key_s2[126], key_s1[126], key_s0[126]}), .b ({key_s2[62], key_s1[62], key_s0[62]}), .c ({new_AGEMA_signal_1491, new_AGEMA_signal_1490, wk[62]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U58 ( .a ({key_s2[125], key_s1[125], key_s0[125]}), .b ({key_s2[61], key_s1[61], key_s0[61]}), .c ({new_AGEMA_signal_1497, new_AGEMA_signal_1496, wk[61]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U57 ( .a ({key_s2[124], key_s1[124], key_s0[124]}), .b ({key_s2[60], key_s1[60], key_s0[60]}), .c ({new_AGEMA_signal_1503, new_AGEMA_signal_1502, wk[60]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U56 ( .a ({key_s2[5], key_s1[5], key_s0[5]}), .b ({key_s2[69], key_s1[69], key_s0[69]}), .c ({new_AGEMA_signal_1509, new_AGEMA_signal_1508, wk[5]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U55 ( .a ({key_s2[123], key_s1[123], key_s0[123]}), .b ({key_s2[59], key_s1[59], key_s0[59]}), .c ({new_AGEMA_signal_1515, new_AGEMA_signal_1514, wk[59]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U54 ( .a ({key_s2[122], key_s1[122], key_s0[122]}), .b ({key_s2[58], key_s1[58], key_s0[58]}), .c ({new_AGEMA_signal_1521, new_AGEMA_signal_1520, wk[58]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U53 ( .a ({key_s2[121], key_s1[121], key_s0[121]}), .b ({key_s2[57], key_s1[57], key_s0[57]}), .c ({new_AGEMA_signal_1527, new_AGEMA_signal_1526, wk[57]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U52 ( .a ({key_s2[120], key_s1[120], key_s0[120]}), .b ({key_s2[56], key_s1[56], key_s0[56]}), .c ({new_AGEMA_signal_1533, new_AGEMA_signal_1532, wk[56]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U51 ( .a ({key_s2[119], key_s1[119], key_s0[119]}), .b ({key_s2[55], key_s1[55], key_s0[55]}), .c ({new_AGEMA_signal_1539, new_AGEMA_signal_1538, wk[55]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U50 ( .a ({key_s2[118], key_s1[118], key_s0[118]}), .b ({key_s2[54], key_s1[54], key_s0[54]}), .c ({new_AGEMA_signal_1545, new_AGEMA_signal_1544, wk[54]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U49 ( .a ({key_s2[117], key_s1[117], key_s0[117]}), .b ({key_s2[53], key_s1[53], key_s0[53]}), .c ({new_AGEMA_signal_1551, new_AGEMA_signal_1550, wk[53]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U48 ( .a ({key_s2[116], key_s1[116], key_s0[116]}), .b ({key_s2[52], key_s1[52], key_s0[52]}), .c ({new_AGEMA_signal_1557, new_AGEMA_signal_1556, wk[52]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U47 ( .a ({key_s2[115], key_s1[115], key_s0[115]}), .b ({key_s2[51], key_s1[51], key_s0[51]}), .c ({new_AGEMA_signal_1563, new_AGEMA_signal_1562, wk[51]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U46 ( .a ({key_s2[114], key_s1[114], key_s0[114]}), .b ({key_s2[50], key_s1[50], key_s0[50]}), .c ({new_AGEMA_signal_1569, new_AGEMA_signal_1568, wk[50]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U45 ( .a ({key_s2[4], key_s1[4], key_s0[4]}), .b ({key_s2[68], key_s1[68], key_s0[68]}), .c ({new_AGEMA_signal_1575, new_AGEMA_signal_1574, wk[4]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U44 ( .a ({key_s2[113], key_s1[113], key_s0[113]}), .b ({key_s2[49], key_s1[49], key_s0[49]}), .c ({new_AGEMA_signal_1581, new_AGEMA_signal_1580, wk[49]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U43 ( .a ({key_s2[112], key_s1[112], key_s0[112]}), .b ({key_s2[48], key_s1[48], key_s0[48]}), .c ({new_AGEMA_signal_1587, new_AGEMA_signal_1586, wk[48]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U42 ( .a ({key_s2[111], key_s1[111], key_s0[111]}), .b ({key_s2[47], key_s1[47], key_s0[47]}), .c ({new_AGEMA_signal_1593, new_AGEMA_signal_1592, wk[47]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U41 ( .a ({key_s2[110], key_s1[110], key_s0[110]}), .b ({key_s2[46], key_s1[46], key_s0[46]}), .c ({new_AGEMA_signal_1599, new_AGEMA_signal_1598, wk[46]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U40 ( .a ({key_s2[109], key_s1[109], key_s0[109]}), .b ({key_s2[45], key_s1[45], key_s0[45]}), .c ({new_AGEMA_signal_1605, new_AGEMA_signal_1604, wk[45]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U39 ( .a ({key_s2[108], key_s1[108], key_s0[108]}), .b ({key_s2[44], key_s1[44], key_s0[44]}), .c ({new_AGEMA_signal_1611, new_AGEMA_signal_1610, wk[44]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U38 ( .a ({key_s2[107], key_s1[107], key_s0[107]}), .b ({key_s2[43], key_s1[43], key_s0[43]}), .c ({new_AGEMA_signal_1617, new_AGEMA_signal_1616, wk[43]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U37 ( .a ({key_s2[106], key_s1[106], key_s0[106]}), .b ({key_s2[42], key_s1[42], key_s0[42]}), .c ({new_AGEMA_signal_1623, new_AGEMA_signal_1622, wk[42]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U36 ( .a ({key_s2[105], key_s1[105], key_s0[105]}), .b ({key_s2[41], key_s1[41], key_s0[41]}), .c ({new_AGEMA_signal_1629, new_AGEMA_signal_1628, wk[41]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U35 ( .a ({key_s2[104], key_s1[104], key_s0[104]}), .b ({key_s2[40], key_s1[40], key_s0[40]}), .c ({new_AGEMA_signal_1635, new_AGEMA_signal_1634, wk[40]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U34 ( .a ({key_s2[3], key_s1[3], key_s0[3]}), .b ({key_s2[67], key_s1[67], key_s0[67]}), .c ({new_AGEMA_signal_1641, new_AGEMA_signal_1640, wk[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U33 ( .a ({key_s2[103], key_s1[103], key_s0[103]}), .b ({key_s2[39], key_s1[39], key_s0[39]}), .c ({new_AGEMA_signal_1647, new_AGEMA_signal_1646, wk[39]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U32 ( .a ({key_s2[102], key_s1[102], key_s0[102]}), .b ({key_s2[38], key_s1[38], key_s0[38]}), .c ({new_AGEMA_signal_1653, new_AGEMA_signal_1652, wk[38]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U31 ( .a ({key_s2[101], key_s1[101], key_s0[101]}), .b ({key_s2[37], key_s1[37], key_s0[37]}), .c ({new_AGEMA_signal_1659, new_AGEMA_signal_1658, wk[37]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U30 ( .a ({key_s2[100], key_s1[100], key_s0[100]}), .b ({key_s2[36], key_s1[36], key_s0[36]}), .c ({new_AGEMA_signal_1665, new_AGEMA_signal_1664, wk[36]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U29 ( .a ({key_s2[35], key_s1[35], key_s0[35]}), .b ({key_s2[99], key_s1[99], key_s0[99]}), .c ({new_AGEMA_signal_1671, new_AGEMA_signal_1670, wk[35]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U28 ( .a ({key_s2[34], key_s1[34], key_s0[34]}), .b ({key_s2[98], key_s1[98], key_s0[98]}), .c ({new_AGEMA_signal_1677, new_AGEMA_signal_1676, wk[34]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U27 ( .a ({key_s2[33], key_s1[33], key_s0[33]}), .b ({key_s2[97], key_s1[97], key_s0[97]}), .c ({new_AGEMA_signal_1683, new_AGEMA_signal_1682, wk[33]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U26 ( .a ({key_s2[32], key_s1[32], key_s0[32]}), .b ({key_s2[96], key_s1[96], key_s0[96]}), .c ({new_AGEMA_signal_1689, new_AGEMA_signal_1688, wk[32]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U25 ( .a ({key_s2[31], key_s1[31], key_s0[31]}), .b ({key_s2[95], key_s1[95], key_s0[95]}), .c ({new_AGEMA_signal_1695, new_AGEMA_signal_1694, wk[31]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U24 ( .a ({key_s2[30], key_s1[30], key_s0[30]}), .b ({key_s2[94], key_s1[94], key_s0[94]}), .c ({new_AGEMA_signal_1701, new_AGEMA_signal_1700, wk[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U23 ( .a ({key_s2[2], key_s1[2], key_s0[2]}), .b ({key_s2[66], key_s1[66], key_s0[66]}), .c ({new_AGEMA_signal_1707, new_AGEMA_signal_1706, wk[2]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U22 ( .a ({key_s2[29], key_s1[29], key_s0[29]}), .b ({key_s2[93], key_s1[93], key_s0[93]}), .c ({new_AGEMA_signal_1713, new_AGEMA_signal_1712, wk[29]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U21 ( .a ({key_s2[28], key_s1[28], key_s0[28]}), .b ({key_s2[92], key_s1[92], key_s0[92]}), .c ({new_AGEMA_signal_1719, new_AGEMA_signal_1718, wk[28]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U20 ( .a ({key_s2[27], key_s1[27], key_s0[27]}), .b ({key_s2[91], key_s1[91], key_s0[91]}), .c ({new_AGEMA_signal_1725, new_AGEMA_signal_1724, wk[27]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U19 ( .a ({key_s2[26], key_s1[26], key_s0[26]}), .b ({key_s2[90], key_s1[90], key_s0[90]}), .c ({new_AGEMA_signal_1731, new_AGEMA_signal_1730, wk[26]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U18 ( .a ({key_s2[25], key_s1[25], key_s0[25]}), .b ({key_s2[89], key_s1[89], key_s0[89]}), .c ({new_AGEMA_signal_1737, new_AGEMA_signal_1736, wk[25]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U17 ( .a ({key_s2[24], key_s1[24], key_s0[24]}), .b ({key_s2[88], key_s1[88], key_s0[88]}), .c ({new_AGEMA_signal_1743, new_AGEMA_signal_1742, wk[24]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U16 ( .a ({key_s2[23], key_s1[23], key_s0[23]}), .b ({key_s2[87], key_s1[87], key_s0[87]}), .c ({new_AGEMA_signal_1749, new_AGEMA_signal_1748, wk[23]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U15 ( .a ({key_s2[22], key_s1[22], key_s0[22]}), .b ({key_s2[86], key_s1[86], key_s0[86]}), .c ({new_AGEMA_signal_1755, new_AGEMA_signal_1754, wk[22]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U14 ( .a ({key_s2[21], key_s1[21], key_s0[21]}), .b ({key_s2[85], key_s1[85], key_s0[85]}), .c ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, wk[21]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U13 ( .a ({key_s2[20], key_s1[20], key_s0[20]}), .b ({key_s2[84], key_s1[84], key_s0[84]}), .c ({new_AGEMA_signal_1767, new_AGEMA_signal_1766, wk[20]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U12 ( .a ({key_s2[1], key_s1[1], key_s0[1]}), .b ({key_s2[65], key_s1[65], key_s0[65]}), .c ({new_AGEMA_signal_1773, new_AGEMA_signal_1772, wk[1]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U11 ( .a ({key_s2[19], key_s1[19], key_s0[19]}), .b ({key_s2[83], key_s1[83], key_s0[83]}), .c ({new_AGEMA_signal_1779, new_AGEMA_signal_1778, wk[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U10 ( .a ({key_s2[18], key_s1[18], key_s0[18]}), .b ({key_s2[82], key_s1[82], key_s0[82]}), .c ({new_AGEMA_signal_1785, new_AGEMA_signal_1784, wk[18]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U9 ( .a ({key_s2[17], key_s1[17], key_s0[17]}), .b ({key_s2[81], key_s1[81], key_s0[81]}), .c ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, wk[17]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U8 ( .a ({key_s2[16], key_s1[16], key_s0[16]}), .b ({key_s2[80], key_s1[80], key_s0[80]}), .c ({new_AGEMA_signal_1797, new_AGEMA_signal_1796, wk[16]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U7 ( .a ({key_s2[15], key_s1[15], key_s0[15]}), .b ({key_s2[79], key_s1[79], key_s0[79]}), .c ({new_AGEMA_signal_1803, new_AGEMA_signal_1802, wk[15]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U6 ( .a ({key_s2[14], key_s1[14], key_s0[14]}), .b ({key_s2[78], key_s1[78], key_s0[78]}), .c ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, wk[14]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U5 ( .a ({key_s2[13], key_s1[13], key_s0[13]}), .b ({key_s2[77], key_s1[77], key_s0[77]}), .c ({new_AGEMA_signal_1815, new_AGEMA_signal_1814, wk[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U4 ( .a ({key_s2[12], key_s1[12], key_s0[12]}), .b ({key_s2[76], key_s1[76], key_s0[76]}), .c ({new_AGEMA_signal_1821, new_AGEMA_signal_1820, wk[12]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U3 ( .a ({key_s2[11], key_s1[11], key_s0[11]}), .b ({key_s2[75], key_s1[75], key_s0[75]}), .c ({new_AGEMA_signal_1827, new_AGEMA_signal_1826, wk[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U2 ( .a ({key_s2[10], key_s1[10], key_s0[10]}), .b ({key_s2[74], key_s1[74], key_s0[74]}), .c ({new_AGEMA_signal_1833, new_AGEMA_signal_1832, wk[10]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) keys_U1 ( .a ({key_s2[0], key_s1[0], key_s0[0]}), .b ({key_s2[64], key_s1[64], key_s0[64]}), .c ({new_AGEMA_signal_1839, new_AGEMA_signal_1838, wk[0]}) ) ;
    NOR2_X1 controller_U3 ( .A1 (controller_n2), .A2 (controller_n1), .ZN (done) ) ;
    NAND2_X1 controller_U2 ( .A1 (round_Signal[0]), .A2 (round_Signal[1]), .ZN (controller_n1) ) ;
    NAND2_X1 controller_U1 ( .A1 (round_Signal[2]), .A2 (round_Signal[3]), .ZN (controller_n2) ) ;
    INV_X1 controller_roundCounter_U14 ( .A (controller_roundCounter_n13), .ZN (controller_roundCounter_n2) ) ;
    MUX2_X1 controller_roundCounter_U13 ( .S (controller_roundCounter_n6), .A (controller_roundCounter_n12), .B (controller_roundCounter_n11), .Z (controller_roundCounter_n13) ) ;
    NOR2_X1 controller_roundCounter_U12 ( .A1 (reset), .A2 (controller_roundCounter_n10), .ZN (controller_roundCounter_N8) ) ;
    XNOR2_X1 controller_roundCounter_U11 ( .A (round_Signal[0]), .B (round_Signal[1]), .ZN (controller_roundCounter_n10) ) ;
    MUX2_X1 controller_roundCounter_U10 ( .S (round_Signal[3]), .A (controller_roundCounter_n9), .B (controller_roundCounter_n8), .Z (controller_roundCounter_N10) ) ;
    NAND2_X1 controller_roundCounter_U9 ( .A1 (controller_roundCounter_n12), .A2 (controller_roundCounter_n7), .ZN (controller_roundCounter_n8) ) ;
    NAND2_X1 controller_roundCounter_U8 ( .A1 (controller_roundCounter_n6), .A2 (controller_roundCounter_n3), .ZN (controller_roundCounter_n7) ) ;
    NOR2_X1 controller_roundCounter_U7 ( .A1 (controller_roundCounter_n5), .A2 (controller_roundCounter_N7), .ZN (controller_roundCounter_n12) ) ;
    NOR2_X1 controller_roundCounter_U6 ( .A1 (round_Signal[1]), .A2 (reset), .ZN (controller_roundCounter_n5) ) ;
    NOR2_X1 controller_roundCounter_U5 ( .A1 (controller_roundCounter_n6), .A2 (controller_roundCounter_n11), .ZN (controller_roundCounter_n9) ) ;
    NAND2_X1 controller_roundCounter_U4 ( .A1 (round_Signal[1]), .A2 (controller_roundCounter_n4), .ZN (controller_roundCounter_n11) ) ;
    NOR2_X1 controller_roundCounter_U3 ( .A1 (reset), .A2 (controller_roundCounter_n1), .ZN (controller_roundCounter_n4) ) ;
    NOR2_X1 controller_roundCounter_U2 ( .A1 (reset), .A2 (round_Signal[0]), .ZN (controller_roundCounter_N7) ) ;
    INV_X1 controller_roundCounter_U1 ( .A (reset), .ZN (controller_roundCounter_n3) ) ;
    INV_X1 controller_roundCounter_count_reg_0__U1 ( .A (round_Signal[0]), .ZN (controller_roundCounter_n1) ) ;
    INV_X1 controller_roundCounter_count_reg_2__U1 ( .A (round_Signal[2]), .ZN (controller_roundCounter_n6) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U64 ( .a ({new_AGEMA_signal_1461, new_AGEMA_signal_1460, wk[9]}), .b ({DataIn_s2[9], DataIn_s1[9], DataIn_s0[9]}), .c ({new_AGEMA_signal_2125, new_AGEMA_signal_2124, Midori_add_Result_Start[9]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U63 ( .a ({new_AGEMA_signal_1467, new_AGEMA_signal_1466, wk[8]}), .b ({DataIn_s2[8], DataIn_s1[8], DataIn_s0[8]}), .c ({new_AGEMA_signal_2129, new_AGEMA_signal_2128, Midori_add_Result_Start[8]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U62 ( .a ({new_AGEMA_signal_1473, new_AGEMA_signal_1472, wk[7]}), .b ({DataIn_s2[7], DataIn_s1[7], DataIn_s0[7]}), .c ({new_AGEMA_signal_2133, new_AGEMA_signal_2132, Midori_add_Result_Start[7]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U61 ( .a ({new_AGEMA_signal_1479, new_AGEMA_signal_1478, wk[6]}), .b ({DataIn_s2[6], DataIn_s1[6], DataIn_s0[6]}), .c ({new_AGEMA_signal_2137, new_AGEMA_signal_2136, Midori_add_Result_Start[6]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U60 ( .a ({new_AGEMA_signal_1485, new_AGEMA_signal_1484, wk[63]}), .b ({DataIn_s2[63], DataIn_s1[63], DataIn_s0[63]}), .c ({new_AGEMA_signal_2141, new_AGEMA_signal_2140, Midori_add_Result_Start[63]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U59 ( .a ({new_AGEMA_signal_1491, new_AGEMA_signal_1490, wk[62]}), .b ({DataIn_s2[62], DataIn_s1[62], DataIn_s0[62]}), .c ({new_AGEMA_signal_2145, new_AGEMA_signal_2144, Midori_add_Result_Start[62]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U58 ( .a ({new_AGEMA_signal_1497, new_AGEMA_signal_1496, wk[61]}), .b ({DataIn_s2[61], DataIn_s1[61], DataIn_s0[61]}), .c ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, Midori_add_Result_Start[61]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U57 ( .a ({new_AGEMA_signal_1503, new_AGEMA_signal_1502, wk[60]}), .b ({DataIn_s2[60], DataIn_s1[60], DataIn_s0[60]}), .c ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, Midori_add_Result_Start[60]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U56 ( .a ({new_AGEMA_signal_1509, new_AGEMA_signal_1508, wk[5]}), .b ({DataIn_s2[5], DataIn_s1[5], DataIn_s0[5]}), .c ({new_AGEMA_signal_2157, new_AGEMA_signal_2156, Midori_add_Result_Start[5]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U55 ( .a ({new_AGEMA_signal_1515, new_AGEMA_signal_1514, wk[59]}), .b ({DataIn_s2[59], DataIn_s1[59], DataIn_s0[59]}), .c ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, Midori_add_Result_Start[59]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U54 ( .a ({new_AGEMA_signal_1521, new_AGEMA_signal_1520, wk[58]}), .b ({DataIn_s2[58], DataIn_s1[58], DataIn_s0[58]}), .c ({new_AGEMA_signal_2165, new_AGEMA_signal_2164, Midori_add_Result_Start[58]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U53 ( .a ({new_AGEMA_signal_1527, new_AGEMA_signal_1526, wk[57]}), .b ({DataIn_s2[57], DataIn_s1[57], DataIn_s0[57]}), .c ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, Midori_add_Result_Start[57]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U52 ( .a ({new_AGEMA_signal_1533, new_AGEMA_signal_1532, wk[56]}), .b ({DataIn_s2[56], DataIn_s1[56], DataIn_s0[56]}), .c ({new_AGEMA_signal_2173, new_AGEMA_signal_2172, Midori_add_Result_Start[56]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U51 ( .a ({new_AGEMA_signal_1539, new_AGEMA_signal_1538, wk[55]}), .b ({DataIn_s2[55], DataIn_s1[55], DataIn_s0[55]}), .c ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, Midori_add_Result_Start[55]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U50 ( .a ({new_AGEMA_signal_1545, new_AGEMA_signal_1544, wk[54]}), .b ({DataIn_s2[54], DataIn_s1[54], DataIn_s0[54]}), .c ({new_AGEMA_signal_2181, new_AGEMA_signal_2180, Midori_add_Result_Start[54]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U49 ( .a ({new_AGEMA_signal_1551, new_AGEMA_signal_1550, wk[53]}), .b ({DataIn_s2[53], DataIn_s1[53], DataIn_s0[53]}), .c ({new_AGEMA_signal_2185, new_AGEMA_signal_2184, Midori_add_Result_Start[53]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U48 ( .a ({new_AGEMA_signal_1557, new_AGEMA_signal_1556, wk[52]}), .b ({DataIn_s2[52], DataIn_s1[52], DataIn_s0[52]}), .c ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, Midori_add_Result_Start[52]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U47 ( .a ({new_AGEMA_signal_1563, new_AGEMA_signal_1562, wk[51]}), .b ({DataIn_s2[51], DataIn_s1[51], DataIn_s0[51]}), .c ({new_AGEMA_signal_2193, new_AGEMA_signal_2192, Midori_add_Result_Start[51]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U46 ( .a ({new_AGEMA_signal_1569, new_AGEMA_signal_1568, wk[50]}), .b ({DataIn_s2[50], DataIn_s1[50], DataIn_s0[50]}), .c ({new_AGEMA_signal_2197, new_AGEMA_signal_2196, Midori_add_Result_Start[50]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U45 ( .a ({new_AGEMA_signal_1575, new_AGEMA_signal_1574, wk[4]}), .b ({DataIn_s2[4], DataIn_s1[4], DataIn_s0[4]}), .c ({new_AGEMA_signal_2201, new_AGEMA_signal_2200, Midori_add_Result_Start[4]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U44 ( .a ({new_AGEMA_signal_1581, new_AGEMA_signal_1580, wk[49]}), .b ({DataIn_s2[49], DataIn_s1[49], DataIn_s0[49]}), .c ({new_AGEMA_signal_2205, new_AGEMA_signal_2204, Midori_add_Result_Start[49]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U43 ( .a ({new_AGEMA_signal_1587, new_AGEMA_signal_1586, wk[48]}), .b ({DataIn_s2[48], DataIn_s1[48], DataIn_s0[48]}), .c ({new_AGEMA_signal_2209, new_AGEMA_signal_2208, Midori_add_Result_Start[48]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U42 ( .a ({new_AGEMA_signal_1593, new_AGEMA_signal_1592, wk[47]}), .b ({DataIn_s2[47], DataIn_s1[47], DataIn_s0[47]}), .c ({new_AGEMA_signal_2213, new_AGEMA_signal_2212, Midori_add_Result_Start[47]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U41 ( .a ({new_AGEMA_signal_1599, new_AGEMA_signal_1598, wk[46]}), .b ({DataIn_s2[46], DataIn_s1[46], DataIn_s0[46]}), .c ({new_AGEMA_signal_2217, new_AGEMA_signal_2216, Midori_add_Result_Start[46]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U40 ( .a ({new_AGEMA_signal_1605, new_AGEMA_signal_1604, wk[45]}), .b ({DataIn_s2[45], DataIn_s1[45], DataIn_s0[45]}), .c ({new_AGEMA_signal_2221, new_AGEMA_signal_2220, Midori_add_Result_Start[45]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U39 ( .a ({new_AGEMA_signal_1611, new_AGEMA_signal_1610, wk[44]}), .b ({DataIn_s2[44], DataIn_s1[44], DataIn_s0[44]}), .c ({new_AGEMA_signal_2225, new_AGEMA_signal_2224, Midori_add_Result_Start[44]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U38 ( .a ({new_AGEMA_signal_1617, new_AGEMA_signal_1616, wk[43]}), .b ({DataIn_s2[43], DataIn_s1[43], DataIn_s0[43]}), .c ({new_AGEMA_signal_2229, new_AGEMA_signal_2228, Midori_add_Result_Start[43]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U37 ( .a ({new_AGEMA_signal_1623, new_AGEMA_signal_1622, wk[42]}), .b ({DataIn_s2[42], DataIn_s1[42], DataIn_s0[42]}), .c ({new_AGEMA_signal_2233, new_AGEMA_signal_2232, Midori_add_Result_Start[42]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U36 ( .a ({new_AGEMA_signal_1629, new_AGEMA_signal_1628, wk[41]}), .b ({DataIn_s2[41], DataIn_s1[41], DataIn_s0[41]}), .c ({new_AGEMA_signal_2237, new_AGEMA_signal_2236, Midori_add_Result_Start[41]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U35 ( .a ({new_AGEMA_signal_1635, new_AGEMA_signal_1634, wk[40]}), .b ({DataIn_s2[40], DataIn_s1[40], DataIn_s0[40]}), .c ({new_AGEMA_signal_2241, new_AGEMA_signal_2240, Midori_add_Result_Start[40]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U34 ( .a ({new_AGEMA_signal_1641, new_AGEMA_signal_1640, wk[3]}), .b ({DataIn_s2[3], DataIn_s1[3], DataIn_s0[3]}), .c ({new_AGEMA_signal_2245, new_AGEMA_signal_2244, Midori_add_Result_Start[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U33 ( .a ({new_AGEMA_signal_1647, new_AGEMA_signal_1646, wk[39]}), .b ({DataIn_s2[39], DataIn_s1[39], DataIn_s0[39]}), .c ({new_AGEMA_signal_2249, new_AGEMA_signal_2248, Midori_add_Result_Start[39]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U32 ( .a ({new_AGEMA_signal_1653, new_AGEMA_signal_1652, wk[38]}), .b ({DataIn_s2[38], DataIn_s1[38], DataIn_s0[38]}), .c ({new_AGEMA_signal_2253, new_AGEMA_signal_2252, Midori_add_Result_Start[38]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U31 ( .a ({new_AGEMA_signal_1659, new_AGEMA_signal_1658, wk[37]}), .b ({DataIn_s2[37], DataIn_s1[37], DataIn_s0[37]}), .c ({new_AGEMA_signal_2257, new_AGEMA_signal_2256, Midori_add_Result_Start[37]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U30 ( .a ({new_AGEMA_signal_1665, new_AGEMA_signal_1664, wk[36]}), .b ({DataIn_s2[36], DataIn_s1[36], DataIn_s0[36]}), .c ({new_AGEMA_signal_2261, new_AGEMA_signal_2260, Midori_add_Result_Start[36]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U29 ( .a ({new_AGEMA_signal_1671, new_AGEMA_signal_1670, wk[35]}), .b ({DataIn_s2[35], DataIn_s1[35], DataIn_s0[35]}), .c ({new_AGEMA_signal_2265, new_AGEMA_signal_2264, Midori_add_Result_Start[35]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U28 ( .a ({new_AGEMA_signal_1677, new_AGEMA_signal_1676, wk[34]}), .b ({DataIn_s2[34], DataIn_s1[34], DataIn_s0[34]}), .c ({new_AGEMA_signal_2269, new_AGEMA_signal_2268, Midori_add_Result_Start[34]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U27 ( .a ({new_AGEMA_signal_1683, new_AGEMA_signal_1682, wk[33]}), .b ({DataIn_s2[33], DataIn_s1[33], DataIn_s0[33]}), .c ({new_AGEMA_signal_2273, new_AGEMA_signal_2272, Midori_add_Result_Start[33]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U26 ( .a ({new_AGEMA_signal_1689, new_AGEMA_signal_1688, wk[32]}), .b ({DataIn_s2[32], DataIn_s1[32], DataIn_s0[32]}), .c ({new_AGEMA_signal_2277, new_AGEMA_signal_2276, Midori_add_Result_Start[32]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U25 ( .a ({new_AGEMA_signal_1695, new_AGEMA_signal_1694, wk[31]}), .b ({DataIn_s2[31], DataIn_s1[31], DataIn_s0[31]}), .c ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, Midori_add_Result_Start[31]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U24 ( .a ({new_AGEMA_signal_1701, new_AGEMA_signal_1700, wk[30]}), .b ({DataIn_s2[30], DataIn_s1[30], DataIn_s0[30]}), .c ({new_AGEMA_signal_2285, new_AGEMA_signal_2284, Midori_add_Result_Start[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U23 ( .a ({new_AGEMA_signal_1707, new_AGEMA_signal_1706, wk[2]}), .b ({DataIn_s2[2], DataIn_s1[2], DataIn_s0[2]}), .c ({new_AGEMA_signal_2289, new_AGEMA_signal_2288, Midori_add_Result_Start[2]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U22 ( .a ({new_AGEMA_signal_1713, new_AGEMA_signal_1712, wk[29]}), .b ({DataIn_s2[29], DataIn_s1[29], DataIn_s0[29]}), .c ({new_AGEMA_signal_2293, new_AGEMA_signal_2292, Midori_add_Result_Start[29]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U21 ( .a ({new_AGEMA_signal_1719, new_AGEMA_signal_1718, wk[28]}), .b ({DataIn_s2[28], DataIn_s1[28], DataIn_s0[28]}), .c ({new_AGEMA_signal_2297, new_AGEMA_signal_2296, Midori_add_Result_Start[28]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U20 ( .a ({new_AGEMA_signal_1725, new_AGEMA_signal_1724, wk[27]}), .b ({DataIn_s2[27], DataIn_s1[27], DataIn_s0[27]}), .c ({new_AGEMA_signal_2301, new_AGEMA_signal_2300, Midori_add_Result_Start[27]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U19 ( .a ({new_AGEMA_signal_1731, new_AGEMA_signal_1730, wk[26]}), .b ({DataIn_s2[26], DataIn_s1[26], DataIn_s0[26]}), .c ({new_AGEMA_signal_2305, new_AGEMA_signal_2304, Midori_add_Result_Start[26]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U18 ( .a ({new_AGEMA_signal_1737, new_AGEMA_signal_1736, wk[25]}), .b ({DataIn_s2[25], DataIn_s1[25], DataIn_s0[25]}), .c ({new_AGEMA_signal_2309, new_AGEMA_signal_2308, Midori_add_Result_Start[25]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U17 ( .a ({new_AGEMA_signal_1743, new_AGEMA_signal_1742, wk[24]}), .b ({DataIn_s2[24], DataIn_s1[24], DataIn_s0[24]}), .c ({new_AGEMA_signal_2313, new_AGEMA_signal_2312, Midori_add_Result_Start[24]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U16 ( .a ({new_AGEMA_signal_1749, new_AGEMA_signal_1748, wk[23]}), .b ({DataIn_s2[23], DataIn_s1[23], DataIn_s0[23]}), .c ({new_AGEMA_signal_2317, new_AGEMA_signal_2316, Midori_add_Result_Start[23]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U15 ( .a ({new_AGEMA_signal_1755, new_AGEMA_signal_1754, wk[22]}), .b ({DataIn_s2[22], DataIn_s1[22], DataIn_s0[22]}), .c ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, Midori_add_Result_Start[22]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U14 ( .a ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, wk[21]}), .b ({DataIn_s2[21], DataIn_s1[21], DataIn_s0[21]}), .c ({new_AGEMA_signal_2325, new_AGEMA_signal_2324, Midori_add_Result_Start[21]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U13 ( .a ({new_AGEMA_signal_1767, new_AGEMA_signal_1766, wk[20]}), .b ({DataIn_s2[20], DataIn_s1[20], DataIn_s0[20]}), .c ({new_AGEMA_signal_2329, new_AGEMA_signal_2328, Midori_add_Result_Start[20]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U12 ( .a ({new_AGEMA_signal_1773, new_AGEMA_signal_1772, wk[1]}), .b ({DataIn_s2[1], DataIn_s1[1], DataIn_s0[1]}), .c ({new_AGEMA_signal_2333, new_AGEMA_signal_2332, Midori_add_Result_Start[1]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U11 ( .a ({new_AGEMA_signal_1779, new_AGEMA_signal_1778, wk[19]}), .b ({DataIn_s2[19], DataIn_s1[19], DataIn_s0[19]}), .c ({new_AGEMA_signal_2337, new_AGEMA_signal_2336, Midori_add_Result_Start[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U10 ( .a ({new_AGEMA_signal_1785, new_AGEMA_signal_1784, wk[18]}), .b ({DataIn_s2[18], DataIn_s1[18], DataIn_s0[18]}), .c ({new_AGEMA_signal_2341, new_AGEMA_signal_2340, Midori_add_Result_Start[18]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U9 ( .a ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, wk[17]}), .b ({DataIn_s2[17], DataIn_s1[17], DataIn_s0[17]}), .c ({new_AGEMA_signal_2345, new_AGEMA_signal_2344, Midori_add_Result_Start[17]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U8 ( .a ({new_AGEMA_signal_1797, new_AGEMA_signal_1796, wk[16]}), .b ({DataIn_s2[16], DataIn_s1[16], DataIn_s0[16]}), .c ({new_AGEMA_signal_2349, new_AGEMA_signal_2348, Midori_add_Result_Start[16]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U7 ( .a ({new_AGEMA_signal_1803, new_AGEMA_signal_1802, wk[15]}), .b ({DataIn_s2[15], DataIn_s1[15], DataIn_s0[15]}), .c ({new_AGEMA_signal_2353, new_AGEMA_signal_2352, Midori_add_Result_Start[15]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U6 ( .a ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, wk[14]}), .b ({DataIn_s2[14], DataIn_s1[14], DataIn_s0[14]}), .c ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, Midori_add_Result_Start[14]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U5 ( .a ({new_AGEMA_signal_1815, new_AGEMA_signal_1814, wk[13]}), .b ({DataIn_s2[13], DataIn_s1[13], DataIn_s0[13]}), .c ({new_AGEMA_signal_2361, new_AGEMA_signal_2360, Midori_add_Result_Start[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U4 ( .a ({new_AGEMA_signal_1821, new_AGEMA_signal_1820, wk[12]}), .b ({DataIn_s2[12], DataIn_s1[12], DataIn_s0[12]}), .c ({new_AGEMA_signal_2365, new_AGEMA_signal_2364, Midori_add_Result_Start[12]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U3 ( .a ({new_AGEMA_signal_1827, new_AGEMA_signal_1826, wk[11]}), .b ({DataIn_s2[11], DataIn_s1[11], DataIn_s0[11]}), .c ({new_AGEMA_signal_2369, new_AGEMA_signal_2368, Midori_add_Result_Start[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U2 ( .a ({new_AGEMA_signal_1833, new_AGEMA_signal_1832, wk[10]}), .b ({DataIn_s2[10], DataIn_s1[10], DataIn_s0[10]}), .c ({new_AGEMA_signal_2373, new_AGEMA_signal_2372, Midori_add_Result_Start[10]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U1 ( .a ({new_AGEMA_signal_1839, new_AGEMA_signal_1838, wk[0]}), .b ({DataIn_s2[0], DataIn_s1[0], DataIn_s0[0]}), .c ({new_AGEMA_signal_2377, new_AGEMA_signal_2376, Midori_add_Result_Start[0]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U78 ( .a ({new_AGEMA_signal_1851, new_AGEMA_signal_1850, Midori_rounds_SelectedKey_8_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[2]}), .c ({new_AGEMA_signal_3427, new_AGEMA_signal_3426, Midori_rounds_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U71 ( .a ({new_AGEMA_signal_2665, new_AGEMA_signal_2664, Midori_rounds_SelectedKey_60_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[15]}), .c ({new_AGEMA_signal_3537, new_AGEMA_signal_3536, Midori_rounds_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U65 ( .a ({new_AGEMA_signal_2657, new_AGEMA_signal_2656, Midori_rounds_SelectedKey_56_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[14]}), .c ({new_AGEMA_signal_3539, new_AGEMA_signal_3538, Midori_rounds_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U60 ( .a ({new_AGEMA_signal_2649, new_AGEMA_signal_2648, Midori_rounds_SelectedKey_52_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[13]}), .c ({new_AGEMA_signal_3541, new_AGEMA_signal_3540, Midori_rounds_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U56 ( .a ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, Midori_rounds_SelectedKey_4_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[1]}), .c ({new_AGEMA_signal_3543, new_AGEMA_signal_3542, Midori_rounds_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U53 ( .a ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, Midori_rounds_SelectedKey_48_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[12]}), .c ({new_AGEMA_signal_3781, new_AGEMA_signal_3780, Midori_rounds_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U48 ( .a ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, Midori_rounds_SelectedKey_44_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[11]}), .c ({new_AGEMA_signal_3465, new_AGEMA_signal_3464, Midori_rounds_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U43 ( .a ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, Midori_rounds_SelectedKey_40_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[10]}), .c ({new_AGEMA_signal_3545, new_AGEMA_signal_3544, Midori_rounds_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U37 ( .a ({new_AGEMA_signal_2617, new_AGEMA_signal_2616, Midori_rounds_SelectedKey_36_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[9]}), .c ({new_AGEMA_signal_3481, new_AGEMA_signal_3480, Midori_rounds_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U32 ( .a ({new_AGEMA_signal_2609, new_AGEMA_signal_2608, Midori_rounds_SelectedKey_32_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[8]}), .c ({new_AGEMA_signal_3547, new_AGEMA_signal_3546, Midori_rounds_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U26 ( .a ({new_AGEMA_signal_2601, new_AGEMA_signal_2600, Midori_rounds_SelectedKey_28_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[7]}), .c ({new_AGEMA_signal_3673, new_AGEMA_signal_3672, Midori_rounds_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U21 ( .a ({new_AGEMA_signal_2595, new_AGEMA_signal_2594, Midori_rounds_SelectedKey_24_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[6]}), .c ({new_AGEMA_signal_3549, new_AGEMA_signal_3548, Midori_rounds_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U16 ( .a ({new_AGEMA_signal_2587, new_AGEMA_signal_2586, Midori_rounds_SelectedKey_20_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[5]}), .c ({new_AGEMA_signal_3509, new_AGEMA_signal_3508, Midori_rounds_n4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U10 ( .a ({new_AGEMA_signal_2579, new_AGEMA_signal_2578, Midori_rounds_SelectedKey_16_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[4]}), .c ({new_AGEMA_signal_3551, new_AGEMA_signal_3550, Midori_rounds_n3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U5 ( .a ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, Midori_rounds_SelectedKey_12_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[3]}), .c ({new_AGEMA_signal_3553, new_AGEMA_signal_3552, Midori_rounds_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U1 ( .a ({new_AGEMA_signal_1841, new_AGEMA_signal_1840, Midori_rounds_SelectedKey_0_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[0]}), .c ({new_AGEMA_signal_3555, new_AGEMA_signal_3554, Midori_rounds_n1}) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U106 ( .A1 (Midori_rounds_constant_MUX_n217), .A2 (Midori_rounds_constant_MUX_n216), .ZN (Midori_rounds_round_Constant[9]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U105 ( .A1 (Midori_rounds_constant_MUX_n215), .A2 (Midori_rounds_constant_MUX_n214), .ZN (Midori_rounds_constant_MUX_n217) ) ;
    OR2_X1 Midori_rounds_constant_MUX_U104 ( .A1 (Midori_rounds_constant_MUX_n213), .A2 (Midori_rounds_constant_MUX_n212), .ZN (Midori_rounds_constant_MUX_n214) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U103 ( .A1 (Midori_rounds_constant_MUX_n211), .A2 (Midori_rounds_constant_MUX_n210), .ZN (Midori_rounds_round_Constant[8]) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U102 ( .A1 (Midori_rounds_constant_MUX_n209), .A2 (Midori_rounds_constant_MUX_n208), .ZN (Midori_rounds_round_Constant[7]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U101 ( .A1 (Midori_rounds_round_Constant[11]), .A2 (Midori_rounds_constant_MUX_n207), .ZN (Midori_rounds_constant_MUX_n208) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U100 ( .A1 (Midori_rounds_constant_MUX_n206), .A2 (Midori_rounds_constant_MUX_n205), .ZN (Midori_rounds_constant_MUX_n207) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U99 ( .A1 (Midori_rounds_constant_MUX_n204), .A2 (Midori_rounds_constant_MUX_n203), .ZN (Midori_rounds_constant_MUX_n206) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U98 ( .A1 (Midori_rounds_constant_MUX_n202), .A2 (Midori_rounds_constant_MUX_n201), .ZN (Midori_rounds_round_Constant[6]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U97 ( .A1 (Midori_rounds_constant_MUX_n200), .A2 (Midori_rounds_constant_MUX_n199), .ZN (Midori_rounds_constant_MUX_n201) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U96 ( .A1 (Midori_rounds_constant_MUX_n198), .A2 (Midori_rounds_constant_MUX_n197), .ZN (Midori_rounds_round_Constant[5]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U95 ( .A1 (Midori_rounds_constant_MUX_n212), .A2 (Midori_rounds_constant_MUX_n196), .ZN (Midori_rounds_constant_MUX_n197) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U94 ( .A1 (Midori_rounds_constant_MUX_n195), .A2 (Midori_rounds_constant_MUX_n205), .ZN (Midori_rounds_constant_MUX_n196) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U93 ( .A1 (Midori_rounds_constant_MUX_n194), .A2 (Midori_rounds_constant_MUX_n195), .ZN (Midori_rounds_round_Constant[4]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U92 ( .A1 (Midori_rounds_constant_MUX_n193), .A2 (Midori_rounds_constant_MUX_n192), .ZN (Midori_rounds_constant_MUX_n195) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U91 ( .A1 (Midori_rounds_constant_MUX_n191), .A2 (Midori_rounds_constant_MUX_n190), .ZN (Midori_rounds_round_Constant[3]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U90 ( .A1 (Midori_rounds_constant_MUX_n215), .A2 (Midori_rounds_constant_MUX_n189), .ZN (Midori_rounds_constant_MUX_n191) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U89 ( .A1 (Midori_rounds_constant_MUX_n188), .A2 (Midori_rounds_constant_MUX_n205), .ZN (Midori_rounds_constant_MUX_n189) ) ;
    INV_X1 Midori_rounds_constant_MUX_U88 ( .A (Midori_rounds_constant_MUX_n187), .ZN (Midori_rounds_constant_MUX_n188) ) ;
    OR2_X1 Midori_rounds_constant_MUX_U87 ( .A1 (Midori_rounds_constant_MUX_n215), .A2 (Midori_rounds_constant_MUX_n186), .ZN (Midori_rounds_round_Constant[2]) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U86 ( .A1 (Midori_rounds_constant_MUX_n202), .A2 (Midori_rounds_constant_MUX_n185), .ZN (Midori_rounds_constant_MUX_n186) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U85 ( .A1 (Midori_rounds_constant_MUX_n184), .A2 (Midori_rounds_constant_MUX_n212), .ZN (Midori_rounds_constant_MUX_n202) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U84 ( .A1 (Midori_rounds_constant_MUX_n183), .A2 (Midori_rounds_constant_MUX_n210), .ZN (Midori_rounds_constant_MUX_n215) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U83 ( .A1 (Midori_rounds_constant_MUX_n182), .A2 (Midori_rounds_constant_MUX_n181), .ZN (Midori_rounds_round_Constant[1]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U82 ( .A1 (Midori_rounds_constant_MUX_n187), .A2 (Midori_rounds_constant_MUX_n180), .ZN (Midori_rounds_constant_MUX_n181) ) ;
    OR2_X1 Midori_rounds_constant_MUX_U81 ( .A1 (Midori_rounds_constant_MUX_n212), .A2 (Midori_rounds_constant_MUX_n204), .ZN (Midori_rounds_constant_MUX_n180) ) ;
    INV_X1 Midori_rounds_constant_MUX_U80 ( .A (Midori_rounds_constant_MUX_n183), .ZN (Midori_rounds_constant_MUX_n204) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U79 ( .A1 (Midori_rounds_constant_MUX_n179), .A2 (Midori_rounds_constant_MUX_n178), .ZN (Midori_rounds_constant_MUX_n183) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U78 ( .A1 (Midori_rounds_constant_MUX_n177), .A2 (Midori_rounds_constant_MUX_n176), .ZN (Midori_rounds_constant_MUX_n178) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U77 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n175), .ZN (Midori_rounds_constant_MUX_n212) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U76 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n174), .B (Midori_rounds_constant_MUX_n173), .Z (Midori_rounds_constant_MUX_n175) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U75 ( .A1 (Midori_rounds_constant_MUX_n172), .A2 (Midori_rounds_constant_MUX_n171), .ZN (Midori_rounds_round_Constant[15]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U74 ( .A1 (Midori_rounds_constant_MUX_n200), .A2 (Midori_rounds_constant_MUX_n187), .ZN (Midori_rounds_constant_MUX_n172) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U73 ( .A1 (Midori_rounds_constant_MUX_n170), .A2 (Midori_rounds_constant_MUX_n194), .ZN (Midori_rounds_round_Constant[14]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U72 ( .A1 (Midori_rounds_constant_MUX_n169), .A2 (Midori_rounds_constant_MUX_n168), .ZN (Midori_rounds_constant_MUX_n194) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U71 ( .A1 (Midori_rounds_constant_MUX_n216), .A2 (Midori_rounds_constant_MUX_n205), .ZN (Midori_rounds_constant_MUX_n168) ) ;
    OR2_X1 Midori_rounds_constant_MUX_U70 ( .A1 (Midori_rounds_constant_MUX_n129), .A2 (Midori_rounds_constant_MUX_n167), .ZN (Midori_rounds_constant_MUX_n205) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U69 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n166), .B (Midori_rounds_constant_MUX_n165), .Z (Midori_rounds_constant_MUX_n167) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U68 ( .A1 (Midori_rounds_constant_MUX_n185), .A2 (Midori_rounds_constant_MUX_n164), .ZN (Midori_rounds_round_Constant[13]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U67 ( .A1 (Midori_rounds_constant_MUX_n163), .A2 (Midori_rounds_constant_MUX_n162), .ZN (Midori_rounds_constant_MUX_n164) ) ;
    INV_X1 Midori_rounds_constant_MUX_U66 ( .A (Midori_rounds_constant_MUX_n170), .ZN (Midori_rounds_constant_MUX_n162) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U65 ( .A1 (Midori_rounds_constant_MUX_n161), .A2 (Midori_rounds_constant_MUX_n192), .ZN (Midori_rounds_constant_MUX_n185) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U64 ( .A1 (Midori_rounds_constant_MUX_n160), .A2 (Midori_rounds_constant_MUX_n190), .ZN (Midori_rounds_round_Constant[12]) ) ;
    INV_X1 Midori_rounds_constant_MUX_U63 ( .A (Midori_rounds_constant_MUX_n184), .ZN (Midori_rounds_constant_MUX_n190) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U62 ( .A1 (Midori_rounds_constant_MUX_n203), .A2 (Midori_rounds_constant_MUX_n159), .ZN (Midori_rounds_constant_MUX_n160) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U61 ( .A1 (Midori_rounds_constant_MUX_n211), .A2 (Midori_rounds_constant_MUX_n170), .ZN (Midori_rounds_constant_MUX_n159) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U60 ( .A1 (Midori_rounds_constant_MUX_n193), .A2 (Midori_rounds_constant_MUX_n169), .ZN (Midori_rounds_constant_MUX_n211) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U59 ( .A1 (Midori_rounds_constant_MUX_n198), .A2 (Midori_rounds_constant_MUX_n158), .ZN (Midori_rounds_constant_MUX_n169) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U58 ( .A1 (Midori_rounds_constant_MUX_n129), .A2 (Midori_rounds_constant_MUX_n157), .ZN (Midori_rounds_constant_MUX_n158) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U57 ( .A1 (Midori_rounds_constant_MUX_n165), .A2 (Midori_rounds_constant_MUX_n177), .ZN (Midori_rounds_constant_MUX_n157) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U56 ( .A1 (Midori_rounds_constant_MUX_n200), .A2 (Midori_rounds_constant_MUX_n156), .ZN (Midori_rounds_constant_MUX_n198) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U55 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n155), .ZN (Midori_rounds_constant_MUX_n156) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U54 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n176), .B (Midori_rounds_constant_MUX_n166), .Z (Midori_rounds_constant_MUX_n155) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U53 ( .A1 (Midori_rounds_constant_MUX_n129), .A2 (Midori_rounds_constant_MUX_n154), .ZN (Midori_rounds_constant_MUX_n200) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U52 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n174), .B (Midori_rounds_constant_MUX_n153), .Z (Midori_rounds_constant_MUX_n154) ) ;
    OR2_X1 Midori_rounds_constant_MUX_U51 ( .A1 (Midori_rounds_constant_MUX_n199), .A2 (Midori_rounds_constant_MUX_n213), .ZN (Midori_rounds_round_Constant[11]) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U50 ( .A1 (Midori_rounds_constant_MUX_n170), .A2 (Midori_rounds_constant_MUX_n210), .ZN (Midori_rounds_constant_MUX_n199) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U49 ( .A1 (Midori_rounds_constant_MUX_n152), .A2 (Midori_rounds_constant_MUX_n151), .ZN (Midori_rounds_constant_MUX_n210) ) ;
    AND2_X1 Midori_rounds_constant_MUX_U48 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (round_Signal[2]), .ZN (Midori_rounds_constant_MUX_n151) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U47 ( .A1 (Midori_rounds_constant_MUX_n150), .A2 (Midori_rounds_constant_MUX_n187), .ZN (Midori_rounds_constant_MUX_n170) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U46 ( .A1 (Midori_rounds_constant_MUX_n129), .A2 (Midori_rounds_constant_MUX_n149), .ZN (Midori_rounds_constant_MUX_n187) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U45 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n165), .B (Midori_rounds_constant_MUX_n166), .Z (Midori_rounds_constant_MUX_n149) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U44 ( .A1 (Midori_rounds_constant_MUX_n129), .A2 (Midori_rounds_constant_MUX_n148), .ZN (Midori_rounds_constant_MUX_n150) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U43 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n153), .B (Midori_rounds_constant_MUX_n174), .Z (Midori_rounds_constant_MUX_n148) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U42 ( .A1 (Midori_rounds_constant_MUX_n147), .A2 (Midori_rounds_constant_MUX_n171), .ZN (Midori_rounds_round_Constant[10]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U41 ( .A1 (Midori_rounds_constant_MUX_n146), .A2 (Midori_rounds_constant_MUX_n213), .ZN (Midori_rounds_constant_MUX_n171) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U40 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n145), .ZN (Midori_rounds_constant_MUX_n213) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U39 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n165), .B (Midori_rounds_constant_MUX_n177), .Z (Midori_rounds_constant_MUX_n145) ) ;
    INV_X1 Midori_rounds_constant_MUX_U38 ( .A (Midori_rounds_constant_MUX_n144), .ZN (Midori_rounds_constant_MUX_n146) ) ;
    INV_X1 Midori_rounds_constant_MUX_U37 ( .A (Midori_rounds_constant_MUX_n193), .ZN (Midori_rounds_constant_MUX_n147) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U36 ( .A1 (Midori_rounds_constant_MUX_n182), .A2 (Midori_rounds_constant_MUX_n144), .ZN (Midori_rounds_round_Constant[0]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U35 ( .A1 (Midori_rounds_constant_MUX_n203), .A2 (Midori_rounds_constant_MUX_n192), .ZN (Midori_rounds_constant_MUX_n144) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U34 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n143), .ZN (Midori_rounds_constant_MUX_n192) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U33 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n173), .B (Midori_rounds_constant_MUX_n174), .Z (Midori_rounds_constant_MUX_n143) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U32 ( .A1 (Midori_rounds_constant_MUX_n142), .A2 (Midori_rounds_constant_MUX_n141), .ZN (Midori_rounds_constant_MUX_n174) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U31 ( .A1 (Midori_rounds_constant_MUX_n140), .A2 (round_Signal[1]), .ZN (Midori_rounds_constant_MUX_n173) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U30 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n139), .ZN (Midori_rounds_constant_MUX_n203) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U29 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n166), .B (Midori_rounds_constant_MUX_n176), .Z (Midori_rounds_constant_MUX_n139) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U28 ( .A1 (enc_dec), .A2 (Midori_rounds_constant_MUX_n152), .ZN (Midori_rounds_constant_MUX_n176) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U27 ( .A1 (round_Signal[3]), .A2 (Midori_rounds_constant_MUX_n141), .ZN (Midori_rounds_constant_MUX_n152) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U26 ( .A1 (Midori_rounds_constant_MUX_n138), .A2 (Midori_rounds_constant_MUX_n141), .ZN (Midori_rounds_constant_MUX_n166) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U25 ( .A1 (Midori_rounds_constant_MUX_n184), .A2 (Midori_rounds_constant_MUX_n137), .ZN (Midori_rounds_constant_MUX_n182) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U24 ( .A1 (Midori_rounds_constant_MUX_n209), .A2 (Midori_rounds_constant_MUX_n216), .ZN (Midori_rounds_constant_MUX_n137) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U23 ( .A1 (Midori_rounds_constant_MUX_n163), .A2 (Midori_rounds_constant_MUX_n136), .ZN (Midori_rounds_constant_MUX_n216) ) ;
    OR2_X1 Midori_rounds_constant_MUX_U22 ( .A1 (Midori_rounds_constant_MUX_n140), .A2 (Midori_rounds_constant_MUX_n142), .ZN (Midori_rounds_constant_MUX_n136) ) ;
    AND2_X1 Midori_rounds_constant_MUX_U21 ( .A1 (round_Signal[1]), .A2 (Midori_rounds_constant_MUX_n179), .ZN (Midori_rounds_constant_MUX_n163) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U20 ( .A1 (Midori_rounds_constant_MUX_n129), .A2 (round_Signal[2]), .ZN (Midori_rounds_constant_MUX_n179) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U19 ( .A1 (Midori_rounds_constant_MUX_n193), .A2 (Midori_rounds_constant_MUX_n161), .ZN (Midori_rounds_constant_MUX_n209) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U18 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n135), .ZN (Midori_rounds_constant_MUX_n161) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U17 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n177), .B (Midori_rounds_constant_MUX_n165), .Z (Midori_rounds_constant_MUX_n135) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U16 ( .A1 (enc_dec), .A2 (Midori_rounds_constant_MUX_n134), .ZN (Midori_rounds_constant_MUX_n165) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U15 ( .A1 (round_Signal[3]), .A2 (round_Signal[1]), .ZN (Midori_rounds_constant_MUX_n134) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U14 ( .A1 (round_Signal[1]), .A2 (Midori_rounds_constant_MUX_n138), .ZN (Midori_rounds_constant_MUX_n177) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U13 ( .A1 (enc_dec), .A2 (Midori_rounds_constant_MUX_n133), .ZN (Midori_rounds_constant_MUX_n138) ) ;
    INV_X1 Midori_rounds_constant_MUX_U12 ( .A (round_Signal[3]), .ZN (Midori_rounds_constant_MUX_n133) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U11 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n132), .ZN (Midori_rounds_constant_MUX_n193) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U10 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n153), .B (Midori_rounds_constant_MUX_n131), .Z (Midori_rounds_constant_MUX_n132) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U9 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n130), .ZN (Midori_rounds_constant_MUX_n184) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U8 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n131), .B (Midori_rounds_constant_MUX_n153), .Z (Midori_rounds_constant_MUX_n130) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U7 ( .A1 (Midori_rounds_constant_MUX_n140), .A2 (Midori_rounds_constant_MUX_n141), .ZN (Midori_rounds_constant_MUX_n153) ) ;
    INV_X1 Midori_rounds_constant_MUX_U6 ( .A (round_Signal[1]), .ZN (Midori_rounds_constant_MUX_n141) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U5 ( .A1 (enc_dec), .A2 (round_Signal[3]), .ZN (Midori_rounds_constant_MUX_n140) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U4 ( .A1 (Midori_rounds_constant_MUX_n142), .A2 (round_Signal[1]), .ZN (Midori_rounds_constant_MUX_n131) ) ;
    AND2_X1 Midori_rounds_constant_MUX_U3 ( .A1 (enc_dec), .A2 (round_Signal[3]), .ZN (Midori_rounds_constant_MUX_n142) ) ;
    INV_X1 Midori_rounds_constant_MUX_U2 ( .A (Midori_rounds_constant_MUX_n129), .ZN (Midori_rounds_constant_MUX_n128) ) ;
    INV_X1 Midori_rounds_constant_MUX_U1 ( .A (round_Signal[0]), .ZN (Midori_rounds_constant_MUX_n129) ) ;
    INV_X1 Midori_rounds_MUXInst_U4 ( .A (round_Signal[0]), .ZN (Midori_rounds_MUXInst_n11) ) ;
    INV_X1 Midori_rounds_MUXInst_U3 ( .A (Midori_rounds_MUXInst_n11), .ZN (Midori_rounds_MUXInst_n8) ) ;
    INV_X1 Midori_rounds_MUXInst_U2 ( .A (Midori_rounds_MUXInst_n11), .ZN (Midori_rounds_MUXInst_n9) ) ;
    INV_X1 Midori_rounds_MUXInst_U1 ( .A (Midori_rounds_MUXInst_n11), .ZN (Midori_rounds_MUXInst_n10) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_0_U1 ( .s (round_Signal[0]), .b ({key_s2[64], key_s1[64], key_s0[64]}), .a ({key_s2[0], key_s1[0], key_s0[0]}), .c ({new_AGEMA_signal_1841, new_AGEMA_signal_1840, Midori_rounds_SelectedKey_0_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_1_U1 ( .s (round_Signal[0]), .b ({key_s2[65], key_s1[65], key_s0[65]}), .a ({key_s2[1], key_s1[1], key_s0[1]}), .c ({new_AGEMA_signal_1843, new_AGEMA_signal_1842, Midori_rounds_SelectedKey_1_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_2_U1 ( .s (round_Signal[0]), .b ({key_s2[66], key_s1[66], key_s0[66]}), .a ({key_s2[2], key_s1[2], key_s0[2]}), .c ({new_AGEMA_signal_1845, new_AGEMA_signal_1844, Midori_rounds_SelectedKey_2_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_3_U1 ( .s (round_Signal[0]), .b ({key_s2[67], key_s1[67], key_s0[67]}), .a ({key_s2[3], key_s1[3], key_s0[3]}), .c ({new_AGEMA_signal_1847, new_AGEMA_signal_1846, Midori_rounds_SelectedKey_3_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_4_U1 ( .s (round_Signal[0]), .b ({key_s2[68], key_s1[68], key_s0[68]}), .a ({key_s2[4], key_s1[4], key_s0[4]}), .c ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, Midori_rounds_SelectedKey_4_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_5_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[69], key_s1[69], key_s0[69]}), .a ({key_s2[5], key_s1[5], key_s0[5]}), .c ({new_AGEMA_signal_2571, new_AGEMA_signal_2570, Midori_rounds_SelectedKey_5_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_6_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[70], key_s1[70], key_s0[70]}), .a ({key_s2[6], key_s1[6], key_s0[6]}), .c ({new_AGEMA_signal_2573, new_AGEMA_signal_2572, Midori_rounds_SelectedKey_6_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_7_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[71], key_s1[71], key_s0[71]}), .a ({key_s2[7], key_s1[7], key_s0[7]}), .c ({new_AGEMA_signal_2575, new_AGEMA_signal_2574, Midori_rounds_SelectedKey_7_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_8_U1 ( .s (round_Signal[0]), .b ({key_s2[72], key_s1[72], key_s0[72]}), .a ({key_s2[8], key_s1[8], key_s0[8]}), .c ({new_AGEMA_signal_1851, new_AGEMA_signal_1850, Midori_rounds_SelectedKey_8_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_9_U1 ( .s (round_Signal[0]), .b ({key_s2[73], key_s1[73], key_s0[73]}), .a ({key_s2[9], key_s1[9], key_s0[9]}), .c ({new_AGEMA_signal_1853, new_AGEMA_signal_1852, Midori_rounds_SelectedKey_9_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_10_U1 ( .s (round_Signal[0]), .b ({key_s2[74], key_s1[74], key_s0[74]}), .a ({key_s2[10], key_s1[10], key_s0[10]}), .c ({new_AGEMA_signal_1855, new_AGEMA_signal_1854, Midori_rounds_SelectedKey_10_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_11_U1 ( .s (round_Signal[0]), .b ({key_s2[75], key_s1[75], key_s0[75]}), .a ({key_s2[11], key_s1[11], key_s0[11]}), .c ({new_AGEMA_signal_1857, new_AGEMA_signal_1856, Midori_rounds_SelectedKey_11_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_12_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[76], key_s1[76], key_s0[76]}), .a ({key_s2[12], key_s1[12], key_s0[12]}), .c ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, Midori_rounds_SelectedKey_12_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_13_U1 ( .s (round_Signal[0]), .b ({key_s2[77], key_s1[77], key_s0[77]}), .a ({key_s2[13], key_s1[13], key_s0[13]}), .c ({new_AGEMA_signal_1859, new_AGEMA_signal_1858, Midori_rounds_SelectedKey_13_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_14_U1 ( .s (round_Signal[0]), .b ({key_s2[78], key_s1[78], key_s0[78]}), .a ({key_s2[14], key_s1[14], key_s0[14]}), .c ({new_AGEMA_signal_1861, new_AGEMA_signal_1860, Midori_rounds_SelectedKey_14_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_15_U1 ( .s (round_Signal[0]), .b ({key_s2[79], key_s1[79], key_s0[79]}), .a ({key_s2[15], key_s1[15], key_s0[15]}), .c ({new_AGEMA_signal_1863, new_AGEMA_signal_1862, Midori_rounds_SelectedKey_15_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_16_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[80], key_s1[80], key_s0[80]}), .a ({key_s2[16], key_s1[16], key_s0[16]}), .c ({new_AGEMA_signal_2579, new_AGEMA_signal_2578, Midori_rounds_SelectedKey_16_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_17_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[81], key_s1[81], key_s0[81]}), .a ({key_s2[17], key_s1[17], key_s0[17]}), .c ({new_AGEMA_signal_2581, new_AGEMA_signal_2580, Midori_rounds_SelectedKey_17_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_18_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[82], key_s1[82], key_s0[82]}), .a ({key_s2[18], key_s1[18], key_s0[18]}), .c ({new_AGEMA_signal_2583, new_AGEMA_signal_2582, Midori_rounds_SelectedKey_18_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_19_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[83], key_s1[83], key_s0[83]}), .a ({key_s2[19], key_s1[19], key_s0[19]}), .c ({new_AGEMA_signal_2585, new_AGEMA_signal_2584, Midori_rounds_SelectedKey_19_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_20_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[84], key_s1[84], key_s0[84]}), .a ({key_s2[20], key_s1[20], key_s0[20]}), .c ({new_AGEMA_signal_2587, new_AGEMA_signal_2586, Midori_rounds_SelectedKey_20_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_21_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[85], key_s1[85], key_s0[85]}), .a ({key_s2[21], key_s1[21], key_s0[21]}), .c ({new_AGEMA_signal_2589, new_AGEMA_signal_2588, Midori_rounds_SelectedKey_21_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_22_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[86], key_s1[86], key_s0[86]}), .a ({key_s2[22], key_s1[22], key_s0[22]}), .c ({new_AGEMA_signal_2591, new_AGEMA_signal_2590, Midori_rounds_SelectedKey_22_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_23_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[87], key_s1[87], key_s0[87]}), .a ({key_s2[23], key_s1[23], key_s0[23]}), .c ({new_AGEMA_signal_2593, new_AGEMA_signal_2592, Midori_rounds_SelectedKey_23_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_24_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[88], key_s1[88], key_s0[88]}), .a ({key_s2[24], key_s1[24], key_s0[24]}), .c ({new_AGEMA_signal_2595, new_AGEMA_signal_2594, Midori_rounds_SelectedKey_24_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_25_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[89], key_s1[89], key_s0[89]}), .a ({key_s2[25], key_s1[25], key_s0[25]}), .c ({new_AGEMA_signal_2597, new_AGEMA_signal_2596, Midori_rounds_SelectedKey_25_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_26_U1 ( .s (round_Signal[0]), .b ({key_s2[90], key_s1[90], key_s0[90]}), .a ({key_s2[26], key_s1[26], key_s0[26]}), .c ({new_AGEMA_signal_1865, new_AGEMA_signal_1864, Midori_rounds_SelectedKey_26_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_27_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[91], key_s1[91], key_s0[91]}), .a ({key_s2[27], key_s1[27], key_s0[27]}), .c ({new_AGEMA_signal_2599, new_AGEMA_signal_2598, Midori_rounds_SelectedKey_27_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_28_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[92], key_s1[92], key_s0[92]}), .a ({key_s2[28], key_s1[28], key_s0[28]}), .c ({new_AGEMA_signal_2601, new_AGEMA_signal_2600, Midori_rounds_SelectedKey_28_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_29_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[93], key_s1[93], key_s0[93]}), .a ({key_s2[29], key_s1[29], key_s0[29]}), .c ({new_AGEMA_signal_2603, new_AGEMA_signal_2602, Midori_rounds_SelectedKey_29_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_30_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[94], key_s1[94], key_s0[94]}), .a ({key_s2[30], key_s1[30], key_s0[30]}), .c ({new_AGEMA_signal_2605, new_AGEMA_signal_2604, Midori_rounds_SelectedKey_30_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_31_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[95], key_s1[95], key_s0[95]}), .a ({key_s2[31], key_s1[31], key_s0[31]}), .c ({new_AGEMA_signal_2607, new_AGEMA_signal_2606, Midori_rounds_SelectedKey_31_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_32_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[96], key_s1[96], key_s0[96]}), .a ({key_s2[32], key_s1[32], key_s0[32]}), .c ({new_AGEMA_signal_2609, new_AGEMA_signal_2608, Midori_rounds_SelectedKey_32_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_33_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[97], key_s1[97], key_s0[97]}), .a ({key_s2[33], key_s1[33], key_s0[33]}), .c ({new_AGEMA_signal_2611, new_AGEMA_signal_2610, Midori_rounds_SelectedKey_33_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_34_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[98], key_s1[98], key_s0[98]}), .a ({key_s2[34], key_s1[34], key_s0[34]}), .c ({new_AGEMA_signal_2613, new_AGEMA_signal_2612, Midori_rounds_SelectedKey_34_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_35_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[99], key_s1[99], key_s0[99]}), .a ({key_s2[35], key_s1[35], key_s0[35]}), .c ({new_AGEMA_signal_2615, new_AGEMA_signal_2614, Midori_rounds_SelectedKey_35_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_36_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[100], key_s1[100], key_s0[100]}), .a ({key_s2[36], key_s1[36], key_s0[36]}), .c ({new_AGEMA_signal_2617, new_AGEMA_signal_2616, Midori_rounds_SelectedKey_36_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_37_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[101], key_s1[101], key_s0[101]}), .a ({key_s2[37], key_s1[37], key_s0[37]}), .c ({new_AGEMA_signal_2619, new_AGEMA_signal_2618, Midori_rounds_SelectedKey_37_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_38_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[102], key_s1[102], key_s0[102]}), .a ({key_s2[38], key_s1[38], key_s0[38]}), .c ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, Midori_rounds_SelectedKey_38_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_39_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[103], key_s1[103], key_s0[103]}), .a ({key_s2[39], key_s1[39], key_s0[39]}), .c ({new_AGEMA_signal_2623, new_AGEMA_signal_2622, Midori_rounds_SelectedKey_39_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_40_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[104], key_s1[104], key_s0[104]}), .a ({key_s2[40], key_s1[40], key_s0[40]}), .c ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, Midori_rounds_SelectedKey_40_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_41_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[105], key_s1[105], key_s0[105]}), .a ({key_s2[41], key_s1[41], key_s0[41]}), .c ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, Midori_rounds_SelectedKey_41_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_42_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[106], key_s1[106], key_s0[106]}), .a ({key_s2[42], key_s1[42], key_s0[42]}), .c ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, Midori_rounds_SelectedKey_42_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_43_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[107], key_s1[107], key_s0[107]}), .a ({key_s2[43], key_s1[43], key_s0[43]}), .c ({new_AGEMA_signal_2631, new_AGEMA_signal_2630, Midori_rounds_SelectedKey_43_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_44_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[108], key_s1[108], key_s0[108]}), .a ({key_s2[44], key_s1[44], key_s0[44]}), .c ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, Midori_rounds_SelectedKey_44_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_45_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[109], key_s1[109], key_s0[109]}), .a ({key_s2[45], key_s1[45], key_s0[45]}), .c ({new_AGEMA_signal_2635, new_AGEMA_signal_2634, Midori_rounds_SelectedKey_45_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_46_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[110], key_s1[110], key_s0[110]}), .a ({key_s2[46], key_s1[46], key_s0[46]}), .c ({new_AGEMA_signal_2637, new_AGEMA_signal_2636, Midori_rounds_SelectedKey_46_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_47_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[111], key_s1[111], key_s0[111]}), .a ({key_s2[47], key_s1[47], key_s0[47]}), .c ({new_AGEMA_signal_2639, new_AGEMA_signal_2638, Midori_rounds_SelectedKey_47_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_48_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[112], key_s1[112], key_s0[112]}), .a ({key_s2[48], key_s1[48], key_s0[48]}), .c ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, Midori_rounds_SelectedKey_48_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_49_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[113], key_s1[113], key_s0[113]}), .a ({key_s2[49], key_s1[49], key_s0[49]}), .c ({new_AGEMA_signal_2643, new_AGEMA_signal_2642, Midori_rounds_SelectedKey_49_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_50_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[114], key_s1[114], key_s0[114]}), .a ({key_s2[50], key_s1[50], key_s0[50]}), .c ({new_AGEMA_signal_2645, new_AGEMA_signal_2644, Midori_rounds_SelectedKey_50_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_51_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[115], key_s1[115], key_s0[115]}), .a ({key_s2[51], key_s1[51], key_s0[51]}), .c ({new_AGEMA_signal_2647, new_AGEMA_signal_2646, Midori_rounds_SelectedKey_51_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_52_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[116], key_s1[116], key_s0[116]}), .a ({key_s2[52], key_s1[52], key_s0[52]}), .c ({new_AGEMA_signal_2649, new_AGEMA_signal_2648, Midori_rounds_SelectedKey_52_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_53_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[117], key_s1[117], key_s0[117]}), .a ({key_s2[53], key_s1[53], key_s0[53]}), .c ({new_AGEMA_signal_2651, new_AGEMA_signal_2650, Midori_rounds_SelectedKey_53_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_54_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[118], key_s1[118], key_s0[118]}), .a ({key_s2[54], key_s1[54], key_s0[54]}), .c ({new_AGEMA_signal_2653, new_AGEMA_signal_2652, Midori_rounds_SelectedKey_54_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_55_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[119], key_s1[119], key_s0[119]}), .a ({key_s2[55], key_s1[55], key_s0[55]}), .c ({new_AGEMA_signal_2655, new_AGEMA_signal_2654, Midori_rounds_SelectedKey_55_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_56_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[120], key_s1[120], key_s0[120]}), .a ({key_s2[56], key_s1[56], key_s0[56]}), .c ({new_AGEMA_signal_2657, new_AGEMA_signal_2656, Midori_rounds_SelectedKey_56_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_57_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[121], key_s1[121], key_s0[121]}), .a ({key_s2[57], key_s1[57], key_s0[57]}), .c ({new_AGEMA_signal_2659, new_AGEMA_signal_2658, Midori_rounds_SelectedKey_57_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_58_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[122], key_s1[122], key_s0[122]}), .a ({key_s2[58], key_s1[58], key_s0[58]}), .c ({new_AGEMA_signal_2661, new_AGEMA_signal_2660, Midori_rounds_SelectedKey_58_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_59_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[123], key_s1[123], key_s0[123]}), .a ({key_s2[59], key_s1[59], key_s0[59]}), .c ({new_AGEMA_signal_2663, new_AGEMA_signal_2662, Midori_rounds_SelectedKey_59_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_60_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[124], key_s1[124], key_s0[124]}), .a ({key_s2[60], key_s1[60], key_s0[60]}), .c ({new_AGEMA_signal_2665, new_AGEMA_signal_2664, Midori_rounds_SelectedKey_60_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_61_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[125], key_s1[125], key_s0[125]}), .a ({key_s2[61], key_s1[61], key_s0[61]}), .c ({new_AGEMA_signal_2667, new_AGEMA_signal_2666, Midori_rounds_SelectedKey_61_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_62_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[126], key_s1[126], key_s0[126]}), .a ({key_s2[62], key_s1[62], key_s0[62]}), .c ({new_AGEMA_signal_2669, new_AGEMA_signal_2668, Midori_rounds_SelectedKey_62_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_MUXInst_mux_inst_63_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[127], key_s1[127], key_s0[127]}), .a ({key_s2[63], key_s1[63], key_s0[63]}), .c ({new_AGEMA_signal_2671, new_AGEMA_signal_2670, Midori_rounds_SelectedKey_63_}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U4 ( .a ({new_AGEMA_signal_1867, new_AGEMA_signal_1866, Midori_rounds_roundReg_out[0]}), .b ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, Midori_rounds_sub_sBox_PRINCE_0_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U2 ( .a ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, Midori_rounds_roundReg_out[3]}), .b ({new_AGEMA_signal_1879, new_AGEMA_signal_1878, Midori_rounds_sub_sBox_PRINCE_0_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U1 ( .a ({new_AGEMA_signal_1873, new_AGEMA_signal_1872, Midori_rounds_roundReg_out[2]}), .b ({new_AGEMA_signal_1881, new_AGEMA_signal_1880, Midori_rounds_sub_sBox_PRINCE_0_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U4 ( .a ({new_AGEMA_signal_1883, new_AGEMA_signal_1882, Midori_rounds_roundReg_out[4]}), .b ({new_AGEMA_signal_1893, new_AGEMA_signal_1892, Midori_rounds_sub_sBox_PRINCE_1_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U2 ( .a ({new_AGEMA_signal_1885, new_AGEMA_signal_1884, Midori_rounds_roundReg_out[7]}), .b ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, Midori_rounds_sub_sBox_PRINCE_1_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U1 ( .a ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, Midori_rounds_roundReg_out[6]}), .b ({new_AGEMA_signal_1897, new_AGEMA_signal_1896, Midori_rounds_sub_sBox_PRINCE_1_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U4 ( .a ({new_AGEMA_signal_1899, new_AGEMA_signal_1898, Midori_rounds_roundReg_out[8]}), .b ({new_AGEMA_signal_1909, new_AGEMA_signal_1908, Midori_rounds_sub_sBox_PRINCE_2_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U2 ( .a ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, Midori_rounds_roundReg_out[11]}), .b ({new_AGEMA_signal_1911, new_AGEMA_signal_1910, Midori_rounds_sub_sBox_PRINCE_2_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U1 ( .a ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, Midori_rounds_roundReg_out[10]}), .b ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, Midori_rounds_sub_sBox_PRINCE_2_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U4 ( .a ({new_AGEMA_signal_1915, new_AGEMA_signal_1914, Midori_rounds_roundReg_out[12]}), .b ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, Midori_rounds_sub_sBox_PRINCE_3_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U2 ( .a ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, Midori_rounds_roundReg_out[15]}), .b ({new_AGEMA_signal_1927, new_AGEMA_signal_1926, Midori_rounds_sub_sBox_PRINCE_3_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U1 ( .a ({new_AGEMA_signal_1921, new_AGEMA_signal_1920, Midori_rounds_roundReg_out[14]}), .b ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, Midori_rounds_sub_sBox_PRINCE_3_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U4 ( .a ({new_AGEMA_signal_1931, new_AGEMA_signal_1930, Midori_rounds_roundReg_out[16]}), .b ({new_AGEMA_signal_1941, new_AGEMA_signal_1940, Midori_rounds_sub_sBox_PRINCE_4_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U2 ( .a ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, Midori_rounds_roundReg_out[19]}), .b ({new_AGEMA_signal_1943, new_AGEMA_signal_1942, Midori_rounds_sub_sBox_PRINCE_4_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U1 ( .a ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, Midori_rounds_roundReg_out[18]}), .b ({new_AGEMA_signal_1945, new_AGEMA_signal_1944, Midori_rounds_sub_sBox_PRINCE_4_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U4 ( .a ({new_AGEMA_signal_1947, new_AGEMA_signal_1946, Midori_rounds_roundReg_out[20]}), .b ({new_AGEMA_signal_1957, new_AGEMA_signal_1956, Midori_rounds_sub_sBox_PRINCE_5_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U2 ( .a ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, Midori_rounds_roundReg_out[23]}), .b ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, Midori_rounds_sub_sBox_PRINCE_5_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U1 ( .a ({new_AGEMA_signal_1953, new_AGEMA_signal_1952, Midori_rounds_roundReg_out[22]}), .b ({new_AGEMA_signal_1961, new_AGEMA_signal_1960, Midori_rounds_sub_sBox_PRINCE_5_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U4 ( .a ({new_AGEMA_signal_1963, new_AGEMA_signal_1962, Midori_rounds_roundReg_out[24]}), .b ({new_AGEMA_signal_1973, new_AGEMA_signal_1972, Midori_rounds_sub_sBox_PRINCE_6_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U2 ( .a ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, Midori_rounds_roundReg_out[27]}), .b ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, Midori_rounds_sub_sBox_PRINCE_6_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U1 ( .a ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, Midori_rounds_roundReg_out[26]}), .b ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, Midori_rounds_sub_sBox_PRINCE_6_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U4 ( .a ({new_AGEMA_signal_1979, new_AGEMA_signal_1978, Midori_rounds_roundReg_out[28]}), .b ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, Midori_rounds_sub_sBox_PRINCE_7_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U2 ( .a ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, Midori_rounds_roundReg_out[31]}), .b ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, Midori_rounds_sub_sBox_PRINCE_7_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U1 ( .a ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, Midori_rounds_roundReg_out[30]}), .b ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, Midori_rounds_sub_sBox_PRINCE_7_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U4 ( .a ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, Midori_rounds_roundReg_out[32]}), .b ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, Midori_rounds_sub_sBox_PRINCE_8_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U2 ( .a ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, Midori_rounds_roundReg_out[35]}), .b ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, Midori_rounds_sub_sBox_PRINCE_8_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U1 ( .a ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, Midori_rounds_roundReg_out[34]}), .b ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, Midori_rounds_sub_sBox_PRINCE_8_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U4 ( .a ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, Midori_rounds_roundReg_out[36]}), .b ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, Midori_rounds_sub_sBox_PRINCE_9_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U2 ( .a ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, Midori_rounds_roundReg_out[39]}), .b ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, Midori_rounds_sub_sBox_PRINCE_9_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U1 ( .a ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, Midori_rounds_roundReg_out[38]}), .b ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, Midori_rounds_sub_sBox_PRINCE_9_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U4 ( .a ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, Midori_rounds_roundReg_out[40]}), .b ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, Midori_rounds_sub_sBox_PRINCE_10_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U2 ( .a ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, Midori_rounds_roundReg_out[43]}), .b ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, Midori_rounds_sub_sBox_PRINCE_10_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U1 ( .a ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, Midori_rounds_roundReg_out[42]}), .b ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, Midori_rounds_sub_sBox_PRINCE_10_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U4 ( .a ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, Midori_rounds_roundReg_out[44]}), .b ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, Midori_rounds_sub_sBox_PRINCE_11_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U2 ( .a ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, Midori_rounds_roundReg_out[47]}), .b ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, Midori_rounds_sub_sBox_PRINCE_11_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U1 ( .a ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, Midori_rounds_roundReg_out[46]}), .b ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, Midori_rounds_sub_sBox_PRINCE_11_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U4 ( .a ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, Midori_rounds_roundReg_out[48]}), .b ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, Midori_rounds_sub_sBox_PRINCE_12_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U2 ( .a ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, Midori_rounds_roundReg_out[51]}), .b ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, Midori_rounds_sub_sBox_PRINCE_12_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U1 ( .a ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, Midori_rounds_roundReg_out[50]}), .b ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, Midori_rounds_sub_sBox_PRINCE_12_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U4 ( .a ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, Midori_rounds_roundReg_out[52]}), .b ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, Midori_rounds_sub_sBox_PRINCE_13_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U2 ( .a ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, Midori_rounds_roundReg_out[55]}), .b ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, Midori_rounds_sub_sBox_PRINCE_13_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U1 ( .a ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, Midori_rounds_roundReg_out[54]}), .b ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, Midori_rounds_sub_sBox_PRINCE_13_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U4 ( .a ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, Midori_rounds_roundReg_out[56]}), .b ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, Midori_rounds_sub_sBox_PRINCE_14_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U2 ( .a ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, Midori_rounds_roundReg_out[59]}), .b ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, Midori_rounds_sub_sBox_PRINCE_14_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U1 ( .a ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, Midori_rounds_roundReg_out[58]}), .b ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, Midori_rounds_sub_sBox_PRINCE_14_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U4 ( .a ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, Midori_rounds_roundReg_out[60]}), .b ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, Midori_rounds_sub_sBox_PRINCE_15_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U2 ( .a ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, Midori_rounds_roundReg_out[63]}), .b ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, Midori_rounds_sub_sBox_PRINCE_15_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U1 ( .a ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, Midori_rounds_roundReg_out[62]}), .b ({new_AGEMA_signal_2121, new_AGEMA_signal_2120, Midori_rounds_sub_sBox_PRINCE_15_n9}) ) ;
    ClockGatingController #(9) ClockGatingInst ( .clk (clk), .rst (reset), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U14 ( .a ({new_AGEMA_signal_1867, new_AGEMA_signal_1866, Midori_rounds_roundReg_out[0]}), .b ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, Midori_rounds_roundReg_out[3]}), .clk (clk), .r ({Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_1871, new_AGEMA_signal_1870, Midori_rounds_sub_sBox_PRINCE_0_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U13 ( .a ({new_AGEMA_signal_1879, new_AGEMA_signal_1878, Midori_rounds_sub_sBox_PRINCE_0_n8}), .b ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, Midori_rounds_sub_sBox_PRINCE_0_n7}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3]}), .c ({new_AGEMA_signal_2381, new_AGEMA_signal_2380, Midori_rounds_sub_sBox_PRINCE_0_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U10 ( .a ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, Midori_rounds_roundReg_out[3]}), .b ({new_AGEMA_signal_1881, new_AGEMA_signal_1880, Midori_rounds_sub_sBox_PRINCE_0_n9}), .clk (clk), .r ({Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, Midori_rounds_sub_sBox_PRINCE_0_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U9 ( .a ({new_AGEMA_signal_1873, new_AGEMA_signal_1872, Midori_rounds_roundReg_out[2]}), .b ({new_AGEMA_signal_1879, new_AGEMA_signal_1878, Midori_rounds_sub_sBox_PRINCE_0_n8}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9]}), .c ({new_AGEMA_signal_2385, new_AGEMA_signal_2384, Midori_rounds_sub_sBox_PRINCE_0_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U5 ( .a ({new_AGEMA_signal_1873, new_AGEMA_signal_1872, Midori_rounds_roundReg_out[2]}), .b ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, Midori_rounds_roundReg_out[3]}), .clk (clk), .r ({Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_1875, new_AGEMA_signal_1874, Midori_rounds_sub_sBox_PRINCE_0_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U3 ( .a ({new_AGEMA_signal_1881, new_AGEMA_signal_1880, Midori_rounds_sub_sBox_PRINCE_0_n9}), .b ({new_AGEMA_signal_1879, new_AGEMA_signal_1878, Midori_rounds_sub_sBox_PRINCE_0_n8}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15]}), .c ({new_AGEMA_signal_2389, new_AGEMA_signal_2388, Midori_rounds_sub_sBox_PRINCE_0_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U14 ( .a ({new_AGEMA_signal_1883, new_AGEMA_signal_1882, Midori_rounds_roundReg_out[4]}), .b ({new_AGEMA_signal_1885, new_AGEMA_signal_1884, Midori_rounds_roundReg_out[7]}), .clk (clk), .r ({Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_1887, new_AGEMA_signal_1886, Midori_rounds_sub_sBox_PRINCE_1_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U13 ( .a ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, Midori_rounds_sub_sBox_PRINCE_1_n8}), .b ({new_AGEMA_signal_1893, new_AGEMA_signal_1892, Midori_rounds_sub_sBox_PRINCE_1_n7}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21]}), .c ({new_AGEMA_signal_2393, new_AGEMA_signal_2392, Midori_rounds_sub_sBox_PRINCE_1_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U10 ( .a ({new_AGEMA_signal_1885, new_AGEMA_signal_1884, Midori_rounds_roundReg_out[7]}), .b ({new_AGEMA_signal_1897, new_AGEMA_signal_1896, Midori_rounds_sub_sBox_PRINCE_1_n9}), .clk (clk), .r ({Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_2395, new_AGEMA_signal_2394, Midori_rounds_sub_sBox_PRINCE_1_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U9 ( .a ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, Midori_rounds_roundReg_out[6]}), .b ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, Midori_rounds_sub_sBox_PRINCE_1_n8}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27]}), .c ({new_AGEMA_signal_2397, new_AGEMA_signal_2396, Midori_rounds_sub_sBox_PRINCE_1_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U5 ( .a ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, Midori_rounds_roundReg_out[6]}), .b ({new_AGEMA_signal_1885, new_AGEMA_signal_1884, Midori_rounds_roundReg_out[7]}), .clk (clk), .r ({Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_1891, new_AGEMA_signal_1890, Midori_rounds_sub_sBox_PRINCE_1_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U3 ( .a ({new_AGEMA_signal_1897, new_AGEMA_signal_1896, Midori_rounds_sub_sBox_PRINCE_1_n9}), .b ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, Midori_rounds_sub_sBox_PRINCE_1_n8}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33]}), .c ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, Midori_rounds_sub_sBox_PRINCE_1_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U14 ( .a ({new_AGEMA_signal_1899, new_AGEMA_signal_1898, Midori_rounds_roundReg_out[8]}), .b ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, Midori_rounds_roundReg_out[11]}), .clk (clk), .r ({Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_1903, new_AGEMA_signal_1902, Midori_rounds_sub_sBox_PRINCE_2_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U13 ( .a ({new_AGEMA_signal_1911, new_AGEMA_signal_1910, Midori_rounds_sub_sBox_PRINCE_2_n8}), .b ({new_AGEMA_signal_1909, new_AGEMA_signal_1908, Midori_rounds_sub_sBox_PRINCE_2_n7}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39]}), .c ({new_AGEMA_signal_2405, new_AGEMA_signal_2404, Midori_rounds_sub_sBox_PRINCE_2_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U10 ( .a ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, Midori_rounds_roundReg_out[11]}), .b ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, Midori_rounds_sub_sBox_PRINCE_2_n9}), .clk (clk), .r ({Fresh[44], Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_2407, new_AGEMA_signal_2406, Midori_rounds_sub_sBox_PRINCE_2_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U9 ( .a ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, Midori_rounds_roundReg_out[10]}), .b ({new_AGEMA_signal_1911, new_AGEMA_signal_1910, Midori_rounds_sub_sBox_PRINCE_2_n8}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45]}), .c ({new_AGEMA_signal_2409, new_AGEMA_signal_2408, Midori_rounds_sub_sBox_PRINCE_2_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U5 ( .a ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, Midori_rounds_roundReg_out[10]}), .b ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, Midori_rounds_roundReg_out[11]}), .clk (clk), .r ({Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, Midori_rounds_sub_sBox_PRINCE_2_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U3 ( .a ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, Midori_rounds_sub_sBox_PRINCE_2_n9}), .b ({new_AGEMA_signal_1911, new_AGEMA_signal_1910, Midori_rounds_sub_sBox_PRINCE_2_n8}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51]}), .c ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, Midori_rounds_sub_sBox_PRINCE_2_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U14 ( .a ({new_AGEMA_signal_1915, new_AGEMA_signal_1914, Midori_rounds_roundReg_out[12]}), .b ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, Midori_rounds_roundReg_out[15]}), .clk (clk), .r ({Fresh[56], Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_1919, new_AGEMA_signal_1918, Midori_rounds_sub_sBox_PRINCE_3_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U13 ( .a ({new_AGEMA_signal_1927, new_AGEMA_signal_1926, Midori_rounds_sub_sBox_PRINCE_3_n8}), .b ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, Midori_rounds_sub_sBox_PRINCE_3_n7}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57]}), .c ({new_AGEMA_signal_2417, new_AGEMA_signal_2416, Midori_rounds_sub_sBox_PRINCE_3_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U10 ( .a ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, Midori_rounds_roundReg_out[15]}), .b ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, Midori_rounds_sub_sBox_PRINCE_3_n9}), .clk (clk), .r ({Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_2419, new_AGEMA_signal_2418, Midori_rounds_sub_sBox_PRINCE_3_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U9 ( .a ({new_AGEMA_signal_1921, new_AGEMA_signal_1920, Midori_rounds_roundReg_out[14]}), .b ({new_AGEMA_signal_1927, new_AGEMA_signal_1926, Midori_rounds_sub_sBox_PRINCE_3_n8}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63]}), .c ({new_AGEMA_signal_2421, new_AGEMA_signal_2420, Midori_rounds_sub_sBox_PRINCE_3_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U5 ( .a ({new_AGEMA_signal_1921, new_AGEMA_signal_1920, Midori_rounds_roundReg_out[14]}), .b ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, Midori_rounds_roundReg_out[15]}), .clk (clk), .r ({Fresh[68], Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_1923, new_AGEMA_signal_1922, Midori_rounds_sub_sBox_PRINCE_3_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U3 ( .a ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, Midori_rounds_sub_sBox_PRINCE_3_n9}), .b ({new_AGEMA_signal_1927, new_AGEMA_signal_1926, Midori_rounds_sub_sBox_PRINCE_3_n8}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69]}), .c ({new_AGEMA_signal_2425, new_AGEMA_signal_2424, Midori_rounds_sub_sBox_PRINCE_3_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U14 ( .a ({new_AGEMA_signal_1931, new_AGEMA_signal_1930, Midori_rounds_roundReg_out[16]}), .b ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, Midori_rounds_roundReg_out[19]}), .clk (clk), .r ({Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_1935, new_AGEMA_signal_1934, Midori_rounds_sub_sBox_PRINCE_4_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U13 ( .a ({new_AGEMA_signal_1943, new_AGEMA_signal_1942, Midori_rounds_sub_sBox_PRINCE_4_n8}), .b ({new_AGEMA_signal_1941, new_AGEMA_signal_1940, Midori_rounds_sub_sBox_PRINCE_4_n7}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75]}), .c ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, Midori_rounds_sub_sBox_PRINCE_4_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U10 ( .a ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, Midori_rounds_roundReg_out[19]}), .b ({new_AGEMA_signal_1945, new_AGEMA_signal_1944, Midori_rounds_sub_sBox_PRINCE_4_n9}), .clk (clk), .r ({Fresh[80], Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_2431, new_AGEMA_signal_2430, Midori_rounds_sub_sBox_PRINCE_4_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U9 ( .a ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, Midori_rounds_roundReg_out[18]}), .b ({new_AGEMA_signal_1943, new_AGEMA_signal_1942, Midori_rounds_sub_sBox_PRINCE_4_n8}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81]}), .c ({new_AGEMA_signal_2433, new_AGEMA_signal_2432, Midori_rounds_sub_sBox_PRINCE_4_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U5 ( .a ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, Midori_rounds_roundReg_out[18]}), .b ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, Midori_rounds_roundReg_out[19]}), .clk (clk), .r ({Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_1939, new_AGEMA_signal_1938, Midori_rounds_sub_sBox_PRINCE_4_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U3 ( .a ({new_AGEMA_signal_1945, new_AGEMA_signal_1944, Midori_rounds_sub_sBox_PRINCE_4_n9}), .b ({new_AGEMA_signal_1943, new_AGEMA_signal_1942, Midori_rounds_sub_sBox_PRINCE_4_n8}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87]}), .c ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, Midori_rounds_sub_sBox_PRINCE_4_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U14 ( .a ({new_AGEMA_signal_1947, new_AGEMA_signal_1946, Midori_rounds_roundReg_out[20]}), .b ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, Midori_rounds_roundReg_out[23]}), .clk (clk), .r ({Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_1951, new_AGEMA_signal_1950, Midori_rounds_sub_sBox_PRINCE_5_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U13 ( .a ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, Midori_rounds_sub_sBox_PRINCE_5_n8}), .b ({new_AGEMA_signal_1957, new_AGEMA_signal_1956, Midori_rounds_sub_sBox_PRINCE_5_n7}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93]}), .c ({new_AGEMA_signal_2441, new_AGEMA_signal_2440, Midori_rounds_sub_sBox_PRINCE_5_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U10 ( .a ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, Midori_rounds_roundReg_out[23]}), .b ({new_AGEMA_signal_1961, new_AGEMA_signal_1960, Midori_rounds_sub_sBox_PRINCE_5_n9}), .clk (clk), .r ({Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_2443, new_AGEMA_signal_2442, Midori_rounds_sub_sBox_PRINCE_5_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U9 ( .a ({new_AGEMA_signal_1953, new_AGEMA_signal_1952, Midori_rounds_roundReg_out[22]}), .b ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, Midori_rounds_sub_sBox_PRINCE_5_n8}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99]}), .c ({new_AGEMA_signal_2445, new_AGEMA_signal_2444, Midori_rounds_sub_sBox_PRINCE_5_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U5 ( .a ({new_AGEMA_signal_1953, new_AGEMA_signal_1952, Midori_rounds_roundReg_out[22]}), .b ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, Midori_rounds_roundReg_out[23]}), .clk (clk), .r ({Fresh[104], Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_1955, new_AGEMA_signal_1954, Midori_rounds_sub_sBox_PRINCE_5_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U3 ( .a ({new_AGEMA_signal_1961, new_AGEMA_signal_1960, Midori_rounds_sub_sBox_PRINCE_5_n9}), .b ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, Midori_rounds_sub_sBox_PRINCE_5_n8}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105]}), .c ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, Midori_rounds_sub_sBox_PRINCE_5_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U14 ( .a ({new_AGEMA_signal_1963, new_AGEMA_signal_1962, Midori_rounds_roundReg_out[24]}), .b ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, Midori_rounds_roundReg_out[27]}), .clk (clk), .r ({Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_1967, new_AGEMA_signal_1966, Midori_rounds_sub_sBox_PRINCE_6_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U13 ( .a ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, Midori_rounds_sub_sBox_PRINCE_6_n8}), .b ({new_AGEMA_signal_1973, new_AGEMA_signal_1972, Midori_rounds_sub_sBox_PRINCE_6_n7}), .clk (clk), .r ({Fresh[113], Fresh[112], Fresh[111]}), .c ({new_AGEMA_signal_2453, new_AGEMA_signal_2452, Midori_rounds_sub_sBox_PRINCE_6_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U10 ( .a ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, Midori_rounds_roundReg_out[27]}), .b ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, Midori_rounds_sub_sBox_PRINCE_6_n9}), .clk (clk), .r ({Fresh[116], Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_2455, new_AGEMA_signal_2454, Midori_rounds_sub_sBox_PRINCE_6_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U9 ( .a ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, Midori_rounds_roundReg_out[26]}), .b ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, Midori_rounds_sub_sBox_PRINCE_6_n8}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117]}), .c ({new_AGEMA_signal_2457, new_AGEMA_signal_2456, Midori_rounds_sub_sBox_PRINCE_6_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U5 ( .a ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, Midori_rounds_roundReg_out[26]}), .b ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, Midori_rounds_roundReg_out[27]}), .clk (clk), .r ({Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_1971, new_AGEMA_signal_1970, Midori_rounds_sub_sBox_PRINCE_6_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U3 ( .a ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, Midori_rounds_sub_sBox_PRINCE_6_n9}), .b ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, Midori_rounds_sub_sBox_PRINCE_6_n8}), .clk (clk), .r ({Fresh[125], Fresh[124], Fresh[123]}), .c ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, Midori_rounds_sub_sBox_PRINCE_6_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U14 ( .a ({new_AGEMA_signal_1979, new_AGEMA_signal_1978, Midori_rounds_roundReg_out[28]}), .b ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, Midori_rounds_roundReg_out[31]}), .clk (clk), .r ({Fresh[128], Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, Midori_rounds_sub_sBox_PRINCE_7_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U13 ( .a ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, Midori_rounds_sub_sBox_PRINCE_7_n8}), .b ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, Midori_rounds_sub_sBox_PRINCE_7_n7}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129]}), .c ({new_AGEMA_signal_2465, new_AGEMA_signal_2464, Midori_rounds_sub_sBox_PRINCE_7_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U10 ( .a ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, Midori_rounds_roundReg_out[31]}), .b ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, Midori_rounds_sub_sBox_PRINCE_7_n9}), .clk (clk), .r ({Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_2467, new_AGEMA_signal_2466, Midori_rounds_sub_sBox_PRINCE_7_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U9 ( .a ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, Midori_rounds_roundReg_out[30]}), .b ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, Midori_rounds_sub_sBox_PRINCE_7_n8}), .clk (clk), .r ({Fresh[137], Fresh[136], Fresh[135]}), .c ({new_AGEMA_signal_2469, new_AGEMA_signal_2468, Midori_rounds_sub_sBox_PRINCE_7_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U5 ( .a ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, Midori_rounds_roundReg_out[30]}), .b ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, Midori_rounds_roundReg_out[31]}), .clk (clk), .r ({Fresh[140], Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, Midori_rounds_sub_sBox_PRINCE_7_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U3 ( .a ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, Midori_rounds_sub_sBox_PRINCE_7_n9}), .b ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, Midori_rounds_sub_sBox_PRINCE_7_n8}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141]}), .c ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, Midori_rounds_sub_sBox_PRINCE_7_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U14 ( .a ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, Midori_rounds_roundReg_out[32]}), .b ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, Midori_rounds_roundReg_out[35]}), .clk (clk), .r ({Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, Midori_rounds_sub_sBox_PRINCE_8_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U13 ( .a ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, Midori_rounds_sub_sBox_PRINCE_8_n8}), .b ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, Midori_rounds_sub_sBox_PRINCE_8_n7}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147]}), .c ({new_AGEMA_signal_2477, new_AGEMA_signal_2476, Midori_rounds_sub_sBox_PRINCE_8_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U10 ( .a ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, Midori_rounds_roundReg_out[35]}), .b ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, Midori_rounds_sub_sBox_PRINCE_8_n9}), .clk (clk), .r ({Fresh[152], Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, Midori_rounds_sub_sBox_PRINCE_8_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U9 ( .a ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, Midori_rounds_roundReg_out[34]}), .b ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, Midori_rounds_sub_sBox_PRINCE_8_n8}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153]}), .c ({new_AGEMA_signal_2481, new_AGEMA_signal_2480, Midori_rounds_sub_sBox_PRINCE_8_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U5 ( .a ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, Midori_rounds_roundReg_out[34]}), .b ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, Midori_rounds_roundReg_out[35]}), .clk (clk), .r ({Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_2003, new_AGEMA_signal_2002, Midori_rounds_sub_sBox_PRINCE_8_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U3 ( .a ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, Midori_rounds_sub_sBox_PRINCE_8_n9}), .b ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, Midori_rounds_sub_sBox_PRINCE_8_n8}), .clk (clk), .r ({Fresh[161], Fresh[160], Fresh[159]}), .c ({new_AGEMA_signal_2485, new_AGEMA_signal_2484, Midori_rounds_sub_sBox_PRINCE_8_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U14 ( .a ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, Midori_rounds_roundReg_out[36]}), .b ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, Midori_rounds_roundReg_out[39]}), .clk (clk), .r ({Fresh[164], Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, Midori_rounds_sub_sBox_PRINCE_9_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U13 ( .a ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, Midori_rounds_sub_sBox_PRINCE_9_n8}), .b ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, Midori_rounds_sub_sBox_PRINCE_9_n7}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165]}), .c ({new_AGEMA_signal_2489, new_AGEMA_signal_2488, Midori_rounds_sub_sBox_PRINCE_9_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U10 ( .a ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, Midori_rounds_roundReg_out[39]}), .b ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, Midori_rounds_sub_sBox_PRINCE_9_n9}), .clk (clk), .r ({Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, Midori_rounds_sub_sBox_PRINCE_9_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U9 ( .a ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, Midori_rounds_roundReg_out[38]}), .b ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, Midori_rounds_sub_sBox_PRINCE_9_n8}), .clk (clk), .r ({Fresh[173], Fresh[172], Fresh[171]}), .c ({new_AGEMA_signal_2493, new_AGEMA_signal_2492, Midori_rounds_sub_sBox_PRINCE_9_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U5 ( .a ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, Midori_rounds_roundReg_out[38]}), .b ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, Midori_rounds_roundReg_out[39]}), .clk (clk), .r ({Fresh[176], Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, Midori_rounds_sub_sBox_PRINCE_9_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U3 ( .a ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, Midori_rounds_sub_sBox_PRINCE_9_n9}), .b ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, Midori_rounds_sub_sBox_PRINCE_9_n8}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177]}), .c ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, Midori_rounds_sub_sBox_PRINCE_9_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U14 ( .a ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, Midori_rounds_roundReg_out[40]}), .b ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, Midori_rounds_roundReg_out[43]}), .clk (clk), .r ({Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, Midori_rounds_sub_sBox_PRINCE_10_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U13 ( .a ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, Midori_rounds_sub_sBox_PRINCE_10_n8}), .b ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, Midori_rounds_sub_sBox_PRINCE_10_n7}), .clk (clk), .r ({Fresh[185], Fresh[184], Fresh[183]}), .c ({new_AGEMA_signal_2501, new_AGEMA_signal_2500, Midori_rounds_sub_sBox_PRINCE_10_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U10 ( .a ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, Midori_rounds_roundReg_out[43]}), .b ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, Midori_rounds_sub_sBox_PRINCE_10_n9}), .clk (clk), .r ({Fresh[188], Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_2503, new_AGEMA_signal_2502, Midori_rounds_sub_sBox_PRINCE_10_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U9 ( .a ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, Midori_rounds_roundReg_out[42]}), .b ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, Midori_rounds_sub_sBox_PRINCE_10_n8}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189]}), .c ({new_AGEMA_signal_2505, new_AGEMA_signal_2504, Midori_rounds_sub_sBox_PRINCE_10_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U5 ( .a ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, Midori_rounds_roundReg_out[42]}), .b ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, Midori_rounds_roundReg_out[43]}), .clk (clk), .r ({Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, Midori_rounds_sub_sBox_PRINCE_10_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U3 ( .a ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, Midori_rounds_sub_sBox_PRINCE_10_n9}), .b ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, Midori_rounds_sub_sBox_PRINCE_10_n8}), .clk (clk), .r ({Fresh[197], Fresh[196], Fresh[195]}), .c ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, Midori_rounds_sub_sBox_PRINCE_10_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U14 ( .a ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, Midori_rounds_roundReg_out[44]}), .b ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, Midori_rounds_roundReg_out[47]}), .clk (clk), .r ({Fresh[200], Fresh[199], Fresh[198]}), .c ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, Midori_rounds_sub_sBox_PRINCE_11_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U13 ( .a ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, Midori_rounds_sub_sBox_PRINCE_11_n8}), .b ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, Midori_rounds_sub_sBox_PRINCE_11_n7}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201]}), .c ({new_AGEMA_signal_2513, new_AGEMA_signal_2512, Midori_rounds_sub_sBox_PRINCE_11_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U10 ( .a ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, Midori_rounds_roundReg_out[47]}), .b ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, Midori_rounds_sub_sBox_PRINCE_11_n9}), .clk (clk), .r ({Fresh[206], Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_2515, new_AGEMA_signal_2514, Midori_rounds_sub_sBox_PRINCE_11_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U9 ( .a ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, Midori_rounds_roundReg_out[46]}), .b ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, Midori_rounds_sub_sBox_PRINCE_11_n8}), .clk (clk), .r ({Fresh[209], Fresh[208], Fresh[207]}), .c ({new_AGEMA_signal_2517, new_AGEMA_signal_2516, Midori_rounds_sub_sBox_PRINCE_11_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U5 ( .a ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, Midori_rounds_roundReg_out[46]}), .b ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, Midori_rounds_roundReg_out[47]}), .clk (clk), .r ({Fresh[212], Fresh[211], Fresh[210]}), .c ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, Midori_rounds_sub_sBox_PRINCE_11_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U3 ( .a ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, Midori_rounds_sub_sBox_PRINCE_11_n9}), .b ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, Midori_rounds_sub_sBox_PRINCE_11_n8}), .clk (clk), .r ({Fresh[215], Fresh[214], Fresh[213]}), .c ({new_AGEMA_signal_2521, new_AGEMA_signal_2520, Midori_rounds_sub_sBox_PRINCE_11_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U14 ( .a ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, Midori_rounds_roundReg_out[48]}), .b ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, Midori_rounds_roundReg_out[51]}), .clk (clk), .r ({Fresh[218], Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, Midori_rounds_sub_sBox_PRINCE_12_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U13 ( .a ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, Midori_rounds_sub_sBox_PRINCE_12_n8}), .b ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, Midori_rounds_sub_sBox_PRINCE_12_n7}), .clk (clk), .r ({Fresh[221], Fresh[220], Fresh[219]}), .c ({new_AGEMA_signal_2525, new_AGEMA_signal_2524, Midori_rounds_sub_sBox_PRINCE_12_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U10 ( .a ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, Midori_rounds_roundReg_out[51]}), .b ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, Midori_rounds_sub_sBox_PRINCE_12_n9}), .clk (clk), .r ({Fresh[224], Fresh[223], Fresh[222]}), .c ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, Midori_rounds_sub_sBox_PRINCE_12_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U9 ( .a ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, Midori_rounds_roundReg_out[50]}), .b ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, Midori_rounds_sub_sBox_PRINCE_12_n8}), .clk (clk), .r ({Fresh[227], Fresh[226], Fresh[225]}), .c ({new_AGEMA_signal_2529, new_AGEMA_signal_2528, Midori_rounds_sub_sBox_PRINCE_12_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U5 ( .a ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, Midori_rounds_roundReg_out[50]}), .b ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, Midori_rounds_roundReg_out[51]}), .clk (clk), .r ({Fresh[230], Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, Midori_rounds_sub_sBox_PRINCE_12_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U3 ( .a ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, Midori_rounds_sub_sBox_PRINCE_12_n9}), .b ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, Midori_rounds_sub_sBox_PRINCE_12_n8}), .clk (clk), .r ({Fresh[233], Fresh[232], Fresh[231]}), .c ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, Midori_rounds_sub_sBox_PRINCE_12_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U14 ( .a ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, Midori_rounds_roundReg_out[52]}), .b ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, Midori_rounds_roundReg_out[55]}), .clk (clk), .r ({Fresh[236], Fresh[235], Fresh[234]}), .c ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, Midori_rounds_sub_sBox_PRINCE_13_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U13 ( .a ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, Midori_rounds_sub_sBox_PRINCE_13_n8}), .b ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, Midori_rounds_sub_sBox_PRINCE_13_n7}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237]}), .c ({new_AGEMA_signal_2537, new_AGEMA_signal_2536, Midori_rounds_sub_sBox_PRINCE_13_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U10 ( .a ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, Midori_rounds_roundReg_out[55]}), .b ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, Midori_rounds_sub_sBox_PRINCE_13_n9}), .clk (clk), .r ({Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_2539, new_AGEMA_signal_2538, Midori_rounds_sub_sBox_PRINCE_13_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U9 ( .a ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, Midori_rounds_roundReg_out[54]}), .b ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, Midori_rounds_sub_sBox_PRINCE_13_n8}), .clk (clk), .r ({Fresh[245], Fresh[244], Fresh[243]}), .c ({new_AGEMA_signal_2541, new_AGEMA_signal_2540, Midori_rounds_sub_sBox_PRINCE_13_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U5 ( .a ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, Midori_rounds_roundReg_out[54]}), .b ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, Midori_rounds_roundReg_out[55]}), .clk (clk), .r ({Fresh[248], Fresh[247], Fresh[246]}), .c ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, Midori_rounds_sub_sBox_PRINCE_13_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U3 ( .a ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, Midori_rounds_sub_sBox_PRINCE_13_n9}), .b ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, Midori_rounds_sub_sBox_PRINCE_13_n8}), .clk (clk), .r ({Fresh[251], Fresh[250], Fresh[249]}), .c ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, Midori_rounds_sub_sBox_PRINCE_13_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U14 ( .a ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, Midori_rounds_roundReg_out[56]}), .b ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, Midori_rounds_roundReg_out[59]}), .clk (clk), .r ({Fresh[254], Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, Midori_rounds_sub_sBox_PRINCE_14_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U13 ( .a ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, Midori_rounds_sub_sBox_PRINCE_14_n8}), .b ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, Midori_rounds_sub_sBox_PRINCE_14_n7}), .clk (clk), .r ({Fresh[257], Fresh[256], Fresh[255]}), .c ({new_AGEMA_signal_2549, new_AGEMA_signal_2548, Midori_rounds_sub_sBox_PRINCE_14_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U10 ( .a ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, Midori_rounds_roundReg_out[59]}), .b ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, Midori_rounds_sub_sBox_PRINCE_14_n9}), .clk (clk), .r ({Fresh[260], Fresh[259], Fresh[258]}), .c ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, Midori_rounds_sub_sBox_PRINCE_14_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U9 ( .a ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, Midori_rounds_roundReg_out[58]}), .b ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, Midori_rounds_sub_sBox_PRINCE_14_n8}), .clk (clk), .r ({Fresh[263], Fresh[262], Fresh[261]}), .c ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, Midori_rounds_sub_sBox_PRINCE_14_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U5 ( .a ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, Midori_rounds_roundReg_out[58]}), .b ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, Midori_rounds_roundReg_out[59]}), .clk (clk), .r ({Fresh[266], Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_2099, new_AGEMA_signal_2098, Midori_rounds_sub_sBox_PRINCE_14_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U3 ( .a ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, Midori_rounds_sub_sBox_PRINCE_14_n9}), .b ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, Midori_rounds_sub_sBox_PRINCE_14_n8}), .clk (clk), .r ({Fresh[269], Fresh[268], Fresh[267]}), .c ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, Midori_rounds_sub_sBox_PRINCE_14_n13}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U14 ( .a ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, Midori_rounds_roundReg_out[60]}), .b ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, Midori_rounds_roundReg_out[63]}), .clk (clk), .r ({Fresh[272], Fresh[271], Fresh[270]}), .c ({new_AGEMA_signal_2111, new_AGEMA_signal_2110, Midori_rounds_sub_sBox_PRINCE_15_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U13 ( .a ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, Midori_rounds_sub_sBox_PRINCE_15_n8}), .b ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, Midori_rounds_sub_sBox_PRINCE_15_n7}), .clk (clk), .r ({Fresh[275], Fresh[274], Fresh[273]}), .c ({new_AGEMA_signal_2561, new_AGEMA_signal_2560, Midori_rounds_sub_sBox_PRINCE_15_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U10 ( .a ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, Midori_rounds_roundReg_out[63]}), .b ({new_AGEMA_signal_2121, new_AGEMA_signal_2120, Midori_rounds_sub_sBox_PRINCE_15_n9}), .clk (clk), .r ({Fresh[278], Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, Midori_rounds_sub_sBox_PRINCE_15_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U9 ( .a ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, Midori_rounds_roundReg_out[62]}), .b ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, Midori_rounds_sub_sBox_PRINCE_15_n8}), .clk (clk), .r ({Fresh[281], Fresh[280], Fresh[279]}), .c ({new_AGEMA_signal_2565, new_AGEMA_signal_2564, Midori_rounds_sub_sBox_PRINCE_15_n6}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U5 ( .a ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, Midori_rounds_roundReg_out[62]}), .b ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, Midori_rounds_roundReg_out[63]}), .clk (clk), .r ({Fresh[284], Fresh[283], Fresh[282]}), .c ({new_AGEMA_signal_2115, new_AGEMA_signal_2114, Midori_rounds_sub_sBox_PRINCE_15_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U3 ( .a ({new_AGEMA_signal_2121, new_AGEMA_signal_2120, Midori_rounds_sub_sBox_PRINCE_15_n9}), .b ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, Midori_rounds_sub_sBox_PRINCE_15_n8}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285]}), .c ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, Midori_rounds_sub_sBox_PRINCE_15_n13}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    or_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U18 ( .a ({new_AGEMA_signal_2389, new_AGEMA_signal_2388, Midori_rounds_sub_sBox_PRINCE_0_n13}), .b ({new_AGEMA_signal_2673, new_AGEMA_signal_2672, Midori_rounds_roundReg_out[1]}), .clk (clk), .r ({Fresh[290], Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_2675, new_AGEMA_signal_2674, Midori_rounds_sub_sBox_PRINCE_0_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U15 ( .a ({new_AGEMA_signal_1871, new_AGEMA_signal_1870, Midori_rounds_sub_sBox_PRINCE_0_n10}), .b ({new_AGEMA_signal_1881, new_AGEMA_signal_1880, Midori_rounds_sub_sBox_PRINCE_0_n9}), .clk (clk), .r ({Fresh[293], Fresh[292], Fresh[291]}), .c ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, Midori_rounds_sub_sBox_PRINCE_0_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U11 ( .a ({new_AGEMA_signal_1867, new_AGEMA_signal_1866, Midori_rounds_roundReg_out[0]}), .b ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, Midori_rounds_sub_sBox_PRINCE_0_n4}), .clk (clk), .r ({Fresh[296], Fresh[295], Fresh[294]}), .c ({new_AGEMA_signal_2679, new_AGEMA_signal_2678, Midori_rounds_sub_sBox_PRINCE_0_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U6 ( .a ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, Midori_rounds_sub_sBox_PRINCE_0_n7}), .b ({new_AGEMA_signal_1875, new_AGEMA_signal_1874, Midori_rounds_sub_sBox_PRINCE_0_n1}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297]}), .c ({new_AGEMA_signal_2387, new_AGEMA_signal_2386, Midori_rounds_sub_sBox_PRINCE_0_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U18 ( .a ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, Midori_rounds_sub_sBox_PRINCE_1_n13}), .b ({new_AGEMA_signal_2683, new_AGEMA_signal_2682, Midori_rounds_roundReg_out[5]}), .clk (clk), .r ({Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_2685, new_AGEMA_signal_2684, Midori_rounds_sub_sBox_PRINCE_1_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U15 ( .a ({new_AGEMA_signal_1887, new_AGEMA_signal_1886, Midori_rounds_sub_sBox_PRINCE_1_n10}), .b ({new_AGEMA_signal_1897, new_AGEMA_signal_1896, Midori_rounds_sub_sBox_PRINCE_1_n9}), .clk (clk), .r ({Fresh[305], Fresh[304], Fresh[303]}), .c ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, Midori_rounds_sub_sBox_PRINCE_1_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U11 ( .a ({new_AGEMA_signal_1883, new_AGEMA_signal_1882, Midori_rounds_roundReg_out[4]}), .b ({new_AGEMA_signal_2395, new_AGEMA_signal_2394, Midori_rounds_sub_sBox_PRINCE_1_n4}), .clk (clk), .r ({Fresh[308], Fresh[307], Fresh[306]}), .c ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, Midori_rounds_sub_sBox_PRINCE_1_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U6 ( .a ({new_AGEMA_signal_1893, new_AGEMA_signal_1892, Midori_rounds_sub_sBox_PRINCE_1_n7}), .b ({new_AGEMA_signal_1891, new_AGEMA_signal_1890, Midori_rounds_sub_sBox_PRINCE_1_n1}), .clk (clk), .r ({Fresh[311], Fresh[310], Fresh[309]}), .c ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, Midori_rounds_sub_sBox_PRINCE_1_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U18 ( .a ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, Midori_rounds_sub_sBox_PRINCE_2_n13}), .b ({new_AGEMA_signal_2693, new_AGEMA_signal_2692, Midori_rounds_roundReg_out[9]}), .clk (clk), .r ({Fresh[314], Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_2695, new_AGEMA_signal_2694, Midori_rounds_sub_sBox_PRINCE_2_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U15 ( .a ({new_AGEMA_signal_1903, new_AGEMA_signal_1902, Midori_rounds_sub_sBox_PRINCE_2_n10}), .b ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, Midori_rounds_sub_sBox_PRINCE_2_n9}), .clk (clk), .r ({Fresh[317], Fresh[316], Fresh[315]}), .c ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, Midori_rounds_sub_sBox_PRINCE_2_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U11 ( .a ({new_AGEMA_signal_1899, new_AGEMA_signal_1898, Midori_rounds_roundReg_out[8]}), .b ({new_AGEMA_signal_2407, new_AGEMA_signal_2406, Midori_rounds_sub_sBox_PRINCE_2_n4}), .clk (clk), .r ({Fresh[320], Fresh[319], Fresh[318]}), .c ({new_AGEMA_signal_2699, new_AGEMA_signal_2698, Midori_rounds_sub_sBox_PRINCE_2_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U6 ( .a ({new_AGEMA_signal_1909, new_AGEMA_signal_1908, Midori_rounds_sub_sBox_PRINCE_2_n7}), .b ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, Midori_rounds_sub_sBox_PRINCE_2_n1}), .clk (clk), .r ({Fresh[323], Fresh[322], Fresh[321]}), .c ({new_AGEMA_signal_2411, new_AGEMA_signal_2410, Midori_rounds_sub_sBox_PRINCE_2_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U18 ( .a ({new_AGEMA_signal_2425, new_AGEMA_signal_2424, Midori_rounds_sub_sBox_PRINCE_3_n13}), .b ({new_AGEMA_signal_2703, new_AGEMA_signal_2702, Midori_rounds_roundReg_out[13]}), .clk (clk), .r ({Fresh[326], Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, Midori_rounds_sub_sBox_PRINCE_3_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U15 ( .a ({new_AGEMA_signal_1919, new_AGEMA_signal_1918, Midori_rounds_sub_sBox_PRINCE_3_n10}), .b ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, Midori_rounds_sub_sBox_PRINCE_3_n9}), .clk (clk), .r ({Fresh[329], Fresh[328], Fresh[327]}), .c ({new_AGEMA_signal_2415, new_AGEMA_signal_2414, Midori_rounds_sub_sBox_PRINCE_3_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U11 ( .a ({new_AGEMA_signal_1915, new_AGEMA_signal_1914, Midori_rounds_roundReg_out[12]}), .b ({new_AGEMA_signal_2419, new_AGEMA_signal_2418, Midori_rounds_sub_sBox_PRINCE_3_n4}), .clk (clk), .r ({Fresh[332], Fresh[331], Fresh[330]}), .c ({new_AGEMA_signal_2709, new_AGEMA_signal_2708, Midori_rounds_sub_sBox_PRINCE_3_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U6 ( .a ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, Midori_rounds_sub_sBox_PRINCE_3_n7}), .b ({new_AGEMA_signal_1923, new_AGEMA_signal_1922, Midori_rounds_sub_sBox_PRINCE_3_n1}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333]}), .c ({new_AGEMA_signal_2423, new_AGEMA_signal_2422, Midori_rounds_sub_sBox_PRINCE_3_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U18 ( .a ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, Midori_rounds_sub_sBox_PRINCE_4_n13}), .b ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, Midori_rounds_roundReg_out[17]}), .clk (clk), .r ({Fresh[338], Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_2715, new_AGEMA_signal_2714, Midori_rounds_sub_sBox_PRINCE_4_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U15 ( .a ({new_AGEMA_signal_1935, new_AGEMA_signal_1934, Midori_rounds_sub_sBox_PRINCE_4_n10}), .b ({new_AGEMA_signal_1945, new_AGEMA_signal_1944, Midori_rounds_sub_sBox_PRINCE_4_n9}), .clk (clk), .r ({Fresh[341], Fresh[340], Fresh[339]}), .c ({new_AGEMA_signal_2427, new_AGEMA_signal_2426, Midori_rounds_sub_sBox_PRINCE_4_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U11 ( .a ({new_AGEMA_signal_1931, new_AGEMA_signal_1930, Midori_rounds_roundReg_out[16]}), .b ({new_AGEMA_signal_2431, new_AGEMA_signal_2430, Midori_rounds_sub_sBox_PRINCE_4_n4}), .clk (clk), .r ({Fresh[344], Fresh[343], Fresh[342]}), .c ({new_AGEMA_signal_2719, new_AGEMA_signal_2718, Midori_rounds_sub_sBox_PRINCE_4_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U6 ( .a ({new_AGEMA_signal_1941, new_AGEMA_signal_1940, Midori_rounds_sub_sBox_PRINCE_4_n7}), .b ({new_AGEMA_signal_1939, new_AGEMA_signal_1938, Midori_rounds_sub_sBox_PRINCE_4_n1}), .clk (clk), .r ({Fresh[347], Fresh[346], Fresh[345]}), .c ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, Midori_rounds_sub_sBox_PRINCE_4_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U18 ( .a ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, Midori_rounds_sub_sBox_PRINCE_5_n13}), .b ({new_AGEMA_signal_2723, new_AGEMA_signal_2722, Midori_rounds_roundReg_out[21]}), .clk (clk), .r ({Fresh[350], Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, Midori_rounds_sub_sBox_PRINCE_5_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U15 ( .a ({new_AGEMA_signal_1951, new_AGEMA_signal_1950, Midori_rounds_sub_sBox_PRINCE_5_n10}), .b ({new_AGEMA_signal_1961, new_AGEMA_signal_1960, Midori_rounds_sub_sBox_PRINCE_5_n9}), .clk (clk), .r ({Fresh[353], Fresh[352], Fresh[351]}), .c ({new_AGEMA_signal_2439, new_AGEMA_signal_2438, Midori_rounds_sub_sBox_PRINCE_5_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U11 ( .a ({new_AGEMA_signal_1947, new_AGEMA_signal_1946, Midori_rounds_roundReg_out[20]}), .b ({new_AGEMA_signal_2443, new_AGEMA_signal_2442, Midori_rounds_sub_sBox_PRINCE_5_n4}), .clk (clk), .r ({Fresh[356], Fresh[355], Fresh[354]}), .c ({new_AGEMA_signal_2729, new_AGEMA_signal_2728, Midori_rounds_sub_sBox_PRINCE_5_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U6 ( .a ({new_AGEMA_signal_1957, new_AGEMA_signal_1956, Midori_rounds_sub_sBox_PRINCE_5_n7}), .b ({new_AGEMA_signal_1955, new_AGEMA_signal_1954, Midori_rounds_sub_sBox_PRINCE_5_n1}), .clk (clk), .r ({Fresh[359], Fresh[358], Fresh[357]}), .c ({new_AGEMA_signal_2447, new_AGEMA_signal_2446, Midori_rounds_sub_sBox_PRINCE_5_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U18 ( .a ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, Midori_rounds_sub_sBox_PRINCE_6_n13}), .b ({new_AGEMA_signal_2733, new_AGEMA_signal_2732, Midori_rounds_roundReg_out[25]}), .clk (clk), .r ({Fresh[362], Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_2735, new_AGEMA_signal_2734, Midori_rounds_sub_sBox_PRINCE_6_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U15 ( .a ({new_AGEMA_signal_1967, new_AGEMA_signal_1966, Midori_rounds_sub_sBox_PRINCE_6_n10}), .b ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, Midori_rounds_sub_sBox_PRINCE_6_n9}), .clk (clk), .r ({Fresh[365], Fresh[364], Fresh[363]}), .c ({new_AGEMA_signal_2451, new_AGEMA_signal_2450, Midori_rounds_sub_sBox_PRINCE_6_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U11 ( .a ({new_AGEMA_signal_1963, new_AGEMA_signal_1962, Midori_rounds_roundReg_out[24]}), .b ({new_AGEMA_signal_2455, new_AGEMA_signal_2454, Midori_rounds_sub_sBox_PRINCE_6_n4}), .clk (clk), .r ({Fresh[368], Fresh[367], Fresh[366]}), .c ({new_AGEMA_signal_2739, new_AGEMA_signal_2738, Midori_rounds_sub_sBox_PRINCE_6_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U6 ( .a ({new_AGEMA_signal_1973, new_AGEMA_signal_1972, Midori_rounds_sub_sBox_PRINCE_6_n7}), .b ({new_AGEMA_signal_1971, new_AGEMA_signal_1970, Midori_rounds_sub_sBox_PRINCE_6_n1}), .clk (clk), .r ({Fresh[371], Fresh[370], Fresh[369]}), .c ({new_AGEMA_signal_2459, new_AGEMA_signal_2458, Midori_rounds_sub_sBox_PRINCE_6_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U18 ( .a ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, Midori_rounds_sub_sBox_PRINCE_7_n13}), .b ({new_AGEMA_signal_2743, new_AGEMA_signal_2742, Midori_rounds_roundReg_out[29]}), .clk (clk), .r ({Fresh[374], Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_2745, new_AGEMA_signal_2744, Midori_rounds_sub_sBox_PRINCE_7_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U15 ( .a ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, Midori_rounds_sub_sBox_PRINCE_7_n10}), .b ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, Midori_rounds_sub_sBox_PRINCE_7_n9}), .clk (clk), .r ({Fresh[377], Fresh[376], Fresh[375]}), .c ({new_AGEMA_signal_2463, new_AGEMA_signal_2462, Midori_rounds_sub_sBox_PRINCE_7_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U11 ( .a ({new_AGEMA_signal_1979, new_AGEMA_signal_1978, Midori_rounds_roundReg_out[28]}), .b ({new_AGEMA_signal_2467, new_AGEMA_signal_2466, Midori_rounds_sub_sBox_PRINCE_7_n4}), .clk (clk), .r ({Fresh[380], Fresh[379], Fresh[378]}), .c ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, Midori_rounds_sub_sBox_PRINCE_7_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U6 ( .a ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, Midori_rounds_sub_sBox_PRINCE_7_n7}), .b ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, Midori_rounds_sub_sBox_PRINCE_7_n1}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381]}), .c ({new_AGEMA_signal_2471, new_AGEMA_signal_2470, Midori_rounds_sub_sBox_PRINCE_7_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U18 ( .a ({new_AGEMA_signal_2485, new_AGEMA_signal_2484, Midori_rounds_sub_sBox_PRINCE_8_n13}), .b ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, Midori_rounds_roundReg_out[33]}), .clk (clk), .r ({Fresh[386], Fresh[385], Fresh[384]}), .c ({new_AGEMA_signal_2755, new_AGEMA_signal_2754, Midori_rounds_sub_sBox_PRINCE_8_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U15 ( .a ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, Midori_rounds_sub_sBox_PRINCE_8_n10}), .b ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, Midori_rounds_sub_sBox_PRINCE_8_n9}), .clk (clk), .r ({Fresh[389], Fresh[388], Fresh[387]}), .c ({new_AGEMA_signal_2475, new_AGEMA_signal_2474, Midori_rounds_sub_sBox_PRINCE_8_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U11 ( .a ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, Midori_rounds_roundReg_out[32]}), .b ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, Midori_rounds_sub_sBox_PRINCE_8_n4}), .clk (clk), .r ({Fresh[392], Fresh[391], Fresh[390]}), .c ({new_AGEMA_signal_2759, new_AGEMA_signal_2758, Midori_rounds_sub_sBox_PRINCE_8_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U6 ( .a ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, Midori_rounds_sub_sBox_PRINCE_8_n7}), .b ({new_AGEMA_signal_2003, new_AGEMA_signal_2002, Midori_rounds_sub_sBox_PRINCE_8_n1}), .clk (clk), .r ({Fresh[395], Fresh[394], Fresh[393]}), .c ({new_AGEMA_signal_2483, new_AGEMA_signal_2482, Midori_rounds_sub_sBox_PRINCE_8_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U18 ( .a ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, Midori_rounds_sub_sBox_PRINCE_9_n13}), .b ({new_AGEMA_signal_2763, new_AGEMA_signal_2762, Midori_rounds_roundReg_out[37]}), .clk (clk), .r ({Fresh[398], Fresh[397], Fresh[396]}), .c ({new_AGEMA_signal_2765, new_AGEMA_signal_2764, Midori_rounds_sub_sBox_PRINCE_9_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U15 ( .a ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, Midori_rounds_sub_sBox_PRINCE_9_n10}), .b ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, Midori_rounds_sub_sBox_PRINCE_9_n9}), .clk (clk), .r ({Fresh[401], Fresh[400], Fresh[399]}), .c ({new_AGEMA_signal_2487, new_AGEMA_signal_2486, Midori_rounds_sub_sBox_PRINCE_9_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U11 ( .a ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, Midori_rounds_roundReg_out[36]}), .b ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, Midori_rounds_sub_sBox_PRINCE_9_n4}), .clk (clk), .r ({Fresh[404], Fresh[403], Fresh[402]}), .c ({new_AGEMA_signal_2769, new_AGEMA_signal_2768, Midori_rounds_sub_sBox_PRINCE_9_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U6 ( .a ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, Midori_rounds_sub_sBox_PRINCE_9_n7}), .b ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, Midori_rounds_sub_sBox_PRINCE_9_n1}), .clk (clk), .r ({Fresh[407], Fresh[406], Fresh[405]}), .c ({new_AGEMA_signal_2495, new_AGEMA_signal_2494, Midori_rounds_sub_sBox_PRINCE_9_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U18 ( .a ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, Midori_rounds_sub_sBox_PRINCE_10_n13}), .b ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, Midori_rounds_roundReg_out[41]}), .clk (clk), .r ({Fresh[410], Fresh[409], Fresh[408]}), .c ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, Midori_rounds_sub_sBox_PRINCE_10_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U15 ( .a ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, Midori_rounds_sub_sBox_PRINCE_10_n10}), .b ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, Midori_rounds_sub_sBox_PRINCE_10_n9}), .clk (clk), .r ({Fresh[413], Fresh[412], Fresh[411]}), .c ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, Midori_rounds_sub_sBox_PRINCE_10_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U11 ( .a ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, Midori_rounds_roundReg_out[40]}), .b ({new_AGEMA_signal_2503, new_AGEMA_signal_2502, Midori_rounds_sub_sBox_PRINCE_10_n4}), .clk (clk), .r ({Fresh[416], Fresh[415], Fresh[414]}), .c ({new_AGEMA_signal_2779, new_AGEMA_signal_2778, Midori_rounds_sub_sBox_PRINCE_10_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U6 ( .a ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, Midori_rounds_sub_sBox_PRINCE_10_n7}), .b ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, Midori_rounds_sub_sBox_PRINCE_10_n1}), .clk (clk), .r ({Fresh[419], Fresh[418], Fresh[417]}), .c ({new_AGEMA_signal_2507, new_AGEMA_signal_2506, Midori_rounds_sub_sBox_PRINCE_10_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U18 ( .a ({new_AGEMA_signal_2521, new_AGEMA_signal_2520, Midori_rounds_sub_sBox_PRINCE_11_n13}), .b ({new_AGEMA_signal_2783, new_AGEMA_signal_2782, Midori_rounds_roundReg_out[45]}), .clk (clk), .r ({Fresh[422], Fresh[421], Fresh[420]}), .c ({new_AGEMA_signal_2785, new_AGEMA_signal_2784, Midori_rounds_sub_sBox_PRINCE_11_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U15 ( .a ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, Midori_rounds_sub_sBox_PRINCE_11_n10}), .b ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, Midori_rounds_sub_sBox_PRINCE_11_n9}), .clk (clk), .r ({Fresh[425], Fresh[424], Fresh[423]}), .c ({new_AGEMA_signal_2511, new_AGEMA_signal_2510, Midori_rounds_sub_sBox_PRINCE_11_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U11 ( .a ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, Midori_rounds_roundReg_out[44]}), .b ({new_AGEMA_signal_2515, new_AGEMA_signal_2514, Midori_rounds_sub_sBox_PRINCE_11_n4}), .clk (clk), .r ({Fresh[428], Fresh[427], Fresh[426]}), .c ({new_AGEMA_signal_2789, new_AGEMA_signal_2788, Midori_rounds_sub_sBox_PRINCE_11_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U6 ( .a ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, Midori_rounds_sub_sBox_PRINCE_11_n7}), .b ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, Midori_rounds_sub_sBox_PRINCE_11_n1}), .clk (clk), .r ({Fresh[431], Fresh[430], Fresh[429]}), .c ({new_AGEMA_signal_2519, new_AGEMA_signal_2518, Midori_rounds_sub_sBox_PRINCE_11_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U18 ( .a ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, Midori_rounds_sub_sBox_PRINCE_12_n13}), .b ({new_AGEMA_signal_2793, new_AGEMA_signal_2792, Midori_rounds_roundReg_out[49]}), .clk (clk), .r ({Fresh[434], Fresh[433], Fresh[432]}), .c ({new_AGEMA_signal_2795, new_AGEMA_signal_2794, Midori_rounds_sub_sBox_PRINCE_12_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U15 ( .a ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, Midori_rounds_sub_sBox_PRINCE_12_n10}), .b ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, Midori_rounds_sub_sBox_PRINCE_12_n9}), .clk (clk), .r ({Fresh[437], Fresh[436], Fresh[435]}), .c ({new_AGEMA_signal_2523, new_AGEMA_signal_2522, Midori_rounds_sub_sBox_PRINCE_12_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U11 ( .a ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, Midori_rounds_roundReg_out[48]}), .b ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, Midori_rounds_sub_sBox_PRINCE_12_n4}), .clk (clk), .r ({Fresh[440], Fresh[439], Fresh[438]}), .c ({new_AGEMA_signal_2799, new_AGEMA_signal_2798, Midori_rounds_sub_sBox_PRINCE_12_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U6 ( .a ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, Midori_rounds_sub_sBox_PRINCE_12_n7}), .b ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, Midori_rounds_sub_sBox_PRINCE_12_n1}), .clk (clk), .r ({Fresh[443], Fresh[442], Fresh[441]}), .c ({new_AGEMA_signal_2531, new_AGEMA_signal_2530, Midori_rounds_sub_sBox_PRINCE_12_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U18 ( .a ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, Midori_rounds_sub_sBox_PRINCE_13_n13}), .b ({new_AGEMA_signal_2803, new_AGEMA_signal_2802, Midori_rounds_roundReg_out[53]}), .clk (clk), .r ({Fresh[446], Fresh[445], Fresh[444]}), .c ({new_AGEMA_signal_2805, new_AGEMA_signal_2804, Midori_rounds_sub_sBox_PRINCE_13_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U15 ( .a ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, Midori_rounds_sub_sBox_PRINCE_13_n10}), .b ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, Midori_rounds_sub_sBox_PRINCE_13_n9}), .clk (clk), .r ({Fresh[449], Fresh[448], Fresh[447]}), .c ({new_AGEMA_signal_2535, new_AGEMA_signal_2534, Midori_rounds_sub_sBox_PRINCE_13_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U11 ( .a ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, Midori_rounds_roundReg_out[52]}), .b ({new_AGEMA_signal_2539, new_AGEMA_signal_2538, Midori_rounds_sub_sBox_PRINCE_13_n4}), .clk (clk), .r ({Fresh[452], Fresh[451], Fresh[450]}), .c ({new_AGEMA_signal_2809, new_AGEMA_signal_2808, Midori_rounds_sub_sBox_PRINCE_13_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U6 ( .a ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, Midori_rounds_sub_sBox_PRINCE_13_n7}), .b ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, Midori_rounds_sub_sBox_PRINCE_13_n1}), .clk (clk), .r ({Fresh[455], Fresh[454], Fresh[453]}), .c ({new_AGEMA_signal_2543, new_AGEMA_signal_2542, Midori_rounds_sub_sBox_PRINCE_13_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U18 ( .a ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, Midori_rounds_sub_sBox_PRINCE_14_n13}), .b ({new_AGEMA_signal_2813, new_AGEMA_signal_2812, Midori_rounds_roundReg_out[57]}), .clk (clk), .r ({Fresh[458], Fresh[457], Fresh[456]}), .c ({new_AGEMA_signal_2815, new_AGEMA_signal_2814, Midori_rounds_sub_sBox_PRINCE_14_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U15 ( .a ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, Midori_rounds_sub_sBox_PRINCE_14_n10}), .b ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, Midori_rounds_sub_sBox_PRINCE_14_n9}), .clk (clk), .r ({Fresh[461], Fresh[460], Fresh[459]}), .c ({new_AGEMA_signal_2547, new_AGEMA_signal_2546, Midori_rounds_sub_sBox_PRINCE_14_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U11 ( .a ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, Midori_rounds_roundReg_out[56]}), .b ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, Midori_rounds_sub_sBox_PRINCE_14_n4}), .clk (clk), .r ({Fresh[464], Fresh[463], Fresh[462]}), .c ({new_AGEMA_signal_2819, new_AGEMA_signal_2818, Midori_rounds_sub_sBox_PRINCE_14_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U6 ( .a ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, Midori_rounds_sub_sBox_PRINCE_14_n7}), .b ({new_AGEMA_signal_2099, new_AGEMA_signal_2098, Midori_rounds_sub_sBox_PRINCE_14_n1}), .clk (clk), .r ({Fresh[467], Fresh[466], Fresh[465]}), .c ({new_AGEMA_signal_2555, new_AGEMA_signal_2554, Midori_rounds_sub_sBox_PRINCE_14_n2}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U18 ( .a ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, Midori_rounds_sub_sBox_PRINCE_15_n13}), .b ({new_AGEMA_signal_2823, new_AGEMA_signal_2822, Midori_rounds_roundReg_out[61]}), .clk (clk), .r ({Fresh[470], Fresh[469], Fresh[468]}), .c ({new_AGEMA_signal_2825, new_AGEMA_signal_2824, Midori_rounds_sub_sBox_PRINCE_15_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U15 ( .a ({new_AGEMA_signal_2111, new_AGEMA_signal_2110, Midori_rounds_sub_sBox_PRINCE_15_n10}), .b ({new_AGEMA_signal_2121, new_AGEMA_signal_2120, Midori_rounds_sub_sBox_PRINCE_15_n9}), .clk (clk), .r ({Fresh[473], Fresh[472], Fresh[471]}), .c ({new_AGEMA_signal_2559, new_AGEMA_signal_2558, Midori_rounds_sub_sBox_PRINCE_15_n11}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U11 ( .a ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, Midori_rounds_roundReg_out[60]}), .b ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, Midori_rounds_sub_sBox_PRINCE_15_n4}), .clk (clk), .r ({Fresh[476], Fresh[475], Fresh[474]}), .c ({new_AGEMA_signal_2829, new_AGEMA_signal_2828, Midori_rounds_sub_sBox_PRINCE_15_n5}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U6 ( .a ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, Midori_rounds_sub_sBox_PRINCE_15_n7}), .b ({new_AGEMA_signal_2115, new_AGEMA_signal_2114, Midori_rounds_sub_sBox_PRINCE_15_n1}), .clk (clk), .r ({Fresh[479], Fresh[478], Fresh[477]}), .c ({new_AGEMA_signal_2567, new_AGEMA_signal_2566, Midori_rounds_sub_sBox_PRINCE_15_n2}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U128 ( .a ({new_AGEMA_signal_1461, new_AGEMA_signal_1460, wk[9]}), .b ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, Midori_rounds_SR_Result[9]}), .c ({DataOut_s2[9], DataOut_s1[9], DataOut_s0[9]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U126 ( .a ({new_AGEMA_signal_1473, new_AGEMA_signal_1472, wk[7]}), .b ({new_AGEMA_signal_2841, new_AGEMA_signal_2840, Midori_rounds_SR_Result[47]}), .c ({DataOut_s2[7], DataOut_s1[7], DataOut_s0[7]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U124 ( .a ({new_AGEMA_signal_1485, new_AGEMA_signal_1484, wk[63]}), .b ({new_AGEMA_signal_2953, new_AGEMA_signal_2952, Midori_rounds_SR_Result[63]}), .c ({DataOut_s2[63], DataOut_s1[63], DataOut_s0[63]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U122 ( .a ({new_AGEMA_signal_1497, new_AGEMA_signal_1496, wk[61]}), .b ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, Midori_rounds_SR_Result[61]}), .c ({DataOut_s2[61], DataOut_s1[61], DataOut_s0[61]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U120 ( .a ({new_AGEMA_signal_1509, new_AGEMA_signal_1508, wk[5]}), .b ({new_AGEMA_signal_2845, new_AGEMA_signal_2844, Midori_rounds_SR_Result[45]}), .c ({DataOut_s2[5], DataOut_s1[5], DataOut_s0[5]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U119 ( .a ({new_AGEMA_signal_1515, new_AGEMA_signal_1514, wk[59]}), .b ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, Midori_rounds_SR_Result[35]}), .c ({DataOut_s2[59], DataOut_s1[59], DataOut_s0[59]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U117 ( .a ({new_AGEMA_signal_1527, new_AGEMA_signal_1526, wk[57]}), .b ({new_AGEMA_signal_2949, new_AGEMA_signal_2948, Midori_rounds_SR_Result[33]}), .c ({DataOut_s2[57], DataOut_s1[57], DataOut_s0[57]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U115 ( .a ({new_AGEMA_signal_1539, new_AGEMA_signal_1538, wk[55]}), .b ({new_AGEMA_signal_2937, new_AGEMA_signal_2936, Midori_rounds_SR_Result[7]}), .c ({DataOut_s2[55], DataOut_s1[55], DataOut_s0[55]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U113 ( .a ({new_AGEMA_signal_1551, new_AGEMA_signal_1550, wk[53]}), .b ({new_AGEMA_signal_2941, new_AGEMA_signal_2940, Midori_rounds_SR_Result[5]}), .c ({DataOut_s2[53], DataOut_s1[53], DataOut_s0[53]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U111 ( .a ({new_AGEMA_signal_1563, new_AGEMA_signal_1562, wk[51]}), .b ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, Midori_rounds_SR_Result[27]}), .c ({DataOut_s2[51], DataOut_s1[51], DataOut_s0[51]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U108 ( .a ({new_AGEMA_signal_1581, new_AGEMA_signal_1580, wk[49]}), .b ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, Midori_rounds_SR_Result[25]}), .c ({DataOut_s2[49], DataOut_s1[49], DataOut_s0[49]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U106 ( .a ({new_AGEMA_signal_1593, new_AGEMA_signal_1592, wk[47]}), .b ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, Midori_rounds_SR_Result[43]}), .c ({DataOut_s2[47], DataOut_s1[47], DataOut_s0[47]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U104 ( .a ({new_AGEMA_signal_1605, new_AGEMA_signal_1604, wk[45]}), .b ({new_AGEMA_signal_2925, new_AGEMA_signal_2924, Midori_rounds_SR_Result[41]}), .c ({DataOut_s2[45], DataOut_s1[45], DataOut_s0[45]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U102 ( .a ({new_AGEMA_signal_1617, new_AGEMA_signal_1616, wk[43]}), .b ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, Midori_rounds_SR_Result[55]}), .c ({DataOut_s2[43], DataOut_s1[43], DataOut_s0[43]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U100 ( .a ({new_AGEMA_signal_1629, new_AGEMA_signal_1628, wk[41]}), .b ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, Midori_rounds_SR_Result[53]}), .c ({DataOut_s2[41], DataOut_s1[41], DataOut_s0[41]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U98 ( .a ({new_AGEMA_signal_1641, new_AGEMA_signal_1640, wk[3]}), .b ({new_AGEMA_signal_2833, new_AGEMA_signal_2832, Midori_rounds_SR_Result[51]}), .c ({DataOut_s2[3], DataOut_s1[3], DataOut_s0[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U97 ( .a ({new_AGEMA_signal_1647, new_AGEMA_signal_1646, wk[39]}), .b ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, Midori_rounds_SR_Result[19]}), .c ({DataOut_s2[39], DataOut_s1[39], DataOut_s0[39]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U95 ( .a ({new_AGEMA_signal_1659, new_AGEMA_signal_1658, wk[37]}), .b ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, Midori_rounds_SR_Result[17]}), .c ({DataOut_s2[37], DataOut_s1[37], DataOut_s0[37]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U93 ( .a ({new_AGEMA_signal_1671, new_AGEMA_signal_1670, wk[35]}), .b ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, Midori_rounds_SR_Result[15]}), .c ({DataOut_s2[35], DataOut_s1[35], DataOut_s0[35]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U91 ( .a ({new_AGEMA_signal_1683, new_AGEMA_signal_1682, wk[33]}), .b ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, Midori_rounds_SR_Result[13]}), .c ({DataOut_s2[33], DataOut_s1[33], DataOut_s0[33]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U89 ( .a ({new_AGEMA_signal_1695, new_AGEMA_signal_1694, wk[31]}), .b ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, Midori_rounds_SR_Result[3]}), .c ({DataOut_s2[31], DataOut_s1[31], DataOut_s0[31]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U86 ( .a ({new_AGEMA_signal_1713, new_AGEMA_signal_1712, wk[29]}), .b ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, Midori_rounds_SR_Result[1]}), .c ({DataOut_s2[29], DataOut_s1[29], DataOut_s0[29]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U84 ( .a ({new_AGEMA_signal_1725, new_AGEMA_signal_1724, wk[27]}), .b ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, Midori_rounds_SR_Result[31]}), .c ({DataOut_s2[27], DataOut_s1[27], DataOut_s0[27]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U82 ( .a ({new_AGEMA_signal_1737, new_AGEMA_signal_1736, wk[25]}), .b ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, Midori_rounds_SR_Result[29]}), .c ({DataOut_s2[25], DataOut_s1[25], DataOut_s0[25]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U80 ( .a ({new_AGEMA_signal_1749, new_AGEMA_signal_1748, wk[23]}), .b ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, Midori_rounds_SR_Result[59]}), .c ({DataOut_s2[23], DataOut_s1[23], DataOut_s0[23]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U78 ( .a ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, wk[21]}), .b ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, Midori_rounds_SR_Result[57]}), .c ({DataOut_s2[21], DataOut_s1[21], DataOut_s0[21]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U76 ( .a ({new_AGEMA_signal_1773, new_AGEMA_signal_1772, wk[1]}), .b ({new_AGEMA_signal_2837, new_AGEMA_signal_2836, Midori_rounds_SR_Result[49]}), .c ({DataOut_s2[1], DataOut_s1[1], DataOut_s0[1]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U75 ( .a ({new_AGEMA_signal_1779, new_AGEMA_signal_1778, wk[19]}), .b ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, Midori_rounds_SR_Result[39]}), .c ({DataOut_s2[19], DataOut_s1[19], DataOut_s0[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U73 ( .a ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, wk[17]}), .b ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, Midori_rounds_SR_Result[37]}), .c ({DataOut_s2[17], DataOut_s1[17], DataOut_s0[17]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U71 ( .a ({new_AGEMA_signal_1803, new_AGEMA_signal_1802, wk[15]}), .b ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, Midori_rounds_SR_Result[23]}), .c ({DataOut_s2[15], DataOut_s1[15], DataOut_s0[15]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U69 ( .a ({new_AGEMA_signal_1815, new_AGEMA_signal_1814, wk[13]}), .b ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, Midori_rounds_SR_Result[21]}), .c ({DataOut_s2[13], DataOut_s1[13], DataOut_s0[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U67 ( .a ({new_AGEMA_signal_1827, new_AGEMA_signal_1826, wk[11]}), .b ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, Midori_rounds_SR_Result[11]}), .c ({DataOut_s2[11], DataOut_s1[11], DataOut_s0[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U144 ( .a ({new_AGEMA_signal_1853, new_AGEMA_signal_1852, Midori_rounds_SelectedKey_9_}), .b ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, Midori_rounds_SR_Result[9]}), .c ({new_AGEMA_signal_3089, new_AGEMA_signal_3088, Midori_rounds_sub_ResultXORkey[9]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U142 ( .a ({new_AGEMA_signal_2575, new_AGEMA_signal_2574, Midori_rounds_SelectedKey_7_}), .b ({new_AGEMA_signal_2841, new_AGEMA_signal_2840, Midori_rounds_SR_Result[47]}), .c ({new_AGEMA_signal_3091, new_AGEMA_signal_3090, Midori_rounds_sub_ResultXORkey[7]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U140 ( .a ({new_AGEMA_signal_2671, new_AGEMA_signal_2670, Midori_rounds_SelectedKey_63_}), .b ({new_AGEMA_signal_2953, new_AGEMA_signal_2952, Midori_rounds_SR_Result[63]}), .c ({new_AGEMA_signal_3095, new_AGEMA_signal_3094, Midori_rounds_sub_ResultXORkey[63]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U138 ( .a ({new_AGEMA_signal_2667, new_AGEMA_signal_2666, Midori_rounds_SelectedKey_61_}), .b ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, Midori_rounds_SR_Result[61]}), .c ({new_AGEMA_signal_3099, new_AGEMA_signal_3098, Midori_rounds_sub_ResultXORkey[61]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U136 ( .a ({new_AGEMA_signal_2571, new_AGEMA_signal_2570, Midori_rounds_SelectedKey_5_}), .b ({new_AGEMA_signal_2845, new_AGEMA_signal_2844, Midori_rounds_SR_Result[45]}), .c ({new_AGEMA_signal_3101, new_AGEMA_signal_3100, Midori_rounds_sub_ResultXORkey[5]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U135 ( .a ({new_AGEMA_signal_2663, new_AGEMA_signal_2662, Midori_rounds_SelectedKey_59_}), .b ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, Midori_rounds_SR_Result[35]}), .c ({new_AGEMA_signal_3103, new_AGEMA_signal_3102, Midori_rounds_sub_ResultXORkey[59]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U133 ( .a ({new_AGEMA_signal_2659, new_AGEMA_signal_2658, Midori_rounds_SelectedKey_57_}), .b ({new_AGEMA_signal_2949, new_AGEMA_signal_2948, Midori_rounds_SR_Result[33]}), .c ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, Midori_rounds_sub_ResultXORkey[57]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U131 ( .a ({new_AGEMA_signal_2655, new_AGEMA_signal_2654, Midori_rounds_SelectedKey_55_}), .b ({new_AGEMA_signal_2937, new_AGEMA_signal_2936, Midori_rounds_SR_Result[7]}), .c ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, Midori_rounds_sub_ResultXORkey[55]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U129 ( .a ({new_AGEMA_signal_2651, new_AGEMA_signal_2650, Midori_rounds_SelectedKey_53_}), .b ({new_AGEMA_signal_2941, new_AGEMA_signal_2940, Midori_rounds_SR_Result[5]}), .c ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, Midori_rounds_sub_ResultXORkey[53]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U127 ( .a ({new_AGEMA_signal_2647, new_AGEMA_signal_2646, Midori_rounds_SelectedKey_51_}), .b ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, Midori_rounds_SR_Result[27]}), .c ({new_AGEMA_signal_3115, new_AGEMA_signal_3114, Midori_rounds_sub_ResultXORkey[51]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U124 ( .a ({new_AGEMA_signal_2643, new_AGEMA_signal_2642, Midori_rounds_SelectedKey_49_}), .b ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, Midori_rounds_SR_Result[25]}), .c ({new_AGEMA_signal_3119, new_AGEMA_signal_3118, Midori_rounds_sub_ResultXORkey[49]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U122 ( .a ({new_AGEMA_signal_2639, new_AGEMA_signal_2638, Midori_rounds_SelectedKey_47_}), .b ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, Midori_rounds_SR_Result[43]}), .c ({new_AGEMA_signal_3121, new_AGEMA_signal_3120, Midori_rounds_sub_ResultXORkey[47]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U120 ( .a ({new_AGEMA_signal_2635, new_AGEMA_signal_2634, Midori_rounds_SelectedKey_45_}), .b ({new_AGEMA_signal_2925, new_AGEMA_signal_2924, Midori_rounds_SR_Result[41]}), .c ({new_AGEMA_signal_3125, new_AGEMA_signal_3124, Midori_rounds_sub_ResultXORkey[45]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U118 ( .a ({new_AGEMA_signal_2631, new_AGEMA_signal_2630, Midori_rounds_SelectedKey_43_}), .b ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, Midori_rounds_SR_Result[55]}), .c ({new_AGEMA_signal_3127, new_AGEMA_signal_3126, Midori_rounds_sub_ResultXORkey[43]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U116 ( .a ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, Midori_rounds_SelectedKey_41_}), .b ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, Midori_rounds_SR_Result[53]}), .c ({new_AGEMA_signal_3131, new_AGEMA_signal_3130, Midori_rounds_sub_ResultXORkey[41]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U114 ( .a ({new_AGEMA_signal_1847, new_AGEMA_signal_1846, Midori_rounds_SelectedKey_3_}), .b ({new_AGEMA_signal_2833, new_AGEMA_signal_2832, Midori_rounds_SR_Result[51]}), .c ({new_AGEMA_signal_3133, new_AGEMA_signal_3132, Midori_rounds_sub_ResultXORkey[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U113 ( .a ({new_AGEMA_signal_2623, new_AGEMA_signal_2622, Midori_rounds_SelectedKey_39_}), .b ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, Midori_rounds_SR_Result[19]}), .c ({new_AGEMA_signal_3135, new_AGEMA_signal_3134, Midori_rounds_sub_ResultXORkey[39]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U111 ( .a ({new_AGEMA_signal_2619, new_AGEMA_signal_2618, Midori_rounds_SelectedKey_37_}), .b ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, Midori_rounds_SR_Result[17]}), .c ({new_AGEMA_signal_3139, new_AGEMA_signal_3138, Midori_rounds_sub_ResultXORkey[37]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U109 ( .a ({new_AGEMA_signal_2615, new_AGEMA_signal_2614, Midori_rounds_SelectedKey_35_}), .b ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, Midori_rounds_SR_Result[15]}), .c ({new_AGEMA_signal_3141, new_AGEMA_signal_3140, Midori_rounds_sub_ResultXORkey[35]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U107 ( .a ({new_AGEMA_signal_2611, new_AGEMA_signal_2610, Midori_rounds_SelectedKey_33_}), .b ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, Midori_rounds_SR_Result[13]}), .c ({new_AGEMA_signal_3145, new_AGEMA_signal_3144, Midori_rounds_sub_ResultXORkey[33]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U105 ( .a ({new_AGEMA_signal_2607, new_AGEMA_signal_2606, Midori_rounds_SelectedKey_31_}), .b ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, Midori_rounds_SR_Result[3]}), .c ({new_AGEMA_signal_3147, new_AGEMA_signal_3146, Midori_rounds_sub_ResultXORkey[31]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U102 ( .a ({new_AGEMA_signal_2603, new_AGEMA_signal_2602, Midori_rounds_SelectedKey_29_}), .b ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, Midori_rounds_SR_Result[1]}), .c ({new_AGEMA_signal_3153, new_AGEMA_signal_3152, Midori_rounds_sub_ResultXORkey[29]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U100 ( .a ({new_AGEMA_signal_2599, new_AGEMA_signal_2598, Midori_rounds_SelectedKey_27_}), .b ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, Midori_rounds_SR_Result[31]}), .c ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, Midori_rounds_sub_ResultXORkey[27]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U98 ( .a ({new_AGEMA_signal_2597, new_AGEMA_signal_2596, Midori_rounds_SelectedKey_25_}), .b ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, Midori_rounds_SR_Result[29]}), .c ({new_AGEMA_signal_3159, new_AGEMA_signal_3158, Midori_rounds_sub_ResultXORkey[25]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U96 ( .a ({new_AGEMA_signal_2593, new_AGEMA_signal_2592, Midori_rounds_SelectedKey_23_}), .b ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, Midori_rounds_SR_Result[59]}), .c ({new_AGEMA_signal_3161, new_AGEMA_signal_3160, Midori_rounds_sub_ResultXORkey[23]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U94 ( .a ({new_AGEMA_signal_2589, new_AGEMA_signal_2588, Midori_rounds_SelectedKey_21_}), .b ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, Midori_rounds_SR_Result[57]}), .c ({new_AGEMA_signal_3165, new_AGEMA_signal_3164, Midori_rounds_sub_ResultXORkey[21]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U92 ( .a ({new_AGEMA_signal_1843, new_AGEMA_signal_1842, Midori_rounds_SelectedKey_1_}), .b ({new_AGEMA_signal_2837, new_AGEMA_signal_2836, Midori_rounds_SR_Result[49]}), .c ({new_AGEMA_signal_3167, new_AGEMA_signal_3166, Midori_rounds_sub_ResultXORkey[1]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U91 ( .a ({new_AGEMA_signal_2585, new_AGEMA_signal_2584, Midori_rounds_SelectedKey_19_}), .b ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, Midori_rounds_SR_Result[39]}), .c ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, Midori_rounds_sub_ResultXORkey[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U89 ( .a ({new_AGEMA_signal_2581, new_AGEMA_signal_2580, Midori_rounds_SelectedKey_17_}), .b ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, Midori_rounds_SR_Result[37]}), .c ({new_AGEMA_signal_3173, new_AGEMA_signal_3172, Midori_rounds_sub_ResultXORkey[17]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U87 ( .a ({new_AGEMA_signal_1863, new_AGEMA_signal_1862, Midori_rounds_SelectedKey_15_}), .b ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, Midori_rounds_SR_Result[23]}), .c ({new_AGEMA_signal_3175, new_AGEMA_signal_3174, Midori_rounds_sub_ResultXORkey[15]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U85 ( .a ({new_AGEMA_signal_1859, new_AGEMA_signal_1858, Midori_rounds_SelectedKey_13_}), .b ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, Midori_rounds_SR_Result[21]}), .c ({new_AGEMA_signal_3179, new_AGEMA_signal_3178, Midori_rounds_sub_ResultXORkey[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U83 ( .a ({new_AGEMA_signal_1857, new_AGEMA_signal_1856, Midori_rounds_SelectedKey_11_}), .b ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, Midori_rounds_SR_Result[11]}), .c ({new_AGEMA_signal_3181, new_AGEMA_signal_3180, Midori_rounds_sub_ResultXORkey[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U80 ( .a ({new_AGEMA_signal_1853, new_AGEMA_signal_1852, Midori_rounds_SelectedKey_9_}), .b ({new_AGEMA_signal_3401, new_AGEMA_signal_3400, Midori_rounds_SR_Inv_Result[9]}), .c ({new_AGEMA_signal_3425, new_AGEMA_signal_3424, Midori_rounds_mul_ResultXORkey[9]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U77 ( .a ({new_AGEMA_signal_2575, new_AGEMA_signal_2574, Midori_rounds_SelectedKey_7_}), .b ({new_AGEMA_signal_3403, new_AGEMA_signal_3402, Midori_rounds_SR_Inv_Result[55]}), .c ({new_AGEMA_signal_3429, new_AGEMA_signal_3428, Midori_rounds_mul_ResultXORkey[7]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U75 ( .a ({new_AGEMA_signal_2671, new_AGEMA_signal_2670, Midori_rounds_SelectedKey_63_}), .b ({new_AGEMA_signal_3343, new_AGEMA_signal_3342, Midori_rounds_SR_Inv_Result[63]}), .c ({new_AGEMA_signal_3433, new_AGEMA_signal_3432, Midori_rounds_mul_ResultXORkey[63]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U73 ( .a ({new_AGEMA_signal_2667, new_AGEMA_signal_2666, Midori_rounds_SelectedKey_61_}), .b ({new_AGEMA_signal_3347, new_AGEMA_signal_3346, Midori_rounds_SR_Inv_Result[61]}), .c ({new_AGEMA_signal_3437, new_AGEMA_signal_3436, Midori_rounds_mul_ResultXORkey[61]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U70 ( .a ({new_AGEMA_signal_2571, new_AGEMA_signal_2570, Midori_rounds_SelectedKey_5_}), .b ({new_AGEMA_signal_3407, new_AGEMA_signal_3406, Midori_rounds_SR_Inv_Result[53]}), .c ({new_AGEMA_signal_3439, new_AGEMA_signal_3438, Midori_rounds_mul_ResultXORkey[5]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U69 ( .a ({new_AGEMA_signal_2663, new_AGEMA_signal_2662, Midori_rounds_SelectedKey_59_}), .b ({new_AGEMA_signal_3349, new_AGEMA_signal_3348, Midori_rounds_SR_Inv_Result[23]}), .c ({new_AGEMA_signal_3441, new_AGEMA_signal_3440, Midori_rounds_mul_ResultXORkey[59]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U67 ( .a ({new_AGEMA_signal_2659, new_AGEMA_signal_2658, Midori_rounds_SelectedKey_57_}), .b ({new_AGEMA_signal_3329, new_AGEMA_signal_3328, Midori_rounds_SR_Inv_Result[21]}), .c ({new_AGEMA_signal_3445, new_AGEMA_signal_3444, Midori_rounds_mul_ResultXORkey[57]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U64 ( .a ({new_AGEMA_signal_2655, new_AGEMA_signal_2654, Midori_rounds_SelectedKey_55_}), .b ({new_AGEMA_signal_3331, new_AGEMA_signal_3330, Midori_rounds_SR_Inv_Result[43]}), .c ({new_AGEMA_signal_3447, new_AGEMA_signal_3446, Midori_rounds_mul_ResultXORkey[55]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U62 ( .a ({new_AGEMA_signal_2651, new_AGEMA_signal_2650, Midori_rounds_SelectedKey_53_}), .b ({new_AGEMA_signal_3335, new_AGEMA_signal_3334, Midori_rounds_SR_Inv_Result[41]}), .c ({new_AGEMA_signal_3451, new_AGEMA_signal_3450, Midori_rounds_mul_ResultXORkey[53]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U59 ( .a ({new_AGEMA_signal_2647, new_AGEMA_signal_2646, Midori_rounds_SelectedKey_51_}), .b ({new_AGEMA_signal_3337, new_AGEMA_signal_3336, Midori_rounds_SR_Inv_Result[3]}), .c ({new_AGEMA_signal_3453, new_AGEMA_signal_3452, Midori_rounds_mul_ResultXORkey[51]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U55 ( .a ({new_AGEMA_signal_2643, new_AGEMA_signal_2642, Midori_rounds_SelectedKey_49_}), .b ({new_AGEMA_signal_3341, new_AGEMA_signal_3340, Midori_rounds_SR_Inv_Result[1]}), .c ({new_AGEMA_signal_3457, new_AGEMA_signal_3456, Midori_rounds_mul_ResultXORkey[49]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U52 ( .a ({new_AGEMA_signal_2639, new_AGEMA_signal_2638, Midori_rounds_SelectedKey_47_}), .b ({new_AGEMA_signal_3367, new_AGEMA_signal_3366, Midori_rounds_SR_Inv_Result[7]}), .c ({new_AGEMA_signal_3459, new_AGEMA_signal_3458, Midori_rounds_mul_ResultXORkey[47]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U50 ( .a ({new_AGEMA_signal_2635, new_AGEMA_signal_2634, Midori_rounds_SelectedKey_45_}), .b ({new_AGEMA_signal_3371, new_AGEMA_signal_3370, Midori_rounds_SR_Inv_Result[5]}), .c ({new_AGEMA_signal_3463, new_AGEMA_signal_3462, Midori_rounds_mul_ResultXORkey[45]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U47 ( .a ({new_AGEMA_signal_2631, new_AGEMA_signal_2630, Midori_rounds_SelectedKey_43_}), .b ({new_AGEMA_signal_3373, new_AGEMA_signal_3372, Midori_rounds_SR_Inv_Result[47]}), .c ({new_AGEMA_signal_3467, new_AGEMA_signal_3466, Midori_rounds_mul_ResultXORkey[43]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U45 ( .a ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, Midori_rounds_SelectedKey_41_}), .b ({new_AGEMA_signal_3353, new_AGEMA_signal_3352, Midori_rounds_SR_Inv_Result[45]}), .c ({new_AGEMA_signal_3471, new_AGEMA_signal_3470, Midori_rounds_mul_ResultXORkey[41]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U42 ( .a ({new_AGEMA_signal_1847, new_AGEMA_signal_1846, Midori_rounds_SelectedKey_3_}), .b ({new_AGEMA_signal_3409, new_AGEMA_signal_3408, Midori_rounds_SR_Inv_Result[31]}), .c ({new_AGEMA_signal_3473, new_AGEMA_signal_3472, Midori_rounds_mul_ResultXORkey[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U41 ( .a ({new_AGEMA_signal_2623, new_AGEMA_signal_2622, Midori_rounds_SelectedKey_39_}), .b ({new_AGEMA_signal_3355, new_AGEMA_signal_3354, Midori_rounds_SR_Inv_Result[19]}), .c ({new_AGEMA_signal_3475, new_AGEMA_signal_3474, Midori_rounds_mul_ResultXORkey[39]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U39 ( .a ({new_AGEMA_signal_2619, new_AGEMA_signal_2618, Midori_rounds_SelectedKey_37_}), .b ({new_AGEMA_signal_3359, new_AGEMA_signal_3358, Midori_rounds_SR_Inv_Result[17]}), .c ({new_AGEMA_signal_3479, new_AGEMA_signal_3478, Midori_rounds_mul_ResultXORkey[37]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U36 ( .a ({new_AGEMA_signal_2615, new_AGEMA_signal_2614, Midori_rounds_SelectedKey_35_}), .b ({new_AGEMA_signal_3361, new_AGEMA_signal_3360, Midori_rounds_SR_Inv_Result[59]}), .c ({new_AGEMA_signal_3483, new_AGEMA_signal_3482, Midori_rounds_mul_ResultXORkey[35]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U34 ( .a ({new_AGEMA_signal_2611, new_AGEMA_signal_2610, Midori_rounds_SelectedKey_33_}), .b ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, Midori_rounds_SR_Inv_Result[57]}), .c ({new_AGEMA_signal_3487, new_AGEMA_signal_3486, Midori_rounds_mul_ResultXORkey[33]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U31 ( .a ({new_AGEMA_signal_2607, new_AGEMA_signal_2606, Midori_rounds_SelectedKey_31_}), .b ({new_AGEMA_signal_3391, new_AGEMA_signal_3390, Midori_rounds_SR_Inv_Result[27]}), .c ({new_AGEMA_signal_3489, new_AGEMA_signal_3488, Midori_rounds_mul_ResultXORkey[31]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U28 ( .a ({new_AGEMA_signal_2603, new_AGEMA_signal_2602, Midori_rounds_SelectedKey_29_}), .b ({new_AGEMA_signal_3395, new_AGEMA_signal_3394, Midori_rounds_SR_Inv_Result[25]}), .c ({new_AGEMA_signal_3495, new_AGEMA_signal_3494, Midori_rounds_mul_ResultXORkey[29]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U25 ( .a ({new_AGEMA_signal_2599, new_AGEMA_signal_2598, Midori_rounds_SelectedKey_27_}), .b ({new_AGEMA_signal_3397, new_AGEMA_signal_3396, Midori_rounds_SR_Inv_Result[51]}), .c ({new_AGEMA_signal_3497, new_AGEMA_signal_3496, Midori_rounds_mul_ResultXORkey[27]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U23 ( .a ({new_AGEMA_signal_2597, new_AGEMA_signal_2596, Midori_rounds_SelectedKey_25_}), .b ({new_AGEMA_signal_3377, new_AGEMA_signal_3376, Midori_rounds_SR_Inv_Result[49]}), .c ({new_AGEMA_signal_3501, new_AGEMA_signal_3500, Midori_rounds_mul_ResultXORkey[25]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U20 ( .a ({new_AGEMA_signal_2593, new_AGEMA_signal_2592, Midori_rounds_SelectedKey_23_}), .b ({new_AGEMA_signal_3379, new_AGEMA_signal_3378, Midori_rounds_SR_Inv_Result[15]}), .c ({new_AGEMA_signal_3503, new_AGEMA_signal_3502, Midori_rounds_mul_ResultXORkey[23]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U18 ( .a ({new_AGEMA_signal_2589, new_AGEMA_signal_2588, Midori_rounds_SelectedKey_21_}), .b ({new_AGEMA_signal_3383, new_AGEMA_signal_3382, Midori_rounds_SR_Inv_Result[13]}), .c ({new_AGEMA_signal_3507, new_AGEMA_signal_3506, Midori_rounds_mul_ResultXORkey[21]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U15 ( .a ({new_AGEMA_signal_1843, new_AGEMA_signal_1842, Midori_rounds_SelectedKey_1_}), .b ({new_AGEMA_signal_3413, new_AGEMA_signal_3412, Midori_rounds_SR_Inv_Result[29]}), .c ({new_AGEMA_signal_3511, new_AGEMA_signal_3510, Midori_rounds_mul_ResultXORkey[1]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U14 ( .a ({new_AGEMA_signal_2585, new_AGEMA_signal_2584, Midori_rounds_SelectedKey_19_}), .b ({new_AGEMA_signal_3385, new_AGEMA_signal_3384, Midori_rounds_SR_Inv_Result[39]}), .c ({new_AGEMA_signal_3513, new_AGEMA_signal_3512, Midori_rounds_mul_ResultXORkey[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U12 ( .a ({new_AGEMA_signal_2581, new_AGEMA_signal_2580, Midori_rounds_SelectedKey_17_}), .b ({new_AGEMA_signal_3389, new_AGEMA_signal_3388, Midori_rounds_SR_Inv_Result[37]}), .c ({new_AGEMA_signal_3517, new_AGEMA_signal_3516, Midori_rounds_mul_ResultXORkey[17]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U9 ( .a ({new_AGEMA_signal_1863, new_AGEMA_signal_1862, Midori_rounds_SelectedKey_15_}), .b ({new_AGEMA_signal_3415, new_AGEMA_signal_3414, Midori_rounds_SR_Inv_Result[35]}), .c ({new_AGEMA_signal_3519, new_AGEMA_signal_3518, Midori_rounds_mul_ResultXORkey[15]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U7 ( .a ({new_AGEMA_signal_1859, new_AGEMA_signal_1858, Midori_rounds_SelectedKey_13_}), .b ({new_AGEMA_signal_3419, new_AGEMA_signal_3418, Midori_rounds_SR_Inv_Result[33]}), .c ({new_AGEMA_signal_3523, new_AGEMA_signal_3522, Midori_rounds_mul_ResultXORkey[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U4 ( .a ({new_AGEMA_signal_1857, new_AGEMA_signal_1856, Midori_rounds_SelectedKey_11_}), .b ({new_AGEMA_signal_3421, new_AGEMA_signal_3420, Midori_rounds_SR_Inv_Result[11]}), .c ({new_AGEMA_signal_3525, new_AGEMA_signal_3524, Midori_rounds_mul_ResultXORkey[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_1_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3557, new_AGEMA_signal_3556, Midori_rounds_round_Result[1]}), .a ({new_AGEMA_signal_2333, new_AGEMA_signal_2332, Midori_add_Result_Start[1]}), .c ({new_AGEMA_signal_3675, new_AGEMA_signal_3674, Midori_rounds_roundResult_Reg_SFF_1_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_3_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, Midori_rounds_round_Result[3]}), .a ({new_AGEMA_signal_2245, new_AGEMA_signal_2244, Midori_add_Result_Start[3]}), .c ({new_AGEMA_signal_3679, new_AGEMA_signal_3678, Midori_rounds_roundResult_Reg_SFF_3_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_5_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3563, new_AGEMA_signal_3562, Midori_rounds_round_Result[5]}), .a ({new_AGEMA_signal_2157, new_AGEMA_signal_2156, Midori_add_Result_Start[5]}), .c ({new_AGEMA_signal_3681, new_AGEMA_signal_3680, Midori_rounds_roundResult_Reg_SFF_5_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_7_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3567, new_AGEMA_signal_3566, Midori_rounds_round_Result[7]}), .a ({new_AGEMA_signal_2133, new_AGEMA_signal_2132, Midori_add_Result_Start[7]}), .c ({new_AGEMA_signal_3685, new_AGEMA_signal_3684, Midori_rounds_roundResult_Reg_SFF_7_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_9_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3569, new_AGEMA_signal_3568, Midori_rounds_round_Result[9]}), .a ({new_AGEMA_signal_2125, new_AGEMA_signal_2124, Midori_add_Result_Start[9]}), .c ({new_AGEMA_signal_3687, new_AGEMA_signal_3686, Midori_rounds_roundResult_Reg_SFF_9_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_11_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3573, new_AGEMA_signal_3572, Midori_rounds_round_Result[11]}), .a ({new_AGEMA_signal_2369, new_AGEMA_signal_2368, Midori_add_Result_Start[11]}), .c ({new_AGEMA_signal_3691, new_AGEMA_signal_3690, Midori_rounds_roundResult_Reg_SFF_11_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_13_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3575, new_AGEMA_signal_3574, Midori_rounds_round_Result[13]}), .a ({new_AGEMA_signal_2361, new_AGEMA_signal_2360, Midori_add_Result_Start[13]}), .c ({new_AGEMA_signal_3693, new_AGEMA_signal_3692, Midori_rounds_roundResult_Reg_SFF_13_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_15_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3579, new_AGEMA_signal_3578, Midori_rounds_round_Result[15]}), .a ({new_AGEMA_signal_2353, new_AGEMA_signal_2352, Midori_add_Result_Start[15]}), .c ({new_AGEMA_signal_3697, new_AGEMA_signal_3696, Midori_rounds_roundResult_Reg_SFF_15_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_17_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3581, new_AGEMA_signal_3580, Midori_rounds_round_Result[17]}), .a ({new_AGEMA_signal_2345, new_AGEMA_signal_2344, Midori_add_Result_Start[17]}), .c ({new_AGEMA_signal_3699, new_AGEMA_signal_3698, Midori_rounds_roundResult_Reg_SFF_17_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_19_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3585, new_AGEMA_signal_3584, Midori_rounds_round_Result[19]}), .a ({new_AGEMA_signal_2337, new_AGEMA_signal_2336, Midori_add_Result_Start[19]}), .c ({new_AGEMA_signal_3703, new_AGEMA_signal_3702, Midori_rounds_roundResult_Reg_SFF_19_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_21_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3587, new_AGEMA_signal_3586, Midori_rounds_round_Result[21]}), .a ({new_AGEMA_signal_2325, new_AGEMA_signal_2324, Midori_add_Result_Start[21]}), .c ({new_AGEMA_signal_3705, new_AGEMA_signal_3704, Midori_rounds_roundResult_Reg_SFF_21_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_23_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3591, new_AGEMA_signal_3590, Midori_rounds_round_Result[23]}), .a ({new_AGEMA_signal_2317, new_AGEMA_signal_2316, Midori_add_Result_Start[23]}), .c ({new_AGEMA_signal_3709, new_AGEMA_signal_3708, Midori_rounds_roundResult_Reg_SFF_23_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_25_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3593, new_AGEMA_signal_3592, Midori_rounds_round_Result[25]}), .a ({new_AGEMA_signal_2309, new_AGEMA_signal_2308, Midori_add_Result_Start[25]}), .c ({new_AGEMA_signal_3711, new_AGEMA_signal_3710, Midori_rounds_roundResult_Reg_SFF_25_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_27_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3597, new_AGEMA_signal_3596, Midori_rounds_round_Result[27]}), .a ({new_AGEMA_signal_2301, new_AGEMA_signal_2300, Midori_add_Result_Start[27]}), .c ({new_AGEMA_signal_3715, new_AGEMA_signal_3714, Midori_rounds_roundResult_Reg_SFF_27_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_29_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3599, new_AGEMA_signal_3598, Midori_rounds_round_Result[29]}), .a ({new_AGEMA_signal_2293, new_AGEMA_signal_2292, Midori_add_Result_Start[29]}), .c ({new_AGEMA_signal_3717, new_AGEMA_signal_3716, Midori_rounds_roundResult_Reg_SFF_29_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_31_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3603, new_AGEMA_signal_3602, Midori_rounds_round_Result[31]}), .a ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, Midori_add_Result_Start[31]}), .c ({new_AGEMA_signal_3721, new_AGEMA_signal_3720, Midori_rounds_roundResult_Reg_SFF_31_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_33_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3605, new_AGEMA_signal_3604, Midori_rounds_round_Result[33]}), .a ({new_AGEMA_signal_2273, new_AGEMA_signal_2272, Midori_add_Result_Start[33]}), .c ({new_AGEMA_signal_3723, new_AGEMA_signal_3722, Midori_rounds_roundResult_Reg_SFF_33_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_35_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3609, new_AGEMA_signal_3608, Midori_rounds_round_Result[35]}), .a ({new_AGEMA_signal_2265, new_AGEMA_signal_2264, Midori_add_Result_Start[35]}), .c ({new_AGEMA_signal_3727, new_AGEMA_signal_3726, Midori_rounds_roundResult_Reg_SFF_35_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_37_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3611, new_AGEMA_signal_3610, Midori_rounds_round_Result[37]}), .a ({new_AGEMA_signal_2257, new_AGEMA_signal_2256, Midori_add_Result_Start[37]}), .c ({new_AGEMA_signal_3729, new_AGEMA_signal_3728, Midori_rounds_roundResult_Reg_SFF_37_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_39_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3615, new_AGEMA_signal_3614, Midori_rounds_round_Result[39]}), .a ({new_AGEMA_signal_2249, new_AGEMA_signal_2248, Midori_add_Result_Start[39]}), .c ({new_AGEMA_signal_3733, new_AGEMA_signal_3732, Midori_rounds_roundResult_Reg_SFF_39_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_41_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3617, new_AGEMA_signal_3616, Midori_rounds_round_Result[41]}), .a ({new_AGEMA_signal_2237, new_AGEMA_signal_2236, Midori_add_Result_Start[41]}), .c ({new_AGEMA_signal_3735, new_AGEMA_signal_3734, Midori_rounds_roundResult_Reg_SFF_41_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_43_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3621, new_AGEMA_signal_3620, Midori_rounds_round_Result[43]}), .a ({new_AGEMA_signal_2229, new_AGEMA_signal_2228, Midori_add_Result_Start[43]}), .c ({new_AGEMA_signal_3739, new_AGEMA_signal_3738, Midori_rounds_roundResult_Reg_SFF_43_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_45_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3623, new_AGEMA_signal_3622, Midori_rounds_round_Result[45]}), .a ({new_AGEMA_signal_2221, new_AGEMA_signal_2220, Midori_add_Result_Start[45]}), .c ({new_AGEMA_signal_3741, new_AGEMA_signal_3740, Midori_rounds_roundResult_Reg_SFF_45_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_47_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3627, new_AGEMA_signal_3626, Midori_rounds_round_Result[47]}), .a ({new_AGEMA_signal_2213, new_AGEMA_signal_2212, Midori_add_Result_Start[47]}), .c ({new_AGEMA_signal_3745, new_AGEMA_signal_3744, Midori_rounds_roundResult_Reg_SFF_47_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_49_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3629, new_AGEMA_signal_3628, Midori_rounds_round_Result[49]}), .a ({new_AGEMA_signal_2205, new_AGEMA_signal_2204, Midori_add_Result_Start[49]}), .c ({new_AGEMA_signal_3747, new_AGEMA_signal_3746, Midori_rounds_roundResult_Reg_SFF_49_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_51_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3633, new_AGEMA_signal_3632, Midori_rounds_round_Result[51]}), .a ({new_AGEMA_signal_2193, new_AGEMA_signal_2192, Midori_add_Result_Start[51]}), .c ({new_AGEMA_signal_3751, new_AGEMA_signal_3750, Midori_rounds_roundResult_Reg_SFF_51_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_53_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3635, new_AGEMA_signal_3634, Midori_rounds_round_Result[53]}), .a ({new_AGEMA_signal_2185, new_AGEMA_signal_2184, Midori_add_Result_Start[53]}), .c ({new_AGEMA_signal_3753, new_AGEMA_signal_3752, Midori_rounds_roundResult_Reg_SFF_53_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_55_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3639, new_AGEMA_signal_3638, Midori_rounds_round_Result[55]}), .a ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, Midori_add_Result_Start[55]}), .c ({new_AGEMA_signal_3757, new_AGEMA_signal_3756, Midori_rounds_roundResult_Reg_SFF_55_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_57_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3641, new_AGEMA_signal_3640, Midori_rounds_round_Result[57]}), .a ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, Midori_add_Result_Start[57]}), .c ({new_AGEMA_signal_3759, new_AGEMA_signal_3758, Midori_rounds_roundResult_Reg_SFF_57_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_59_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3645, new_AGEMA_signal_3644, Midori_rounds_round_Result[59]}), .a ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, Midori_add_Result_Start[59]}), .c ({new_AGEMA_signal_3763, new_AGEMA_signal_3762, Midori_rounds_roundResult_Reg_SFF_59_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_61_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3647, new_AGEMA_signal_3646, Midori_rounds_round_Result[61]}), .a ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, Midori_add_Result_Start[61]}), .c ({new_AGEMA_signal_3765, new_AGEMA_signal_3764, Midori_rounds_roundResult_Reg_SFF_61_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_63_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3651, new_AGEMA_signal_3650, Midori_rounds_round_Result[63]}), .a ({new_AGEMA_signal_2141, new_AGEMA_signal_2140, Midori_add_Result_Start[63]}), .c ({new_AGEMA_signal_3769, new_AGEMA_signal_3768, Midori_rounds_roundResult_Reg_SFF_63_DQ}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U19 ( .a ({new_AGEMA_signal_2381, new_AGEMA_signal_2380, Midori_rounds_sub_sBox_PRINCE_0_n15}), .b ({new_AGEMA_signal_2675, new_AGEMA_signal_2674, Midori_rounds_sub_sBox_PRINCE_0_n14}), .clk (clk), .r ({Fresh[482], Fresh[481], Fresh[480]}), .c ({new_AGEMA_signal_2833, new_AGEMA_signal_2832, Midori_rounds_SR_Result[51]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U16 ( .a ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, Midori_rounds_sub_sBox_PRINCE_0_n11}), .b ({new_AGEMA_signal_2673, new_AGEMA_signal_2672, Midori_rounds_roundReg_out[1]}), .clk (clk), .r ({Fresh[485], Fresh[484], Fresh[483]}), .c ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, Midori_rounds_sub_sBox_PRINCE_0_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U12 ( .a ({new_AGEMA_signal_2385, new_AGEMA_signal_2384, Midori_rounds_sub_sBox_PRINCE_0_n6}), .b ({new_AGEMA_signal_2679, new_AGEMA_signal_2678, Midori_rounds_sub_sBox_PRINCE_0_n5}), .clk (clk), .r ({Fresh[488], Fresh[487], Fresh[486]}), .c ({new_AGEMA_signal_2837, new_AGEMA_signal_2836, Midori_rounds_SR_Result[49]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U7 ( .a ({new_AGEMA_signal_2673, new_AGEMA_signal_2672, Midori_rounds_roundReg_out[1]}), .b ({new_AGEMA_signal_2387, new_AGEMA_signal_2386, Midori_rounds_sub_sBox_PRINCE_0_n2}), .clk (clk), .r ({Fresh[491], Fresh[490], Fresh[489]}), .c ({new_AGEMA_signal_2681, new_AGEMA_signal_2680, Midori_rounds_sub_sBox_PRINCE_0_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U19 ( .a ({new_AGEMA_signal_2393, new_AGEMA_signal_2392, Midori_rounds_sub_sBox_PRINCE_1_n15}), .b ({new_AGEMA_signal_2685, new_AGEMA_signal_2684, Midori_rounds_sub_sBox_PRINCE_1_n14}), .clk (clk), .r ({Fresh[494], Fresh[493], Fresh[492]}), .c ({new_AGEMA_signal_2841, new_AGEMA_signal_2840, Midori_rounds_SR_Result[47]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U16 ( .a ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, Midori_rounds_sub_sBox_PRINCE_1_n11}), .b ({new_AGEMA_signal_2683, new_AGEMA_signal_2682, Midori_rounds_roundReg_out[5]}), .clk (clk), .r ({Fresh[497], Fresh[496], Fresh[495]}), .c ({new_AGEMA_signal_2687, new_AGEMA_signal_2686, Midori_rounds_sub_sBox_PRINCE_1_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U12 ( .a ({new_AGEMA_signal_2397, new_AGEMA_signal_2396, Midori_rounds_sub_sBox_PRINCE_1_n6}), .b ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, Midori_rounds_sub_sBox_PRINCE_1_n5}), .clk (clk), .r ({Fresh[500], Fresh[499], Fresh[498]}), .c ({new_AGEMA_signal_2845, new_AGEMA_signal_2844, Midori_rounds_SR_Result[45]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U7 ( .a ({new_AGEMA_signal_2683, new_AGEMA_signal_2682, Midori_rounds_roundReg_out[5]}), .b ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, Midori_rounds_sub_sBox_PRINCE_1_n2}), .clk (clk), .r ({Fresh[503], Fresh[502], Fresh[501]}), .c ({new_AGEMA_signal_2691, new_AGEMA_signal_2690, Midori_rounds_sub_sBox_PRINCE_1_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U19 ( .a ({new_AGEMA_signal_2405, new_AGEMA_signal_2404, Midori_rounds_sub_sBox_PRINCE_2_n15}), .b ({new_AGEMA_signal_2695, new_AGEMA_signal_2694, Midori_rounds_sub_sBox_PRINCE_2_n14}), .clk (clk), .r ({Fresh[506], Fresh[505], Fresh[504]}), .c ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, Midori_rounds_SR_Result[11]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U16 ( .a ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, Midori_rounds_sub_sBox_PRINCE_2_n11}), .b ({new_AGEMA_signal_2693, new_AGEMA_signal_2692, Midori_rounds_roundReg_out[9]}), .clk (clk), .r ({Fresh[509], Fresh[508], Fresh[507]}), .c ({new_AGEMA_signal_2697, new_AGEMA_signal_2696, Midori_rounds_sub_sBox_PRINCE_2_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U12 ( .a ({new_AGEMA_signal_2409, new_AGEMA_signal_2408, Midori_rounds_sub_sBox_PRINCE_2_n6}), .b ({new_AGEMA_signal_2699, new_AGEMA_signal_2698, Midori_rounds_sub_sBox_PRINCE_2_n5}), .clk (clk), .r ({Fresh[512], Fresh[511], Fresh[510]}), .c ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, Midori_rounds_SR_Result[9]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U7 ( .a ({new_AGEMA_signal_2693, new_AGEMA_signal_2692, Midori_rounds_roundReg_out[9]}), .b ({new_AGEMA_signal_2411, new_AGEMA_signal_2410, Midori_rounds_sub_sBox_PRINCE_2_n2}), .clk (clk), .r ({Fresh[515], Fresh[514], Fresh[513]}), .c ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, Midori_rounds_sub_sBox_PRINCE_2_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U19 ( .a ({new_AGEMA_signal_2417, new_AGEMA_signal_2416, Midori_rounds_sub_sBox_PRINCE_3_n15}), .b ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, Midori_rounds_sub_sBox_PRINCE_3_n14}), .clk (clk), .r ({Fresh[518], Fresh[517], Fresh[516]}), .c ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, Midori_rounds_SR_Result[23]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U16 ( .a ({new_AGEMA_signal_2415, new_AGEMA_signal_2414, Midori_rounds_sub_sBox_PRINCE_3_n11}), .b ({new_AGEMA_signal_2703, new_AGEMA_signal_2702, Midori_rounds_roundReg_out[13]}), .clk (clk), .r ({Fresh[521], Fresh[520], Fresh[519]}), .c ({new_AGEMA_signal_2707, new_AGEMA_signal_2706, Midori_rounds_sub_sBox_PRINCE_3_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U12 ( .a ({new_AGEMA_signal_2421, new_AGEMA_signal_2420, Midori_rounds_sub_sBox_PRINCE_3_n6}), .b ({new_AGEMA_signal_2709, new_AGEMA_signal_2708, Midori_rounds_sub_sBox_PRINCE_3_n5}), .clk (clk), .r ({Fresh[524], Fresh[523], Fresh[522]}), .c ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, Midori_rounds_SR_Result[21]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U7 ( .a ({new_AGEMA_signal_2703, new_AGEMA_signal_2702, Midori_rounds_roundReg_out[13]}), .b ({new_AGEMA_signal_2423, new_AGEMA_signal_2422, Midori_rounds_sub_sBox_PRINCE_3_n2}), .clk (clk), .r ({Fresh[527], Fresh[526], Fresh[525]}), .c ({new_AGEMA_signal_2711, new_AGEMA_signal_2710, Midori_rounds_sub_sBox_PRINCE_3_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U19 ( .a ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, Midori_rounds_sub_sBox_PRINCE_4_n15}), .b ({new_AGEMA_signal_2715, new_AGEMA_signal_2714, Midori_rounds_sub_sBox_PRINCE_4_n14}), .clk (clk), .r ({Fresh[530], Fresh[529], Fresh[528]}), .c ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, Midori_rounds_SR_Result[39]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U16 ( .a ({new_AGEMA_signal_2427, new_AGEMA_signal_2426, Midori_rounds_sub_sBox_PRINCE_4_n11}), .b ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, Midori_rounds_roundReg_out[17]}), .clk (clk), .r ({Fresh[533], Fresh[532], Fresh[531]}), .c ({new_AGEMA_signal_2717, new_AGEMA_signal_2716, Midori_rounds_sub_sBox_PRINCE_4_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U12 ( .a ({new_AGEMA_signal_2433, new_AGEMA_signal_2432, Midori_rounds_sub_sBox_PRINCE_4_n6}), .b ({new_AGEMA_signal_2719, new_AGEMA_signal_2718, Midori_rounds_sub_sBox_PRINCE_4_n5}), .clk (clk), .r ({Fresh[536], Fresh[535], Fresh[534]}), .c ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, Midori_rounds_SR_Result[37]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U7 ( .a ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, Midori_rounds_roundReg_out[17]}), .b ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, Midori_rounds_sub_sBox_PRINCE_4_n2}), .clk (clk), .r ({Fresh[539], Fresh[538], Fresh[537]}), .c ({new_AGEMA_signal_2721, new_AGEMA_signal_2720, Midori_rounds_sub_sBox_PRINCE_4_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U19 ( .a ({new_AGEMA_signal_2441, new_AGEMA_signal_2440, Midori_rounds_sub_sBox_PRINCE_5_n15}), .b ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, Midori_rounds_sub_sBox_PRINCE_5_n14}), .clk (clk), .r ({Fresh[542], Fresh[541], Fresh[540]}), .c ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, Midori_rounds_SR_Result[59]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U16 ( .a ({new_AGEMA_signal_2439, new_AGEMA_signal_2438, Midori_rounds_sub_sBox_PRINCE_5_n11}), .b ({new_AGEMA_signal_2723, new_AGEMA_signal_2722, Midori_rounds_roundReg_out[21]}), .clk (clk), .r ({Fresh[545], Fresh[544], Fresh[543]}), .c ({new_AGEMA_signal_2727, new_AGEMA_signal_2726, Midori_rounds_sub_sBox_PRINCE_5_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U12 ( .a ({new_AGEMA_signal_2445, new_AGEMA_signal_2444, Midori_rounds_sub_sBox_PRINCE_5_n6}), .b ({new_AGEMA_signal_2729, new_AGEMA_signal_2728, Midori_rounds_sub_sBox_PRINCE_5_n5}), .clk (clk), .r ({Fresh[548], Fresh[547], Fresh[546]}), .c ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, Midori_rounds_SR_Result[57]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U7 ( .a ({new_AGEMA_signal_2723, new_AGEMA_signal_2722, Midori_rounds_roundReg_out[21]}), .b ({new_AGEMA_signal_2447, new_AGEMA_signal_2446, Midori_rounds_sub_sBox_PRINCE_5_n2}), .clk (clk), .r ({Fresh[551], Fresh[550], Fresh[549]}), .c ({new_AGEMA_signal_2731, new_AGEMA_signal_2730, Midori_rounds_sub_sBox_PRINCE_5_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U19 ( .a ({new_AGEMA_signal_2453, new_AGEMA_signal_2452, Midori_rounds_sub_sBox_PRINCE_6_n15}), .b ({new_AGEMA_signal_2735, new_AGEMA_signal_2734, Midori_rounds_sub_sBox_PRINCE_6_n14}), .clk (clk), .r ({Fresh[554], Fresh[553], Fresh[552]}), .c ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, Midori_rounds_SR_Result[31]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U16 ( .a ({new_AGEMA_signal_2451, new_AGEMA_signal_2450, Midori_rounds_sub_sBox_PRINCE_6_n11}), .b ({new_AGEMA_signal_2733, new_AGEMA_signal_2732, Midori_rounds_roundReg_out[25]}), .clk (clk), .r ({Fresh[557], Fresh[556], Fresh[555]}), .c ({new_AGEMA_signal_2737, new_AGEMA_signal_2736, Midori_rounds_sub_sBox_PRINCE_6_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U12 ( .a ({new_AGEMA_signal_2457, new_AGEMA_signal_2456, Midori_rounds_sub_sBox_PRINCE_6_n6}), .b ({new_AGEMA_signal_2739, new_AGEMA_signal_2738, Midori_rounds_sub_sBox_PRINCE_6_n5}), .clk (clk), .r ({Fresh[560], Fresh[559], Fresh[558]}), .c ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, Midori_rounds_SR_Result[29]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U7 ( .a ({new_AGEMA_signal_2733, new_AGEMA_signal_2732, Midori_rounds_roundReg_out[25]}), .b ({new_AGEMA_signal_2459, new_AGEMA_signal_2458, Midori_rounds_sub_sBox_PRINCE_6_n2}), .clk (clk), .r ({Fresh[563], Fresh[562], Fresh[561]}), .c ({new_AGEMA_signal_2741, new_AGEMA_signal_2740, Midori_rounds_sub_sBox_PRINCE_6_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U19 ( .a ({new_AGEMA_signal_2465, new_AGEMA_signal_2464, Midori_rounds_sub_sBox_PRINCE_7_n15}), .b ({new_AGEMA_signal_2745, new_AGEMA_signal_2744, Midori_rounds_sub_sBox_PRINCE_7_n14}), .clk (clk), .r ({Fresh[566], Fresh[565], Fresh[564]}), .c ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, Midori_rounds_SR_Result[3]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U16 ( .a ({new_AGEMA_signal_2463, new_AGEMA_signal_2462, Midori_rounds_sub_sBox_PRINCE_7_n11}), .b ({new_AGEMA_signal_2743, new_AGEMA_signal_2742, Midori_rounds_roundReg_out[29]}), .clk (clk), .r ({Fresh[569], Fresh[568], Fresh[567]}), .c ({new_AGEMA_signal_2747, new_AGEMA_signal_2746, Midori_rounds_sub_sBox_PRINCE_7_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U12 ( .a ({new_AGEMA_signal_2469, new_AGEMA_signal_2468, Midori_rounds_sub_sBox_PRINCE_7_n6}), .b ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, Midori_rounds_sub_sBox_PRINCE_7_n5}), .clk (clk), .r ({Fresh[572], Fresh[571], Fresh[570]}), .c ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, Midori_rounds_SR_Result[1]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U7 ( .a ({new_AGEMA_signal_2743, new_AGEMA_signal_2742, Midori_rounds_roundReg_out[29]}), .b ({new_AGEMA_signal_2471, new_AGEMA_signal_2470, Midori_rounds_sub_sBox_PRINCE_7_n2}), .clk (clk), .r ({Fresh[575], Fresh[574], Fresh[573]}), .c ({new_AGEMA_signal_2751, new_AGEMA_signal_2750, Midori_rounds_sub_sBox_PRINCE_7_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U19 ( .a ({new_AGEMA_signal_2477, new_AGEMA_signal_2476, Midori_rounds_sub_sBox_PRINCE_8_n15}), .b ({new_AGEMA_signal_2755, new_AGEMA_signal_2754, Midori_rounds_sub_sBox_PRINCE_8_n14}), .clk (clk), .r ({Fresh[578], Fresh[577], Fresh[576]}), .c ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, Midori_rounds_SR_Result[15]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U16 ( .a ({new_AGEMA_signal_2475, new_AGEMA_signal_2474, Midori_rounds_sub_sBox_PRINCE_8_n11}), .b ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, Midori_rounds_roundReg_out[33]}), .clk (clk), .r ({Fresh[581], Fresh[580], Fresh[579]}), .c ({new_AGEMA_signal_2757, new_AGEMA_signal_2756, Midori_rounds_sub_sBox_PRINCE_8_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U12 ( .a ({new_AGEMA_signal_2481, new_AGEMA_signal_2480, Midori_rounds_sub_sBox_PRINCE_8_n6}), .b ({new_AGEMA_signal_2759, new_AGEMA_signal_2758, Midori_rounds_sub_sBox_PRINCE_8_n5}), .clk (clk), .r ({Fresh[584], Fresh[583], Fresh[582]}), .c ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, Midori_rounds_SR_Result[13]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U7 ( .a ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, Midori_rounds_roundReg_out[33]}), .b ({new_AGEMA_signal_2483, new_AGEMA_signal_2482, Midori_rounds_sub_sBox_PRINCE_8_n2}), .clk (clk), .r ({Fresh[587], Fresh[586], Fresh[585]}), .c ({new_AGEMA_signal_2761, new_AGEMA_signal_2760, Midori_rounds_sub_sBox_PRINCE_8_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U19 ( .a ({new_AGEMA_signal_2489, new_AGEMA_signal_2488, Midori_rounds_sub_sBox_PRINCE_9_n15}), .b ({new_AGEMA_signal_2765, new_AGEMA_signal_2764, Midori_rounds_sub_sBox_PRINCE_9_n14}), .clk (clk), .r ({Fresh[590], Fresh[589], Fresh[588]}), .c ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, Midori_rounds_SR_Result[19]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U16 ( .a ({new_AGEMA_signal_2487, new_AGEMA_signal_2486, Midori_rounds_sub_sBox_PRINCE_9_n11}), .b ({new_AGEMA_signal_2763, new_AGEMA_signal_2762, Midori_rounds_roundReg_out[37]}), .clk (clk), .r ({Fresh[593], Fresh[592], Fresh[591]}), .c ({new_AGEMA_signal_2767, new_AGEMA_signal_2766, Midori_rounds_sub_sBox_PRINCE_9_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U12 ( .a ({new_AGEMA_signal_2493, new_AGEMA_signal_2492, Midori_rounds_sub_sBox_PRINCE_9_n6}), .b ({new_AGEMA_signal_2769, new_AGEMA_signal_2768, Midori_rounds_sub_sBox_PRINCE_9_n5}), .clk (clk), .r ({Fresh[596], Fresh[595], Fresh[594]}), .c ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, Midori_rounds_SR_Result[17]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U7 ( .a ({new_AGEMA_signal_2763, new_AGEMA_signal_2762, Midori_rounds_roundReg_out[37]}), .b ({new_AGEMA_signal_2495, new_AGEMA_signal_2494, Midori_rounds_sub_sBox_PRINCE_9_n2}), .clk (clk), .r ({Fresh[599], Fresh[598], Fresh[597]}), .c ({new_AGEMA_signal_2771, new_AGEMA_signal_2770, Midori_rounds_sub_sBox_PRINCE_9_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U19 ( .a ({new_AGEMA_signal_2501, new_AGEMA_signal_2500, Midori_rounds_sub_sBox_PRINCE_10_n15}), .b ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, Midori_rounds_sub_sBox_PRINCE_10_n14}), .clk (clk), .r ({Fresh[602], Fresh[601], Fresh[600]}), .c ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, Midori_rounds_SR_Result[55]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U16 ( .a ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, Midori_rounds_sub_sBox_PRINCE_10_n11}), .b ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, Midori_rounds_roundReg_out[41]}), .clk (clk), .r ({Fresh[605], Fresh[604], Fresh[603]}), .c ({new_AGEMA_signal_2777, new_AGEMA_signal_2776, Midori_rounds_sub_sBox_PRINCE_10_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U12 ( .a ({new_AGEMA_signal_2505, new_AGEMA_signal_2504, Midori_rounds_sub_sBox_PRINCE_10_n6}), .b ({new_AGEMA_signal_2779, new_AGEMA_signal_2778, Midori_rounds_sub_sBox_PRINCE_10_n5}), .clk (clk), .r ({Fresh[608], Fresh[607], Fresh[606]}), .c ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, Midori_rounds_SR_Result[53]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U7 ( .a ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, Midori_rounds_roundReg_out[41]}), .b ({new_AGEMA_signal_2507, new_AGEMA_signal_2506, Midori_rounds_sub_sBox_PRINCE_10_n2}), .clk (clk), .r ({Fresh[611], Fresh[610], Fresh[609]}), .c ({new_AGEMA_signal_2781, new_AGEMA_signal_2780, Midori_rounds_sub_sBox_PRINCE_10_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U19 ( .a ({new_AGEMA_signal_2513, new_AGEMA_signal_2512, Midori_rounds_sub_sBox_PRINCE_11_n15}), .b ({new_AGEMA_signal_2785, new_AGEMA_signal_2784, Midori_rounds_sub_sBox_PRINCE_11_n14}), .clk (clk), .r ({Fresh[614], Fresh[613], Fresh[612]}), .c ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, Midori_rounds_SR_Result[43]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U16 ( .a ({new_AGEMA_signal_2511, new_AGEMA_signal_2510, Midori_rounds_sub_sBox_PRINCE_11_n11}), .b ({new_AGEMA_signal_2783, new_AGEMA_signal_2782, Midori_rounds_roundReg_out[45]}), .clk (clk), .r ({Fresh[617], Fresh[616], Fresh[615]}), .c ({new_AGEMA_signal_2787, new_AGEMA_signal_2786, Midori_rounds_sub_sBox_PRINCE_11_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U12 ( .a ({new_AGEMA_signal_2517, new_AGEMA_signal_2516, Midori_rounds_sub_sBox_PRINCE_11_n6}), .b ({new_AGEMA_signal_2789, new_AGEMA_signal_2788, Midori_rounds_sub_sBox_PRINCE_11_n5}), .clk (clk), .r ({Fresh[620], Fresh[619], Fresh[618]}), .c ({new_AGEMA_signal_2925, new_AGEMA_signal_2924, Midori_rounds_SR_Result[41]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U7 ( .a ({new_AGEMA_signal_2783, new_AGEMA_signal_2782, Midori_rounds_roundReg_out[45]}), .b ({new_AGEMA_signal_2519, new_AGEMA_signal_2518, Midori_rounds_sub_sBox_PRINCE_11_n2}), .clk (clk), .r ({Fresh[623], Fresh[622], Fresh[621]}), .c ({new_AGEMA_signal_2791, new_AGEMA_signal_2790, Midori_rounds_sub_sBox_PRINCE_11_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U19 ( .a ({new_AGEMA_signal_2525, new_AGEMA_signal_2524, Midori_rounds_sub_sBox_PRINCE_12_n15}), .b ({new_AGEMA_signal_2795, new_AGEMA_signal_2794, Midori_rounds_sub_sBox_PRINCE_12_n14}), .clk (clk), .r ({Fresh[626], Fresh[625], Fresh[624]}), .c ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, Midori_rounds_SR_Result[27]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U16 ( .a ({new_AGEMA_signal_2523, new_AGEMA_signal_2522, Midori_rounds_sub_sBox_PRINCE_12_n11}), .b ({new_AGEMA_signal_2793, new_AGEMA_signal_2792, Midori_rounds_roundReg_out[49]}), .clk (clk), .r ({Fresh[629], Fresh[628], Fresh[627]}), .c ({new_AGEMA_signal_2797, new_AGEMA_signal_2796, Midori_rounds_sub_sBox_PRINCE_12_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U12 ( .a ({new_AGEMA_signal_2529, new_AGEMA_signal_2528, Midori_rounds_sub_sBox_PRINCE_12_n6}), .b ({new_AGEMA_signal_2799, new_AGEMA_signal_2798, Midori_rounds_sub_sBox_PRINCE_12_n5}), .clk (clk), .r ({Fresh[632], Fresh[631], Fresh[630]}), .c ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, Midori_rounds_SR_Result[25]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U7 ( .a ({new_AGEMA_signal_2793, new_AGEMA_signal_2792, Midori_rounds_roundReg_out[49]}), .b ({new_AGEMA_signal_2531, new_AGEMA_signal_2530, Midori_rounds_sub_sBox_PRINCE_12_n2}), .clk (clk), .r ({Fresh[635], Fresh[634], Fresh[633]}), .c ({new_AGEMA_signal_2801, new_AGEMA_signal_2800, Midori_rounds_sub_sBox_PRINCE_12_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U19 ( .a ({new_AGEMA_signal_2537, new_AGEMA_signal_2536, Midori_rounds_sub_sBox_PRINCE_13_n15}), .b ({new_AGEMA_signal_2805, new_AGEMA_signal_2804, Midori_rounds_sub_sBox_PRINCE_13_n14}), .clk (clk), .r ({Fresh[638], Fresh[637], Fresh[636]}), .c ({new_AGEMA_signal_2937, new_AGEMA_signal_2936, Midori_rounds_SR_Result[7]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U16 ( .a ({new_AGEMA_signal_2535, new_AGEMA_signal_2534, Midori_rounds_sub_sBox_PRINCE_13_n11}), .b ({new_AGEMA_signal_2803, new_AGEMA_signal_2802, Midori_rounds_roundReg_out[53]}), .clk (clk), .r ({Fresh[641], Fresh[640], Fresh[639]}), .c ({new_AGEMA_signal_2807, new_AGEMA_signal_2806, Midori_rounds_sub_sBox_PRINCE_13_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U12 ( .a ({new_AGEMA_signal_2541, new_AGEMA_signal_2540, Midori_rounds_sub_sBox_PRINCE_13_n6}), .b ({new_AGEMA_signal_2809, new_AGEMA_signal_2808, Midori_rounds_sub_sBox_PRINCE_13_n5}), .clk (clk), .r ({Fresh[644], Fresh[643], Fresh[642]}), .c ({new_AGEMA_signal_2941, new_AGEMA_signal_2940, Midori_rounds_SR_Result[5]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U7 ( .a ({new_AGEMA_signal_2803, new_AGEMA_signal_2802, Midori_rounds_roundReg_out[53]}), .b ({new_AGEMA_signal_2543, new_AGEMA_signal_2542, Midori_rounds_sub_sBox_PRINCE_13_n2}), .clk (clk), .r ({Fresh[647], Fresh[646], Fresh[645]}), .c ({new_AGEMA_signal_2811, new_AGEMA_signal_2810, Midori_rounds_sub_sBox_PRINCE_13_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U19 ( .a ({new_AGEMA_signal_2549, new_AGEMA_signal_2548, Midori_rounds_sub_sBox_PRINCE_14_n15}), .b ({new_AGEMA_signal_2815, new_AGEMA_signal_2814, Midori_rounds_sub_sBox_PRINCE_14_n14}), .clk (clk), .r ({Fresh[650], Fresh[649], Fresh[648]}), .c ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, Midori_rounds_SR_Result[35]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U16 ( .a ({new_AGEMA_signal_2547, new_AGEMA_signal_2546, Midori_rounds_sub_sBox_PRINCE_14_n11}), .b ({new_AGEMA_signal_2813, new_AGEMA_signal_2812, Midori_rounds_roundReg_out[57]}), .clk (clk), .r ({Fresh[653], Fresh[652], Fresh[651]}), .c ({new_AGEMA_signal_2817, new_AGEMA_signal_2816, Midori_rounds_sub_sBox_PRINCE_14_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U12 ( .a ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, Midori_rounds_sub_sBox_PRINCE_14_n6}), .b ({new_AGEMA_signal_2819, new_AGEMA_signal_2818, Midori_rounds_sub_sBox_PRINCE_14_n5}), .clk (clk), .r ({Fresh[656], Fresh[655], Fresh[654]}), .c ({new_AGEMA_signal_2949, new_AGEMA_signal_2948, Midori_rounds_SR_Result[33]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U7 ( .a ({new_AGEMA_signal_2813, new_AGEMA_signal_2812, Midori_rounds_roundReg_out[57]}), .b ({new_AGEMA_signal_2555, new_AGEMA_signal_2554, Midori_rounds_sub_sBox_PRINCE_14_n2}), .clk (clk), .r ({Fresh[659], Fresh[658], Fresh[657]}), .c ({new_AGEMA_signal_2821, new_AGEMA_signal_2820, Midori_rounds_sub_sBox_PRINCE_14_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U19 ( .a ({new_AGEMA_signal_2561, new_AGEMA_signal_2560, Midori_rounds_sub_sBox_PRINCE_15_n15}), .b ({new_AGEMA_signal_2825, new_AGEMA_signal_2824, Midori_rounds_sub_sBox_PRINCE_15_n14}), .clk (clk), .r ({Fresh[662], Fresh[661], Fresh[660]}), .c ({new_AGEMA_signal_2953, new_AGEMA_signal_2952, Midori_rounds_SR_Result[63]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U16 ( .a ({new_AGEMA_signal_2559, new_AGEMA_signal_2558, Midori_rounds_sub_sBox_PRINCE_15_n11}), .b ({new_AGEMA_signal_2823, new_AGEMA_signal_2822, Midori_rounds_roundReg_out[61]}), .clk (clk), .r ({Fresh[665], Fresh[664], Fresh[663]}), .c ({new_AGEMA_signal_2827, new_AGEMA_signal_2826, Midori_rounds_sub_sBox_PRINCE_15_n12}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U12 ( .a ({new_AGEMA_signal_2565, new_AGEMA_signal_2564, Midori_rounds_sub_sBox_PRINCE_15_n6}), .b ({new_AGEMA_signal_2829, new_AGEMA_signal_2828, Midori_rounds_sub_sBox_PRINCE_15_n5}), .clk (clk), .r ({Fresh[668], Fresh[667], Fresh[666]}), .c ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, Midori_rounds_SR_Result[61]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U7 ( .a ({new_AGEMA_signal_2823, new_AGEMA_signal_2822, Midori_rounds_roundReg_out[61]}), .b ({new_AGEMA_signal_2567, new_AGEMA_signal_2566, Midori_rounds_sub_sBox_PRINCE_15_n2}), .clk (clk), .r ({Fresh[671], Fresh[670], Fresh[669]}), .c ({new_AGEMA_signal_2831, new_AGEMA_signal_2830, Midori_rounds_sub_sBox_PRINCE_15_n3}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_1_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, Midori_rounds_SR_Result[1]}), .a ({new_AGEMA_signal_3167, new_AGEMA_signal_3166, Midori_rounds_sub_ResultXORkey[1]}), .c ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, Midori_rounds_mul_input[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_3_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, Midori_rounds_SR_Result[3]}), .a ({new_AGEMA_signal_3133, new_AGEMA_signal_3132, Midori_rounds_sub_ResultXORkey[3]}), .c ({new_AGEMA_signal_3189, new_AGEMA_signal_3188, Midori_rounds_mul_input[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_5_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2941, new_AGEMA_signal_2940, Midori_rounds_SR_Result[5]}), .a ({new_AGEMA_signal_3101, new_AGEMA_signal_3100, Midori_rounds_sub_ResultXORkey[5]}), .c ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, Midori_rounds_mul_input[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_7_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2937, new_AGEMA_signal_2936, Midori_rounds_SR_Result[7]}), .a ({new_AGEMA_signal_3091, new_AGEMA_signal_3090, Midori_rounds_sub_ResultXORkey[7]}), .c ({new_AGEMA_signal_3195, new_AGEMA_signal_3194, Midori_rounds_mul_input[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_9_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, Midori_rounds_SR_Result[9]}), .a ({new_AGEMA_signal_3089, new_AGEMA_signal_3088, Midori_rounds_sub_ResultXORkey[9]}), .c ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, Midori_rounds_mul_input[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_11_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, Midori_rounds_SR_Result[11]}), .a ({new_AGEMA_signal_3181, new_AGEMA_signal_3180, Midori_rounds_sub_ResultXORkey[11]}), .c ({new_AGEMA_signal_3201, new_AGEMA_signal_3200, Midori_rounds_mul_input[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_13_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, Midori_rounds_SR_Result[13]}), .a ({new_AGEMA_signal_3179, new_AGEMA_signal_3178, Midori_rounds_sub_ResultXORkey[13]}), .c ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, Midori_rounds_mul_input[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_15_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, Midori_rounds_SR_Result[15]}), .a ({new_AGEMA_signal_3175, new_AGEMA_signal_3174, Midori_rounds_sub_ResultXORkey[15]}), .c ({new_AGEMA_signal_3207, new_AGEMA_signal_3206, Midori_rounds_mul_input[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_17_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, Midori_rounds_SR_Result[17]}), .a ({new_AGEMA_signal_3173, new_AGEMA_signal_3172, Midori_rounds_sub_ResultXORkey[17]}), .c ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, Midori_rounds_mul_input[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_19_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, Midori_rounds_SR_Result[19]}), .a ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, Midori_rounds_sub_ResultXORkey[19]}), .c ({new_AGEMA_signal_3213, new_AGEMA_signal_3212, Midori_rounds_mul_input[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_21_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, Midori_rounds_SR_Result[21]}), .a ({new_AGEMA_signal_3165, new_AGEMA_signal_3164, Midori_rounds_sub_ResultXORkey[21]}), .c ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, Midori_rounds_mul_input[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_23_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, Midori_rounds_SR_Result[23]}), .a ({new_AGEMA_signal_3161, new_AGEMA_signal_3160, Midori_rounds_sub_ResultXORkey[23]}), .c ({new_AGEMA_signal_3219, new_AGEMA_signal_3218, Midori_rounds_mul_input[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_25_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, Midori_rounds_SR_Result[25]}), .a ({new_AGEMA_signal_3159, new_AGEMA_signal_3158, Midori_rounds_sub_ResultXORkey[25]}), .c ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, Midori_rounds_mul_input[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_27_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, Midori_rounds_SR_Result[27]}), .a ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, Midori_rounds_sub_ResultXORkey[27]}), .c ({new_AGEMA_signal_3225, new_AGEMA_signal_3224, Midori_rounds_mul_input[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_29_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, Midori_rounds_SR_Result[29]}), .a ({new_AGEMA_signal_3153, new_AGEMA_signal_3152, Midori_rounds_sub_ResultXORkey[29]}), .c ({new_AGEMA_signal_3227, new_AGEMA_signal_3226, Midori_rounds_mul_input[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_31_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, Midori_rounds_SR_Result[31]}), .a ({new_AGEMA_signal_3147, new_AGEMA_signal_3146, Midori_rounds_sub_ResultXORkey[31]}), .c ({new_AGEMA_signal_3231, new_AGEMA_signal_3230, Midori_rounds_mul_input[31]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_33_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2949, new_AGEMA_signal_2948, Midori_rounds_SR_Result[33]}), .a ({new_AGEMA_signal_3145, new_AGEMA_signal_3144, Midori_rounds_sub_ResultXORkey[33]}), .c ({new_AGEMA_signal_3233, new_AGEMA_signal_3232, Midori_rounds_mul_input[33]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_35_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, Midori_rounds_SR_Result[35]}), .a ({new_AGEMA_signal_3141, new_AGEMA_signal_3140, Midori_rounds_sub_ResultXORkey[35]}), .c ({new_AGEMA_signal_3237, new_AGEMA_signal_3236, Midori_rounds_mul_input[35]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_37_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, Midori_rounds_SR_Result[37]}), .a ({new_AGEMA_signal_3139, new_AGEMA_signal_3138, Midori_rounds_sub_ResultXORkey[37]}), .c ({new_AGEMA_signal_3239, new_AGEMA_signal_3238, Midori_rounds_mul_input[37]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_39_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, Midori_rounds_SR_Result[39]}), .a ({new_AGEMA_signal_3135, new_AGEMA_signal_3134, Midori_rounds_sub_ResultXORkey[39]}), .c ({new_AGEMA_signal_3243, new_AGEMA_signal_3242, Midori_rounds_mul_input[39]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_41_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2925, new_AGEMA_signal_2924, Midori_rounds_SR_Result[41]}), .a ({new_AGEMA_signal_3131, new_AGEMA_signal_3130, Midori_rounds_sub_ResultXORkey[41]}), .c ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, Midori_rounds_mul_input[41]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_43_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, Midori_rounds_SR_Result[43]}), .a ({new_AGEMA_signal_3127, new_AGEMA_signal_3126, Midori_rounds_sub_ResultXORkey[43]}), .c ({new_AGEMA_signal_3249, new_AGEMA_signal_3248, Midori_rounds_mul_input[43]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_45_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2845, new_AGEMA_signal_2844, Midori_rounds_SR_Result[45]}), .a ({new_AGEMA_signal_3125, new_AGEMA_signal_3124, Midori_rounds_sub_ResultXORkey[45]}), .c ({new_AGEMA_signal_3251, new_AGEMA_signal_3250, Midori_rounds_mul_input[45]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_47_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2841, new_AGEMA_signal_2840, Midori_rounds_SR_Result[47]}), .a ({new_AGEMA_signal_3121, new_AGEMA_signal_3120, Midori_rounds_sub_ResultXORkey[47]}), .c ({new_AGEMA_signal_3255, new_AGEMA_signal_3254, Midori_rounds_mul_input[47]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_49_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2837, new_AGEMA_signal_2836, Midori_rounds_SR_Result[49]}), .a ({new_AGEMA_signal_3119, new_AGEMA_signal_3118, Midori_rounds_sub_ResultXORkey[49]}), .c ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, Midori_rounds_mul_input[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_51_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2833, new_AGEMA_signal_2832, Midori_rounds_SR_Result[51]}), .a ({new_AGEMA_signal_3115, new_AGEMA_signal_3114, Midori_rounds_sub_ResultXORkey[51]}), .c ({new_AGEMA_signal_3261, new_AGEMA_signal_3260, Midori_rounds_mul_input[51]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_53_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, Midori_rounds_SR_Result[53]}), .a ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, Midori_rounds_sub_ResultXORkey[53]}), .c ({new_AGEMA_signal_3263, new_AGEMA_signal_3262, Midori_rounds_mul_input[53]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_55_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, Midori_rounds_SR_Result[55]}), .a ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, Midori_rounds_sub_ResultXORkey[55]}), .c ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, Midori_rounds_mul_input[55]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_57_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, Midori_rounds_SR_Result[57]}), .a ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, Midori_rounds_sub_ResultXORkey[57]}), .c ({new_AGEMA_signal_3269, new_AGEMA_signal_3268, Midori_rounds_mul_input[57]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_59_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, Midori_rounds_SR_Result[59]}), .a ({new_AGEMA_signal_3103, new_AGEMA_signal_3102, Midori_rounds_sub_ResultXORkey[59]}), .c ({new_AGEMA_signal_3273, new_AGEMA_signal_3272, Midori_rounds_mul_input[59]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_61_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, Midori_rounds_SR_Result[61]}), .a ({new_AGEMA_signal_3099, new_AGEMA_signal_3098, Midori_rounds_sub_ResultXORkey[61]}), .c ({new_AGEMA_signal_3275, new_AGEMA_signal_3274, Midori_rounds_mul_input[61]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_63_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2953, new_AGEMA_signal_2952, Midori_rounds_SR_Result[63]}), .a ({new_AGEMA_signal_3095, new_AGEMA_signal_3094, Midori_rounds_sub_ResultXORkey[63]}), .c ({new_AGEMA_signal_3279, new_AGEMA_signal_3278, Midori_rounds_mul_input[63]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC1_U24 ( .a ({new_AGEMA_signal_3275, new_AGEMA_signal_3274, Midori_rounds_mul_input[61]}), .b ({new_AGEMA_signal_3287, new_AGEMA_signal_3286, Midori_rounds_mul_MC1_n8}), .c ({new_AGEMA_signal_3329, new_AGEMA_signal_3328, Midori_rounds_SR_Inv_Result[21]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC1_U22 ( .a ({new_AGEMA_signal_3261, new_AGEMA_signal_3260, Midori_rounds_mul_input[51]}), .b ({new_AGEMA_signal_3281, new_AGEMA_signal_3280, Midori_rounds_mul_MC1_n6}), .c ({new_AGEMA_signal_3331, new_AGEMA_signal_3330, Midori_rounds_SR_Inv_Result[43]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC1_U20 ( .a ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, Midori_rounds_mul_input[49]}), .b ({new_AGEMA_signal_3285, new_AGEMA_signal_3284, Midori_rounds_mul_MC1_n4}), .c ({new_AGEMA_signal_3335, new_AGEMA_signal_3334, Midori_rounds_SR_Inv_Result[41]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC1_U18 ( .a ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, Midori_rounds_mul_input[55]}), .b ({new_AGEMA_signal_3281, new_AGEMA_signal_3280, Midori_rounds_mul_MC1_n6}), .c ({new_AGEMA_signal_3337, new_AGEMA_signal_3336, Midori_rounds_SR_Inv_Result[3]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC1_U17 ( .a ({new_AGEMA_signal_3279, new_AGEMA_signal_3278, Midori_rounds_mul_input[63]}), .b ({new_AGEMA_signal_3273, new_AGEMA_signal_3272, Midori_rounds_mul_input[59]}), .c ({new_AGEMA_signal_3281, new_AGEMA_signal_3280, Midori_rounds_mul_MC1_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC1_U14 ( .a ({new_AGEMA_signal_3263, new_AGEMA_signal_3262, Midori_rounds_mul_input[53]}), .b ({new_AGEMA_signal_3285, new_AGEMA_signal_3284, Midori_rounds_mul_MC1_n4}), .c ({new_AGEMA_signal_3341, new_AGEMA_signal_3340, Midori_rounds_SR_Inv_Result[1]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC1_U13 ( .a ({new_AGEMA_signal_3269, new_AGEMA_signal_3268, Midori_rounds_mul_input[57]}), .b ({new_AGEMA_signal_3275, new_AGEMA_signal_3274, Midori_rounds_mul_input[61]}), .c ({new_AGEMA_signal_3285, new_AGEMA_signal_3284, Midori_rounds_mul_MC1_n4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC1_U12 ( .a ({new_AGEMA_signal_3273, new_AGEMA_signal_3272, Midori_rounds_mul_input[59]}), .b ({new_AGEMA_signal_3289, new_AGEMA_signal_3288, Midori_rounds_mul_MC1_n2}), .c ({new_AGEMA_signal_3343, new_AGEMA_signal_3342, Midori_rounds_SR_Inv_Result[63]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC1_U10 ( .a ({new_AGEMA_signal_3269, new_AGEMA_signal_3268, Midori_rounds_mul_input[57]}), .b ({new_AGEMA_signal_3287, new_AGEMA_signal_3286, Midori_rounds_mul_MC1_n8}), .c ({new_AGEMA_signal_3347, new_AGEMA_signal_3346, Midori_rounds_SR_Inv_Result[61]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC1_U9 ( .a ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, Midori_rounds_mul_input[49]}), .b ({new_AGEMA_signal_3263, new_AGEMA_signal_3262, Midori_rounds_mul_input[53]}), .c ({new_AGEMA_signal_3287, new_AGEMA_signal_3286, Midori_rounds_mul_MC1_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC1_U6 ( .a ({new_AGEMA_signal_3279, new_AGEMA_signal_3278, Midori_rounds_mul_input[63]}), .b ({new_AGEMA_signal_3289, new_AGEMA_signal_3288, Midori_rounds_mul_MC1_n2}), .c ({new_AGEMA_signal_3349, new_AGEMA_signal_3348, Midori_rounds_SR_Inv_Result[23]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC1_U5 ( .a ({new_AGEMA_signal_3261, new_AGEMA_signal_3260, Midori_rounds_mul_input[51]}), .b ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, Midori_rounds_mul_input[55]}), .c ({new_AGEMA_signal_3289, new_AGEMA_signal_3288, Midori_rounds_mul_MC1_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC2_U24 ( .a ({new_AGEMA_signal_3251, new_AGEMA_signal_3250, Midori_rounds_mul_input[45]}), .b ({new_AGEMA_signal_3299, new_AGEMA_signal_3298, Midori_rounds_mul_MC2_n8}), .c ({new_AGEMA_signal_3353, new_AGEMA_signal_3352, Midori_rounds_SR_Inv_Result[45]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC2_U22 ( .a ({new_AGEMA_signal_3237, new_AGEMA_signal_3236, Midori_rounds_mul_input[35]}), .b ({new_AGEMA_signal_3293, new_AGEMA_signal_3292, Midori_rounds_mul_MC2_n6}), .c ({new_AGEMA_signal_3355, new_AGEMA_signal_3354, Midori_rounds_SR_Inv_Result[19]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC2_U20 ( .a ({new_AGEMA_signal_3233, new_AGEMA_signal_3232, Midori_rounds_mul_input[33]}), .b ({new_AGEMA_signal_3297, new_AGEMA_signal_3296, Midori_rounds_mul_MC2_n4}), .c ({new_AGEMA_signal_3359, new_AGEMA_signal_3358, Midori_rounds_SR_Inv_Result[17]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC2_U18 ( .a ({new_AGEMA_signal_3243, new_AGEMA_signal_3242, Midori_rounds_mul_input[39]}), .b ({new_AGEMA_signal_3293, new_AGEMA_signal_3292, Midori_rounds_mul_MC2_n6}), .c ({new_AGEMA_signal_3361, new_AGEMA_signal_3360, Midori_rounds_SR_Inv_Result[59]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC2_U17 ( .a ({new_AGEMA_signal_3255, new_AGEMA_signal_3254, Midori_rounds_mul_input[47]}), .b ({new_AGEMA_signal_3249, new_AGEMA_signal_3248, Midori_rounds_mul_input[43]}), .c ({new_AGEMA_signal_3293, new_AGEMA_signal_3292, Midori_rounds_mul_MC2_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC2_U14 ( .a ({new_AGEMA_signal_3239, new_AGEMA_signal_3238, Midori_rounds_mul_input[37]}), .b ({new_AGEMA_signal_3297, new_AGEMA_signal_3296, Midori_rounds_mul_MC2_n4}), .c ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, Midori_rounds_SR_Inv_Result[57]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC2_U13 ( .a ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, Midori_rounds_mul_input[41]}), .b ({new_AGEMA_signal_3251, new_AGEMA_signal_3250, Midori_rounds_mul_input[45]}), .c ({new_AGEMA_signal_3297, new_AGEMA_signal_3296, Midori_rounds_mul_MC2_n4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC2_U12 ( .a ({new_AGEMA_signal_3249, new_AGEMA_signal_3248, Midori_rounds_mul_input[43]}), .b ({new_AGEMA_signal_3301, new_AGEMA_signal_3300, Midori_rounds_mul_MC2_n2}), .c ({new_AGEMA_signal_3367, new_AGEMA_signal_3366, Midori_rounds_SR_Inv_Result[7]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC2_U10 ( .a ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, Midori_rounds_mul_input[41]}), .b ({new_AGEMA_signal_3299, new_AGEMA_signal_3298, Midori_rounds_mul_MC2_n8}), .c ({new_AGEMA_signal_3371, new_AGEMA_signal_3370, Midori_rounds_SR_Inv_Result[5]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC2_U9 ( .a ({new_AGEMA_signal_3233, new_AGEMA_signal_3232, Midori_rounds_mul_input[33]}), .b ({new_AGEMA_signal_3239, new_AGEMA_signal_3238, Midori_rounds_mul_input[37]}), .c ({new_AGEMA_signal_3299, new_AGEMA_signal_3298, Midori_rounds_mul_MC2_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC2_U6 ( .a ({new_AGEMA_signal_3255, new_AGEMA_signal_3254, Midori_rounds_mul_input[47]}), .b ({new_AGEMA_signal_3301, new_AGEMA_signal_3300, Midori_rounds_mul_MC2_n2}), .c ({new_AGEMA_signal_3373, new_AGEMA_signal_3372, Midori_rounds_SR_Inv_Result[47]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC2_U5 ( .a ({new_AGEMA_signal_3237, new_AGEMA_signal_3236, Midori_rounds_mul_input[35]}), .b ({new_AGEMA_signal_3243, new_AGEMA_signal_3242, Midori_rounds_mul_input[39]}), .c ({new_AGEMA_signal_3301, new_AGEMA_signal_3300, Midori_rounds_mul_MC2_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC3_U24 ( .a ({new_AGEMA_signal_3227, new_AGEMA_signal_3226, Midori_rounds_mul_input[29]}), .b ({new_AGEMA_signal_3311, new_AGEMA_signal_3310, Midori_rounds_mul_MC3_n8}), .c ({new_AGEMA_signal_3377, new_AGEMA_signal_3376, Midori_rounds_SR_Inv_Result[49]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC3_U22 ( .a ({new_AGEMA_signal_3213, new_AGEMA_signal_3212, Midori_rounds_mul_input[19]}), .b ({new_AGEMA_signal_3305, new_AGEMA_signal_3304, Midori_rounds_mul_MC3_n6}), .c ({new_AGEMA_signal_3379, new_AGEMA_signal_3378, Midori_rounds_SR_Inv_Result[15]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC3_U20 ( .a ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, Midori_rounds_mul_input[17]}), .b ({new_AGEMA_signal_3309, new_AGEMA_signal_3308, Midori_rounds_mul_MC3_n4}), .c ({new_AGEMA_signal_3383, new_AGEMA_signal_3382, Midori_rounds_SR_Inv_Result[13]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC3_U18 ( .a ({new_AGEMA_signal_3219, new_AGEMA_signal_3218, Midori_rounds_mul_input[23]}), .b ({new_AGEMA_signal_3305, new_AGEMA_signal_3304, Midori_rounds_mul_MC3_n6}), .c ({new_AGEMA_signal_3385, new_AGEMA_signal_3384, Midori_rounds_SR_Inv_Result[39]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC3_U17 ( .a ({new_AGEMA_signal_3231, new_AGEMA_signal_3230, Midori_rounds_mul_input[31]}), .b ({new_AGEMA_signal_3225, new_AGEMA_signal_3224, Midori_rounds_mul_input[27]}), .c ({new_AGEMA_signal_3305, new_AGEMA_signal_3304, Midori_rounds_mul_MC3_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC3_U14 ( .a ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, Midori_rounds_mul_input[21]}), .b ({new_AGEMA_signal_3309, new_AGEMA_signal_3308, Midori_rounds_mul_MC3_n4}), .c ({new_AGEMA_signal_3389, new_AGEMA_signal_3388, Midori_rounds_SR_Inv_Result[37]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC3_U13 ( .a ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, Midori_rounds_mul_input[25]}), .b ({new_AGEMA_signal_3227, new_AGEMA_signal_3226, Midori_rounds_mul_input[29]}), .c ({new_AGEMA_signal_3309, new_AGEMA_signal_3308, Midori_rounds_mul_MC3_n4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC3_U12 ( .a ({new_AGEMA_signal_3225, new_AGEMA_signal_3224, Midori_rounds_mul_input[27]}), .b ({new_AGEMA_signal_3313, new_AGEMA_signal_3312, Midori_rounds_mul_MC3_n2}), .c ({new_AGEMA_signal_3391, new_AGEMA_signal_3390, Midori_rounds_SR_Inv_Result[27]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC3_U10 ( .a ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, Midori_rounds_mul_input[25]}), .b ({new_AGEMA_signal_3311, new_AGEMA_signal_3310, Midori_rounds_mul_MC3_n8}), .c ({new_AGEMA_signal_3395, new_AGEMA_signal_3394, Midori_rounds_SR_Inv_Result[25]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC3_U9 ( .a ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, Midori_rounds_mul_input[17]}), .b ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, Midori_rounds_mul_input[21]}), .c ({new_AGEMA_signal_3311, new_AGEMA_signal_3310, Midori_rounds_mul_MC3_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC3_U6 ( .a ({new_AGEMA_signal_3231, new_AGEMA_signal_3230, Midori_rounds_mul_input[31]}), .b ({new_AGEMA_signal_3313, new_AGEMA_signal_3312, Midori_rounds_mul_MC3_n2}), .c ({new_AGEMA_signal_3397, new_AGEMA_signal_3396, Midori_rounds_SR_Inv_Result[51]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC3_U5 ( .a ({new_AGEMA_signal_3213, new_AGEMA_signal_3212, Midori_rounds_mul_input[19]}), .b ({new_AGEMA_signal_3219, new_AGEMA_signal_3218, Midori_rounds_mul_input[23]}), .c ({new_AGEMA_signal_3313, new_AGEMA_signal_3312, Midori_rounds_mul_MC3_n2}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC4_U24 ( .a ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, Midori_rounds_mul_input[13]}), .b ({new_AGEMA_signal_3323, new_AGEMA_signal_3322, Midori_rounds_mul_MC4_n8}), .c ({new_AGEMA_signal_3401, new_AGEMA_signal_3400, Midori_rounds_SR_Inv_Result[9]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC4_U22 ( .a ({new_AGEMA_signal_3189, new_AGEMA_signal_3188, Midori_rounds_mul_input[3]}), .b ({new_AGEMA_signal_3317, new_AGEMA_signal_3316, Midori_rounds_mul_MC4_n6}), .c ({new_AGEMA_signal_3403, new_AGEMA_signal_3402, Midori_rounds_SR_Inv_Result[55]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC4_U20 ( .a ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, Midori_rounds_mul_input[1]}), .b ({new_AGEMA_signal_3321, new_AGEMA_signal_3320, Midori_rounds_mul_MC4_n4}), .c ({new_AGEMA_signal_3407, new_AGEMA_signal_3406, Midori_rounds_SR_Inv_Result[53]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC4_U18 ( .a ({new_AGEMA_signal_3195, new_AGEMA_signal_3194, Midori_rounds_mul_input[7]}), .b ({new_AGEMA_signal_3317, new_AGEMA_signal_3316, Midori_rounds_mul_MC4_n6}), .c ({new_AGEMA_signal_3409, new_AGEMA_signal_3408, Midori_rounds_SR_Inv_Result[31]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC4_U17 ( .a ({new_AGEMA_signal_3207, new_AGEMA_signal_3206, Midori_rounds_mul_input[15]}), .b ({new_AGEMA_signal_3201, new_AGEMA_signal_3200, Midori_rounds_mul_input[11]}), .c ({new_AGEMA_signal_3317, new_AGEMA_signal_3316, Midori_rounds_mul_MC4_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC4_U14 ( .a ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, Midori_rounds_mul_input[5]}), .b ({new_AGEMA_signal_3321, new_AGEMA_signal_3320, Midori_rounds_mul_MC4_n4}), .c ({new_AGEMA_signal_3413, new_AGEMA_signal_3412, Midori_rounds_SR_Inv_Result[29]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC4_U13 ( .a ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, Midori_rounds_mul_input[9]}), .b ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, Midori_rounds_mul_input[13]}), .c ({new_AGEMA_signal_3321, new_AGEMA_signal_3320, Midori_rounds_mul_MC4_n4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC4_U12 ( .a ({new_AGEMA_signal_3201, new_AGEMA_signal_3200, Midori_rounds_mul_input[11]}), .b ({new_AGEMA_signal_3325, new_AGEMA_signal_3324, Midori_rounds_mul_MC4_n2}), .c ({new_AGEMA_signal_3415, new_AGEMA_signal_3414, Midori_rounds_SR_Inv_Result[35]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC4_U10 ( .a ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, Midori_rounds_mul_input[9]}), .b ({new_AGEMA_signal_3323, new_AGEMA_signal_3322, Midori_rounds_mul_MC4_n8}), .c ({new_AGEMA_signal_3419, new_AGEMA_signal_3418, Midori_rounds_SR_Inv_Result[33]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC4_U9 ( .a ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, Midori_rounds_mul_input[1]}), .b ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, Midori_rounds_mul_input[5]}), .c ({new_AGEMA_signal_3323, new_AGEMA_signal_3322, Midori_rounds_mul_MC4_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC4_U6 ( .a ({new_AGEMA_signal_3207, new_AGEMA_signal_3206, Midori_rounds_mul_input[15]}), .b ({new_AGEMA_signal_3325, new_AGEMA_signal_3324, Midori_rounds_mul_MC4_n2}), .c ({new_AGEMA_signal_3421, new_AGEMA_signal_3420, Midori_rounds_SR_Inv_Result[11]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC4_U5 ( .a ({new_AGEMA_signal_3189, new_AGEMA_signal_3188, Midori_rounds_mul_input[3]}), .b ({new_AGEMA_signal_3195, new_AGEMA_signal_3194, Midori_rounds_mul_input[7]}), .c ({new_AGEMA_signal_3325, new_AGEMA_signal_3324, Midori_rounds_mul_MC4_n2}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_1_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3511, new_AGEMA_signal_3510, Midori_rounds_mul_ResultXORkey[1]}), .a ({new_AGEMA_signal_3341, new_AGEMA_signal_3340, Midori_rounds_SR_Inv_Result[1]}), .c ({new_AGEMA_signal_3557, new_AGEMA_signal_3556, Midori_rounds_round_Result[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_3_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3473, new_AGEMA_signal_3472, Midori_rounds_mul_ResultXORkey[3]}), .a ({new_AGEMA_signal_3337, new_AGEMA_signal_3336, Midori_rounds_SR_Inv_Result[3]}), .c ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, Midori_rounds_round_Result[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_5_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3439, new_AGEMA_signal_3438, Midori_rounds_mul_ResultXORkey[5]}), .a ({new_AGEMA_signal_3371, new_AGEMA_signal_3370, Midori_rounds_SR_Inv_Result[5]}), .c ({new_AGEMA_signal_3563, new_AGEMA_signal_3562, Midori_rounds_round_Result[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_7_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3429, new_AGEMA_signal_3428, Midori_rounds_mul_ResultXORkey[7]}), .a ({new_AGEMA_signal_3367, new_AGEMA_signal_3366, Midori_rounds_SR_Inv_Result[7]}), .c ({new_AGEMA_signal_3567, new_AGEMA_signal_3566, Midori_rounds_round_Result[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_9_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3425, new_AGEMA_signal_3424, Midori_rounds_mul_ResultXORkey[9]}), .a ({new_AGEMA_signal_3401, new_AGEMA_signal_3400, Midori_rounds_SR_Inv_Result[9]}), .c ({new_AGEMA_signal_3569, new_AGEMA_signal_3568, Midori_rounds_round_Result[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_11_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3525, new_AGEMA_signal_3524, Midori_rounds_mul_ResultXORkey[11]}), .a ({new_AGEMA_signal_3421, new_AGEMA_signal_3420, Midori_rounds_SR_Inv_Result[11]}), .c ({new_AGEMA_signal_3573, new_AGEMA_signal_3572, Midori_rounds_round_Result[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_13_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3523, new_AGEMA_signal_3522, Midori_rounds_mul_ResultXORkey[13]}), .a ({new_AGEMA_signal_3383, new_AGEMA_signal_3382, Midori_rounds_SR_Inv_Result[13]}), .c ({new_AGEMA_signal_3575, new_AGEMA_signal_3574, Midori_rounds_round_Result[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_15_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3519, new_AGEMA_signal_3518, Midori_rounds_mul_ResultXORkey[15]}), .a ({new_AGEMA_signal_3379, new_AGEMA_signal_3378, Midori_rounds_SR_Inv_Result[15]}), .c ({new_AGEMA_signal_3579, new_AGEMA_signal_3578, Midori_rounds_round_Result[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_17_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3517, new_AGEMA_signal_3516, Midori_rounds_mul_ResultXORkey[17]}), .a ({new_AGEMA_signal_3359, new_AGEMA_signal_3358, Midori_rounds_SR_Inv_Result[17]}), .c ({new_AGEMA_signal_3581, new_AGEMA_signal_3580, Midori_rounds_round_Result[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_19_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3513, new_AGEMA_signal_3512, Midori_rounds_mul_ResultXORkey[19]}), .a ({new_AGEMA_signal_3355, new_AGEMA_signal_3354, Midori_rounds_SR_Inv_Result[19]}), .c ({new_AGEMA_signal_3585, new_AGEMA_signal_3584, Midori_rounds_round_Result[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_21_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3507, new_AGEMA_signal_3506, Midori_rounds_mul_ResultXORkey[21]}), .a ({new_AGEMA_signal_3329, new_AGEMA_signal_3328, Midori_rounds_SR_Inv_Result[21]}), .c ({new_AGEMA_signal_3587, new_AGEMA_signal_3586, Midori_rounds_round_Result[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_23_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3503, new_AGEMA_signal_3502, Midori_rounds_mul_ResultXORkey[23]}), .a ({new_AGEMA_signal_3349, new_AGEMA_signal_3348, Midori_rounds_SR_Inv_Result[23]}), .c ({new_AGEMA_signal_3591, new_AGEMA_signal_3590, Midori_rounds_round_Result[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_25_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3501, new_AGEMA_signal_3500, Midori_rounds_mul_ResultXORkey[25]}), .a ({new_AGEMA_signal_3395, new_AGEMA_signal_3394, Midori_rounds_SR_Inv_Result[25]}), .c ({new_AGEMA_signal_3593, new_AGEMA_signal_3592, Midori_rounds_round_Result[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_27_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3497, new_AGEMA_signal_3496, Midori_rounds_mul_ResultXORkey[27]}), .a ({new_AGEMA_signal_3391, new_AGEMA_signal_3390, Midori_rounds_SR_Inv_Result[27]}), .c ({new_AGEMA_signal_3597, new_AGEMA_signal_3596, Midori_rounds_round_Result[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_29_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3495, new_AGEMA_signal_3494, Midori_rounds_mul_ResultXORkey[29]}), .a ({new_AGEMA_signal_3413, new_AGEMA_signal_3412, Midori_rounds_SR_Inv_Result[29]}), .c ({new_AGEMA_signal_3599, new_AGEMA_signal_3598, Midori_rounds_round_Result[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_31_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3489, new_AGEMA_signal_3488, Midori_rounds_mul_ResultXORkey[31]}), .a ({new_AGEMA_signal_3409, new_AGEMA_signal_3408, Midori_rounds_SR_Inv_Result[31]}), .c ({new_AGEMA_signal_3603, new_AGEMA_signal_3602, Midori_rounds_round_Result[31]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_33_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3487, new_AGEMA_signal_3486, Midori_rounds_mul_ResultXORkey[33]}), .a ({new_AGEMA_signal_3419, new_AGEMA_signal_3418, Midori_rounds_SR_Inv_Result[33]}), .c ({new_AGEMA_signal_3605, new_AGEMA_signal_3604, Midori_rounds_round_Result[33]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_35_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3483, new_AGEMA_signal_3482, Midori_rounds_mul_ResultXORkey[35]}), .a ({new_AGEMA_signal_3415, new_AGEMA_signal_3414, Midori_rounds_SR_Inv_Result[35]}), .c ({new_AGEMA_signal_3609, new_AGEMA_signal_3608, Midori_rounds_round_Result[35]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_37_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3479, new_AGEMA_signal_3478, Midori_rounds_mul_ResultXORkey[37]}), .a ({new_AGEMA_signal_3389, new_AGEMA_signal_3388, Midori_rounds_SR_Inv_Result[37]}), .c ({new_AGEMA_signal_3611, new_AGEMA_signal_3610, Midori_rounds_round_Result[37]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_39_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3475, new_AGEMA_signal_3474, Midori_rounds_mul_ResultXORkey[39]}), .a ({new_AGEMA_signal_3385, new_AGEMA_signal_3384, Midori_rounds_SR_Inv_Result[39]}), .c ({new_AGEMA_signal_3615, new_AGEMA_signal_3614, Midori_rounds_round_Result[39]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_41_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3471, new_AGEMA_signal_3470, Midori_rounds_mul_ResultXORkey[41]}), .a ({new_AGEMA_signal_3335, new_AGEMA_signal_3334, Midori_rounds_SR_Inv_Result[41]}), .c ({new_AGEMA_signal_3617, new_AGEMA_signal_3616, Midori_rounds_round_Result[41]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_43_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3467, new_AGEMA_signal_3466, Midori_rounds_mul_ResultXORkey[43]}), .a ({new_AGEMA_signal_3331, new_AGEMA_signal_3330, Midori_rounds_SR_Inv_Result[43]}), .c ({new_AGEMA_signal_3621, new_AGEMA_signal_3620, Midori_rounds_round_Result[43]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_45_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3463, new_AGEMA_signal_3462, Midori_rounds_mul_ResultXORkey[45]}), .a ({new_AGEMA_signal_3353, new_AGEMA_signal_3352, Midori_rounds_SR_Inv_Result[45]}), .c ({new_AGEMA_signal_3623, new_AGEMA_signal_3622, Midori_rounds_round_Result[45]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_47_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3459, new_AGEMA_signal_3458, Midori_rounds_mul_ResultXORkey[47]}), .a ({new_AGEMA_signal_3373, new_AGEMA_signal_3372, Midori_rounds_SR_Inv_Result[47]}), .c ({new_AGEMA_signal_3627, new_AGEMA_signal_3626, Midori_rounds_round_Result[47]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_49_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3457, new_AGEMA_signal_3456, Midori_rounds_mul_ResultXORkey[49]}), .a ({new_AGEMA_signal_3377, new_AGEMA_signal_3376, Midori_rounds_SR_Inv_Result[49]}), .c ({new_AGEMA_signal_3629, new_AGEMA_signal_3628, Midori_rounds_round_Result[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_51_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3453, new_AGEMA_signal_3452, Midori_rounds_mul_ResultXORkey[51]}), .a ({new_AGEMA_signal_3397, new_AGEMA_signal_3396, Midori_rounds_SR_Inv_Result[51]}), .c ({new_AGEMA_signal_3633, new_AGEMA_signal_3632, Midori_rounds_round_Result[51]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_53_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3451, new_AGEMA_signal_3450, Midori_rounds_mul_ResultXORkey[53]}), .a ({new_AGEMA_signal_3407, new_AGEMA_signal_3406, Midori_rounds_SR_Inv_Result[53]}), .c ({new_AGEMA_signal_3635, new_AGEMA_signal_3634, Midori_rounds_round_Result[53]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_55_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3447, new_AGEMA_signal_3446, Midori_rounds_mul_ResultXORkey[55]}), .a ({new_AGEMA_signal_3403, new_AGEMA_signal_3402, Midori_rounds_SR_Inv_Result[55]}), .c ({new_AGEMA_signal_3639, new_AGEMA_signal_3638, Midori_rounds_round_Result[55]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_57_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3445, new_AGEMA_signal_3444, Midori_rounds_mul_ResultXORkey[57]}), .a ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, Midori_rounds_SR_Inv_Result[57]}), .c ({new_AGEMA_signal_3641, new_AGEMA_signal_3640, Midori_rounds_round_Result[57]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_59_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3441, new_AGEMA_signal_3440, Midori_rounds_mul_ResultXORkey[59]}), .a ({new_AGEMA_signal_3361, new_AGEMA_signal_3360, Midori_rounds_SR_Inv_Result[59]}), .c ({new_AGEMA_signal_3645, new_AGEMA_signal_3644, Midori_rounds_round_Result[59]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_61_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3437, new_AGEMA_signal_3436, Midori_rounds_mul_ResultXORkey[61]}), .a ({new_AGEMA_signal_3347, new_AGEMA_signal_3346, Midori_rounds_SR_Inv_Result[61]}), .c ({new_AGEMA_signal_3647, new_AGEMA_signal_3646, Midori_rounds_round_Result[61]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_63_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3433, new_AGEMA_signal_3432, Midori_rounds_mul_ResultXORkey[63]}), .a ({new_AGEMA_signal_3343, new_AGEMA_signal_3342, Midori_rounds_SR_Inv_Result[63]}), .c ({new_AGEMA_signal_3651, new_AGEMA_signal_3650, Midori_rounds_round_Result[63]}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U127 ( .a ({new_AGEMA_signal_1467, new_AGEMA_signal_1466, wk[8]}), .b ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, Midori_rounds_SR_Result[8]}), .c ({DataOut_s2[8], DataOut_s1[8], DataOut_s0[8]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U125 ( .a ({new_AGEMA_signal_1479, new_AGEMA_signal_1478, wk[6]}), .b ({new_AGEMA_signal_2843, new_AGEMA_signal_2842, Midori_rounds_SR_Result[46]}), .c ({DataOut_s2[6], DataOut_s1[6], DataOut_s0[6]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U123 ( .a ({new_AGEMA_signal_1491, new_AGEMA_signal_1490, wk[62]}), .b ({new_AGEMA_signal_2955, new_AGEMA_signal_2954, Midori_rounds_SR_Result[62]}), .c ({DataOut_s2[62], DataOut_s1[62], DataOut_s0[62]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U121 ( .a ({new_AGEMA_signal_1503, new_AGEMA_signal_1502, wk[60]}), .b ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, Midori_rounds_SR_Result[60]}), .c ({DataOut_s2[60], DataOut_s1[60], DataOut_s0[60]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U118 ( .a ({new_AGEMA_signal_1521, new_AGEMA_signal_1520, wk[58]}), .b ({new_AGEMA_signal_2947, new_AGEMA_signal_2946, Midori_rounds_SR_Result[34]}), .c ({DataOut_s2[58], DataOut_s1[58], DataOut_s0[58]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U116 ( .a ({new_AGEMA_signal_1533, new_AGEMA_signal_1532, wk[56]}), .b ({new_AGEMA_signal_2951, new_AGEMA_signal_2950, Midori_rounds_SR_Result[32]}), .c ({DataOut_s2[56], DataOut_s1[56], DataOut_s0[56]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U114 ( .a ({new_AGEMA_signal_1545, new_AGEMA_signal_1544, wk[54]}), .b ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, Midori_rounds_SR_Result[6]}), .c ({DataOut_s2[54], DataOut_s1[54], DataOut_s0[54]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U112 ( .a ({new_AGEMA_signal_1557, new_AGEMA_signal_1556, wk[52]}), .b ({new_AGEMA_signal_2943, new_AGEMA_signal_2942, Midori_rounds_SR_Result[4]}), .c ({DataOut_s2[52], DataOut_s1[52], DataOut_s0[52]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U110 ( .a ({new_AGEMA_signal_1569, new_AGEMA_signal_1568, wk[50]}), .b ({new_AGEMA_signal_2931, new_AGEMA_signal_2930, Midori_rounds_SR_Result[26]}), .c ({DataOut_s2[50], DataOut_s1[50], DataOut_s0[50]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U109 ( .a ({new_AGEMA_signal_1575, new_AGEMA_signal_1574, wk[4]}), .b ({new_AGEMA_signal_2847, new_AGEMA_signal_2846, Midori_rounds_SR_Result[44]}), .c ({DataOut_s2[4], DataOut_s1[4], DataOut_s0[4]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U107 ( .a ({new_AGEMA_signal_1587, new_AGEMA_signal_1586, wk[48]}), .b ({new_AGEMA_signal_2935, new_AGEMA_signal_2934, Midori_rounds_SR_Result[24]}), .c ({DataOut_s2[48], DataOut_s1[48], DataOut_s0[48]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U105 ( .a ({new_AGEMA_signal_1599, new_AGEMA_signal_1598, wk[46]}), .b ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, Midori_rounds_SR_Result[42]}), .c ({DataOut_s2[46], DataOut_s1[46], DataOut_s0[46]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U103 ( .a ({new_AGEMA_signal_1611, new_AGEMA_signal_1610, wk[44]}), .b ({new_AGEMA_signal_2927, new_AGEMA_signal_2926, Midori_rounds_SR_Result[40]}), .c ({DataOut_s2[44], DataOut_s1[44], DataOut_s0[44]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U101 ( .a ({new_AGEMA_signal_1623, new_AGEMA_signal_1622, wk[42]}), .b ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, Midori_rounds_SR_Result[54]}), .c ({DataOut_s2[42], DataOut_s1[42], DataOut_s0[42]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U99 ( .a ({new_AGEMA_signal_1635, new_AGEMA_signal_1634, wk[40]}), .b ({new_AGEMA_signal_2919, new_AGEMA_signal_2918, Midori_rounds_SR_Result[52]}), .c ({DataOut_s2[40], DataOut_s1[40], DataOut_s0[40]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U96 ( .a ({new_AGEMA_signal_1653, new_AGEMA_signal_1652, wk[38]}), .b ({new_AGEMA_signal_2907, new_AGEMA_signal_2906, Midori_rounds_SR_Result[18]}), .c ({DataOut_s2[38], DataOut_s1[38], DataOut_s0[38]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U94 ( .a ({new_AGEMA_signal_1665, new_AGEMA_signal_1664, wk[36]}), .b ({new_AGEMA_signal_2911, new_AGEMA_signal_2910, Midori_rounds_SR_Result[16]}), .c ({DataOut_s2[36], DataOut_s1[36], DataOut_s0[36]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U92 ( .a ({new_AGEMA_signal_1677, new_AGEMA_signal_1676, wk[34]}), .b ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, Midori_rounds_SR_Result[14]}), .c ({DataOut_s2[34], DataOut_s1[34], DataOut_s0[34]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U90 ( .a ({new_AGEMA_signal_1689, new_AGEMA_signal_1688, wk[32]}), .b ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, Midori_rounds_SR_Result[12]}), .c ({DataOut_s2[32], DataOut_s1[32], DataOut_s0[32]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U88 ( .a ({new_AGEMA_signal_1701, new_AGEMA_signal_1700, wk[30]}), .b ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, Midori_rounds_SR_Result[2]}), .c ({DataOut_s2[30], DataOut_s1[30], DataOut_s0[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U87 ( .a ({new_AGEMA_signal_1707, new_AGEMA_signal_1706, wk[2]}), .b ({new_AGEMA_signal_2835, new_AGEMA_signal_2834, Midori_rounds_SR_Result[50]}), .c ({DataOut_s2[2], DataOut_s1[2], DataOut_s0[2]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U85 ( .a ({new_AGEMA_signal_1719, new_AGEMA_signal_1718, wk[28]}), .b ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, Midori_rounds_SR_Result[0]}), .c ({DataOut_s2[28], DataOut_s1[28], DataOut_s0[28]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U83 ( .a ({new_AGEMA_signal_1731, new_AGEMA_signal_1730, wk[26]}), .b ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, Midori_rounds_SR_Result[30]}), .c ({DataOut_s2[26], DataOut_s1[26], DataOut_s0[26]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U81 ( .a ({new_AGEMA_signal_1743, new_AGEMA_signal_1742, wk[24]}), .b ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, Midori_rounds_SR_Result[28]}), .c ({DataOut_s2[24], DataOut_s1[24], DataOut_s0[24]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U79 ( .a ({new_AGEMA_signal_1755, new_AGEMA_signal_1754, wk[22]}), .b ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, Midori_rounds_SR_Result[58]}), .c ({DataOut_s2[22], DataOut_s1[22], DataOut_s0[22]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U77 ( .a ({new_AGEMA_signal_1767, new_AGEMA_signal_1766, wk[20]}), .b ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, Midori_rounds_SR_Result[56]}), .c ({DataOut_s2[20], DataOut_s1[20], DataOut_s0[20]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U74 ( .a ({new_AGEMA_signal_1785, new_AGEMA_signal_1784, wk[18]}), .b ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, Midori_rounds_SR_Result[38]}), .c ({DataOut_s2[18], DataOut_s1[18], DataOut_s0[18]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U72 ( .a ({new_AGEMA_signal_1797, new_AGEMA_signal_1796, wk[16]}), .b ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, Midori_rounds_SR_Result[36]}), .c ({DataOut_s2[16], DataOut_s1[16], DataOut_s0[16]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U70 ( .a ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, wk[14]}), .b ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, Midori_rounds_SR_Result[22]}), .c ({DataOut_s2[14], DataOut_s1[14], DataOut_s0[14]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U68 ( .a ({new_AGEMA_signal_1821, new_AGEMA_signal_1820, wk[12]}), .b ({new_AGEMA_signal_2863, new_AGEMA_signal_2862, Midori_rounds_SR_Result[20]}), .c ({DataOut_s2[12], DataOut_s1[12], DataOut_s0[12]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U66 ( .a ({new_AGEMA_signal_1833, new_AGEMA_signal_1832, wk[10]}), .b ({new_AGEMA_signal_2851, new_AGEMA_signal_2850, Midori_rounds_SR_Result[10]}), .c ({DataOut_s2[10], DataOut_s1[10], DataOut_s0[10]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_U65 ( .a ({new_AGEMA_signal_1839, new_AGEMA_signal_1838, wk[0]}), .b ({new_AGEMA_signal_2839, new_AGEMA_signal_2838, Midori_rounds_SR_Result[48]}), .c ({DataOut_s2[0], DataOut_s1[0], DataOut_s0[0]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U143 ( .a ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, Midori_rounds_SR_Result[8]}), .b ({new_AGEMA_signal_3427, new_AGEMA_signal_3426, Midori_rounds_n16}), .c ({new_AGEMA_signal_3529, new_AGEMA_signal_3528, Midori_rounds_sub_ResultXORkey[8]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U141 ( .a ({new_AGEMA_signal_2573, new_AGEMA_signal_2572, Midori_rounds_SelectedKey_6_}), .b ({new_AGEMA_signal_2843, new_AGEMA_signal_2842, Midori_rounds_SR_Result[46]}), .c ({new_AGEMA_signal_3093, new_AGEMA_signal_3092, Midori_rounds_sub_ResultXORkey[6]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U139 ( .a ({new_AGEMA_signal_2669, new_AGEMA_signal_2668, Midori_rounds_SelectedKey_62_}), .b ({new_AGEMA_signal_2955, new_AGEMA_signal_2954, Midori_rounds_SR_Result[62]}), .c ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, Midori_rounds_sub_ResultXORkey[62]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U137 ( .a ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, Midori_rounds_SR_Result[60]}), .b ({new_AGEMA_signal_3537, new_AGEMA_signal_3536, Midori_rounds_n15}), .c ({new_AGEMA_signal_3653, new_AGEMA_signal_3652, Midori_rounds_sub_ResultXORkey[60]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U134 ( .a ({new_AGEMA_signal_2661, new_AGEMA_signal_2660, Midori_rounds_SelectedKey_58_}), .b ({new_AGEMA_signal_2947, new_AGEMA_signal_2946, Midori_rounds_SR_Result[34]}), .c ({new_AGEMA_signal_3105, new_AGEMA_signal_3104, Midori_rounds_sub_ResultXORkey[58]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U132 ( .a ({new_AGEMA_signal_2951, new_AGEMA_signal_2950, Midori_rounds_SR_Result[32]}), .b ({new_AGEMA_signal_3539, new_AGEMA_signal_3538, Midori_rounds_n14}), .c ({new_AGEMA_signal_3655, new_AGEMA_signal_3654, Midori_rounds_sub_ResultXORkey[56]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U130 ( .a ({new_AGEMA_signal_2653, new_AGEMA_signal_2652, Midori_rounds_SelectedKey_54_}), .b ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, Midori_rounds_SR_Result[6]}), .c ({new_AGEMA_signal_3111, new_AGEMA_signal_3110, Midori_rounds_sub_ResultXORkey[54]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U128 ( .a ({new_AGEMA_signal_2943, new_AGEMA_signal_2942, Midori_rounds_SR_Result[4]}), .b ({new_AGEMA_signal_3541, new_AGEMA_signal_3540, Midori_rounds_n13}), .c ({new_AGEMA_signal_3657, new_AGEMA_signal_3656, Midori_rounds_sub_ResultXORkey[52]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U126 ( .a ({new_AGEMA_signal_2645, new_AGEMA_signal_2644, Midori_rounds_SelectedKey_50_}), .b ({new_AGEMA_signal_2931, new_AGEMA_signal_2930, Midori_rounds_SR_Result[26]}), .c ({new_AGEMA_signal_3117, new_AGEMA_signal_3116, Midori_rounds_sub_ResultXORkey[50]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U125 ( .a ({new_AGEMA_signal_2847, new_AGEMA_signal_2846, Midori_rounds_SR_Result[44]}), .b ({new_AGEMA_signal_3543, new_AGEMA_signal_3542, Midori_rounds_n12}), .c ({new_AGEMA_signal_3659, new_AGEMA_signal_3658, Midori_rounds_sub_ResultXORkey[4]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U123 ( .a ({new_AGEMA_signal_2935, new_AGEMA_signal_2934, Midori_rounds_SR_Result[24]}), .b ({new_AGEMA_signal_3781, new_AGEMA_signal_3780, Midori_rounds_n11}), .c ({new_AGEMA_signal_3803, new_AGEMA_signal_3802, Midori_rounds_sub_ResultXORkey[48]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U121 ( .a ({new_AGEMA_signal_2637, new_AGEMA_signal_2636, Midori_rounds_SelectedKey_46_}), .b ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, Midori_rounds_SR_Result[42]}), .c ({new_AGEMA_signal_3123, new_AGEMA_signal_3122, Midori_rounds_sub_ResultXORkey[46]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U119 ( .a ({new_AGEMA_signal_2927, new_AGEMA_signal_2926, Midori_rounds_SR_Result[40]}), .b ({new_AGEMA_signal_3465, new_AGEMA_signal_3464, Midori_rounds_n10}), .c ({new_AGEMA_signal_3531, new_AGEMA_signal_3530, Midori_rounds_sub_ResultXORkey[44]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U117 ( .a ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, Midori_rounds_SelectedKey_42_}), .b ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, Midori_rounds_SR_Result[54]}), .c ({new_AGEMA_signal_3129, new_AGEMA_signal_3128, Midori_rounds_sub_ResultXORkey[42]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U115 ( .a ({new_AGEMA_signal_2919, new_AGEMA_signal_2918, Midori_rounds_SR_Result[52]}), .b ({new_AGEMA_signal_3545, new_AGEMA_signal_3544, Midori_rounds_n9}), .c ({new_AGEMA_signal_3661, new_AGEMA_signal_3660, Midori_rounds_sub_ResultXORkey[40]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U112 ( .a ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, Midori_rounds_SelectedKey_38_}), .b ({new_AGEMA_signal_2907, new_AGEMA_signal_2906, Midori_rounds_SR_Result[18]}), .c ({new_AGEMA_signal_3137, new_AGEMA_signal_3136, Midori_rounds_sub_ResultXORkey[38]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U110 ( .a ({new_AGEMA_signal_2911, new_AGEMA_signal_2910, Midori_rounds_SR_Result[16]}), .b ({new_AGEMA_signal_3481, new_AGEMA_signal_3480, Midori_rounds_n8}), .c ({new_AGEMA_signal_3533, new_AGEMA_signal_3532, Midori_rounds_sub_ResultXORkey[36]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U108 ( .a ({new_AGEMA_signal_2613, new_AGEMA_signal_2612, Midori_rounds_SelectedKey_34_}), .b ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, Midori_rounds_SR_Result[14]}), .c ({new_AGEMA_signal_3143, new_AGEMA_signal_3142, Midori_rounds_sub_ResultXORkey[34]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U106 ( .a ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, Midori_rounds_SR_Result[12]}), .b ({new_AGEMA_signal_3547, new_AGEMA_signal_3546, Midori_rounds_n7}), .c ({new_AGEMA_signal_3663, new_AGEMA_signal_3662, Midori_rounds_sub_ResultXORkey[32]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U104 ( .a ({new_AGEMA_signal_2605, new_AGEMA_signal_2604, Midori_rounds_SelectedKey_30_}), .b ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, Midori_rounds_SR_Result[2]}), .c ({new_AGEMA_signal_3149, new_AGEMA_signal_3148, Midori_rounds_sub_ResultXORkey[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U103 ( .a ({new_AGEMA_signal_1845, new_AGEMA_signal_1844, Midori_rounds_SelectedKey_2_}), .b ({new_AGEMA_signal_2835, new_AGEMA_signal_2834, Midori_rounds_SR_Result[50]}), .c ({new_AGEMA_signal_3151, new_AGEMA_signal_3150, Midori_rounds_sub_ResultXORkey[2]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U101 ( .a ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, Midori_rounds_SR_Result[0]}), .b ({new_AGEMA_signal_3673, new_AGEMA_signal_3672, Midori_rounds_n6}), .c ({new_AGEMA_signal_3779, new_AGEMA_signal_3778, Midori_rounds_sub_ResultXORkey[28]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U99 ( .a ({new_AGEMA_signal_1865, new_AGEMA_signal_1864, Midori_rounds_SelectedKey_26_}), .b ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, Midori_rounds_SR_Result[30]}), .c ({new_AGEMA_signal_3157, new_AGEMA_signal_3156, Midori_rounds_sub_ResultXORkey[26]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U97 ( .a ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, Midori_rounds_SR_Result[28]}), .b ({new_AGEMA_signal_3549, new_AGEMA_signal_3548, Midori_rounds_n5}), .c ({new_AGEMA_signal_3665, new_AGEMA_signal_3664, Midori_rounds_sub_ResultXORkey[24]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U95 ( .a ({new_AGEMA_signal_2591, new_AGEMA_signal_2590, Midori_rounds_SelectedKey_22_}), .b ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, Midori_rounds_SR_Result[58]}), .c ({new_AGEMA_signal_3163, new_AGEMA_signal_3162, Midori_rounds_sub_ResultXORkey[22]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U93 ( .a ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, Midori_rounds_SR_Result[56]}), .b ({new_AGEMA_signal_3509, new_AGEMA_signal_3508, Midori_rounds_n4}), .c ({new_AGEMA_signal_3535, new_AGEMA_signal_3534, Midori_rounds_sub_ResultXORkey[20]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U90 ( .a ({new_AGEMA_signal_2583, new_AGEMA_signal_2582, Midori_rounds_SelectedKey_18_}), .b ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, Midori_rounds_SR_Result[38]}), .c ({new_AGEMA_signal_3171, new_AGEMA_signal_3170, Midori_rounds_sub_ResultXORkey[18]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U88 ( .a ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, Midori_rounds_SR_Result[36]}), .b ({new_AGEMA_signal_3551, new_AGEMA_signal_3550, Midori_rounds_n3}), .c ({new_AGEMA_signal_3667, new_AGEMA_signal_3666, Midori_rounds_sub_ResultXORkey[16]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U86 ( .a ({new_AGEMA_signal_1861, new_AGEMA_signal_1860, Midori_rounds_SelectedKey_14_}), .b ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, Midori_rounds_SR_Result[22]}), .c ({new_AGEMA_signal_3177, new_AGEMA_signal_3176, Midori_rounds_sub_ResultXORkey[14]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U84 ( .a ({new_AGEMA_signal_2863, new_AGEMA_signal_2862, Midori_rounds_SR_Result[20]}), .b ({new_AGEMA_signal_3553, new_AGEMA_signal_3552, Midori_rounds_n2}), .c ({new_AGEMA_signal_3669, new_AGEMA_signal_3668, Midori_rounds_sub_ResultXORkey[12]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U82 ( .a ({new_AGEMA_signal_1855, new_AGEMA_signal_1854, Midori_rounds_SelectedKey_10_}), .b ({new_AGEMA_signal_2851, new_AGEMA_signal_2850, Midori_rounds_SR_Result[10]}), .c ({new_AGEMA_signal_3183, new_AGEMA_signal_3182, Midori_rounds_sub_ResultXORkey[10]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U81 ( .a ({new_AGEMA_signal_2839, new_AGEMA_signal_2838, Midori_rounds_SR_Result[48]}), .b ({new_AGEMA_signal_3555, new_AGEMA_signal_3554, Midori_rounds_n1}), .c ({new_AGEMA_signal_3671, new_AGEMA_signal_3670, Midori_rounds_sub_ResultXORkey[0]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U79 ( .a ({new_AGEMA_signal_3837, new_AGEMA_signal_3836, Midori_rounds_SR_Inv_Result[8]}), .b ({new_AGEMA_signal_3427, new_AGEMA_signal_3426, Midori_rounds_n16}), .c ({new_AGEMA_signal_3845, new_AGEMA_signal_3844, Midori_rounds_mul_ResultXORkey[8]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U76 ( .a ({new_AGEMA_signal_2573, new_AGEMA_signal_2572, Midori_rounds_SelectedKey_6_}), .b ({new_AGEMA_signal_3405, new_AGEMA_signal_3404, Midori_rounds_SR_Inv_Result[54]}), .c ({new_AGEMA_signal_3431, new_AGEMA_signal_3430, Midori_rounds_mul_ResultXORkey[6]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U74 ( .a ({new_AGEMA_signal_2669, new_AGEMA_signal_2668, Midori_rounds_SelectedKey_62_}), .b ({new_AGEMA_signal_3345, new_AGEMA_signal_3344, Midori_rounds_SR_Inv_Result[62]}), .c ({new_AGEMA_signal_3435, new_AGEMA_signal_3434, Midori_rounds_mul_ResultXORkey[62]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U72 ( .a ({new_AGEMA_signal_3883, new_AGEMA_signal_3882, Midori_rounds_SR_Inv_Result[60]}), .b ({new_AGEMA_signal_3537, new_AGEMA_signal_3536, Midori_rounds_n15}), .c ({new_AGEMA_signal_3907, new_AGEMA_signal_3906, Midori_rounds_mul_ResultXORkey[60]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U68 ( .a ({new_AGEMA_signal_2661, new_AGEMA_signal_2660, Midori_rounds_SelectedKey_58_}), .b ({new_AGEMA_signal_3351, new_AGEMA_signal_3350, Midori_rounds_SR_Inv_Result[22]}), .c ({new_AGEMA_signal_3443, new_AGEMA_signal_3442, Midori_rounds_mul_ResultXORkey[58]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U66 ( .a ({new_AGEMA_signal_3881, new_AGEMA_signal_3880, Midori_rounds_SR_Inv_Result[20]}), .b ({new_AGEMA_signal_3539, new_AGEMA_signal_3538, Midori_rounds_n14}), .c ({new_AGEMA_signal_3909, new_AGEMA_signal_3908, Midori_rounds_mul_ResultXORkey[56]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U63 ( .a ({new_AGEMA_signal_2653, new_AGEMA_signal_2652, Midori_rounds_SelectedKey_54_}), .b ({new_AGEMA_signal_3333, new_AGEMA_signal_3332, Midori_rounds_SR_Inv_Result[42]}), .c ({new_AGEMA_signal_3449, new_AGEMA_signal_3448, Midori_rounds_mul_ResultXORkey[54]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U61 ( .a ({new_AGEMA_signal_3867, new_AGEMA_signal_3866, Midori_rounds_SR_Inv_Result[40]}), .b ({new_AGEMA_signal_3541, new_AGEMA_signal_3540, Midori_rounds_n13}), .c ({new_AGEMA_signal_3875, new_AGEMA_signal_3874, Midori_rounds_mul_ResultXORkey[52]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U58 ( .a ({new_AGEMA_signal_2645, new_AGEMA_signal_2644, Midori_rounds_SelectedKey_50_}), .b ({new_AGEMA_signal_3339, new_AGEMA_signal_3338, Midori_rounds_SR_Inv_Result[2]}), .c ({new_AGEMA_signal_3455, new_AGEMA_signal_3454, Midori_rounds_mul_ResultXORkey[50]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U57 ( .a ({new_AGEMA_signal_3839, new_AGEMA_signal_3838, Midori_rounds_SR_Inv_Result[52]}), .b ({new_AGEMA_signal_3543, new_AGEMA_signal_3542, Midori_rounds_n12}), .c ({new_AGEMA_signal_3847, new_AGEMA_signal_3846, Midori_rounds_mul_ResultXORkey[4]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U54 ( .a ({new_AGEMA_signal_3821, new_AGEMA_signal_3820, Midori_rounds_SR_Inv_Result[0]}), .b ({new_AGEMA_signal_3781, new_AGEMA_signal_3780, Midori_rounds_n11}), .c ({new_AGEMA_signal_3849, new_AGEMA_signal_3848, Midori_rounds_mul_ResultXORkey[48]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U51 ( .a ({new_AGEMA_signal_2637, new_AGEMA_signal_2636, Midori_rounds_SelectedKey_46_}), .b ({new_AGEMA_signal_3369, new_AGEMA_signal_3368, Midori_rounds_SR_Inv_Result[6]}), .c ({new_AGEMA_signal_3461, new_AGEMA_signal_3460, Midori_rounds_mul_ResultXORkey[46]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U49 ( .a ({new_AGEMA_signal_3827, new_AGEMA_signal_3826, Midori_rounds_SR_Inv_Result[4]}), .b ({new_AGEMA_signal_3465, new_AGEMA_signal_3464, Midori_rounds_n10}), .c ({new_AGEMA_signal_3851, new_AGEMA_signal_3850, Midori_rounds_mul_ResultXORkey[44]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U46 ( .a ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, Midori_rounds_SelectedKey_42_}), .b ({new_AGEMA_signal_3375, new_AGEMA_signal_3374, Midori_rounds_SR_Inv_Result[46]}), .c ({new_AGEMA_signal_3469, new_AGEMA_signal_3468, Midori_rounds_mul_ResultXORkey[42]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U44 ( .a ({new_AGEMA_signal_3823, new_AGEMA_signal_3822, Midori_rounds_SR_Inv_Result[44]}), .b ({new_AGEMA_signal_3545, new_AGEMA_signal_3544, Midori_rounds_n9}), .c ({new_AGEMA_signal_3853, new_AGEMA_signal_3852, Midori_rounds_mul_ResultXORkey[40]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U40 ( .a ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, Midori_rounds_SelectedKey_38_}), .b ({new_AGEMA_signal_3357, new_AGEMA_signal_3356, Midori_rounds_SR_Inv_Result[18]}), .c ({new_AGEMA_signal_3477, new_AGEMA_signal_3476, Midori_rounds_mul_ResultXORkey[38]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U38 ( .a ({new_AGEMA_signal_3825, new_AGEMA_signal_3824, Midori_rounds_SR_Inv_Result[16]}), .b ({new_AGEMA_signal_3481, new_AGEMA_signal_3480, Midori_rounds_n8}), .c ({new_AGEMA_signal_3855, new_AGEMA_signal_3854, Midori_rounds_mul_ResultXORkey[36]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U35 ( .a ({new_AGEMA_signal_2613, new_AGEMA_signal_2612, Midori_rounds_SelectedKey_34_}), .b ({new_AGEMA_signal_3363, new_AGEMA_signal_3362, Midori_rounds_SR_Inv_Result[58]}), .c ({new_AGEMA_signal_3485, new_AGEMA_signal_3484, Midori_rounds_mul_ResultXORkey[34]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U33 ( .a ({new_AGEMA_signal_3829, new_AGEMA_signal_3828, Midori_rounds_SR_Inv_Result[56]}), .b ({new_AGEMA_signal_3547, new_AGEMA_signal_3546, Midori_rounds_n7}), .c ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, Midori_rounds_mul_ResultXORkey[32]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U30 ( .a ({new_AGEMA_signal_2605, new_AGEMA_signal_2604, Midori_rounds_SelectedKey_30_}), .b ({new_AGEMA_signal_3393, new_AGEMA_signal_3392, Midori_rounds_SR_Inv_Result[26]}), .c ({new_AGEMA_signal_3491, new_AGEMA_signal_3490, Midori_rounds_mul_ResultXORkey[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U29 ( .a ({new_AGEMA_signal_1845, new_AGEMA_signal_1844, Midori_rounds_SelectedKey_2_}), .b ({new_AGEMA_signal_3411, new_AGEMA_signal_3410, Midori_rounds_SR_Inv_Result[30]}), .c ({new_AGEMA_signal_3493, new_AGEMA_signal_3492, Midori_rounds_mul_ResultXORkey[2]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U27 ( .a ({new_AGEMA_signal_3833, new_AGEMA_signal_3832, Midori_rounds_SR_Inv_Result[24]}), .b ({new_AGEMA_signal_3673, new_AGEMA_signal_3672, Midori_rounds_n6}), .c ({new_AGEMA_signal_3859, new_AGEMA_signal_3858, Midori_rounds_mul_ResultXORkey[28]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U24 ( .a ({new_AGEMA_signal_1865, new_AGEMA_signal_1864, Midori_rounds_SelectedKey_26_}), .b ({new_AGEMA_signal_3399, new_AGEMA_signal_3398, Midori_rounds_SR_Inv_Result[50]}), .c ({new_AGEMA_signal_3499, new_AGEMA_signal_3498, Midori_rounds_mul_ResultXORkey[26]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U22 ( .a ({new_AGEMA_signal_3831, new_AGEMA_signal_3830, Midori_rounds_SR_Inv_Result[48]}), .b ({new_AGEMA_signal_3549, new_AGEMA_signal_3548, Midori_rounds_n5}), .c ({new_AGEMA_signal_3861, new_AGEMA_signal_3860, Midori_rounds_mul_ResultXORkey[24]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U19 ( .a ({new_AGEMA_signal_2591, new_AGEMA_signal_2590, Midori_rounds_SelectedKey_22_}), .b ({new_AGEMA_signal_3381, new_AGEMA_signal_3380, Midori_rounds_SR_Inv_Result[14]}), .c ({new_AGEMA_signal_3505, new_AGEMA_signal_3504, Midori_rounds_mul_ResultXORkey[22]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U17 ( .a ({new_AGEMA_signal_3871, new_AGEMA_signal_3870, Midori_rounds_SR_Inv_Result[12]}), .b ({new_AGEMA_signal_3509, new_AGEMA_signal_3508, Midori_rounds_n4}), .c ({new_AGEMA_signal_3877, new_AGEMA_signal_3876, Midori_rounds_mul_ResultXORkey[20]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U13 ( .a ({new_AGEMA_signal_2583, new_AGEMA_signal_2582, Midori_rounds_SelectedKey_18_}), .b ({new_AGEMA_signal_3387, new_AGEMA_signal_3386, Midori_rounds_SR_Inv_Result[38]}), .c ({new_AGEMA_signal_3515, new_AGEMA_signal_3514, Midori_rounds_mul_ResultXORkey[18]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U11 ( .a ({new_AGEMA_signal_3873, new_AGEMA_signal_3872, Midori_rounds_SR_Inv_Result[36]}), .b ({new_AGEMA_signal_3551, new_AGEMA_signal_3550, Midori_rounds_n3}), .c ({new_AGEMA_signal_3879, new_AGEMA_signal_3878, Midori_rounds_mul_ResultXORkey[16]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U8 ( .a ({new_AGEMA_signal_1861, new_AGEMA_signal_1860, Midori_rounds_SelectedKey_14_}), .b ({new_AGEMA_signal_3417, new_AGEMA_signal_3416, Midori_rounds_SR_Inv_Result[34]}), .c ({new_AGEMA_signal_3521, new_AGEMA_signal_3520, Midori_rounds_mul_ResultXORkey[14]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U6 ( .a ({new_AGEMA_signal_3841, new_AGEMA_signal_3840, Midori_rounds_SR_Inv_Result[32]}), .b ({new_AGEMA_signal_3553, new_AGEMA_signal_3552, Midori_rounds_n2}), .c ({new_AGEMA_signal_3863, new_AGEMA_signal_3862, Midori_rounds_mul_ResultXORkey[12]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U3 ( .a ({new_AGEMA_signal_1855, new_AGEMA_signal_1854, Midori_rounds_SelectedKey_10_}), .b ({new_AGEMA_signal_3423, new_AGEMA_signal_3422, Midori_rounds_SR_Inv_Result[10]}), .c ({new_AGEMA_signal_3527, new_AGEMA_signal_3526, Midori_rounds_mul_ResultXORkey[10]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_U2 ( .a ({new_AGEMA_signal_3843, new_AGEMA_signal_3842, Midori_rounds_SR_Inv_Result[28]}), .b ({new_AGEMA_signal_3555, new_AGEMA_signal_3554, Midori_rounds_n1}), .c ({new_AGEMA_signal_3865, new_AGEMA_signal_3864, Midori_rounds_mul_ResultXORkey[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_0_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3885, new_AGEMA_signal_3884, Midori_rounds_round_Result[0]}), .a ({new_AGEMA_signal_2377, new_AGEMA_signal_2376, Midori_add_Result_Start[0]}), .c ({new_AGEMA_signal_3911, new_AGEMA_signal_3910, Midori_rounds_roundResult_Reg_SFF_0_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_2_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3559, new_AGEMA_signal_3558, Midori_rounds_round_Result[2]}), .a ({new_AGEMA_signal_2289, new_AGEMA_signal_2288, Midori_add_Result_Start[2]}), .c ({new_AGEMA_signal_3677, new_AGEMA_signal_3676, Midori_rounds_roundResult_Reg_SFF_2_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_4_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3887, new_AGEMA_signal_3886, Midori_rounds_round_Result[4]}), .a ({new_AGEMA_signal_2201, new_AGEMA_signal_2200, Midori_add_Result_Start[4]}), .c ({new_AGEMA_signal_3913, new_AGEMA_signal_3912, Midori_rounds_roundResult_Reg_SFF_4_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_6_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3565, new_AGEMA_signal_3564, Midori_rounds_round_Result[6]}), .a ({new_AGEMA_signal_2137, new_AGEMA_signal_2136, Midori_add_Result_Start[6]}), .c ({new_AGEMA_signal_3683, new_AGEMA_signal_3682, Midori_rounds_roundResult_Reg_SFF_6_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_8_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3889, new_AGEMA_signal_3888, Midori_rounds_round_Result[8]}), .a ({new_AGEMA_signal_2129, new_AGEMA_signal_2128, Midori_add_Result_Start[8]}), .c ({new_AGEMA_signal_3915, new_AGEMA_signal_3914, Midori_rounds_roundResult_Reg_SFF_8_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_10_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3571, new_AGEMA_signal_3570, Midori_rounds_round_Result[10]}), .a ({new_AGEMA_signal_2373, new_AGEMA_signal_2372, Midori_add_Result_Start[10]}), .c ({new_AGEMA_signal_3689, new_AGEMA_signal_3688, Midori_rounds_roundResult_Reg_SFF_10_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_12_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3891, new_AGEMA_signal_3890, Midori_rounds_round_Result[12]}), .a ({new_AGEMA_signal_2365, new_AGEMA_signal_2364, Midori_add_Result_Start[12]}), .c ({new_AGEMA_signal_3917, new_AGEMA_signal_3916, Midori_rounds_roundResult_Reg_SFF_12_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_14_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3577, new_AGEMA_signal_3576, Midori_rounds_round_Result[14]}), .a ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, Midori_add_Result_Start[14]}), .c ({new_AGEMA_signal_3695, new_AGEMA_signal_3694, Midori_rounds_roundResult_Reg_SFF_14_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_16_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3933, new_AGEMA_signal_3932, Midori_rounds_round_Result[16]}), .a ({new_AGEMA_signal_2349, new_AGEMA_signal_2348, Midori_add_Result_Start[16]}), .c ({new_AGEMA_signal_3939, new_AGEMA_signal_3938, Midori_rounds_roundResult_Reg_SFF_16_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_18_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3583, new_AGEMA_signal_3582, Midori_rounds_round_Result[18]}), .a ({new_AGEMA_signal_2341, new_AGEMA_signal_2340, Midori_add_Result_Start[18]}), .c ({new_AGEMA_signal_3701, new_AGEMA_signal_3700, Midori_rounds_roundResult_Reg_SFF_18_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_20_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3935, new_AGEMA_signal_3934, Midori_rounds_round_Result[20]}), .a ({new_AGEMA_signal_2329, new_AGEMA_signal_2328, Midori_add_Result_Start[20]}), .c ({new_AGEMA_signal_3941, new_AGEMA_signal_3940, Midori_rounds_roundResult_Reg_SFF_20_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_22_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3589, new_AGEMA_signal_3588, Midori_rounds_round_Result[22]}), .a ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, Midori_add_Result_Start[22]}), .c ({new_AGEMA_signal_3707, new_AGEMA_signal_3706, Midori_rounds_roundResult_Reg_SFF_22_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_24_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3893, new_AGEMA_signal_3892, Midori_rounds_round_Result[24]}), .a ({new_AGEMA_signal_2313, new_AGEMA_signal_2312, Midori_add_Result_Start[24]}), .c ({new_AGEMA_signal_3919, new_AGEMA_signal_3918, Midori_rounds_roundResult_Reg_SFF_24_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_26_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3595, new_AGEMA_signal_3594, Midori_rounds_round_Result[26]}), .a ({new_AGEMA_signal_2305, new_AGEMA_signal_2304, Midori_add_Result_Start[26]}), .c ({new_AGEMA_signal_3713, new_AGEMA_signal_3712, Midori_rounds_roundResult_Reg_SFF_26_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_28_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3895, new_AGEMA_signal_3894, Midori_rounds_round_Result[28]}), .a ({new_AGEMA_signal_2297, new_AGEMA_signal_2296, Midori_add_Result_Start[28]}), .c ({new_AGEMA_signal_3921, new_AGEMA_signal_3920, Midori_rounds_roundResult_Reg_SFF_28_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_30_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3601, new_AGEMA_signal_3600, Midori_rounds_round_Result[30]}), .a ({new_AGEMA_signal_2285, new_AGEMA_signal_2284, Midori_add_Result_Start[30]}), .c ({new_AGEMA_signal_3719, new_AGEMA_signal_3718, Midori_rounds_roundResult_Reg_SFF_30_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_32_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3897, new_AGEMA_signal_3896, Midori_rounds_round_Result[32]}), .a ({new_AGEMA_signal_2277, new_AGEMA_signal_2276, Midori_add_Result_Start[32]}), .c ({new_AGEMA_signal_3923, new_AGEMA_signal_3922, Midori_rounds_roundResult_Reg_SFF_32_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_34_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3607, new_AGEMA_signal_3606, Midori_rounds_round_Result[34]}), .a ({new_AGEMA_signal_2269, new_AGEMA_signal_2268, Midori_add_Result_Start[34]}), .c ({new_AGEMA_signal_3725, new_AGEMA_signal_3724, Midori_rounds_roundResult_Reg_SFF_34_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_36_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3899, new_AGEMA_signal_3898, Midori_rounds_round_Result[36]}), .a ({new_AGEMA_signal_2261, new_AGEMA_signal_2260, Midori_add_Result_Start[36]}), .c ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, Midori_rounds_roundResult_Reg_SFF_36_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_38_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3613, new_AGEMA_signal_3612, Midori_rounds_round_Result[38]}), .a ({new_AGEMA_signal_2253, new_AGEMA_signal_2252, Midori_add_Result_Start[38]}), .c ({new_AGEMA_signal_3731, new_AGEMA_signal_3730, Midori_rounds_roundResult_Reg_SFF_38_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_40_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3901, new_AGEMA_signal_3900, Midori_rounds_round_Result[40]}), .a ({new_AGEMA_signal_2241, new_AGEMA_signal_2240, Midori_add_Result_Start[40]}), .c ({new_AGEMA_signal_3927, new_AGEMA_signal_3926, Midori_rounds_roundResult_Reg_SFF_40_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_42_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3619, new_AGEMA_signal_3618, Midori_rounds_round_Result[42]}), .a ({new_AGEMA_signal_2233, new_AGEMA_signal_2232, Midori_add_Result_Start[42]}), .c ({new_AGEMA_signal_3737, new_AGEMA_signal_3736, Midori_rounds_roundResult_Reg_SFF_42_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_44_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3903, new_AGEMA_signal_3902, Midori_rounds_round_Result[44]}), .a ({new_AGEMA_signal_2225, new_AGEMA_signal_2224, Midori_add_Result_Start[44]}), .c ({new_AGEMA_signal_3929, new_AGEMA_signal_3928, Midori_rounds_roundResult_Reg_SFF_44_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_46_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3625, new_AGEMA_signal_3624, Midori_rounds_round_Result[46]}), .a ({new_AGEMA_signal_2217, new_AGEMA_signal_2216, Midori_add_Result_Start[46]}), .c ({new_AGEMA_signal_3743, new_AGEMA_signal_3742, Midori_rounds_roundResult_Reg_SFF_46_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_48_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3905, new_AGEMA_signal_3904, Midori_rounds_round_Result[48]}), .a ({new_AGEMA_signal_2209, new_AGEMA_signal_2208, Midori_add_Result_Start[48]}), .c ({new_AGEMA_signal_3931, new_AGEMA_signal_3930, Midori_rounds_roundResult_Reg_SFF_48_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_50_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3631, new_AGEMA_signal_3630, Midori_rounds_round_Result[50]}), .a ({new_AGEMA_signal_2197, new_AGEMA_signal_2196, Midori_add_Result_Start[50]}), .c ({new_AGEMA_signal_3749, new_AGEMA_signal_3748, Midori_rounds_roundResult_Reg_SFF_50_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_52_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3937, new_AGEMA_signal_3936, Midori_rounds_round_Result[52]}), .a ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, Midori_add_Result_Start[52]}), .c ({new_AGEMA_signal_3943, new_AGEMA_signal_3942, Midori_rounds_roundResult_Reg_SFF_52_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_54_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3637, new_AGEMA_signal_3636, Midori_rounds_round_Result[54]}), .a ({new_AGEMA_signal_2181, new_AGEMA_signal_2180, Midori_add_Result_Start[54]}), .c ({new_AGEMA_signal_3755, new_AGEMA_signal_3754, Midori_rounds_roundResult_Reg_SFF_54_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_56_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3945, new_AGEMA_signal_3944, Midori_rounds_round_Result[56]}), .a ({new_AGEMA_signal_2173, new_AGEMA_signal_2172, Midori_add_Result_Start[56]}), .c ({new_AGEMA_signal_3949, new_AGEMA_signal_3948, Midori_rounds_roundResult_Reg_SFF_56_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_58_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3643, new_AGEMA_signal_3642, Midori_rounds_round_Result[58]}), .a ({new_AGEMA_signal_2165, new_AGEMA_signal_2164, Midori_add_Result_Start[58]}), .c ({new_AGEMA_signal_3761, new_AGEMA_signal_3760, Midori_rounds_roundResult_Reg_SFF_58_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_60_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3947, new_AGEMA_signal_3946, Midori_rounds_round_Result[60]}), .a ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, Midori_add_Result_Start[60]}), .c ({new_AGEMA_signal_3951, new_AGEMA_signal_3950, Midori_rounds_roundResult_Reg_SFF_60_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_62_MUXInst_U1 ( .s (reset), .b ({new_AGEMA_signal_3649, new_AGEMA_signal_3648, Midori_rounds_round_Result[62]}), .a ({new_AGEMA_signal_2145, new_AGEMA_signal_2144, Midori_add_Result_Start[62]}), .c ({new_AGEMA_signal_3767, new_AGEMA_signal_3766, Midori_rounds_roundResult_Reg_SFF_62_DQ}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U17 ( .a ({new_AGEMA_signal_2381, new_AGEMA_signal_2380, Midori_rounds_sub_sBox_PRINCE_0_n15}), .b ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, Midori_rounds_sub_sBox_PRINCE_0_n12}), .clk (clk), .r ({Fresh[674], Fresh[673], Fresh[672]}), .c ({new_AGEMA_signal_2835, new_AGEMA_signal_2834, Midori_rounds_SR_Result[50]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_0_U8 ( .a ({new_AGEMA_signal_2389, new_AGEMA_signal_2388, Midori_rounds_sub_sBox_PRINCE_0_n13}), .b ({new_AGEMA_signal_2681, new_AGEMA_signal_2680, Midori_rounds_sub_sBox_PRINCE_0_n3}), .clk (clk), .r ({Fresh[677], Fresh[676], Fresh[675]}), .c ({new_AGEMA_signal_2839, new_AGEMA_signal_2838, Midori_rounds_SR_Result[48]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U17 ( .a ({new_AGEMA_signal_2393, new_AGEMA_signal_2392, Midori_rounds_sub_sBox_PRINCE_1_n15}), .b ({new_AGEMA_signal_2687, new_AGEMA_signal_2686, Midori_rounds_sub_sBox_PRINCE_1_n12}), .clk (clk), .r ({Fresh[680], Fresh[679], Fresh[678]}), .c ({new_AGEMA_signal_2843, new_AGEMA_signal_2842, Midori_rounds_SR_Result[46]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_1_U8 ( .a ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, Midori_rounds_sub_sBox_PRINCE_1_n13}), .b ({new_AGEMA_signal_2691, new_AGEMA_signal_2690, Midori_rounds_sub_sBox_PRINCE_1_n3}), .clk (clk), .r ({Fresh[683], Fresh[682], Fresh[681]}), .c ({new_AGEMA_signal_2847, new_AGEMA_signal_2846, Midori_rounds_SR_Result[44]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U17 ( .a ({new_AGEMA_signal_2405, new_AGEMA_signal_2404, Midori_rounds_sub_sBox_PRINCE_2_n15}), .b ({new_AGEMA_signal_2697, new_AGEMA_signal_2696, Midori_rounds_sub_sBox_PRINCE_2_n12}), .clk (clk), .r ({Fresh[686], Fresh[685], Fresh[684]}), .c ({new_AGEMA_signal_2851, new_AGEMA_signal_2850, Midori_rounds_SR_Result[10]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_2_U8 ( .a ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, Midori_rounds_sub_sBox_PRINCE_2_n13}), .b ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, Midori_rounds_sub_sBox_PRINCE_2_n3}), .clk (clk), .r ({Fresh[689], Fresh[688], Fresh[687]}), .c ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, Midori_rounds_SR_Result[8]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U17 ( .a ({new_AGEMA_signal_2417, new_AGEMA_signal_2416, Midori_rounds_sub_sBox_PRINCE_3_n15}), .b ({new_AGEMA_signal_2707, new_AGEMA_signal_2706, Midori_rounds_sub_sBox_PRINCE_3_n12}), .clk (clk), .r ({Fresh[692], Fresh[691], Fresh[690]}), .c ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, Midori_rounds_SR_Result[22]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_3_U8 ( .a ({new_AGEMA_signal_2425, new_AGEMA_signal_2424, Midori_rounds_sub_sBox_PRINCE_3_n13}), .b ({new_AGEMA_signal_2711, new_AGEMA_signal_2710, Midori_rounds_sub_sBox_PRINCE_3_n3}), .clk (clk), .r ({Fresh[695], Fresh[694], Fresh[693]}), .c ({new_AGEMA_signal_2863, new_AGEMA_signal_2862, Midori_rounds_SR_Result[20]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U17 ( .a ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, Midori_rounds_sub_sBox_PRINCE_4_n15}), .b ({new_AGEMA_signal_2717, new_AGEMA_signal_2716, Midori_rounds_sub_sBox_PRINCE_4_n12}), .clk (clk), .r ({Fresh[698], Fresh[697], Fresh[696]}), .c ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, Midori_rounds_SR_Result[38]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_4_U8 ( .a ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, Midori_rounds_sub_sBox_PRINCE_4_n13}), .b ({new_AGEMA_signal_2721, new_AGEMA_signal_2720, Midori_rounds_sub_sBox_PRINCE_4_n3}), .clk (clk), .r ({Fresh[701], Fresh[700], Fresh[699]}), .c ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, Midori_rounds_SR_Result[36]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U17 ( .a ({new_AGEMA_signal_2441, new_AGEMA_signal_2440, Midori_rounds_sub_sBox_PRINCE_5_n15}), .b ({new_AGEMA_signal_2727, new_AGEMA_signal_2726, Midori_rounds_sub_sBox_PRINCE_5_n12}), .clk (clk), .r ({Fresh[704], Fresh[703], Fresh[702]}), .c ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, Midori_rounds_SR_Result[58]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_5_U8 ( .a ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, Midori_rounds_sub_sBox_PRINCE_5_n13}), .b ({new_AGEMA_signal_2731, new_AGEMA_signal_2730, Midori_rounds_sub_sBox_PRINCE_5_n3}), .clk (clk), .r ({Fresh[707], Fresh[706], Fresh[705]}), .c ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, Midori_rounds_SR_Result[56]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U17 ( .a ({new_AGEMA_signal_2453, new_AGEMA_signal_2452, Midori_rounds_sub_sBox_PRINCE_6_n15}), .b ({new_AGEMA_signal_2737, new_AGEMA_signal_2736, Midori_rounds_sub_sBox_PRINCE_6_n12}), .clk (clk), .r ({Fresh[710], Fresh[709], Fresh[708]}), .c ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, Midori_rounds_SR_Result[30]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_6_U8 ( .a ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, Midori_rounds_sub_sBox_PRINCE_6_n13}), .b ({new_AGEMA_signal_2741, new_AGEMA_signal_2740, Midori_rounds_sub_sBox_PRINCE_6_n3}), .clk (clk), .r ({Fresh[713], Fresh[712], Fresh[711]}), .c ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, Midori_rounds_SR_Result[28]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U17 ( .a ({new_AGEMA_signal_2465, new_AGEMA_signal_2464, Midori_rounds_sub_sBox_PRINCE_7_n15}), .b ({new_AGEMA_signal_2747, new_AGEMA_signal_2746, Midori_rounds_sub_sBox_PRINCE_7_n12}), .clk (clk), .r ({Fresh[716], Fresh[715], Fresh[714]}), .c ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, Midori_rounds_SR_Result[2]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_7_U8 ( .a ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, Midori_rounds_sub_sBox_PRINCE_7_n13}), .b ({new_AGEMA_signal_2751, new_AGEMA_signal_2750, Midori_rounds_sub_sBox_PRINCE_7_n3}), .clk (clk), .r ({Fresh[719], Fresh[718], Fresh[717]}), .c ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, Midori_rounds_SR_Result[0]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U17 ( .a ({new_AGEMA_signal_2477, new_AGEMA_signal_2476, Midori_rounds_sub_sBox_PRINCE_8_n15}), .b ({new_AGEMA_signal_2757, new_AGEMA_signal_2756, Midori_rounds_sub_sBox_PRINCE_8_n12}), .clk (clk), .r ({Fresh[722], Fresh[721], Fresh[720]}), .c ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, Midori_rounds_SR_Result[14]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_8_U8 ( .a ({new_AGEMA_signal_2485, new_AGEMA_signal_2484, Midori_rounds_sub_sBox_PRINCE_8_n13}), .b ({new_AGEMA_signal_2761, new_AGEMA_signal_2760, Midori_rounds_sub_sBox_PRINCE_8_n3}), .clk (clk), .r ({Fresh[725], Fresh[724], Fresh[723]}), .c ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, Midori_rounds_SR_Result[12]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U17 ( .a ({new_AGEMA_signal_2489, new_AGEMA_signal_2488, Midori_rounds_sub_sBox_PRINCE_9_n15}), .b ({new_AGEMA_signal_2767, new_AGEMA_signal_2766, Midori_rounds_sub_sBox_PRINCE_9_n12}), .clk (clk), .r ({Fresh[728], Fresh[727], Fresh[726]}), .c ({new_AGEMA_signal_2907, new_AGEMA_signal_2906, Midori_rounds_SR_Result[18]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_9_U8 ( .a ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, Midori_rounds_sub_sBox_PRINCE_9_n13}), .b ({new_AGEMA_signal_2771, new_AGEMA_signal_2770, Midori_rounds_sub_sBox_PRINCE_9_n3}), .clk (clk), .r ({Fresh[731], Fresh[730], Fresh[729]}), .c ({new_AGEMA_signal_2911, new_AGEMA_signal_2910, Midori_rounds_SR_Result[16]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U17 ( .a ({new_AGEMA_signal_2501, new_AGEMA_signal_2500, Midori_rounds_sub_sBox_PRINCE_10_n15}), .b ({new_AGEMA_signal_2777, new_AGEMA_signal_2776, Midori_rounds_sub_sBox_PRINCE_10_n12}), .clk (clk), .r ({Fresh[734], Fresh[733], Fresh[732]}), .c ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, Midori_rounds_SR_Result[54]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_10_U8 ( .a ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, Midori_rounds_sub_sBox_PRINCE_10_n13}), .b ({new_AGEMA_signal_2781, new_AGEMA_signal_2780, Midori_rounds_sub_sBox_PRINCE_10_n3}), .clk (clk), .r ({Fresh[737], Fresh[736], Fresh[735]}), .c ({new_AGEMA_signal_2919, new_AGEMA_signal_2918, Midori_rounds_SR_Result[52]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U17 ( .a ({new_AGEMA_signal_2513, new_AGEMA_signal_2512, Midori_rounds_sub_sBox_PRINCE_11_n15}), .b ({new_AGEMA_signal_2787, new_AGEMA_signal_2786, Midori_rounds_sub_sBox_PRINCE_11_n12}), .clk (clk), .r ({Fresh[740], Fresh[739], Fresh[738]}), .c ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, Midori_rounds_SR_Result[42]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_11_U8 ( .a ({new_AGEMA_signal_2521, new_AGEMA_signal_2520, Midori_rounds_sub_sBox_PRINCE_11_n13}), .b ({new_AGEMA_signal_2791, new_AGEMA_signal_2790, Midori_rounds_sub_sBox_PRINCE_11_n3}), .clk (clk), .r ({Fresh[743], Fresh[742], Fresh[741]}), .c ({new_AGEMA_signal_2927, new_AGEMA_signal_2926, Midori_rounds_SR_Result[40]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U17 ( .a ({new_AGEMA_signal_2525, new_AGEMA_signal_2524, Midori_rounds_sub_sBox_PRINCE_12_n15}), .b ({new_AGEMA_signal_2797, new_AGEMA_signal_2796, Midori_rounds_sub_sBox_PRINCE_12_n12}), .clk (clk), .r ({Fresh[746], Fresh[745], Fresh[744]}), .c ({new_AGEMA_signal_2931, new_AGEMA_signal_2930, Midori_rounds_SR_Result[26]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_12_U8 ( .a ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, Midori_rounds_sub_sBox_PRINCE_12_n13}), .b ({new_AGEMA_signal_2801, new_AGEMA_signal_2800, Midori_rounds_sub_sBox_PRINCE_12_n3}), .clk (clk), .r ({Fresh[749], Fresh[748], Fresh[747]}), .c ({new_AGEMA_signal_2935, new_AGEMA_signal_2934, Midori_rounds_SR_Result[24]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U17 ( .a ({new_AGEMA_signal_2537, new_AGEMA_signal_2536, Midori_rounds_sub_sBox_PRINCE_13_n15}), .b ({new_AGEMA_signal_2807, new_AGEMA_signal_2806, Midori_rounds_sub_sBox_PRINCE_13_n12}), .clk (clk), .r ({Fresh[752], Fresh[751], Fresh[750]}), .c ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, Midori_rounds_SR_Result[6]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_13_U8 ( .a ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, Midori_rounds_sub_sBox_PRINCE_13_n13}), .b ({new_AGEMA_signal_2811, new_AGEMA_signal_2810, Midori_rounds_sub_sBox_PRINCE_13_n3}), .clk (clk), .r ({Fresh[755], Fresh[754], Fresh[753]}), .c ({new_AGEMA_signal_2943, new_AGEMA_signal_2942, Midori_rounds_SR_Result[4]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U17 ( .a ({new_AGEMA_signal_2549, new_AGEMA_signal_2548, Midori_rounds_sub_sBox_PRINCE_14_n15}), .b ({new_AGEMA_signal_2817, new_AGEMA_signal_2816, Midori_rounds_sub_sBox_PRINCE_14_n12}), .clk (clk), .r ({Fresh[758], Fresh[757], Fresh[756]}), .c ({new_AGEMA_signal_2947, new_AGEMA_signal_2946, Midori_rounds_SR_Result[34]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_14_U8 ( .a ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, Midori_rounds_sub_sBox_PRINCE_14_n13}), .b ({new_AGEMA_signal_2821, new_AGEMA_signal_2820, Midori_rounds_sub_sBox_PRINCE_14_n3}), .clk (clk), .r ({Fresh[761], Fresh[760], Fresh[759]}), .c ({new_AGEMA_signal_2951, new_AGEMA_signal_2950, Midori_rounds_SR_Result[32]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U17 ( .a ({new_AGEMA_signal_2561, new_AGEMA_signal_2560, Midori_rounds_sub_sBox_PRINCE_15_n15}), .b ({new_AGEMA_signal_2827, new_AGEMA_signal_2826, Midori_rounds_sub_sBox_PRINCE_15_n12}), .clk (clk), .r ({Fresh[764], Fresh[763], Fresh[762]}), .c ({new_AGEMA_signal_2955, new_AGEMA_signal_2954, Midori_rounds_SR_Result[62]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_sub_sBox_PRINCE_15_U8 ( .a ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, Midori_rounds_sub_sBox_PRINCE_15_n13}), .b ({new_AGEMA_signal_2831, new_AGEMA_signal_2830, Midori_rounds_sub_sBox_PRINCE_15_n3}), .clk (clk), .r ({Fresh[767], Fresh[766], Fresh[765]}), .c ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, Midori_rounds_SR_Result[60]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_0_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, Midori_rounds_SR_Result[0]}), .a ({new_AGEMA_signal_3671, new_AGEMA_signal_3670, Midori_rounds_sub_ResultXORkey[0]}), .c ({new_AGEMA_signal_3783, new_AGEMA_signal_3782, Midori_rounds_mul_input[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_2_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, Midori_rounds_SR_Result[2]}), .a ({new_AGEMA_signal_3151, new_AGEMA_signal_3150, Midori_rounds_sub_ResultXORkey[2]}), .c ({new_AGEMA_signal_3187, new_AGEMA_signal_3186, Midori_rounds_mul_input[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_4_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2943, new_AGEMA_signal_2942, Midori_rounds_SR_Result[4]}), .a ({new_AGEMA_signal_3659, new_AGEMA_signal_3658, Midori_rounds_sub_ResultXORkey[4]}), .c ({new_AGEMA_signal_3785, new_AGEMA_signal_3784, Midori_rounds_mul_input[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_6_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, Midori_rounds_SR_Result[6]}), .a ({new_AGEMA_signal_3093, new_AGEMA_signal_3092, Midori_rounds_sub_ResultXORkey[6]}), .c ({new_AGEMA_signal_3193, new_AGEMA_signal_3192, Midori_rounds_mul_input[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_8_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, Midori_rounds_SR_Result[8]}), .a ({new_AGEMA_signal_3529, new_AGEMA_signal_3528, Midori_rounds_sub_ResultXORkey[8]}), .c ({new_AGEMA_signal_3771, new_AGEMA_signal_3770, Midori_rounds_mul_input[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_10_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2851, new_AGEMA_signal_2850, Midori_rounds_SR_Result[10]}), .a ({new_AGEMA_signal_3183, new_AGEMA_signal_3182, Midori_rounds_sub_ResultXORkey[10]}), .c ({new_AGEMA_signal_3199, new_AGEMA_signal_3198, Midori_rounds_mul_input[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_12_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, Midori_rounds_SR_Result[12]}), .a ({new_AGEMA_signal_3669, new_AGEMA_signal_3668, Midori_rounds_sub_ResultXORkey[12]}), .c ({new_AGEMA_signal_3787, new_AGEMA_signal_3786, Midori_rounds_mul_input[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_14_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, Midori_rounds_SR_Result[14]}), .a ({new_AGEMA_signal_3177, new_AGEMA_signal_3176, Midori_rounds_sub_ResultXORkey[14]}), .c ({new_AGEMA_signal_3205, new_AGEMA_signal_3204, Midori_rounds_mul_input[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_16_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2911, new_AGEMA_signal_2910, Midori_rounds_SR_Result[16]}), .a ({new_AGEMA_signal_3667, new_AGEMA_signal_3666, Midori_rounds_sub_ResultXORkey[16]}), .c ({new_AGEMA_signal_3789, new_AGEMA_signal_3788, Midori_rounds_mul_input[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_18_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2907, new_AGEMA_signal_2906, Midori_rounds_SR_Result[18]}), .a ({new_AGEMA_signal_3171, new_AGEMA_signal_3170, Midori_rounds_sub_ResultXORkey[18]}), .c ({new_AGEMA_signal_3211, new_AGEMA_signal_3210, Midori_rounds_mul_input[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_20_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2863, new_AGEMA_signal_2862, Midori_rounds_SR_Result[20]}), .a ({new_AGEMA_signal_3535, new_AGEMA_signal_3534, Midori_rounds_sub_ResultXORkey[20]}), .c ({new_AGEMA_signal_3773, new_AGEMA_signal_3772, Midori_rounds_mul_input[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_22_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, Midori_rounds_SR_Result[22]}), .a ({new_AGEMA_signal_3163, new_AGEMA_signal_3162, Midori_rounds_sub_ResultXORkey[22]}), .c ({new_AGEMA_signal_3217, new_AGEMA_signal_3216, Midori_rounds_mul_input[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_24_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2935, new_AGEMA_signal_2934, Midori_rounds_SR_Result[24]}), .a ({new_AGEMA_signal_3665, new_AGEMA_signal_3664, Midori_rounds_sub_ResultXORkey[24]}), .c ({new_AGEMA_signal_3791, new_AGEMA_signal_3790, Midori_rounds_mul_input[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_26_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2931, new_AGEMA_signal_2930, Midori_rounds_SR_Result[26]}), .a ({new_AGEMA_signal_3157, new_AGEMA_signal_3156, Midori_rounds_sub_ResultXORkey[26]}), .c ({new_AGEMA_signal_3223, new_AGEMA_signal_3222, Midori_rounds_mul_input[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_28_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, Midori_rounds_SR_Result[28]}), .a ({new_AGEMA_signal_3779, new_AGEMA_signal_3778, Midori_rounds_sub_ResultXORkey[28]}), .c ({new_AGEMA_signal_3805, new_AGEMA_signal_3804, Midori_rounds_mul_input[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_30_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, Midori_rounds_SR_Result[30]}), .a ({new_AGEMA_signal_3149, new_AGEMA_signal_3148, Midori_rounds_sub_ResultXORkey[30]}), .c ({new_AGEMA_signal_3229, new_AGEMA_signal_3228, Midori_rounds_mul_input[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_32_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2951, new_AGEMA_signal_2950, Midori_rounds_SR_Result[32]}), .a ({new_AGEMA_signal_3663, new_AGEMA_signal_3662, Midori_rounds_sub_ResultXORkey[32]}), .c ({new_AGEMA_signal_3793, new_AGEMA_signal_3792, Midori_rounds_mul_input[32]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_34_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2947, new_AGEMA_signal_2946, Midori_rounds_SR_Result[34]}), .a ({new_AGEMA_signal_3143, new_AGEMA_signal_3142, Midori_rounds_sub_ResultXORkey[34]}), .c ({new_AGEMA_signal_3235, new_AGEMA_signal_3234, Midori_rounds_mul_input[34]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_36_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, Midori_rounds_SR_Result[36]}), .a ({new_AGEMA_signal_3533, new_AGEMA_signal_3532, Midori_rounds_sub_ResultXORkey[36]}), .c ({new_AGEMA_signal_3775, new_AGEMA_signal_3774, Midori_rounds_mul_input[36]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_38_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, Midori_rounds_SR_Result[38]}), .a ({new_AGEMA_signal_3137, new_AGEMA_signal_3136, Midori_rounds_sub_ResultXORkey[38]}), .c ({new_AGEMA_signal_3241, new_AGEMA_signal_3240, Midori_rounds_mul_input[38]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_40_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2927, new_AGEMA_signal_2926, Midori_rounds_SR_Result[40]}), .a ({new_AGEMA_signal_3661, new_AGEMA_signal_3660, Midori_rounds_sub_ResultXORkey[40]}), .c ({new_AGEMA_signal_3795, new_AGEMA_signal_3794, Midori_rounds_mul_input[40]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_42_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, Midori_rounds_SR_Result[42]}), .a ({new_AGEMA_signal_3129, new_AGEMA_signal_3128, Midori_rounds_sub_ResultXORkey[42]}), .c ({new_AGEMA_signal_3247, new_AGEMA_signal_3246, Midori_rounds_mul_input[42]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_44_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2847, new_AGEMA_signal_2846, Midori_rounds_SR_Result[44]}), .a ({new_AGEMA_signal_3531, new_AGEMA_signal_3530, Midori_rounds_sub_ResultXORkey[44]}), .c ({new_AGEMA_signal_3777, new_AGEMA_signal_3776, Midori_rounds_mul_input[44]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_46_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2843, new_AGEMA_signal_2842, Midori_rounds_SR_Result[46]}), .a ({new_AGEMA_signal_3123, new_AGEMA_signal_3122, Midori_rounds_sub_ResultXORkey[46]}), .c ({new_AGEMA_signal_3253, new_AGEMA_signal_3252, Midori_rounds_mul_input[46]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_48_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2839, new_AGEMA_signal_2838, Midori_rounds_SR_Result[48]}), .a ({new_AGEMA_signal_3803, new_AGEMA_signal_3802, Midori_rounds_sub_ResultXORkey[48]}), .c ({new_AGEMA_signal_3819, new_AGEMA_signal_3818, Midori_rounds_mul_input[48]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_50_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2835, new_AGEMA_signal_2834, Midori_rounds_SR_Result[50]}), .a ({new_AGEMA_signal_3117, new_AGEMA_signal_3116, Midori_rounds_sub_ResultXORkey[50]}), .c ({new_AGEMA_signal_3259, new_AGEMA_signal_3258, Midori_rounds_mul_input[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_52_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2919, new_AGEMA_signal_2918, Midori_rounds_SR_Result[52]}), .a ({new_AGEMA_signal_3657, new_AGEMA_signal_3656, Midori_rounds_sub_ResultXORkey[52]}), .c ({new_AGEMA_signal_3797, new_AGEMA_signal_3796, Midori_rounds_mul_input[52]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_54_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, Midori_rounds_SR_Result[54]}), .a ({new_AGEMA_signal_3111, new_AGEMA_signal_3110, Midori_rounds_sub_ResultXORkey[54]}), .c ({new_AGEMA_signal_3265, new_AGEMA_signal_3264, Midori_rounds_mul_input[54]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_56_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, Midori_rounds_SR_Result[56]}), .a ({new_AGEMA_signal_3655, new_AGEMA_signal_3654, Midori_rounds_sub_ResultXORkey[56]}), .c ({new_AGEMA_signal_3799, new_AGEMA_signal_3798, Midori_rounds_mul_input[56]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_58_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, Midori_rounds_SR_Result[58]}), .a ({new_AGEMA_signal_3105, new_AGEMA_signal_3104, Midori_rounds_sub_ResultXORkey[58]}), .c ({new_AGEMA_signal_3271, new_AGEMA_signal_3270, Midori_rounds_mul_input[58]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_60_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, Midori_rounds_SR_Result[60]}), .a ({new_AGEMA_signal_3653, new_AGEMA_signal_3652, Midori_rounds_sub_ResultXORkey[60]}), .c ({new_AGEMA_signal_3801, new_AGEMA_signal_3800, Midori_rounds_mul_input[60]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_mul_input_Inst_mux_inst_62_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_2955, new_AGEMA_signal_2954, Midori_rounds_SR_Result[62]}), .a ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, Midori_rounds_sub_ResultXORkey[62]}), .c ({new_AGEMA_signal_3277, new_AGEMA_signal_3276, Midori_rounds_mul_input[62]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC1_U23 ( .a ({new_AGEMA_signal_3801, new_AGEMA_signal_3800, Midori_rounds_mul_input[60]}), .b ({new_AGEMA_signal_3869, new_AGEMA_signal_3868, Midori_rounds_mul_MC1_n7}), .c ({new_AGEMA_signal_3881, new_AGEMA_signal_3880, Midori_rounds_SR_Inv_Result[20]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC1_U21 ( .a ({new_AGEMA_signal_3259, new_AGEMA_signal_3258, Midori_rounds_mul_input[50]}), .b ({new_AGEMA_signal_3283, new_AGEMA_signal_3282, Midori_rounds_mul_MC1_n5}), .c ({new_AGEMA_signal_3333, new_AGEMA_signal_3332, Midori_rounds_SR_Inv_Result[42]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC1_U19 ( .a ({new_AGEMA_signal_3819, new_AGEMA_signal_3818, Midori_rounds_mul_input[48]}), .b ({new_AGEMA_signal_3807, new_AGEMA_signal_3806, Midori_rounds_mul_MC1_n3}), .c ({new_AGEMA_signal_3867, new_AGEMA_signal_3866, Midori_rounds_SR_Inv_Result[40]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC1_U16 ( .a ({new_AGEMA_signal_3265, new_AGEMA_signal_3264, Midori_rounds_mul_input[54]}), .b ({new_AGEMA_signal_3283, new_AGEMA_signal_3282, Midori_rounds_mul_MC1_n5}), .c ({new_AGEMA_signal_3339, new_AGEMA_signal_3338, Midori_rounds_SR_Inv_Result[2]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC1_U15 ( .a ({new_AGEMA_signal_3277, new_AGEMA_signal_3276, Midori_rounds_mul_input[62]}), .b ({new_AGEMA_signal_3271, new_AGEMA_signal_3270, Midori_rounds_mul_input[58]}), .c ({new_AGEMA_signal_3283, new_AGEMA_signal_3282, Midori_rounds_mul_MC1_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC1_U11 ( .a ({new_AGEMA_signal_3271, new_AGEMA_signal_3270, Midori_rounds_mul_input[58]}), .b ({new_AGEMA_signal_3291, new_AGEMA_signal_3290, Midori_rounds_mul_MC1_n1}), .c ({new_AGEMA_signal_3345, new_AGEMA_signal_3344, Midori_rounds_SR_Inv_Result[62]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC1_U8 ( .a ({new_AGEMA_signal_3799, new_AGEMA_signal_3798, Midori_rounds_mul_input[56]}), .b ({new_AGEMA_signal_3869, new_AGEMA_signal_3868, Midori_rounds_mul_MC1_n7}), .c ({new_AGEMA_signal_3883, new_AGEMA_signal_3882, Midori_rounds_SR_Inv_Result[60]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC1_U7 ( .a ({new_AGEMA_signal_3797, new_AGEMA_signal_3796, Midori_rounds_mul_input[52]}), .b ({new_AGEMA_signal_3819, new_AGEMA_signal_3818, Midori_rounds_mul_input[48]}), .c ({new_AGEMA_signal_3869, new_AGEMA_signal_3868, Midori_rounds_mul_MC1_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC1_U4 ( .a ({new_AGEMA_signal_3277, new_AGEMA_signal_3276, Midori_rounds_mul_input[62]}), .b ({new_AGEMA_signal_3291, new_AGEMA_signal_3290, Midori_rounds_mul_MC1_n1}), .c ({new_AGEMA_signal_3351, new_AGEMA_signal_3350, Midori_rounds_SR_Inv_Result[22]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC1_U3 ( .a ({new_AGEMA_signal_3259, new_AGEMA_signal_3258, Midori_rounds_mul_input[50]}), .b ({new_AGEMA_signal_3265, new_AGEMA_signal_3264, Midori_rounds_mul_input[54]}), .c ({new_AGEMA_signal_3291, new_AGEMA_signal_3290, Midori_rounds_mul_MC1_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC1_U2 ( .a ({new_AGEMA_signal_3797, new_AGEMA_signal_3796, Midori_rounds_mul_input[52]}), .b ({new_AGEMA_signal_3807, new_AGEMA_signal_3806, Midori_rounds_mul_MC1_n3}), .c ({new_AGEMA_signal_3821, new_AGEMA_signal_3820, Midori_rounds_SR_Inv_Result[0]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC1_U1 ( .a ({new_AGEMA_signal_3801, new_AGEMA_signal_3800, Midori_rounds_mul_input[60]}), .b ({new_AGEMA_signal_3799, new_AGEMA_signal_3798, Midori_rounds_mul_input[56]}), .c ({new_AGEMA_signal_3807, new_AGEMA_signal_3806, Midori_rounds_mul_MC1_n3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC2_U23 ( .a ({new_AGEMA_signal_3777, new_AGEMA_signal_3776, Midori_rounds_mul_input[44]}), .b ({new_AGEMA_signal_3809, new_AGEMA_signal_3808, Midori_rounds_mul_MC2_n7}), .c ({new_AGEMA_signal_3823, new_AGEMA_signal_3822, Midori_rounds_SR_Inv_Result[44]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC2_U21 ( .a ({new_AGEMA_signal_3235, new_AGEMA_signal_3234, Midori_rounds_mul_input[34]}), .b ({new_AGEMA_signal_3295, new_AGEMA_signal_3294, Midori_rounds_mul_MC2_n5}), .c ({new_AGEMA_signal_3357, new_AGEMA_signal_3356, Midori_rounds_SR_Inv_Result[18]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC2_U19 ( .a ({new_AGEMA_signal_3793, new_AGEMA_signal_3792, Midori_rounds_mul_input[32]}), .b ({new_AGEMA_signal_3811, new_AGEMA_signal_3810, Midori_rounds_mul_MC2_n3}), .c ({new_AGEMA_signal_3825, new_AGEMA_signal_3824, Midori_rounds_SR_Inv_Result[16]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC2_U16 ( .a ({new_AGEMA_signal_3241, new_AGEMA_signal_3240, Midori_rounds_mul_input[38]}), .b ({new_AGEMA_signal_3295, new_AGEMA_signal_3294, Midori_rounds_mul_MC2_n5}), .c ({new_AGEMA_signal_3363, new_AGEMA_signal_3362, Midori_rounds_SR_Inv_Result[58]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC2_U15 ( .a ({new_AGEMA_signal_3253, new_AGEMA_signal_3252, Midori_rounds_mul_input[46]}), .b ({new_AGEMA_signal_3247, new_AGEMA_signal_3246, Midori_rounds_mul_input[42]}), .c ({new_AGEMA_signal_3295, new_AGEMA_signal_3294, Midori_rounds_mul_MC2_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC2_U11 ( .a ({new_AGEMA_signal_3247, new_AGEMA_signal_3246, Midori_rounds_mul_input[42]}), .b ({new_AGEMA_signal_3303, new_AGEMA_signal_3302, Midori_rounds_mul_MC2_n1}), .c ({new_AGEMA_signal_3369, new_AGEMA_signal_3368, Midori_rounds_SR_Inv_Result[6]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC2_U8 ( .a ({new_AGEMA_signal_3795, new_AGEMA_signal_3794, Midori_rounds_mul_input[40]}), .b ({new_AGEMA_signal_3809, new_AGEMA_signal_3808, Midori_rounds_mul_MC2_n7}), .c ({new_AGEMA_signal_3827, new_AGEMA_signal_3826, Midori_rounds_SR_Inv_Result[4]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC2_U7 ( .a ({new_AGEMA_signal_3775, new_AGEMA_signal_3774, Midori_rounds_mul_input[36]}), .b ({new_AGEMA_signal_3793, new_AGEMA_signal_3792, Midori_rounds_mul_input[32]}), .c ({new_AGEMA_signal_3809, new_AGEMA_signal_3808, Midori_rounds_mul_MC2_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC2_U4 ( .a ({new_AGEMA_signal_3253, new_AGEMA_signal_3252, Midori_rounds_mul_input[46]}), .b ({new_AGEMA_signal_3303, new_AGEMA_signal_3302, Midori_rounds_mul_MC2_n1}), .c ({new_AGEMA_signal_3375, new_AGEMA_signal_3374, Midori_rounds_SR_Inv_Result[46]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC2_U3 ( .a ({new_AGEMA_signal_3235, new_AGEMA_signal_3234, Midori_rounds_mul_input[34]}), .b ({new_AGEMA_signal_3241, new_AGEMA_signal_3240, Midori_rounds_mul_input[38]}), .c ({new_AGEMA_signal_3303, new_AGEMA_signal_3302, Midori_rounds_mul_MC2_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC2_U2 ( .a ({new_AGEMA_signal_3775, new_AGEMA_signal_3774, Midori_rounds_mul_input[36]}), .b ({new_AGEMA_signal_3811, new_AGEMA_signal_3810, Midori_rounds_mul_MC2_n3}), .c ({new_AGEMA_signal_3829, new_AGEMA_signal_3828, Midori_rounds_SR_Inv_Result[56]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC2_U1 ( .a ({new_AGEMA_signal_3777, new_AGEMA_signal_3776, Midori_rounds_mul_input[44]}), .b ({new_AGEMA_signal_3795, new_AGEMA_signal_3794, Midori_rounds_mul_input[40]}), .c ({new_AGEMA_signal_3811, new_AGEMA_signal_3810, Midori_rounds_mul_MC2_n3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC3_U23 ( .a ({new_AGEMA_signal_3805, new_AGEMA_signal_3804, Midori_rounds_mul_input[28]}), .b ({new_AGEMA_signal_3813, new_AGEMA_signal_3812, Midori_rounds_mul_MC3_n7}), .c ({new_AGEMA_signal_3831, new_AGEMA_signal_3830, Midori_rounds_SR_Inv_Result[48]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC3_U21 ( .a ({new_AGEMA_signal_3211, new_AGEMA_signal_3210, Midori_rounds_mul_input[18]}), .b ({new_AGEMA_signal_3307, new_AGEMA_signal_3306, Midori_rounds_mul_MC3_n5}), .c ({new_AGEMA_signal_3381, new_AGEMA_signal_3380, Midori_rounds_SR_Inv_Result[14]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC3_U19 ( .a ({new_AGEMA_signal_3789, new_AGEMA_signal_3788, Midori_rounds_mul_input[16]}), .b ({new_AGEMA_signal_3835, new_AGEMA_signal_3834, Midori_rounds_mul_MC3_n3}), .c ({new_AGEMA_signal_3871, new_AGEMA_signal_3870, Midori_rounds_SR_Inv_Result[12]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC3_U16 ( .a ({new_AGEMA_signal_3217, new_AGEMA_signal_3216, Midori_rounds_mul_input[22]}), .b ({new_AGEMA_signal_3307, new_AGEMA_signal_3306, Midori_rounds_mul_MC3_n5}), .c ({new_AGEMA_signal_3387, new_AGEMA_signal_3386, Midori_rounds_SR_Inv_Result[38]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC3_U15 ( .a ({new_AGEMA_signal_3229, new_AGEMA_signal_3228, Midori_rounds_mul_input[30]}), .b ({new_AGEMA_signal_3223, new_AGEMA_signal_3222, Midori_rounds_mul_input[26]}), .c ({new_AGEMA_signal_3307, new_AGEMA_signal_3306, Midori_rounds_mul_MC3_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC3_U11 ( .a ({new_AGEMA_signal_3223, new_AGEMA_signal_3222, Midori_rounds_mul_input[26]}), .b ({new_AGEMA_signal_3315, new_AGEMA_signal_3314, Midori_rounds_mul_MC3_n1}), .c ({new_AGEMA_signal_3393, new_AGEMA_signal_3392, Midori_rounds_SR_Inv_Result[26]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC3_U8 ( .a ({new_AGEMA_signal_3791, new_AGEMA_signal_3790, Midori_rounds_mul_input[24]}), .b ({new_AGEMA_signal_3813, new_AGEMA_signal_3812, Midori_rounds_mul_MC3_n7}), .c ({new_AGEMA_signal_3833, new_AGEMA_signal_3832, Midori_rounds_SR_Inv_Result[24]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC3_U7 ( .a ({new_AGEMA_signal_3773, new_AGEMA_signal_3772, Midori_rounds_mul_input[20]}), .b ({new_AGEMA_signal_3789, new_AGEMA_signal_3788, Midori_rounds_mul_input[16]}), .c ({new_AGEMA_signal_3813, new_AGEMA_signal_3812, Midori_rounds_mul_MC3_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC3_U4 ( .a ({new_AGEMA_signal_3229, new_AGEMA_signal_3228, Midori_rounds_mul_input[30]}), .b ({new_AGEMA_signal_3315, new_AGEMA_signal_3314, Midori_rounds_mul_MC3_n1}), .c ({new_AGEMA_signal_3399, new_AGEMA_signal_3398, Midori_rounds_SR_Inv_Result[50]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC3_U3 ( .a ({new_AGEMA_signal_3211, new_AGEMA_signal_3210, Midori_rounds_mul_input[18]}), .b ({new_AGEMA_signal_3217, new_AGEMA_signal_3216, Midori_rounds_mul_input[22]}), .c ({new_AGEMA_signal_3315, new_AGEMA_signal_3314, Midori_rounds_mul_MC3_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC3_U2 ( .a ({new_AGEMA_signal_3773, new_AGEMA_signal_3772, Midori_rounds_mul_input[20]}), .b ({new_AGEMA_signal_3835, new_AGEMA_signal_3834, Midori_rounds_mul_MC3_n3}), .c ({new_AGEMA_signal_3873, new_AGEMA_signal_3872, Midori_rounds_SR_Inv_Result[36]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC3_U1 ( .a ({new_AGEMA_signal_3805, new_AGEMA_signal_3804, Midori_rounds_mul_input[28]}), .b ({new_AGEMA_signal_3791, new_AGEMA_signal_3790, Midori_rounds_mul_input[24]}), .c ({new_AGEMA_signal_3835, new_AGEMA_signal_3834, Midori_rounds_mul_MC3_n3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC4_U23 ( .a ({new_AGEMA_signal_3787, new_AGEMA_signal_3786, Midori_rounds_mul_input[12]}), .b ({new_AGEMA_signal_3815, new_AGEMA_signal_3814, Midori_rounds_mul_MC4_n7}), .c ({new_AGEMA_signal_3837, new_AGEMA_signal_3836, Midori_rounds_SR_Inv_Result[8]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC4_U21 ( .a ({new_AGEMA_signal_3187, new_AGEMA_signal_3186, Midori_rounds_mul_input[2]}), .b ({new_AGEMA_signal_3319, new_AGEMA_signal_3318, Midori_rounds_mul_MC4_n5}), .c ({new_AGEMA_signal_3405, new_AGEMA_signal_3404, Midori_rounds_SR_Inv_Result[54]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC4_U19 ( .a ({new_AGEMA_signal_3783, new_AGEMA_signal_3782, Midori_rounds_mul_input[0]}), .b ({new_AGEMA_signal_3817, new_AGEMA_signal_3816, Midori_rounds_mul_MC4_n3}), .c ({new_AGEMA_signal_3839, new_AGEMA_signal_3838, Midori_rounds_SR_Inv_Result[52]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC4_U16 ( .a ({new_AGEMA_signal_3193, new_AGEMA_signal_3192, Midori_rounds_mul_input[6]}), .b ({new_AGEMA_signal_3319, new_AGEMA_signal_3318, Midori_rounds_mul_MC4_n5}), .c ({new_AGEMA_signal_3411, new_AGEMA_signal_3410, Midori_rounds_SR_Inv_Result[30]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC4_U15 ( .a ({new_AGEMA_signal_3205, new_AGEMA_signal_3204, Midori_rounds_mul_input[14]}), .b ({new_AGEMA_signal_3199, new_AGEMA_signal_3198, Midori_rounds_mul_input[10]}), .c ({new_AGEMA_signal_3319, new_AGEMA_signal_3318, Midori_rounds_mul_MC4_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC4_U11 ( .a ({new_AGEMA_signal_3199, new_AGEMA_signal_3198, Midori_rounds_mul_input[10]}), .b ({new_AGEMA_signal_3327, new_AGEMA_signal_3326, Midori_rounds_mul_MC4_n1}), .c ({new_AGEMA_signal_3417, new_AGEMA_signal_3416, Midori_rounds_SR_Inv_Result[34]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC4_U8 ( .a ({new_AGEMA_signal_3771, new_AGEMA_signal_3770, Midori_rounds_mul_input[8]}), .b ({new_AGEMA_signal_3815, new_AGEMA_signal_3814, Midori_rounds_mul_MC4_n7}), .c ({new_AGEMA_signal_3841, new_AGEMA_signal_3840, Midori_rounds_SR_Inv_Result[32]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC4_U7 ( .a ({new_AGEMA_signal_3785, new_AGEMA_signal_3784, Midori_rounds_mul_input[4]}), .b ({new_AGEMA_signal_3783, new_AGEMA_signal_3782, Midori_rounds_mul_input[0]}), .c ({new_AGEMA_signal_3815, new_AGEMA_signal_3814, Midori_rounds_mul_MC4_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC4_U4 ( .a ({new_AGEMA_signal_3205, new_AGEMA_signal_3204, Midori_rounds_mul_input[14]}), .b ({new_AGEMA_signal_3327, new_AGEMA_signal_3326, Midori_rounds_mul_MC4_n1}), .c ({new_AGEMA_signal_3423, new_AGEMA_signal_3422, Midori_rounds_SR_Inv_Result[10]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC4_U3 ( .a ({new_AGEMA_signal_3187, new_AGEMA_signal_3186, Midori_rounds_mul_input[2]}), .b ({new_AGEMA_signal_3193, new_AGEMA_signal_3192, Midori_rounds_mul_input[6]}), .c ({new_AGEMA_signal_3327, new_AGEMA_signal_3326, Midori_rounds_mul_MC4_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC4_U2 ( .a ({new_AGEMA_signal_3785, new_AGEMA_signal_3784, Midori_rounds_mul_input[4]}), .b ({new_AGEMA_signal_3817, new_AGEMA_signal_3816, Midori_rounds_mul_MC4_n3}), .c ({new_AGEMA_signal_3843, new_AGEMA_signal_3842, Midori_rounds_SR_Inv_Result[28]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) Midori_rounds_mul_MC4_U1 ( .a ({new_AGEMA_signal_3787, new_AGEMA_signal_3786, Midori_rounds_mul_input[12]}), .b ({new_AGEMA_signal_3771, new_AGEMA_signal_3770, Midori_rounds_mul_input[8]}), .c ({new_AGEMA_signal_3817, new_AGEMA_signal_3816, Midori_rounds_mul_MC4_n3}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_0_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3865, new_AGEMA_signal_3864, Midori_rounds_mul_ResultXORkey[0]}), .a ({new_AGEMA_signal_3821, new_AGEMA_signal_3820, Midori_rounds_SR_Inv_Result[0]}), .c ({new_AGEMA_signal_3885, new_AGEMA_signal_3884, Midori_rounds_round_Result[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_2_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3493, new_AGEMA_signal_3492, Midori_rounds_mul_ResultXORkey[2]}), .a ({new_AGEMA_signal_3339, new_AGEMA_signal_3338, Midori_rounds_SR_Inv_Result[2]}), .c ({new_AGEMA_signal_3559, new_AGEMA_signal_3558, Midori_rounds_round_Result[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_4_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3847, new_AGEMA_signal_3846, Midori_rounds_mul_ResultXORkey[4]}), .a ({new_AGEMA_signal_3827, new_AGEMA_signal_3826, Midori_rounds_SR_Inv_Result[4]}), .c ({new_AGEMA_signal_3887, new_AGEMA_signal_3886, Midori_rounds_round_Result[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_6_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3431, new_AGEMA_signal_3430, Midori_rounds_mul_ResultXORkey[6]}), .a ({new_AGEMA_signal_3369, new_AGEMA_signal_3368, Midori_rounds_SR_Inv_Result[6]}), .c ({new_AGEMA_signal_3565, new_AGEMA_signal_3564, Midori_rounds_round_Result[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_8_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3845, new_AGEMA_signal_3844, Midori_rounds_mul_ResultXORkey[8]}), .a ({new_AGEMA_signal_3837, new_AGEMA_signal_3836, Midori_rounds_SR_Inv_Result[8]}), .c ({new_AGEMA_signal_3889, new_AGEMA_signal_3888, Midori_rounds_round_Result[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_10_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3527, new_AGEMA_signal_3526, Midori_rounds_mul_ResultXORkey[10]}), .a ({new_AGEMA_signal_3423, new_AGEMA_signal_3422, Midori_rounds_SR_Inv_Result[10]}), .c ({new_AGEMA_signal_3571, new_AGEMA_signal_3570, Midori_rounds_round_Result[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_12_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3863, new_AGEMA_signal_3862, Midori_rounds_mul_ResultXORkey[12]}), .a ({new_AGEMA_signal_3871, new_AGEMA_signal_3870, Midori_rounds_SR_Inv_Result[12]}), .c ({new_AGEMA_signal_3891, new_AGEMA_signal_3890, Midori_rounds_round_Result[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_14_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3521, new_AGEMA_signal_3520, Midori_rounds_mul_ResultXORkey[14]}), .a ({new_AGEMA_signal_3381, new_AGEMA_signal_3380, Midori_rounds_SR_Inv_Result[14]}), .c ({new_AGEMA_signal_3577, new_AGEMA_signal_3576, Midori_rounds_round_Result[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_16_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3879, new_AGEMA_signal_3878, Midori_rounds_mul_ResultXORkey[16]}), .a ({new_AGEMA_signal_3825, new_AGEMA_signal_3824, Midori_rounds_SR_Inv_Result[16]}), .c ({new_AGEMA_signal_3933, new_AGEMA_signal_3932, Midori_rounds_round_Result[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_18_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3515, new_AGEMA_signal_3514, Midori_rounds_mul_ResultXORkey[18]}), .a ({new_AGEMA_signal_3357, new_AGEMA_signal_3356, Midori_rounds_SR_Inv_Result[18]}), .c ({new_AGEMA_signal_3583, new_AGEMA_signal_3582, Midori_rounds_round_Result[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_20_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3877, new_AGEMA_signal_3876, Midori_rounds_mul_ResultXORkey[20]}), .a ({new_AGEMA_signal_3881, new_AGEMA_signal_3880, Midori_rounds_SR_Inv_Result[20]}), .c ({new_AGEMA_signal_3935, new_AGEMA_signal_3934, Midori_rounds_round_Result[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_22_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3505, new_AGEMA_signal_3504, Midori_rounds_mul_ResultXORkey[22]}), .a ({new_AGEMA_signal_3351, new_AGEMA_signal_3350, Midori_rounds_SR_Inv_Result[22]}), .c ({new_AGEMA_signal_3589, new_AGEMA_signal_3588, Midori_rounds_round_Result[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_24_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3861, new_AGEMA_signal_3860, Midori_rounds_mul_ResultXORkey[24]}), .a ({new_AGEMA_signal_3833, new_AGEMA_signal_3832, Midori_rounds_SR_Inv_Result[24]}), .c ({new_AGEMA_signal_3893, new_AGEMA_signal_3892, Midori_rounds_round_Result[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_26_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3499, new_AGEMA_signal_3498, Midori_rounds_mul_ResultXORkey[26]}), .a ({new_AGEMA_signal_3393, new_AGEMA_signal_3392, Midori_rounds_SR_Inv_Result[26]}), .c ({new_AGEMA_signal_3595, new_AGEMA_signal_3594, Midori_rounds_round_Result[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_28_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3859, new_AGEMA_signal_3858, Midori_rounds_mul_ResultXORkey[28]}), .a ({new_AGEMA_signal_3843, new_AGEMA_signal_3842, Midori_rounds_SR_Inv_Result[28]}), .c ({new_AGEMA_signal_3895, new_AGEMA_signal_3894, Midori_rounds_round_Result[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_30_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3491, new_AGEMA_signal_3490, Midori_rounds_mul_ResultXORkey[30]}), .a ({new_AGEMA_signal_3411, new_AGEMA_signal_3410, Midori_rounds_SR_Inv_Result[30]}), .c ({new_AGEMA_signal_3601, new_AGEMA_signal_3600, Midori_rounds_round_Result[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_32_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, Midori_rounds_mul_ResultXORkey[32]}), .a ({new_AGEMA_signal_3841, new_AGEMA_signal_3840, Midori_rounds_SR_Inv_Result[32]}), .c ({new_AGEMA_signal_3897, new_AGEMA_signal_3896, Midori_rounds_round_Result[32]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_34_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3485, new_AGEMA_signal_3484, Midori_rounds_mul_ResultXORkey[34]}), .a ({new_AGEMA_signal_3417, new_AGEMA_signal_3416, Midori_rounds_SR_Inv_Result[34]}), .c ({new_AGEMA_signal_3607, new_AGEMA_signal_3606, Midori_rounds_round_Result[34]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_36_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3855, new_AGEMA_signal_3854, Midori_rounds_mul_ResultXORkey[36]}), .a ({new_AGEMA_signal_3873, new_AGEMA_signal_3872, Midori_rounds_SR_Inv_Result[36]}), .c ({new_AGEMA_signal_3899, new_AGEMA_signal_3898, Midori_rounds_round_Result[36]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_38_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3477, new_AGEMA_signal_3476, Midori_rounds_mul_ResultXORkey[38]}), .a ({new_AGEMA_signal_3387, new_AGEMA_signal_3386, Midori_rounds_SR_Inv_Result[38]}), .c ({new_AGEMA_signal_3613, new_AGEMA_signal_3612, Midori_rounds_round_Result[38]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_40_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3853, new_AGEMA_signal_3852, Midori_rounds_mul_ResultXORkey[40]}), .a ({new_AGEMA_signal_3867, new_AGEMA_signal_3866, Midori_rounds_SR_Inv_Result[40]}), .c ({new_AGEMA_signal_3901, new_AGEMA_signal_3900, Midori_rounds_round_Result[40]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_42_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3469, new_AGEMA_signal_3468, Midori_rounds_mul_ResultXORkey[42]}), .a ({new_AGEMA_signal_3333, new_AGEMA_signal_3332, Midori_rounds_SR_Inv_Result[42]}), .c ({new_AGEMA_signal_3619, new_AGEMA_signal_3618, Midori_rounds_round_Result[42]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_44_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3851, new_AGEMA_signal_3850, Midori_rounds_mul_ResultXORkey[44]}), .a ({new_AGEMA_signal_3823, new_AGEMA_signal_3822, Midori_rounds_SR_Inv_Result[44]}), .c ({new_AGEMA_signal_3903, new_AGEMA_signal_3902, Midori_rounds_round_Result[44]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_46_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3461, new_AGEMA_signal_3460, Midori_rounds_mul_ResultXORkey[46]}), .a ({new_AGEMA_signal_3375, new_AGEMA_signal_3374, Midori_rounds_SR_Inv_Result[46]}), .c ({new_AGEMA_signal_3625, new_AGEMA_signal_3624, Midori_rounds_round_Result[46]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_48_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3849, new_AGEMA_signal_3848, Midori_rounds_mul_ResultXORkey[48]}), .a ({new_AGEMA_signal_3831, new_AGEMA_signal_3830, Midori_rounds_SR_Inv_Result[48]}), .c ({new_AGEMA_signal_3905, new_AGEMA_signal_3904, Midori_rounds_round_Result[48]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_50_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3455, new_AGEMA_signal_3454, Midori_rounds_mul_ResultXORkey[50]}), .a ({new_AGEMA_signal_3399, new_AGEMA_signal_3398, Midori_rounds_SR_Inv_Result[50]}), .c ({new_AGEMA_signal_3631, new_AGEMA_signal_3630, Midori_rounds_round_Result[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_52_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3875, new_AGEMA_signal_3874, Midori_rounds_mul_ResultXORkey[52]}), .a ({new_AGEMA_signal_3839, new_AGEMA_signal_3838, Midori_rounds_SR_Inv_Result[52]}), .c ({new_AGEMA_signal_3937, new_AGEMA_signal_3936, Midori_rounds_round_Result[52]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_54_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3449, new_AGEMA_signal_3448, Midori_rounds_mul_ResultXORkey[54]}), .a ({new_AGEMA_signal_3405, new_AGEMA_signal_3404, Midori_rounds_SR_Inv_Result[54]}), .c ({new_AGEMA_signal_3637, new_AGEMA_signal_3636, Midori_rounds_round_Result[54]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_56_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3909, new_AGEMA_signal_3908, Midori_rounds_mul_ResultXORkey[56]}), .a ({new_AGEMA_signal_3829, new_AGEMA_signal_3828, Midori_rounds_SR_Inv_Result[56]}), .c ({new_AGEMA_signal_3945, new_AGEMA_signal_3944, Midori_rounds_round_Result[56]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_58_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3443, new_AGEMA_signal_3442, Midori_rounds_mul_ResultXORkey[58]}), .a ({new_AGEMA_signal_3363, new_AGEMA_signal_3362, Midori_rounds_SR_Inv_Result[58]}), .c ({new_AGEMA_signal_3643, new_AGEMA_signal_3642, Midori_rounds_round_Result[58]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_60_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3907, new_AGEMA_signal_3906, Midori_rounds_mul_ResultXORkey[60]}), .a ({new_AGEMA_signal_3883, new_AGEMA_signal_3882, Midori_rounds_SR_Inv_Result[60]}), .c ({new_AGEMA_signal_3947, new_AGEMA_signal_3946, Midori_rounds_round_Result[60]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) Midori_rounds_Res_Inst_mux_inst_62_U1 ( .s (enc_dec), .b ({new_AGEMA_signal_3435, new_AGEMA_signal_3434, Midori_rounds_mul_ResultXORkey[62]}), .a ({new_AGEMA_signal_3345, new_AGEMA_signal_3344, Midori_rounds_SR_Inv_Result[62]}), .c ({new_AGEMA_signal_3649, new_AGEMA_signal_3648, Midori_rounds_round_Result[62]}) ) ;

    /* register cells */
    DFF_X1 controller_roundCounter_count_reg_0__FF_FF ( .CK (clk_gated), .D (controller_roundCounter_N7), .Q (round_Signal[0]), .QN () ) ;
    DFF_X1 controller_roundCounter_count_reg_1__FF_FF ( .CK (clk_gated), .D (controller_roundCounter_N8), .Q (round_Signal[1]), .QN () ) ;
    DFF_X1 controller_roundCounter_count_reg_2__FF_FF ( .CK (clk_gated), .D (controller_roundCounter_n2), .Q (round_Signal[2]), .QN () ) ;
    DFF_X1 controller_roundCounter_count_reg_3__FF_FF ( .CK (clk_gated), .D (controller_roundCounter_N10), .Q (round_Signal[3]), .QN () ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3911, new_AGEMA_signal_3910, Midori_rounds_roundResult_Reg_SFF_0_DQ}), .Q ({new_AGEMA_signal_1867, new_AGEMA_signal_1866, Midori_rounds_roundReg_out[0]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3675, new_AGEMA_signal_3674, Midori_rounds_roundResult_Reg_SFF_1_DQ}), .Q ({new_AGEMA_signal_2673, new_AGEMA_signal_2672, Midori_rounds_roundReg_out[1]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3677, new_AGEMA_signal_3676, Midori_rounds_roundResult_Reg_SFF_2_DQ}), .Q ({new_AGEMA_signal_1873, new_AGEMA_signal_1872, Midori_rounds_roundReg_out[2]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3679, new_AGEMA_signal_3678, Midori_rounds_roundResult_Reg_SFF_3_DQ}), .Q ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, Midori_rounds_roundReg_out[3]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3913, new_AGEMA_signal_3912, Midori_rounds_roundResult_Reg_SFF_4_DQ}), .Q ({new_AGEMA_signal_1883, new_AGEMA_signal_1882, Midori_rounds_roundReg_out[4]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3681, new_AGEMA_signal_3680, Midori_rounds_roundResult_Reg_SFF_5_DQ}), .Q ({new_AGEMA_signal_2683, new_AGEMA_signal_2682, Midori_rounds_roundReg_out[5]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3683, new_AGEMA_signal_3682, Midori_rounds_roundResult_Reg_SFF_6_DQ}), .Q ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, Midori_rounds_roundReg_out[6]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3685, new_AGEMA_signal_3684, Midori_rounds_roundResult_Reg_SFF_7_DQ}), .Q ({new_AGEMA_signal_1885, new_AGEMA_signal_1884, Midori_rounds_roundReg_out[7]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_8_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3915, new_AGEMA_signal_3914, Midori_rounds_roundResult_Reg_SFF_8_DQ}), .Q ({new_AGEMA_signal_1899, new_AGEMA_signal_1898, Midori_rounds_roundReg_out[8]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_9_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3687, new_AGEMA_signal_3686, Midori_rounds_roundResult_Reg_SFF_9_DQ}), .Q ({new_AGEMA_signal_2693, new_AGEMA_signal_2692, Midori_rounds_roundReg_out[9]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_10_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3689, new_AGEMA_signal_3688, Midori_rounds_roundResult_Reg_SFF_10_DQ}), .Q ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, Midori_rounds_roundReg_out[10]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_11_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3691, new_AGEMA_signal_3690, Midori_rounds_roundResult_Reg_SFF_11_DQ}), .Q ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, Midori_rounds_roundReg_out[11]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_12_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3917, new_AGEMA_signal_3916, Midori_rounds_roundResult_Reg_SFF_12_DQ}), .Q ({new_AGEMA_signal_1915, new_AGEMA_signal_1914, Midori_rounds_roundReg_out[12]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_13_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3693, new_AGEMA_signal_3692, Midori_rounds_roundResult_Reg_SFF_13_DQ}), .Q ({new_AGEMA_signal_2703, new_AGEMA_signal_2702, Midori_rounds_roundReg_out[13]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_14_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3695, new_AGEMA_signal_3694, Midori_rounds_roundResult_Reg_SFF_14_DQ}), .Q ({new_AGEMA_signal_1921, new_AGEMA_signal_1920, Midori_rounds_roundReg_out[14]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_15_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3697, new_AGEMA_signal_3696, Midori_rounds_roundResult_Reg_SFF_15_DQ}), .Q ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, Midori_rounds_roundReg_out[15]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_16_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3939, new_AGEMA_signal_3938, Midori_rounds_roundResult_Reg_SFF_16_DQ}), .Q ({new_AGEMA_signal_1931, new_AGEMA_signal_1930, Midori_rounds_roundReg_out[16]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_17_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3699, new_AGEMA_signal_3698, Midori_rounds_roundResult_Reg_SFF_17_DQ}), .Q ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, Midori_rounds_roundReg_out[17]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_18_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3701, new_AGEMA_signal_3700, Midori_rounds_roundResult_Reg_SFF_18_DQ}), .Q ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, Midori_rounds_roundReg_out[18]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_19_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3703, new_AGEMA_signal_3702, Midori_rounds_roundResult_Reg_SFF_19_DQ}), .Q ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, Midori_rounds_roundReg_out[19]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_20_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3941, new_AGEMA_signal_3940, Midori_rounds_roundResult_Reg_SFF_20_DQ}), .Q ({new_AGEMA_signal_1947, new_AGEMA_signal_1946, Midori_rounds_roundReg_out[20]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_21_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3705, new_AGEMA_signal_3704, Midori_rounds_roundResult_Reg_SFF_21_DQ}), .Q ({new_AGEMA_signal_2723, new_AGEMA_signal_2722, Midori_rounds_roundReg_out[21]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_22_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3707, new_AGEMA_signal_3706, Midori_rounds_roundResult_Reg_SFF_22_DQ}), .Q ({new_AGEMA_signal_1953, new_AGEMA_signal_1952, Midori_rounds_roundReg_out[22]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_23_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3709, new_AGEMA_signal_3708, Midori_rounds_roundResult_Reg_SFF_23_DQ}), .Q ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, Midori_rounds_roundReg_out[23]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_24_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3919, new_AGEMA_signal_3918, Midori_rounds_roundResult_Reg_SFF_24_DQ}), .Q ({new_AGEMA_signal_1963, new_AGEMA_signal_1962, Midori_rounds_roundReg_out[24]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_25_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3711, new_AGEMA_signal_3710, Midori_rounds_roundResult_Reg_SFF_25_DQ}), .Q ({new_AGEMA_signal_2733, new_AGEMA_signal_2732, Midori_rounds_roundReg_out[25]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_26_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3713, new_AGEMA_signal_3712, Midori_rounds_roundResult_Reg_SFF_26_DQ}), .Q ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, Midori_rounds_roundReg_out[26]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_27_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3715, new_AGEMA_signal_3714, Midori_rounds_roundResult_Reg_SFF_27_DQ}), .Q ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, Midori_rounds_roundReg_out[27]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_28_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3921, new_AGEMA_signal_3920, Midori_rounds_roundResult_Reg_SFF_28_DQ}), .Q ({new_AGEMA_signal_1979, new_AGEMA_signal_1978, Midori_rounds_roundReg_out[28]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_29_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3717, new_AGEMA_signal_3716, Midori_rounds_roundResult_Reg_SFF_29_DQ}), .Q ({new_AGEMA_signal_2743, new_AGEMA_signal_2742, Midori_rounds_roundReg_out[29]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_30_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3719, new_AGEMA_signal_3718, Midori_rounds_roundResult_Reg_SFF_30_DQ}), .Q ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, Midori_rounds_roundReg_out[30]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_31_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3721, new_AGEMA_signal_3720, Midori_rounds_roundResult_Reg_SFF_31_DQ}), .Q ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, Midori_rounds_roundReg_out[31]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_32_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3923, new_AGEMA_signal_3922, Midori_rounds_roundResult_Reg_SFF_32_DQ}), .Q ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, Midori_rounds_roundReg_out[32]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_33_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3723, new_AGEMA_signal_3722, Midori_rounds_roundResult_Reg_SFF_33_DQ}), .Q ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, Midori_rounds_roundReg_out[33]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_34_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3725, new_AGEMA_signal_3724, Midori_rounds_roundResult_Reg_SFF_34_DQ}), .Q ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, Midori_rounds_roundReg_out[34]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_35_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3727, new_AGEMA_signal_3726, Midori_rounds_roundResult_Reg_SFF_35_DQ}), .Q ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, Midori_rounds_roundReg_out[35]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_36_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, Midori_rounds_roundResult_Reg_SFF_36_DQ}), .Q ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, Midori_rounds_roundReg_out[36]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_37_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3729, new_AGEMA_signal_3728, Midori_rounds_roundResult_Reg_SFF_37_DQ}), .Q ({new_AGEMA_signal_2763, new_AGEMA_signal_2762, Midori_rounds_roundReg_out[37]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_38_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3731, new_AGEMA_signal_3730, Midori_rounds_roundResult_Reg_SFF_38_DQ}), .Q ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, Midori_rounds_roundReg_out[38]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_39_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3733, new_AGEMA_signal_3732, Midori_rounds_roundResult_Reg_SFF_39_DQ}), .Q ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, Midori_rounds_roundReg_out[39]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_40_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3927, new_AGEMA_signal_3926, Midori_rounds_roundResult_Reg_SFF_40_DQ}), .Q ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, Midori_rounds_roundReg_out[40]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_41_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3735, new_AGEMA_signal_3734, Midori_rounds_roundResult_Reg_SFF_41_DQ}), .Q ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, Midori_rounds_roundReg_out[41]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_42_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3737, new_AGEMA_signal_3736, Midori_rounds_roundResult_Reg_SFF_42_DQ}), .Q ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, Midori_rounds_roundReg_out[42]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_43_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3739, new_AGEMA_signal_3738, Midori_rounds_roundResult_Reg_SFF_43_DQ}), .Q ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, Midori_rounds_roundReg_out[43]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_44_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3929, new_AGEMA_signal_3928, Midori_rounds_roundResult_Reg_SFF_44_DQ}), .Q ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, Midori_rounds_roundReg_out[44]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_45_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3741, new_AGEMA_signal_3740, Midori_rounds_roundResult_Reg_SFF_45_DQ}), .Q ({new_AGEMA_signal_2783, new_AGEMA_signal_2782, Midori_rounds_roundReg_out[45]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_46_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3743, new_AGEMA_signal_3742, Midori_rounds_roundResult_Reg_SFF_46_DQ}), .Q ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, Midori_rounds_roundReg_out[46]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_47_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3745, new_AGEMA_signal_3744, Midori_rounds_roundResult_Reg_SFF_47_DQ}), .Q ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, Midori_rounds_roundReg_out[47]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_48_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3931, new_AGEMA_signal_3930, Midori_rounds_roundResult_Reg_SFF_48_DQ}), .Q ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, Midori_rounds_roundReg_out[48]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_49_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3747, new_AGEMA_signal_3746, Midori_rounds_roundResult_Reg_SFF_49_DQ}), .Q ({new_AGEMA_signal_2793, new_AGEMA_signal_2792, Midori_rounds_roundReg_out[49]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_50_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3749, new_AGEMA_signal_3748, Midori_rounds_roundResult_Reg_SFF_50_DQ}), .Q ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, Midori_rounds_roundReg_out[50]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_51_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3751, new_AGEMA_signal_3750, Midori_rounds_roundResult_Reg_SFF_51_DQ}), .Q ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, Midori_rounds_roundReg_out[51]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_52_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3943, new_AGEMA_signal_3942, Midori_rounds_roundResult_Reg_SFF_52_DQ}), .Q ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, Midori_rounds_roundReg_out[52]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_53_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3753, new_AGEMA_signal_3752, Midori_rounds_roundResult_Reg_SFF_53_DQ}), .Q ({new_AGEMA_signal_2803, new_AGEMA_signal_2802, Midori_rounds_roundReg_out[53]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_54_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3755, new_AGEMA_signal_3754, Midori_rounds_roundResult_Reg_SFF_54_DQ}), .Q ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, Midori_rounds_roundReg_out[54]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_55_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3757, new_AGEMA_signal_3756, Midori_rounds_roundResult_Reg_SFF_55_DQ}), .Q ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, Midori_rounds_roundReg_out[55]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_56_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3949, new_AGEMA_signal_3948, Midori_rounds_roundResult_Reg_SFF_56_DQ}), .Q ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, Midori_rounds_roundReg_out[56]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_57_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3759, new_AGEMA_signal_3758, Midori_rounds_roundResult_Reg_SFF_57_DQ}), .Q ({new_AGEMA_signal_2813, new_AGEMA_signal_2812, Midori_rounds_roundReg_out[57]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_58_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3761, new_AGEMA_signal_3760, Midori_rounds_roundResult_Reg_SFF_58_DQ}), .Q ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, Midori_rounds_roundReg_out[58]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_59_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3763, new_AGEMA_signal_3762, Midori_rounds_roundResult_Reg_SFF_59_DQ}), .Q ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, Midori_rounds_roundReg_out[59]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_60_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3951, new_AGEMA_signal_3950, Midori_rounds_roundResult_Reg_SFF_60_DQ}), .Q ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, Midori_rounds_roundReg_out[60]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_61_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3765, new_AGEMA_signal_3764, Midori_rounds_roundResult_Reg_SFF_61_DQ}), .Q ({new_AGEMA_signal_2823, new_AGEMA_signal_2822, Midori_rounds_roundReg_out[61]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_62_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3767, new_AGEMA_signal_3766, Midori_rounds_roundResult_Reg_SFF_62_DQ}), .Q ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, Midori_rounds_roundReg_out[62]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Midori_rounds_roundResult_Reg_SFF_63_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3769, new_AGEMA_signal_3768, Midori_rounds_roundResult_Reg_SFF_63_DQ}), .Q ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, Midori_rounds_roundReg_out[63]}) ) ;
endmodule
