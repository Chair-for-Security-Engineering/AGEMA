/* modified netlist. Source: module LED in file /LED_round-based/AGEMA/LED.v */
/* 4 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 5 register stage(s) in total */

module LED_HPC2_AIG_Pipeline_d1 (IN_plaintext_s0, IN_key_s0, IN_reset, CLK, IN_key_s1, IN_plaintext_s1, Fresh, OUT_ciphertext_s0, OUT_done, OUT_ciphertext_s1);
    input [63:0] IN_plaintext_s0 ;
    input [127:0] IN_key_s0 ;
    input IN_reset ;
    input CLK ;
    input [127:0] IN_key_s1 ;
    input [63:0] IN_plaintext_s1 ;
    input [63:0] Fresh ;
    output [63:0] OUT_ciphertext_s0 ;
    output OUT_done ;
    output [63:0] OUT_ciphertext_s1 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_285 ;
    wire signal_286 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_295 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_356 ;
    wire signal_375 ;
    wire signal_394 ;
    wire signal_413 ;
    wire signal_432 ;
    wire signal_451 ;
    wire signal_470 ;
    wire signal_489 ;
    wire signal_508 ;
    wire signal_527 ;
    wire signal_546 ;
    wire signal_565 ;
    wire signal_584 ;
    wire signal_603 ;
    wire signal_622 ;
    wire signal_641 ;
    wire signal_656 ;
    wire signal_657 ;
    wire signal_658 ;
    wire signal_659 ;
    wire signal_660 ;
    wire signal_661 ;
    wire signal_662 ;
    wire signal_663 ;
    wire signal_664 ;
    wire signal_665 ;
    wire signal_666 ;
    wire signal_667 ;
    wire signal_668 ;
    wire signal_669 ;
    wire signal_670 ;
    wire signal_671 ;
    wire signal_672 ;
    wire signal_673 ;
    wire signal_674 ;
    wire signal_675 ;
    wire signal_676 ;
    wire signal_677 ;
    wire signal_678 ;
    wire signal_679 ;
    wire signal_680 ;
    wire signal_681 ;
    wire signal_682 ;
    wire signal_683 ;
    wire signal_684 ;
    wire signal_685 ;
    wire signal_686 ;
    wire signal_687 ;
    wire signal_688 ;
    wire signal_689 ;
    wire signal_690 ;
    wire signal_691 ;
    wire signal_692 ;
    wire signal_693 ;
    wire signal_694 ;
    wire signal_695 ;
    wire signal_696 ;
    wire signal_697 ;
    wire signal_698 ;
    wire signal_699 ;
    wire signal_700 ;
    wire signal_701 ;
    wire signal_702 ;
    wire signal_703 ;
    wire signal_704 ;
    wire signal_705 ;
    wire signal_706 ;
    wire signal_707 ;
    wire signal_708 ;
    wire signal_709 ;
    wire signal_710 ;
    wire signal_711 ;
    wire signal_712 ;
    wire signal_713 ;
    wire signal_714 ;
    wire signal_715 ;
    wire signal_716 ;
    wire signal_717 ;
    wire signal_718 ;
    wire signal_719 ;
    wire signal_720 ;
    wire signal_721 ;
    wire signal_722 ;
    wire signal_723 ;
    wire signal_724 ;
    wire signal_725 ;
    wire signal_726 ;
    wire signal_727 ;
    wire signal_728 ;
    wire signal_729 ;
    wire signal_730 ;
    wire signal_731 ;
    wire signal_732 ;
    wire signal_733 ;
    wire signal_734 ;
    wire signal_735 ;
    wire signal_736 ;
    wire signal_737 ;
    wire signal_738 ;
    wire signal_739 ;
    wire signal_740 ;
    wire signal_741 ;
    wire signal_742 ;
    wire signal_743 ;
    wire signal_744 ;
    wire signal_745 ;
    wire signal_746 ;
    wire signal_747 ;
    wire signal_748 ;
    wire signal_749 ;
    wire signal_750 ;
    wire signal_751 ;
    wire signal_752 ;
    wire signal_753 ;
    wire signal_754 ;
    wire signal_755 ;
    wire signal_756 ;
    wire signal_757 ;
    wire signal_758 ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_768 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_771 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_774 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_777 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_780 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_783 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_786 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_789 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_792 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_879 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_885 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_888 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_891 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_894 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_897 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_900 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_903 ;
    wire signal_904 ;
    wire signal_905 ;
    wire signal_906 ;
    wire signal_907 ;
    wire signal_908 ;
    wire signal_909 ;
    wire signal_910 ;
    wire signal_911 ;
    wire signal_912 ;
    wire signal_914 ;
    wire signal_915 ;
    wire signal_916 ;
    wire signal_918 ;
    wire signal_919 ;
    wire signal_920 ;
    wire signal_922 ;
    wire signal_923 ;
    wire signal_924 ;
    wire signal_926 ;
    wire signal_927 ;
    wire signal_928 ;
    wire signal_929 ;
    wire signal_930 ;
    wire signal_932 ;
    wire signal_933 ;
    wire signal_934 ;
    wire signal_936 ;
    wire signal_937 ;
    wire signal_938 ;
    wire signal_940 ;
    wire signal_941 ;
    wire signal_942 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1020 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1023 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1276 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1279 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1282 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1285 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1288 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1294 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1297 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1300 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1303 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1309 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1494 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1499 ;
    wire signal_1500 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1503 ;
    wire signal_1504 ;
    wire signal_1505 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1509 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1512 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1518 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1521 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1527 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1530 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1536 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1539 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1564 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1623 ;
    wire signal_1624 ;
    wire signal_1625 ;
    wire signal_1626 ;
    wire signal_1627 ;
    wire signal_1628 ;
    wire signal_1629 ;
    wire signal_1630 ;
    wire signal_1631 ;
    wire signal_1632 ;
    wire signal_1633 ;
    wire signal_1634 ;
    wire signal_1635 ;
    wire signal_1636 ;
    wire signal_1637 ;
    wire signal_1638 ;
    wire signal_1639 ;
    wire signal_1640 ;
    wire signal_1641 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1658 ;
    wire signal_1661 ;
    wire signal_1664 ;
    wire signal_1667 ;
    wire signal_1670 ;
    wire signal_1673 ;
    wire signal_1676 ;
    wire signal_1679 ;
    wire signal_1682 ;
    wire signal_1685 ;
    wire signal_1688 ;
    wire signal_1691 ;
    wire signal_1694 ;
    wire signal_1696 ;
    wire signal_1698 ;
    wire signal_1700 ;
    wire signal_1702 ;
    wire signal_1704 ;
    wire signal_1706 ;
    wire signal_1708 ;
    wire signal_1710 ;
    wire signal_1712 ;
    wire signal_1714 ;
    wire signal_1716 ;
    wire signal_1718 ;
    wire signal_1720 ;
    wire signal_1723 ;
    wire signal_1726 ;
    wire signal_1729 ;
    wire signal_1732 ;
    wire signal_1735 ;
    wire signal_1738 ;
    wire signal_1741 ;
    wire signal_1744 ;
    wire signal_1747 ;
    wire signal_1750 ;
    wire signal_1753 ;
    wire signal_1756 ;
    wire signal_1759 ;
    wire signal_1762 ;
    wire signal_1765 ;
    wire signal_1768 ;
    wire signal_1771 ;
    wire signal_1774 ;
    wire signal_1777 ;
    wire signal_1780 ;
    wire signal_1783 ;
    wire signal_1786 ;
    wire signal_1789 ;
    wire signal_1792 ;
    wire signal_1795 ;
    wire signal_1798 ;
    wire signal_1801 ;
    wire signal_1804 ;
    wire signal_1807 ;
    wire signal_1810 ;
    wire signal_1813 ;
    wire signal_1816 ;
    wire signal_1819 ;
    wire signal_1822 ;
    wire signal_1825 ;
    wire signal_1828 ;
    wire signal_1831 ;
    wire signal_1834 ;
    wire signal_1837 ;
    wire signal_1840 ;
    wire signal_1843 ;
    wire signal_1846 ;
    wire signal_1849 ;
    wire signal_1852 ;
    wire signal_1855 ;
    wire signal_1858 ;
    wire signal_1861 ;
    wire signal_1864 ;
    wire signal_1867 ;
    wire signal_1870 ;
    wire signal_1873 ;
    wire signal_1874 ;
    wire signal_1875 ;
    wire signal_1876 ;
    wire signal_1877 ;
    wire signal_1878 ;
    wire signal_1879 ;
    wire signal_1880 ;
    wire signal_1882 ;
    wire signal_1884 ;
    wire signal_1886 ;
    wire signal_1888 ;
    wire signal_1890 ;
    wire signal_1892 ;
    wire signal_1894 ;
    wire signal_1896 ;
    wire signal_1898 ;
    wire signal_1900 ;
    wire signal_1902 ;
    wire signal_1904 ;
    wire signal_1906 ;
    wire signal_1908 ;
    wire signal_1910 ;
    wire signal_1912 ;
    wire signal_1914 ;
    wire signal_1916 ;
    wire signal_1918 ;
    wire signal_1920 ;
    wire signal_1922 ;
    wire signal_1924 ;
    wire signal_1926 ;
    wire signal_1928 ;
    wire signal_1930 ;
    wire signal_1932 ;
    wire signal_1934 ;
    wire signal_1936 ;
    wire signal_1938 ;
    wire signal_1940 ;
    wire signal_1942 ;
    wire signal_1944 ;
    wire signal_1946 ;
    wire signal_1948 ;
    wire signal_1950 ;
    wire signal_1952 ;
    wire signal_1954 ;
    wire signal_1956 ;
    wire signal_1958 ;
    wire signal_1960 ;
    wire signal_1962 ;
    wire signal_1964 ;
    wire signal_1966 ;
    wire signal_1968 ;
    wire signal_1970 ;
    wire signal_1972 ;
    wire signal_1974 ;
    wire signal_1976 ;
    wire signal_1978 ;
    wire signal_1980 ;
    wire signal_1982 ;
    wire signal_1983 ;
    wire signal_1984 ;
    wire signal_1985 ;
    wire signal_1986 ;
    wire signal_1987 ;
    wire signal_1988 ;
    wire signal_1989 ;
    wire signal_1990 ;
    wire signal_1991 ;
    wire signal_1992 ;
    wire signal_1993 ;
    wire signal_1994 ;
    wire signal_1995 ;
    wire signal_1996 ;
    wire signal_1997 ;
    wire signal_1998 ;
    wire signal_1999 ;
    wire signal_2000 ;
    wire signal_2001 ;
    wire signal_2002 ;
    wire signal_2003 ;
    wire signal_2004 ;
    wire signal_2005 ;
    wire signal_2006 ;
    wire signal_2007 ;
    wire signal_2008 ;
    wire signal_2009 ;
    wire signal_2010 ;
    wire signal_2011 ;
    wire signal_2012 ;
    wire signal_2013 ;
    wire signal_2014 ;
    wire signal_2015 ;
    wire signal_2016 ;
    wire signal_2017 ;
    wire signal_2018 ;
    wire signal_2019 ;
    wire signal_2020 ;
    wire signal_2021 ;
    wire signal_2022 ;
    wire signal_2023 ;
    wire signal_2024 ;
    wire signal_2025 ;
    wire signal_2026 ;
    wire signal_2027 ;
    wire signal_2028 ;
    wire signal_2029 ;
    wire signal_2030 ;
    wire signal_2031 ;
    wire signal_2032 ;
    wire signal_2033 ;
    wire signal_2034 ;
    wire signal_2035 ;
    wire signal_2036 ;
    wire signal_2037 ;
    wire signal_2038 ;
    wire signal_2039 ;
    wire signal_2040 ;
    wire signal_2041 ;
    wire signal_2042 ;
    wire signal_2043 ;
    wire signal_2044 ;
    wire signal_2045 ;
    wire signal_2046 ;
    wire signal_2047 ;
    wire signal_2048 ;
    wire signal_2049 ;
    wire signal_2050 ;
    wire signal_2051 ;
    wire signal_2052 ;
    wire signal_2053 ;
    wire signal_2054 ;
    wire signal_2055 ;
    wire signal_2056 ;
    wire signal_2057 ;
    wire signal_2058 ;
    wire signal_2059 ;
    wire signal_2060 ;
    wire signal_2061 ;
    wire signal_2062 ;
    wire signal_2063 ;
    wire signal_2064 ;
    wire signal_2065 ;
    wire signal_2066 ;
    wire signal_2067 ;
    wire signal_2068 ;
    wire signal_2069 ;
    wire signal_2070 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2079 ;
    wire signal_2080 ;
    wire signal_2081 ;
    wire signal_2082 ;
    wire signal_2083 ;
    wire signal_2084 ;
    wire signal_2085 ;
    wire signal_2086 ;
    wire signal_2087 ;
    wire signal_2088 ;
    wire signal_2089 ;
    wire signal_2090 ;
    wire signal_2091 ;
    wire signal_2092 ;
    wire signal_2093 ;
    wire signal_2094 ;
    wire signal_2095 ;
    wire signal_2096 ;
    wire signal_2097 ;
    wire signal_2098 ;
    wire signal_2099 ;
    wire signal_2100 ;
    wire signal_2101 ;
    wire signal_2102 ;
    wire signal_2103 ;
    wire signal_2104 ;
    wire signal_2105 ;
    wire signal_2106 ;
    wire signal_2107 ;
    wire signal_2108 ;
    wire signal_2109 ;
    wire signal_2110 ;
    wire signal_2111 ;
    wire signal_2112 ;
    wire signal_2113 ;
    wire signal_2114 ;
    wire signal_2115 ;
    wire signal_2116 ;
    wire signal_2117 ;
    wire signal_2118 ;
    wire signal_2119 ;
    wire signal_2120 ;
    wire signal_2121 ;
    wire signal_2122 ;
    wire signal_2123 ;
    wire signal_2124 ;
    wire signal_2125 ;
    wire signal_2126 ;
    wire signal_2127 ;
    wire signal_2128 ;
    wire signal_2129 ;
    wire signal_2130 ;
    wire signal_2131 ;
    wire signal_2132 ;
    wire signal_2133 ;
    wire signal_2134 ;
    wire signal_2135 ;
    wire signal_2136 ;
    wire signal_2137 ;
    wire signal_2138 ;
    wire signal_2139 ;
    wire signal_2140 ;
    wire signal_2141 ;
    wire signal_2142 ;
    wire signal_2143 ;
    wire signal_2144 ;
    wire signal_2145 ;
    wire signal_2146 ;
    wire signal_2147 ;
    wire signal_2148 ;
    wire signal_2149 ;
    wire signal_2150 ;
    wire signal_2151 ;
    wire signal_2152 ;
    wire signal_2153 ;
    wire signal_2154 ;
    wire signal_2155 ;
    wire signal_2156 ;
    wire signal_2157 ;
    wire signal_2158 ;
    wire signal_2159 ;
    wire signal_2160 ;
    wire signal_2161 ;
    wire signal_2162 ;
    wire signal_2163 ;
    wire signal_2164 ;
    wire signal_2165 ;
    wire signal_2166 ;
    wire signal_2167 ;
    wire signal_2168 ;
    wire signal_2169 ;
    wire signal_2170 ;
    wire signal_2171 ;
    wire signal_2172 ;
    wire signal_2173 ;
    wire signal_2174 ;
    wire signal_2175 ;
    wire signal_2176 ;
    wire signal_2177 ;
    wire signal_2178 ;
    wire signal_2179 ;
    wire signal_2180 ;
    wire signal_2181 ;
    wire signal_2182 ;
    wire signal_2183 ;
    wire signal_2184 ;
    wire signal_2185 ;
    wire signal_2186 ;
    wire signal_2187 ;
    wire signal_2188 ;
    wire signal_2189 ;
    wire signal_2190 ;
    wire signal_2191 ;
    wire signal_2192 ;
    wire signal_2193 ;
    wire signal_2194 ;
    wire signal_2195 ;
    wire signal_2196 ;
    wire signal_2197 ;
    wire signal_2198 ;
    wire signal_2199 ;
    wire signal_2200 ;
    wire signal_2201 ;
    wire signal_2202 ;
    wire signal_2203 ;
    wire signal_2204 ;
    wire signal_2205 ;
    wire signal_2206 ;
    wire signal_2207 ;
    wire signal_2208 ;
    wire signal_2209 ;
    wire signal_2210 ;
    wire signal_2211 ;
    wire signal_2212 ;
    wire signal_2213 ;
    wire signal_2214 ;
    wire signal_2215 ;
    wire signal_2216 ;
    wire signal_2217 ;
    wire signal_2218 ;
    wire signal_2219 ;
    wire signal_2220 ;
    wire signal_2221 ;
    wire signal_2222 ;
    wire signal_2223 ;
    wire signal_2224 ;
    wire signal_2225 ;
    wire signal_2226 ;
    wire signal_2227 ;
    wire signal_2228 ;
    wire signal_2229 ;
    wire signal_2230 ;
    wire signal_2231 ;
    wire signal_2232 ;
    wire signal_2233 ;
    wire signal_2234 ;
    wire signal_2235 ;
    wire signal_2236 ;
    wire signal_2237 ;
    wire signal_2238 ;
    wire signal_2239 ;
    wire signal_2240 ;
    wire signal_2241 ;
    wire signal_2242 ;
    wire signal_2243 ;
    wire signal_2244 ;
    wire signal_2245 ;
    wire signal_2246 ;
    wire signal_2247 ;
    wire signal_2248 ;
    wire signal_2249 ;
    wire signal_2250 ;
    wire signal_2251 ;
    wire signal_2252 ;
    wire signal_2253 ;
    wire signal_2254 ;
    wire signal_2255 ;
    wire signal_2256 ;
    wire signal_2257 ;
    wire signal_2258 ;
    wire signal_2259 ;
    wire signal_2260 ;
    wire signal_2261 ;
    wire signal_2262 ;
    wire signal_2263 ;
    wire signal_2264 ;
    wire signal_2265 ;
    wire signal_2266 ;
    wire signal_2267 ;
    wire signal_2268 ;
    wire signal_2269 ;
    wire signal_2270 ;
    wire signal_2271 ;
    wire signal_2272 ;
    wire signal_2273 ;
    wire signal_2274 ;
    wire signal_2275 ;
    wire signal_2276 ;
    wire signal_2277 ;
    wire signal_2278 ;
    wire signal_2279 ;
    wire signal_2280 ;
    wire signal_2281 ;
    wire signal_2282 ;
    wire signal_2283 ;
    wire signal_2284 ;
    wire signal_2285 ;
    wire signal_2286 ;
    wire signal_2287 ;
    wire signal_2288 ;
    wire signal_2289 ;
    wire signal_2290 ;
    wire signal_2291 ;
    wire signal_2292 ;
    wire signal_2293 ;
    wire signal_2294 ;
    wire signal_2295 ;
    wire signal_2296 ;
    wire signal_2297 ;
    wire signal_2298 ;
    wire signal_2299 ;
    wire signal_2300 ;
    wire signal_2301 ;
    wire signal_2302 ;
    wire signal_2303 ;
    wire signal_2304 ;
    wire signal_2305 ;
    wire signal_2306 ;
    wire signal_2307 ;
    wire signal_2308 ;
    wire signal_2309 ;
    wire signal_2310 ;
    wire signal_2311 ;
    wire signal_2312 ;
    wire signal_2313 ;
    wire signal_2314 ;
    wire signal_2315 ;
    wire signal_2316 ;
    wire signal_2317 ;
    wire signal_2318 ;
    wire signal_2319 ;
    wire signal_2320 ;
    wire signal_2321 ;
    wire signal_2322 ;
    wire signal_2323 ;
    wire signal_2324 ;
    wire signal_2325 ;
    wire signal_2326 ;
    wire signal_2327 ;
    wire signal_2328 ;
    wire signal_2329 ;
    wire signal_2330 ;
    wire signal_2331 ;
    wire signal_2332 ;
    wire signal_2333 ;
    wire signal_2334 ;
    wire signal_2335 ;
    wire signal_2336 ;
    wire signal_2337 ;
    wire signal_2338 ;
    wire signal_2339 ;
    wire signal_2340 ;
    wire signal_2341 ;
    wire signal_2342 ;
    wire signal_2343 ;
    wire signal_2344 ;
    wire signal_2345 ;
    wire signal_2346 ;
    wire signal_2347 ;
    wire signal_2348 ;
    wire signal_2349 ;
    wire signal_2350 ;
    wire signal_2351 ;
    wire signal_2352 ;
    wire signal_2353 ;
    wire signal_2354 ;
    wire signal_2355 ;
    wire signal_2356 ;
    wire signal_2357 ;
    wire signal_2358 ;
    wire signal_2359 ;
    wire signal_2360 ;
    wire signal_2361 ;
    wire signal_2362 ;
    wire signal_2363 ;
    wire signal_2364 ;
    wire signal_2365 ;
    wire signal_2366 ;
    wire signal_2367 ;
    wire signal_2368 ;
    wire signal_2369 ;
    wire signal_2370 ;
    wire signal_2371 ;
    wire signal_2372 ;
    wire signal_2373 ;
    wire signal_2374 ;
    wire signal_2375 ;
    wire signal_2376 ;
    wire signal_2377 ;
    wire signal_2378 ;
    wire signal_2379 ;
    wire signal_2380 ;
    wire signal_2381 ;
    wire signal_2382 ;
    wire signal_2383 ;
    wire signal_2384 ;
    wire signal_2385 ;
    wire signal_2386 ;
    wire signal_2387 ;
    wire signal_2388 ;
    wire signal_2389 ;
    wire signal_2390 ;
    wire signal_2391 ;
    wire signal_2392 ;
    wire signal_2393 ;
    wire signal_2394 ;
    wire signal_2395 ;
    wire signal_2396 ;
    wire signal_2397 ;
    wire signal_2398 ;
    wire signal_2399 ;
    wire signal_2400 ;
    wire signal_2401 ;
    wire signal_2402 ;
    wire signal_2403 ;
    wire signal_2404 ;
    wire signal_2405 ;
    wire signal_2406 ;
    wire signal_2407 ;
    wire signal_2408 ;
    wire signal_2409 ;
    wire signal_2410 ;
    wire signal_2411 ;
    wire signal_2412 ;
    wire signal_2413 ;
    wire signal_2414 ;
    wire signal_2415 ;
    wire signal_2416 ;
    wire signal_2417 ;
    wire signal_2418 ;
    wire signal_2419 ;
    wire signal_2420 ;
    wire signal_2421 ;
    wire signal_2422 ;
    wire signal_2423 ;
    wire signal_2424 ;
    wire signal_2425 ;
    wire signal_2426 ;
    wire signal_2427 ;
    wire signal_2428 ;
    wire signal_2429 ;
    wire signal_2430 ;
    wire signal_2431 ;
    wire signal_2432 ;
    wire signal_2433 ;
    wire signal_2434 ;
    wire signal_2435 ;
    wire signal_2436 ;
    wire signal_2437 ;
    wire signal_2438 ;
    wire signal_2439 ;
    wire signal_2440 ;
    wire signal_2441 ;
    wire signal_2442 ;
    wire signal_2443 ;
    wire signal_2444 ;
    wire signal_2445 ;
    wire signal_2446 ;
    wire signal_2447 ;
    wire signal_2448 ;
    wire signal_2449 ;
    wire signal_2450 ;
    wire signal_2451 ;
    wire signal_2452 ;
    wire signal_2453 ;
    wire signal_2454 ;
    wire signal_2455 ;
    wire signal_2456 ;
    wire signal_2457 ;
    wire signal_2458 ;
    wire signal_2459 ;
    wire signal_2460 ;
    wire signal_2461 ;
    wire signal_2462 ;
    wire signal_2463 ;
    wire signal_2464 ;
    wire signal_2465 ;
    wire signal_2466 ;
    wire signal_2467 ;
    wire signal_2468 ;
    wire signal_2469 ;
    wire signal_2470 ;
    wire signal_2471 ;
    wire signal_2472 ;
    wire signal_2473 ;
    wire signal_2474 ;
    wire signal_2475 ;
    wire signal_2476 ;
    wire signal_2477 ;
    wire signal_2478 ;
    wire signal_2479 ;
    wire signal_2480 ;
    wire signal_2481 ;
    wire signal_2482 ;
    wire signal_2483 ;
    wire signal_2484 ;
    wire signal_2485 ;
    wire signal_2486 ;
    wire signal_2487 ;
    wire signal_2488 ;
    wire signal_2489 ;
    wire signal_2490 ;
    wire signal_2491 ;
    wire signal_2492 ;
    wire signal_2493 ;
    wire signal_2494 ;
    wire signal_2495 ;
    wire signal_2496 ;
    wire signal_2497 ;
    wire signal_2498 ;
    wire signal_2499 ;
    wire signal_2500 ;
    wire signal_2501 ;
    wire signal_2502 ;
    wire signal_2503 ;
    wire signal_2504 ;
    wire signal_2505 ;
    wire signal_2506 ;
    wire signal_2507 ;
    wire signal_2508 ;
    wire signal_2509 ;
    wire signal_2510 ;
    wire signal_2511 ;
    wire signal_2512 ;
    wire signal_2513 ;
    wire signal_2514 ;
    wire signal_2515 ;
    wire signal_2516 ;
    wire signal_2517 ;
    wire signal_2518 ;
    wire signal_2519 ;
    wire signal_2520 ;
    wire signal_2521 ;
    wire signal_2522 ;
    wire signal_2523 ;
    wire signal_2524 ;
    wire signal_2525 ;
    wire signal_2526 ;
    wire signal_2527 ;
    wire signal_2528 ;
    wire signal_2529 ;
    wire signal_2530 ;
    wire signal_2531 ;
    wire signal_2532 ;
    wire signal_2533 ;
    wire signal_2534 ;
    wire signal_2535 ;
    wire signal_2536 ;
    wire signal_2537 ;
    wire signal_2538 ;
    wire signal_2539 ;
    wire signal_2540 ;
    wire signal_2541 ;
    wire signal_2542 ;
    wire signal_2543 ;
    wire signal_2544 ;
    wire signal_2545 ;
    wire signal_2546 ;
    wire signal_2547 ;
    wire signal_2548 ;
    wire signal_2549 ;
    wire signal_2550 ;
    wire signal_2551 ;
    wire signal_2552 ;
    wire signal_2553 ;
    wire signal_2554 ;
    wire signal_2555 ;
    wire signal_2556 ;
    wire signal_2557 ;
    wire signal_2558 ;
    wire signal_2559 ;
    wire signal_2561 ;
    wire signal_2562 ;
    wire signal_2563 ;
    wire signal_2564 ;
    wire signal_2565 ;
    wire signal_2566 ;
    wire signal_2567 ;
    wire signal_2568 ;
    wire signal_2569 ;
    wire signal_2570 ;
    wire signal_2571 ;
    wire signal_2572 ;
    wire signal_2573 ;
    wire signal_2574 ;
    wire signal_2575 ;
    wire signal_2576 ;
    wire signal_2577 ;
    wire signal_2578 ;
    wire signal_2579 ;
    wire signal_2580 ;
    wire signal_2581 ;
    wire signal_2582 ;
    wire signal_2583 ;
    wire signal_2584 ;
    wire signal_2585 ;
    wire signal_2587 ;
    wire signal_2589 ;
    wire signal_2591 ;
    wire signal_2593 ;
    wire signal_2595 ;
    wire signal_2597 ;
    wire signal_2599 ;
    wire signal_2601 ;
    wire signal_2603 ;
    wire signal_2604 ;
    wire signal_2605 ;
    wire signal_2606 ;
    wire signal_2607 ;
    wire signal_2608 ;
    wire signal_2609 ;
    wire signal_2610 ;
    wire signal_2611 ;
    wire signal_2612 ;
    wire signal_2613 ;
    wire signal_2614 ;
    wire signal_2615 ;
    wire signal_2616 ;
    wire signal_2617 ;
    wire signal_2618 ;
    wire signal_2619 ;
    wire signal_2620 ;
    wire signal_2621 ;
    wire signal_2622 ;
    wire signal_2623 ;
    wire signal_2624 ;
    wire signal_2625 ;
    wire signal_2626 ;
    wire signal_2627 ;
    wire signal_2628 ;
    wire signal_2629 ;
    wire signal_2630 ;
    wire signal_2631 ;
    wire signal_2632 ;
    wire signal_2633 ;
    wire signal_2634 ;
    wire signal_2635 ;
    wire signal_2637 ;
    wire signal_2639 ;
    wire signal_2641 ;
    wire signal_2643 ;
    wire signal_2644 ;
    wire signal_2645 ;
    wire signal_2646 ;
    wire signal_2647 ;
    wire signal_2648 ;
    wire signal_2649 ;
    wire signal_2650 ;
    wire signal_2651 ;
    wire signal_2652 ;
    wire signal_2653 ;
    wire signal_2654 ;
    wire signal_2655 ;
    wire signal_2656 ;
    wire signal_2657 ;
    wire signal_2658 ;
    wire signal_2659 ;
    wire signal_2660 ;
    wire signal_2661 ;
    wire signal_2662 ;
    wire signal_2663 ;
    wire signal_2664 ;
    wire signal_2665 ;
    wire signal_2666 ;
    wire signal_2667 ;
    wire signal_2668 ;
    wire signal_2669 ;
    wire signal_2670 ;
    wire signal_2671 ;
    wire signal_2672 ;
    wire signal_2673 ;
    wire signal_2674 ;
    wire signal_2675 ;
    wire signal_2676 ;
    wire signal_2677 ;
    wire signal_2679 ;
    wire signal_2681 ;
    wire signal_2683 ;
    wire signal_2685 ;
    wire signal_2687 ;
    wire signal_2689 ;
    wire signal_2691 ;
    wire signal_2693 ;
    wire signal_2694 ;
    wire signal_2695 ;
    wire signal_2696 ;
    wire signal_2697 ;
    wire signal_2698 ;
    wire signal_2699 ;
    wire signal_2700 ;
    wire signal_2701 ;
    wire signal_2702 ;
    wire signal_2703 ;
    wire signal_2704 ;
    wire signal_2705 ;
    wire signal_2706 ;
    wire signal_2707 ;
    wire signal_2708 ;
    wire signal_2709 ;
    wire signal_2710 ;
    wire signal_2711 ;
    wire signal_2712 ;
    wire signal_2713 ;
    wire signal_2714 ;
    wire signal_2715 ;
    wire signal_2716 ;
    wire signal_2717 ;
    wire signal_2718 ;
    wire signal_2719 ;
    wire signal_2720 ;
    wire signal_2721 ;
    wire signal_2722 ;
    wire signal_2723 ;
    wire signal_2724 ;
    wire signal_2725 ;
    wire signal_2726 ;
    wire signal_2728 ;
    wire signal_2730 ;
    wire signal_2732 ;
    wire signal_2734 ;
    wire signal_2736 ;
    wire signal_2738 ;
    wire signal_2740 ;
    wire signal_2742 ;
    wire signal_2743 ;
    wire signal_2744 ;
    wire signal_2745 ;
    wire signal_2746 ;
    wire signal_2747 ;
    wire signal_2748 ;
    wire signal_2749 ;
    wire signal_2750 ;
    wire signal_2751 ;
    wire signal_2752 ;
    wire signal_2753 ;
    wire signal_2754 ;
    wire signal_2755 ;
    wire signal_2756 ;
    wire signal_2757 ;
    wire signal_2758 ;
    wire signal_2759 ;
    wire signal_2760 ;
    wire signal_2761 ;
    wire signal_2763 ;
    wire signal_2765 ;
    wire signal_2767 ;
    wire signal_2769 ;
    wire signal_2771 ;
    wire signal_2773 ;
    wire signal_2775 ;
    wire signal_2777 ;
    wire signal_2779 ;
    wire signal_2781 ;
    wire signal_2783 ;
    wire signal_2785 ;
    wire signal_2786 ;
    wire signal_2787 ;
    wire signal_2788 ;
    wire signal_2789 ;
    wire signal_2790 ;
    wire signal_2791 ;
    wire signal_2792 ;
    wire signal_2793 ;
    wire signal_2794 ;
    wire signal_2795 ;
    wire signal_2796 ;
    wire signal_2797 ;
    wire signal_2798 ;
    wire signal_2799 ;
    wire signal_2800 ;
    wire signal_2801 ;
    wire signal_2803 ;
    wire signal_2805 ;
    wire signal_2807 ;
    wire signal_2809 ;
    wire signal_2811 ;
    wire signal_2813 ;
    wire signal_2815 ;
    wire signal_2816 ;
    wire signal_2817 ;
    wire signal_2818 ;
    wire signal_2819 ;
    wire signal_2820 ;
    wire signal_2821 ;
    wire signal_2823 ;
    wire signal_2825 ;
    wire signal_2827 ;
    wire signal_2829 ;
    wire signal_2831 ;
    wire signal_2833 ;
    wire signal_2835 ;
    wire signal_2836 ;
    wire signal_2837 ;
    wire signal_2838 ;
    wire signal_2839 ;
    wire signal_2840 ;
    wire signal_2841 ;
    wire signal_2842 ;
    wire signal_2843 ;
    wire signal_2844 ;
    wire signal_2845 ;
    wire signal_2846 ;
    wire signal_2847 ;
    wire signal_2848 ;
    wire signal_2849 ;
    wire signal_2850 ;
    wire signal_2851 ;
    wire signal_2852 ;
    wire signal_2853 ;
    wire signal_2854 ;
    wire signal_2855 ;
    wire signal_2857 ;
    wire signal_2859 ;
    wire signal_2860 ;
    wire signal_2861 ;
    wire signal_2862 ;
    wire signal_2863 ;
    wire signal_2865 ;
    wire signal_2867 ;
    wire signal_2869 ;
    wire signal_2871 ;
    wire signal_2873 ;
    wire signal_2875 ;
    wire signal_2940 ;
    wire signal_2941 ;
    wire signal_2942 ;
    wire signal_2943 ;
    wire signal_2944 ;
    wire signal_2945 ;
    wire signal_2946 ;
    wire signal_2947 ;
    wire signal_2948 ;
    wire signal_2949 ;
    wire signal_2950 ;
    wire signal_2951 ;
    wire signal_2952 ;
    wire signal_2953 ;
    wire signal_2954 ;
    wire signal_2955 ;
    wire signal_2956 ;
    wire signal_2957 ;
    wire signal_2958 ;
    wire signal_2959 ;
    wire signal_2960 ;
    wire signal_2961 ;
    wire signal_2962 ;
    wire signal_2963 ;
    wire signal_2964 ;
    wire signal_2965 ;
    wire signal_2966 ;
    wire signal_2967 ;
    wire signal_2968 ;
    wire signal_2969 ;
    wire signal_2970 ;
    wire signal_2971 ;
    wire signal_2972 ;
    wire signal_2973 ;
    wire signal_2974 ;
    wire signal_2975 ;
    wire signal_2976 ;
    wire signal_2977 ;
    wire signal_2978 ;
    wire signal_2979 ;
    wire signal_2980 ;
    wire signal_2981 ;
    wire signal_2982 ;
    wire signal_2983 ;
    wire signal_2984 ;
    wire signal_2985 ;
    wire signal_2986 ;
    wire signal_2987 ;
    wire signal_2988 ;
    wire signal_2989 ;
    wire signal_2990 ;
    wire signal_2991 ;
    wire signal_2992 ;
    wire signal_2993 ;
    wire signal_2994 ;
    wire signal_2995 ;
    wire signal_2996 ;
    wire signal_2997 ;
    wire signal_2998 ;
    wire signal_2999 ;
    wire signal_3000 ;
    wire signal_3001 ;
    wire signal_3002 ;
    wire signal_3003 ;
    wire signal_3004 ;
    wire signal_3005 ;
    wire signal_3006 ;
    wire signal_3007 ;
    wire signal_3008 ;
    wire signal_3009 ;
    wire signal_3010 ;
    wire signal_3011 ;
    wire signal_3012 ;
    wire signal_3013 ;
    wire signal_3014 ;
    wire signal_3015 ;
    wire signal_3016 ;
    wire signal_3017 ;
    wire signal_3018 ;
    wire signal_3019 ;
    wire signal_3020 ;
    wire signal_3021 ;
    wire signal_3022 ;
    wire signal_3023 ;
    wire signal_3024 ;
    wire signal_3025 ;
    wire signal_3026 ;
    wire signal_3027 ;
    wire signal_3028 ;
    wire signal_3029 ;
    wire signal_3030 ;
    wire signal_3031 ;
    wire signal_3032 ;
    wire signal_3033 ;
    wire signal_3034 ;
    wire signal_3035 ;
    wire signal_3036 ;
    wire signal_3037 ;
    wire signal_3038 ;
    wire signal_3039 ;
    wire signal_3040 ;
    wire signal_3041 ;
    wire signal_3042 ;
    wire signal_3043 ;
    wire signal_3044 ;
    wire signal_3045 ;
    wire signal_3046 ;
    wire signal_3047 ;
    wire signal_3048 ;
    wire signal_3049 ;
    wire signal_3050 ;
    wire signal_3051 ;
    wire signal_3052 ;
    wire signal_3053 ;
    wire signal_3054 ;
    wire signal_3055 ;
    wire signal_3056 ;
    wire signal_3057 ;
    wire signal_3058 ;
    wire signal_3059 ;
    wire signal_3060 ;
    wire signal_3061 ;
    wire signal_3062 ;
    wire signal_3063 ;
    wire signal_3064 ;
    wire signal_3065 ;
    wire signal_3066 ;
    wire signal_3067 ;
    wire signal_3068 ;
    wire signal_3069 ;
    wire signal_3070 ;
    wire signal_3071 ;
    wire signal_3072 ;
    wire signal_3073 ;
    wire signal_3074 ;
    wire signal_3075 ;
    wire signal_3076 ;
    wire signal_3077 ;
    wire signal_3078 ;
    wire signal_3079 ;
    wire signal_3080 ;
    wire signal_3081 ;
    wire signal_3082 ;
    wire signal_3083 ;
    wire signal_3084 ;
    wire signal_3085 ;
    wire signal_3086 ;
    wire signal_3087 ;
    wire signal_3088 ;
    wire signal_3089 ;
    wire signal_3090 ;
    wire signal_3091 ;
    wire signal_3092 ;
    wire signal_3093 ;
    wire signal_3094 ;
    wire signal_3095 ;
    wire signal_3096 ;
    wire signal_3097 ;
    wire signal_3098 ;
    wire signal_3099 ;
    wire signal_3100 ;
    wire signal_3101 ;
    wire signal_3102 ;
    wire signal_3103 ;
    wire signal_3104 ;
    wire signal_3105 ;
    wire signal_3106 ;
    wire signal_3107 ;
    wire signal_3108 ;
    wire signal_3109 ;
    wire signal_3110 ;
    wire signal_3111 ;
    wire signal_3112 ;
    wire signal_3113 ;
    wire signal_3114 ;
    wire signal_3115 ;
    wire signal_3116 ;
    wire signal_3117 ;
    wire signal_3118 ;
    wire signal_3119 ;
    wire signal_3120 ;
    wire signal_3121 ;
    wire signal_3122 ;
    wire signal_3123 ;
    wire signal_3124 ;
    wire signal_3125 ;
    wire signal_3126 ;
    wire signal_3127 ;
    wire signal_3128 ;
    wire signal_3129 ;
    wire signal_3130 ;
    wire signal_3131 ;
    wire signal_3132 ;
    wire signal_3133 ;
    wire signal_3134 ;
    wire signal_3135 ;
    wire signal_3136 ;
    wire signal_3137 ;
    wire signal_3138 ;
    wire signal_3139 ;
    wire signal_3140 ;
    wire signal_3141 ;
    wire signal_3142 ;
    wire signal_3143 ;
    wire signal_3144 ;
    wire signal_3145 ;
    wire signal_3146 ;
    wire signal_3147 ;
    wire signal_3148 ;
    wire signal_3149 ;
    wire signal_3150 ;
    wire signal_3151 ;
    wire signal_3152 ;
    wire signal_3153 ;
    wire signal_3154 ;
    wire signal_3155 ;
    wire signal_3156 ;
    wire signal_3157 ;
    wire signal_3158 ;
    wire signal_3159 ;
    wire signal_3160 ;
    wire signal_3161 ;
    wire signal_3162 ;
    wire signal_3163 ;
    wire signal_3164 ;
    wire signal_3165 ;
    wire signal_3166 ;
    wire signal_3167 ;
    wire signal_3168 ;
    wire signal_3169 ;
    wire signal_3170 ;
    wire signal_3171 ;
    wire signal_3172 ;
    wire signal_3173 ;
    wire signal_3174 ;
    wire signal_3175 ;
    wire signal_3176 ;
    wire signal_3177 ;
    wire signal_3178 ;
    wire signal_3179 ;
    wire signal_3180 ;
    wire signal_3181 ;
    wire signal_3182 ;
    wire signal_3183 ;
    wire signal_3184 ;
    wire signal_3185 ;
    wire signal_3186 ;
    wire signal_3187 ;
    wire signal_3188 ;
    wire signal_3189 ;
    wire signal_3190 ;
    wire signal_3191 ;
    wire signal_3192 ;
    wire signal_3193 ;
    wire signal_3194 ;
    wire signal_3195 ;
    wire signal_3196 ;
    wire signal_3197 ;
    wire signal_3198 ;
    wire signal_3199 ;
    wire signal_3200 ;
    wire signal_3201 ;
    wire signal_3202 ;
    wire signal_3203 ;
    wire signal_3204 ;
    wire signal_3205 ;
    wire signal_3206 ;
    wire signal_3207 ;
    wire signal_3208 ;
    wire signal_3209 ;
    wire signal_3210 ;
    wire signal_3211 ;
    wire signal_3212 ;
    wire signal_3213 ;
    wire signal_3214 ;
    wire signal_3215 ;
    wire signal_3216 ;
    wire signal_3217 ;
    wire signal_3218 ;
    wire signal_3219 ;
    wire signal_3220 ;
    wire signal_3221 ;
    wire signal_3222 ;
    wire signal_3223 ;
    wire signal_3224 ;
    wire signal_3225 ;
    wire signal_3226 ;
    wire signal_3227 ;
    wire signal_3228 ;
    wire signal_3229 ;
    wire signal_3230 ;
    wire signal_3231 ;
    wire signal_3232 ;
    wire signal_3233 ;
    wire signal_3234 ;
    wire signal_3235 ;
    wire signal_3236 ;
    wire signal_3237 ;
    wire signal_3238 ;
    wire signal_3239 ;
    wire signal_3240 ;
    wire signal_3241 ;
    wire signal_3242 ;
    wire signal_3243 ;
    wire signal_3244 ;
    wire signal_3245 ;
    wire signal_3246 ;
    wire signal_3247 ;
    wire signal_3248 ;
    wire signal_3249 ;
    wire signal_3250 ;
    wire signal_3251 ;
    wire signal_3252 ;
    wire signal_3253 ;
    wire signal_3254 ;
    wire signal_3255 ;
    wire signal_3256 ;
    wire signal_3257 ;
    wire signal_3258 ;
    wire signal_3259 ;
    wire signal_3260 ;
    wire signal_3261 ;
    wire signal_3262 ;
    wire signal_3263 ;
    wire signal_3264 ;
    wire signal_3265 ;
    wire signal_3266 ;
    wire signal_3267 ;
    wire signal_3268 ;
    wire signal_3269 ;
    wire signal_3270 ;
    wire signal_3271 ;
    wire signal_3272 ;
    wire signal_3273 ;
    wire signal_3274 ;
    wire signal_3275 ;
    wire signal_3276 ;
    wire signal_3277 ;
    wire signal_3278 ;
    wire signal_3279 ;
    wire signal_3280 ;
    wire signal_3281 ;
    wire signal_3282 ;
    wire signal_3283 ;
    wire signal_3284 ;
    wire signal_3285 ;
    wire signal_3286 ;
    wire signal_3287 ;
    wire signal_3288 ;
    wire signal_3289 ;
    wire signal_3290 ;
    wire signal_3291 ;
    wire signal_3292 ;
    wire signal_3293 ;
    wire signal_3294 ;
    wire signal_3295 ;
    wire signal_3296 ;
    wire signal_3297 ;
    wire signal_3298 ;
    wire signal_3299 ;
    wire signal_3300 ;
    wire signal_3301 ;
    wire signal_3302 ;
    wire signal_3303 ;
    wire signal_3304 ;
    wire signal_3305 ;
    wire signal_3306 ;
    wire signal_3307 ;
    wire signal_3308 ;
    wire signal_3309 ;
    wire signal_3310 ;
    wire signal_3311 ;
    wire signal_3312 ;
    wire signal_3313 ;
    wire signal_3314 ;
    wire signal_3315 ;
    wire signal_3316 ;
    wire signal_3317 ;
    wire signal_3318 ;
    wire signal_3319 ;
    wire signal_3320 ;
    wire signal_3321 ;
    wire signal_3322 ;
    wire signal_3323 ;
    wire signal_3324 ;
    wire signal_3325 ;
    wire signal_3326 ;
    wire signal_3327 ;
    wire signal_3328 ;
    wire signal_3329 ;
    wire signal_3330 ;
    wire signal_3331 ;
    wire signal_3332 ;
    wire signal_3333 ;
    wire signal_3334 ;
    wire signal_3335 ;
    wire signal_3336 ;
    wire signal_3337 ;
    wire signal_3338 ;
    wire signal_3339 ;
    wire signal_3340 ;
    wire signal_3341 ;
    wire signal_3342 ;
    wire signal_3343 ;
    wire signal_3344 ;
    wire signal_3345 ;
    wire signal_3346 ;
    wire signal_3347 ;
    wire signal_3348 ;
    wire signal_3349 ;
    wire signal_3350 ;
    wire signal_3351 ;
    wire signal_3352 ;
    wire signal_3353 ;
    wire signal_3354 ;
    wire signal_3355 ;
    wire signal_3356 ;
    wire signal_3357 ;
    wire signal_3358 ;
    wire signal_3359 ;
    wire signal_3360 ;
    wire signal_3361 ;
    wire signal_3362 ;
    wire signal_3363 ;
    wire signal_3364 ;
    wire signal_3365 ;
    wire signal_3366 ;
    wire signal_3367 ;
    wire signal_3368 ;
    wire signal_3369 ;
    wire signal_3370 ;
    wire signal_3371 ;
    wire signal_3372 ;
    wire signal_3373 ;
    wire signal_3374 ;
    wire signal_3375 ;
    wire signal_3376 ;
    wire signal_3377 ;
    wire signal_3378 ;
    wire signal_3379 ;
    wire signal_3380 ;
    wire signal_3381 ;
    wire signal_3382 ;
    wire signal_3383 ;
    wire signal_3384 ;
    wire signal_3385 ;
    wire signal_3386 ;
    wire signal_3387 ;
    wire signal_3388 ;
    wire signal_3389 ;
    wire signal_3390 ;
    wire signal_3391 ;
    wire signal_3392 ;
    wire signal_3393 ;
    wire signal_3394 ;
    wire signal_3395 ;
    wire signal_3396 ;
    wire signal_3397 ;
    wire signal_3398 ;
    wire signal_3399 ;
    wire signal_3400 ;
    wire signal_3401 ;
    wire signal_3402 ;
    wire signal_3403 ;
    wire signal_3404 ;
    wire signal_3405 ;
    wire signal_3406 ;
    wire signal_3407 ;
    wire signal_3408 ;
    wire signal_3409 ;
    wire signal_3410 ;
    wire signal_3411 ;
    wire signal_3412 ;
    wire signal_3413 ;
    wire signal_3414 ;
    wire signal_3415 ;
    wire signal_3416 ;
    wire signal_3417 ;
    wire signal_3418 ;
    wire signal_3419 ;
    wire signal_3420 ;
    wire signal_3421 ;
    wire signal_3422 ;
    wire signal_3423 ;
    wire signal_3424 ;
    wire signal_3425 ;
    wire signal_3426 ;
    wire signal_3427 ;
    wire signal_3428 ;
    wire signal_3429 ;
    wire signal_3430 ;
    wire signal_3431 ;
    wire signal_3432 ;
    wire signal_3433 ;
    wire signal_3434 ;
    wire signal_3435 ;
    wire signal_3436 ;
    wire signal_3437 ;
    wire signal_3438 ;
    wire signal_3439 ;
    wire signal_3440 ;
    wire signal_3441 ;
    wire signal_3442 ;
    wire signal_3443 ;
    wire signal_3444 ;
    wire signal_3445 ;
    wire signal_3446 ;
    wire signal_3447 ;
    wire signal_3448 ;
    wire signal_3449 ;
    wire signal_3450 ;
    wire signal_3451 ;
    wire signal_3452 ;
    wire signal_3453 ;
    wire signal_3454 ;
    wire signal_3455 ;
    wire signal_3456 ;
    wire signal_3457 ;
    wire signal_3458 ;
    wire signal_3459 ;
    wire signal_3460 ;
    wire signal_3461 ;
    wire signal_3462 ;
    wire signal_3463 ;
    wire signal_3464 ;
    wire signal_3465 ;
    wire signal_3466 ;
    wire signal_3467 ;
    wire signal_3468 ;
    wire signal_3469 ;
    wire signal_3470 ;
    wire signal_3471 ;
    wire signal_3472 ;
    wire signal_3473 ;
    wire signal_3474 ;
    wire signal_3475 ;
    wire signal_3476 ;
    wire signal_3477 ;
    wire signal_3478 ;
    wire signal_3479 ;
    wire signal_3480 ;
    wire signal_3481 ;
    wire signal_3482 ;
    wire signal_3483 ;
    wire signal_3484 ;
    wire signal_3485 ;
    wire signal_3486 ;
    wire signal_3487 ;
    wire signal_3488 ;
    wire signal_3489 ;
    wire signal_3490 ;
    wire signal_3491 ;
    wire signal_3492 ;
    wire signal_3493 ;
    wire signal_3494 ;
    wire signal_3495 ;
    wire signal_3496 ;
    wire signal_3497 ;
    wire signal_3498 ;
    wire signal_3499 ;
    wire signal_3500 ;
    wire signal_3501 ;
    wire signal_3502 ;
    wire signal_3503 ;
    wire signal_3504 ;
    wire signal_3505 ;
    wire signal_3506 ;
    wire signal_3507 ;
    wire signal_3508 ;
    wire signal_3509 ;
    wire signal_3510 ;
    wire signal_3511 ;
    wire signal_3512 ;
    wire signal_3513 ;
    wire signal_3514 ;
    wire signal_3515 ;
    wire signal_3516 ;
    wire signal_3517 ;
    wire signal_3518 ;
    wire signal_3519 ;
    wire signal_3520 ;
    wire signal_3521 ;
    wire signal_3522 ;
    wire signal_3523 ;
    wire signal_3524 ;
    wire signal_3525 ;
    wire signal_3526 ;
    wire signal_3527 ;
    wire signal_3528 ;
    wire signal_3529 ;
    wire signal_3530 ;
    wire signal_3531 ;
    wire signal_3532 ;
    wire signal_3533 ;
    wire signal_3534 ;
    wire signal_3535 ;
    wire signal_3536 ;
    wire signal_3537 ;
    wire signal_3538 ;
    wire signal_3539 ;
    wire signal_3540 ;
    wire signal_3541 ;
    wire signal_3542 ;
    wire signal_3543 ;
    wire signal_3544 ;
    wire signal_3545 ;
    wire signal_3546 ;
    wire signal_3547 ;
    wire signal_3548 ;
    wire signal_3549 ;
    wire signal_3550 ;
    wire signal_3551 ;
    wire signal_3552 ;
    wire signal_3553 ;
    wire signal_3554 ;
    wire signal_3555 ;
    wire signal_3556 ;
    wire signal_3557 ;
    wire signal_3558 ;
    wire signal_3559 ;
    wire signal_3560 ;
    wire signal_3561 ;
    wire signal_3562 ;
    wire signal_3563 ;
    wire signal_3564 ;
    wire signal_3565 ;
    wire signal_3566 ;
    wire signal_3567 ;
    wire signal_3568 ;
    wire signal_3569 ;
    wire signal_3570 ;
    wire signal_3571 ;
    wire signal_3572 ;
    wire signal_3573 ;
    wire signal_3574 ;
    wire signal_3575 ;
    wire signal_3576 ;
    wire signal_3577 ;
    wire signal_3578 ;
    wire signal_3579 ;
    wire signal_3580 ;
    wire signal_3581 ;
    wire signal_3582 ;
    wire signal_3583 ;
    wire signal_3584 ;
    wire signal_3585 ;
    wire signal_3586 ;
    wire signal_3587 ;
    wire signal_3588 ;
    wire signal_3589 ;
    wire signal_3590 ;
    wire signal_3591 ;
    wire signal_3592 ;
    wire signal_3593 ;
    wire signal_3594 ;
    wire signal_3595 ;
    wire signal_3596 ;
    wire signal_3597 ;
    wire signal_3598 ;
    wire signal_3599 ;
    wire signal_3600 ;
    wire signal_3601 ;
    wire signal_3602 ;
    wire signal_3603 ;
    wire signal_3604 ;
    wire signal_3605 ;
    wire signal_3606 ;
    wire signal_3607 ;
    wire signal_3608 ;
    wire signal_3609 ;
    wire signal_3610 ;
    wire signal_3611 ;
    wire signal_3612 ;
    wire signal_3613 ;
    wire signal_3614 ;
    wire signal_3615 ;
    wire signal_3616 ;
    wire signal_3617 ;
    wire signal_3618 ;
    wire signal_3619 ;
    wire signal_3620 ;
    wire signal_3621 ;
    wire signal_3622 ;
    wire signal_3623 ;
    wire signal_3624 ;
    wire signal_3625 ;
    wire signal_3626 ;
    wire signal_3627 ;
    wire signal_3628 ;
    wire signal_3629 ;
    wire signal_3630 ;
    wire signal_3631 ;
    wire signal_3632 ;
    wire signal_3633 ;
    wire signal_3634 ;
    wire signal_3635 ;
    wire signal_3636 ;
    wire signal_3637 ;
    wire signal_3638 ;
    wire signal_3639 ;
    wire signal_3640 ;
    wire signal_3641 ;
    wire signal_3642 ;
    wire signal_3643 ;
    wire signal_3644 ;
    wire signal_3645 ;
    wire signal_3646 ;
    wire signal_3647 ;
    wire signal_3648 ;
    wire signal_3649 ;
    wire signal_3650 ;
    wire signal_3651 ;
    wire signal_3652 ;
    wire signal_3653 ;
    wire signal_3654 ;
    wire signal_3655 ;
    wire signal_3656 ;
    wire signal_3657 ;
    wire signal_3658 ;
    wire signal_3659 ;
    wire signal_3660 ;
    wire signal_3661 ;
    wire signal_3662 ;
    wire signal_3663 ;
    wire signal_3664 ;
    wire signal_3665 ;
    wire signal_3666 ;
    wire signal_3667 ;
    wire signal_3668 ;
    wire signal_3669 ;
    wire signal_3670 ;
    wire signal_3671 ;
    wire signal_3672 ;
    wire signal_3673 ;
    wire signal_3674 ;
    wire signal_3675 ;
    wire signal_3676 ;
    wire signal_3677 ;
    wire signal_3678 ;
    wire signal_3679 ;
    wire signal_3680 ;
    wire signal_3681 ;
    wire signal_3682 ;
    wire signal_3683 ;
    wire signal_3684 ;
    wire signal_3685 ;
    wire signal_3686 ;
    wire signal_3687 ;
    wire signal_3688 ;
    wire signal_3689 ;
    wire signal_3690 ;
    wire signal_3691 ;
    wire signal_3692 ;
    wire signal_3693 ;
    wire signal_3694 ;
    wire signal_3695 ;
    wire signal_3696 ;
    wire signal_3697 ;
    wire signal_3698 ;
    wire signal_3699 ;
    wire signal_3700 ;
    wire signal_3701 ;
    wire signal_3702 ;
    wire signal_3703 ;
    wire signal_3704 ;
    wire signal_3705 ;
    wire signal_3706 ;
    wire signal_3707 ;
    wire signal_3708 ;
    wire signal_3709 ;
    wire signal_3710 ;
    wire signal_3711 ;
    wire signal_3712 ;
    wire signal_3713 ;
    wire signal_3714 ;
    wire signal_3715 ;
    wire signal_3716 ;
    wire signal_3717 ;
    wire signal_3718 ;
    wire signal_3719 ;
    wire signal_3720 ;
    wire signal_3721 ;
    wire signal_3722 ;
    wire signal_3723 ;
    wire signal_3724 ;
    wire signal_3725 ;
    wire signal_3726 ;
    wire signal_3727 ;
    wire signal_3728 ;
    wire signal_3729 ;
    wire signal_3730 ;
    wire signal_3731 ;
    wire signal_3732 ;
    wire signal_3733 ;
    wire signal_3734 ;
    wire signal_3735 ;
    wire signal_3736 ;
    wire signal_3737 ;
    wire signal_3738 ;
    wire signal_3739 ;
    wire signal_3740 ;
    wire signal_3741 ;
    wire signal_3742 ;
    wire signal_3743 ;
    wire signal_3744 ;
    wire signal_3745 ;
    wire signal_3746 ;
    wire signal_3747 ;
    wire signal_3748 ;
    wire signal_3749 ;
    wire signal_3750 ;
    wire signal_3751 ;
    wire signal_3752 ;
    wire signal_3753 ;
    wire signal_3754 ;
    wire signal_3755 ;
    wire signal_3756 ;
    wire signal_3757 ;
    wire signal_3758 ;
    wire signal_3759 ;
    wire signal_3760 ;
    wire signal_3761 ;
    wire signal_3762 ;
    wire signal_3763 ;
    wire signal_3764 ;
    wire signal_3765 ;
    wire signal_3766 ;
    wire signal_3767 ;
    wire signal_3768 ;
    wire signal_3769 ;
    wire signal_3770 ;
    wire signal_3771 ;
    wire signal_3772 ;
    wire signal_3773 ;
    wire signal_3774 ;
    wire signal_3775 ;
    wire signal_3776 ;
    wire signal_3777 ;
    wire signal_3778 ;
    wire signal_3779 ;
    wire signal_3780 ;
    wire signal_3781 ;
    wire signal_3782 ;
    wire signal_3783 ;
    wire signal_3784 ;
    wire signal_3785 ;
    wire signal_3786 ;
    wire signal_3787 ;
    wire signal_3788 ;
    wire signal_3789 ;
    wire signal_3790 ;
    wire signal_3791 ;
    wire signal_3792 ;
    wire signal_3793 ;
    wire signal_3794 ;
    wire signal_3795 ;
    wire signal_3796 ;
    wire signal_3797 ;
    wire signal_3798 ;
    wire signal_3799 ;
    wire signal_3800 ;
    wire signal_3801 ;
    wire signal_3802 ;
    wire signal_3803 ;
    wire signal_3804 ;
    wire signal_3805 ;
    wire signal_3806 ;
    wire signal_3807 ;
    wire signal_3808 ;
    wire signal_3809 ;
    wire signal_3810 ;
    wire signal_3811 ;
    wire signal_3812 ;
    wire signal_3813 ;
    wire signal_3814 ;
    wire signal_3815 ;
    wire signal_3816 ;
    wire signal_3817 ;
    wire signal_3818 ;
    wire signal_3819 ;
    wire signal_3820 ;
    wire signal_3821 ;
    wire signal_3822 ;
    wire signal_3823 ;
    wire signal_3824 ;
    wire signal_3825 ;
    wire signal_3826 ;
    wire signal_3827 ;
    wire signal_3828 ;
    wire signal_3829 ;
    wire signal_3830 ;
    wire signal_3831 ;
    wire signal_3832 ;
    wire signal_3833 ;
    wire signal_3834 ;
    wire signal_3835 ;
    wire signal_3836 ;
    wire signal_3837 ;
    wire signal_3838 ;
    wire signal_3839 ;
    wire signal_3840 ;
    wire signal_3841 ;
    wire signal_3842 ;
    wire signal_3843 ;
    wire signal_3844 ;
    wire signal_3845 ;
    wire signal_3846 ;
    wire signal_3847 ;
    wire signal_3848 ;
    wire signal_3849 ;
    wire signal_3850 ;
    wire signal_3851 ;
    wire signal_3852 ;
    wire signal_3853 ;
    wire signal_3854 ;
    wire signal_3855 ;
    wire signal_3856 ;
    wire signal_3857 ;
    wire signal_3858 ;
    wire signal_3859 ;
    wire signal_3860 ;
    wire signal_3861 ;
    wire signal_3862 ;
    wire signal_3863 ;
    wire signal_3864 ;
    wire signal_3865 ;
    wire signal_3866 ;
    wire signal_3867 ;
    wire signal_3868 ;
    wire signal_3869 ;
    wire signal_3870 ;
    wire signal_3871 ;
    wire signal_3872 ;
    wire signal_3873 ;
    wire signal_3874 ;
    wire signal_3875 ;
    wire signal_3876 ;
    wire signal_3877 ;
    wire signal_3878 ;
    wire signal_3879 ;
    wire signal_3880 ;
    wire signal_3881 ;
    wire signal_3882 ;
    wire signal_3883 ;
    wire signal_3884 ;
    wire signal_3885 ;
    wire signal_3886 ;
    wire signal_3887 ;
    wire signal_3888 ;
    wire signal_3889 ;
    wire signal_3890 ;
    wire signal_3891 ;
    wire signal_3892 ;
    wire signal_3893 ;
    wire signal_3894 ;
    wire signal_3895 ;
    wire signal_3896 ;
    wire signal_3897 ;
    wire signal_3898 ;
    wire signal_3899 ;
    wire signal_3900 ;
    wire signal_3901 ;
    wire signal_3902 ;
    wire signal_3903 ;
    wire signal_3904 ;
    wire signal_3905 ;
    wire signal_3906 ;
    wire signal_3907 ;
    wire signal_3908 ;
    wire signal_3909 ;
    wire signal_3910 ;
    wire signal_3911 ;
    wire signal_3912 ;
    wire signal_3913 ;
    wire signal_3914 ;
    wire signal_3915 ;
    wire signal_3916 ;
    wire signal_3917 ;
    wire signal_3918 ;
    wire signal_3919 ;
    wire signal_3920 ;
    wire signal_3921 ;
    wire signal_3922 ;
    wire signal_3923 ;
    wire signal_3924 ;
    wire signal_3925 ;
    wire signal_3926 ;
    wire signal_3927 ;
    wire signal_3928 ;
    wire signal_3929 ;
    wire signal_3930 ;
    wire signal_3931 ;
    wire signal_3932 ;
    wire signal_3933 ;
    wire signal_3934 ;
    wire signal_3935 ;
    wire signal_3936 ;
    wire signal_3937 ;
    wire signal_3938 ;
    wire signal_3939 ;
    wire signal_3940 ;
    wire signal_3941 ;
    wire signal_3942 ;
    wire signal_3943 ;
    wire signal_3944 ;
    wire signal_3945 ;
    wire signal_3946 ;
    wire signal_3947 ;
    wire signal_3948 ;
    wire signal_3949 ;
    wire signal_3950 ;
    wire signal_3951 ;
    wire signal_3952 ;
    wire signal_3953 ;
    wire signal_3954 ;
    wire signal_3955 ;
    wire signal_3956 ;
    wire signal_3957 ;
    wire signal_3958 ;
    wire signal_3959 ;
    wire signal_3960 ;
    wire signal_3961 ;
    wire signal_3962 ;
    wire signal_3963 ;
    wire signal_3964 ;
    wire signal_3965 ;
    wire signal_3966 ;
    wire signal_3967 ;
    wire signal_3968 ;
    wire signal_3969 ;
    wire signal_3970 ;
    wire signal_3971 ;
    wire signal_3972 ;
    wire signal_3973 ;
    wire signal_3974 ;
    wire signal_3975 ;
    wire signal_3976 ;
    wire signal_3977 ;
    wire signal_3978 ;
    wire signal_3979 ;
    wire signal_3980 ;
    wire signal_3981 ;
    wire signal_3982 ;
    wire signal_3983 ;
    wire signal_3984 ;
    wire signal_3985 ;
    wire signal_3986 ;
    wire signal_3987 ;
    wire signal_3988 ;
    wire signal_3989 ;
    wire signal_3990 ;
    wire signal_3991 ;
    wire signal_3992 ;
    wire signal_3993 ;
    wire signal_3994 ;
    wire signal_3995 ;
    wire signal_3996 ;
    wire signal_3997 ;
    wire signal_3998 ;
    wire signal_3999 ;
    wire signal_4000 ;
    wire signal_4001 ;
    wire signal_4002 ;
    wire signal_4003 ;
    wire signal_4004 ;
    wire signal_4005 ;
    wire signal_4006 ;
    wire signal_4007 ;
    wire signal_4008 ;
    wire signal_4009 ;
    wire signal_4010 ;
    wire signal_4011 ;
    wire signal_4012 ;
    wire signal_4013 ;
    wire signal_4014 ;
    wire signal_4015 ;
    wire signal_4016 ;
    wire signal_4017 ;
    wire signal_4018 ;
    wire signal_4019 ;
    wire signal_4020 ;
    wire signal_4021 ;
    wire signal_4022 ;
    wire signal_4023 ;
    wire signal_4024 ;
    wire signal_4025 ;
    wire signal_4026 ;
    wire signal_4027 ;
    wire signal_4028 ;
    wire signal_4029 ;
    wire signal_4030 ;
    wire signal_4031 ;
    wire signal_4032 ;
    wire signal_4033 ;
    wire signal_4034 ;
    wire signal_4035 ;
    wire signal_4036 ;
    wire signal_4037 ;
    wire signal_4038 ;
    wire signal_4039 ;
    wire signal_4040 ;
    wire signal_4041 ;
    wire signal_4042 ;
    wire signal_4043 ;
    wire signal_4044 ;
    wire signal_4045 ;
    wire signal_4046 ;
    wire signal_4047 ;
    wire signal_4048 ;
    wire signal_4049 ;
    wire signal_4050 ;
    wire signal_4051 ;
    wire signal_4052 ;
    wire signal_4053 ;
    wire signal_4054 ;
    wire signal_4055 ;
    wire signal_4056 ;
    wire signal_4057 ;
    wire signal_4058 ;
    wire signal_4059 ;
    wire signal_4060 ;
    wire signal_4061 ;
    wire signal_4062 ;
    wire signal_4063 ;
    wire signal_4064 ;
    wire signal_4065 ;
    wire signal_4066 ;
    wire signal_4067 ;
    wire signal_4068 ;
    wire signal_4069 ;
    wire signal_4070 ;
    wire signal_4071 ;
    wire signal_4072 ;
    wire signal_4073 ;
    wire signal_4074 ;
    wire signal_4075 ;
    wire signal_4076 ;
    wire signal_4077 ;
    wire signal_4078 ;
    wire signal_4079 ;
    wire signal_4080 ;
    wire signal_4081 ;
    wire signal_4082 ;
    wire signal_4083 ;
    wire signal_4084 ;
    wire signal_4085 ;
    wire signal_4086 ;
    wire signal_4087 ;
    wire signal_4088 ;
    wire signal_4089 ;
    wire signal_4090 ;
    wire signal_4091 ;
    wire signal_4092 ;
    wire signal_4093 ;
    wire signal_4094 ;
    wire signal_4095 ;
    wire signal_4096 ;
    wire signal_4097 ;
    wire signal_4098 ;
    wire signal_4099 ;
    wire signal_4100 ;
    wire signal_4101 ;
    wire signal_4102 ;
    wire signal_4103 ;
    wire signal_4104 ;
    wire signal_4105 ;
    wire signal_4106 ;
    wire signal_4107 ;
    wire signal_4108 ;
    wire signal_4109 ;
    wire signal_4110 ;
    wire signal_4111 ;
    wire signal_4112 ;
    wire signal_4113 ;
    wire signal_4114 ;
    wire signal_4115 ;
    wire signal_4116 ;
    wire signal_4117 ;
    wire signal_4118 ;
    wire signal_4119 ;
    wire signal_4120 ;
    wire signal_4121 ;
    wire signal_4122 ;
    wire signal_4123 ;
    wire signal_4124 ;
    wire signal_4125 ;
    wire signal_4126 ;
    wire signal_4127 ;
    wire signal_4128 ;
    wire signal_4129 ;
    wire signal_4130 ;
    wire signal_4131 ;
    wire signal_4132 ;
    wire signal_4133 ;
    wire signal_4134 ;
    wire signal_4135 ;
    wire signal_4136 ;
    wire signal_4137 ;
    wire signal_4138 ;
    wire signal_4139 ;
    wire signal_4140 ;
    wire signal_4141 ;
    wire signal_4142 ;
    wire signal_4143 ;
    wire signal_4144 ;
    wire signal_4145 ;
    wire signal_4146 ;
    wire signal_4147 ;
    wire signal_4148 ;
    wire signal_4149 ;
    wire signal_4150 ;
    wire signal_4151 ;
    wire signal_4152 ;
    wire signal_4153 ;
    wire signal_4154 ;
    wire signal_4155 ;
    wire signal_4156 ;
    wire signal_4157 ;
    wire signal_4158 ;
    wire signal_4159 ;
    wire signal_4160 ;
    wire signal_4161 ;
    wire signal_4162 ;
    wire signal_4163 ;
    wire signal_4164 ;
    wire signal_4165 ;
    wire signal_4166 ;
    wire signal_4167 ;
    wire signal_4168 ;
    wire signal_4169 ;
    wire signal_4170 ;
    wire signal_4171 ;
    wire signal_4172 ;
    wire signal_4173 ;
    wire signal_4174 ;
    wire signal_4175 ;
    wire signal_4176 ;
    wire signal_4177 ;
    wire signal_4178 ;
    wire signal_4179 ;
    wire signal_4180 ;
    wire signal_4181 ;
    wire signal_4182 ;
    wire signal_4183 ;
    wire signal_4184 ;
    wire signal_4185 ;
    wire signal_4186 ;
    wire signal_4187 ;
    wire signal_4188 ;
    wire signal_4189 ;
    wire signal_4190 ;
    wire signal_4191 ;
    wire signal_4192 ;
    wire signal_4193 ;
    wire signal_4194 ;
    wire signal_4195 ;
    wire signal_4196 ;
    wire signal_4197 ;
    wire signal_4198 ;
    wire signal_4199 ;
    wire signal_4200 ;
    wire signal_4201 ;
    wire signal_4202 ;
    wire signal_4203 ;
    wire signal_4204 ;
    wire signal_4205 ;
    wire signal_4206 ;
    wire signal_4207 ;
    wire signal_4208 ;
    wire signal_4209 ;
    wire signal_4210 ;
    wire signal_4211 ;
    wire signal_4212 ;
    wire signal_4213 ;
    wire signal_4214 ;
    wire signal_4215 ;
    wire signal_4216 ;
    wire signal_4217 ;
    wire signal_4218 ;
    wire signal_4219 ;
    wire signal_4220 ;
    wire signal_4221 ;
    wire signal_4222 ;
    wire signal_4223 ;
    wire signal_4224 ;
    wire signal_4225 ;
    wire signal_4226 ;
    wire signal_4227 ;
    wire signal_4228 ;
    wire signal_4229 ;
    wire signal_4230 ;
    wire signal_4231 ;
    wire signal_4232 ;
    wire signal_4233 ;
    wire signal_4234 ;
    wire signal_4235 ;
    wire signal_4236 ;
    wire signal_4237 ;
    wire signal_4238 ;
    wire signal_4239 ;
    wire signal_4240 ;
    wire signal_4241 ;
    wire signal_4242 ;
    wire signal_4243 ;
    wire signal_4244 ;
    wire signal_4245 ;
    wire signal_4246 ;
    wire signal_4247 ;
    wire signal_4248 ;
    wire signal_4249 ;
    wire signal_4250 ;
    wire signal_4251 ;
    wire signal_4252 ;
    wire signal_4253 ;
    wire signal_4254 ;
    wire signal_4255 ;
    wire signal_4256 ;
    wire signal_4257 ;
    wire signal_4258 ;
    wire signal_4259 ;
    wire signal_4260 ;
    wire signal_4261 ;
    wire signal_4262 ;
    wire signal_4263 ;
    wire signal_4264 ;
    wire signal_4265 ;
    wire signal_4266 ;
    wire signal_4267 ;
    wire signal_4268 ;
    wire signal_4269 ;
    wire signal_4270 ;
    wire signal_4271 ;
    wire signal_4272 ;
    wire signal_4273 ;
    wire signal_4274 ;
    wire signal_4275 ;
    wire signal_4276 ;
    wire signal_4277 ;
    wire signal_4278 ;
    wire signal_4279 ;
    wire signal_4280 ;
    wire signal_4281 ;
    wire signal_4282 ;
    wire signal_4283 ;
    wire signal_4284 ;
    wire signal_4285 ;
    wire signal_4286 ;
    wire signal_4287 ;
    wire signal_4288 ;
    wire signal_4289 ;
    wire signal_4290 ;
    wire signal_4291 ;
    wire signal_4292 ;
    wire signal_4293 ;
    wire signal_4294 ;
    wire signal_4295 ;
    wire signal_4296 ;
    wire signal_4297 ;
    wire signal_4298 ;
    wire signal_4299 ;
    wire signal_4300 ;
    wire signal_4301 ;
    wire signal_4302 ;
    wire signal_4303 ;
    wire signal_4304 ;
    wire signal_4305 ;
    wire signal_4306 ;
    wire signal_4307 ;
    wire signal_4308 ;
    wire signal_4309 ;
    wire signal_4310 ;
    wire signal_4311 ;
    wire signal_4312 ;
    wire signal_4313 ;
    wire signal_4314 ;
    wire signal_4315 ;
    wire signal_4316 ;
    wire signal_4317 ;
    wire signal_4318 ;
    wire signal_4319 ;
    wire signal_4320 ;
    wire signal_4321 ;
    wire signal_4322 ;
    wire signal_4323 ;
    wire signal_4324 ;
    wire signal_4325 ;
    wire signal_4326 ;
    wire signal_4327 ;
    wire signal_4328 ;
    wire signal_4329 ;
    wire signal_4330 ;
    wire signal_4331 ;
    wire signal_4332 ;
    wire signal_4333 ;
    wire signal_4334 ;
    wire signal_4335 ;
    wire signal_4336 ;
    wire signal_4337 ;
    wire signal_4338 ;
    wire signal_4339 ;
    wire signal_4340 ;
    wire signal_4341 ;
    wire signal_4342 ;
    wire signal_4343 ;
    wire signal_4344 ;
    wire signal_4345 ;
    wire signal_4346 ;
    wire signal_4347 ;
    wire signal_4348 ;
    wire signal_4349 ;
    wire signal_4350 ;
    wire signal_4351 ;
    wire signal_4352 ;
    wire signal_4353 ;
    wire signal_4354 ;
    wire signal_4355 ;
    wire signal_4356 ;
    wire signal_4357 ;
    wire signal_4358 ;
    wire signal_4359 ;
    wire signal_4360 ;
    wire signal_4361 ;
    wire signal_4362 ;
    wire signal_4363 ;
    wire signal_4364 ;
    wire signal_4365 ;
    wire signal_4366 ;
    wire signal_4367 ;
    wire signal_4368 ;
    wire signal_4369 ;
    wire signal_4370 ;
    wire signal_4371 ;
    wire signal_4372 ;
    wire signal_4373 ;
    wire signal_4374 ;
    wire signal_4375 ;
    wire signal_4376 ;
    wire signal_4377 ;
    wire signal_4378 ;
    wire signal_4379 ;
    wire signal_4380 ;
    wire signal_4381 ;
    wire signal_4382 ;
    wire signal_4383 ;
    wire signal_4384 ;
    wire signal_4385 ;
    wire signal_4386 ;
    wire signal_4387 ;
    wire signal_4388 ;
    wire signal_4389 ;
    wire signal_4390 ;
    wire signal_4391 ;
    wire signal_4392 ;
    wire signal_4393 ;
    wire signal_4394 ;
    wire signal_4395 ;
    wire signal_4396 ;
    wire signal_4397 ;
    wire signal_4398 ;
    wire signal_4399 ;
    wire signal_4400 ;
    wire signal_4401 ;
    wire signal_4402 ;
    wire signal_4403 ;
    wire signal_4404 ;
    wire signal_4405 ;
    wire signal_4406 ;
    wire signal_4407 ;
    wire signal_4408 ;
    wire signal_4409 ;
    wire signal_4410 ;
    wire signal_4411 ;
    wire signal_4412 ;
    wire signal_4413 ;
    wire signal_4414 ;
    wire signal_4415 ;
    wire signal_4416 ;
    wire signal_4417 ;
    wire signal_4418 ;
    wire signal_4419 ;
    wire signal_4420 ;
    wire signal_4421 ;
    wire signal_4422 ;
    wire signal_4423 ;
    wire signal_4424 ;
    wire signal_4425 ;
    wire signal_4426 ;
    wire signal_4427 ;
    wire signal_4428 ;
    wire signal_4429 ;
    wire signal_4430 ;
    wire signal_4431 ;
    wire signal_4432 ;
    wire signal_4433 ;
    wire signal_4434 ;
    wire signal_4435 ;
    wire signal_4436 ;
    wire signal_4437 ;
    wire signal_4438 ;
    wire signal_4439 ;
    wire signal_4440 ;
    wire signal_4441 ;
    wire signal_4442 ;
    wire signal_4443 ;
    wire signal_4444 ;
    wire signal_4445 ;
    wire signal_4446 ;
    wire signal_4447 ;
    wire signal_4448 ;
    wire signal_4449 ;
    wire signal_4450 ;
    wire signal_4451 ;
    wire signal_4452 ;
    wire signal_4453 ;
    wire signal_4454 ;
    wire signal_4455 ;
    wire signal_4456 ;
    wire signal_4457 ;
    wire signal_4458 ;
    wire signal_4459 ;
    wire signal_4460 ;
    wire signal_4461 ;
    wire signal_4462 ;
    wire signal_4463 ;
    wire signal_4464 ;
    wire signal_4465 ;
    wire signal_4466 ;
    wire signal_4467 ;
    wire signal_4468 ;
    wire signal_4469 ;
    wire signal_4470 ;
    wire signal_4471 ;
    wire signal_4472 ;
    wire signal_4473 ;
    wire signal_4474 ;
    wire signal_4475 ;
    wire signal_4476 ;
    wire signal_4477 ;
    wire signal_4478 ;
    wire signal_4479 ;
    wire signal_4480 ;
    wire signal_4481 ;
    wire signal_4482 ;
    wire signal_4483 ;
    wire signal_4484 ;
    wire signal_4485 ;
    wire signal_4486 ;
    wire signal_4487 ;
    wire signal_4488 ;
    wire signal_4489 ;
    wire signal_4490 ;
    wire signal_4491 ;
    wire signal_4492 ;
    wire signal_4493 ;
    wire signal_4494 ;
    wire signal_4495 ;
    wire signal_4496 ;
    wire signal_4497 ;
    wire signal_4498 ;
    wire signal_4499 ;
    wire signal_4500 ;
    wire signal_4501 ;
    wire signal_4502 ;
    wire signal_4503 ;
    wire signal_4504 ;
    wire signal_4505 ;
    wire signal_4506 ;
    wire signal_4507 ;
    wire signal_4508 ;
    wire signal_4509 ;
    wire signal_4510 ;
    wire signal_4511 ;
    wire signal_4512 ;
    wire signal_4513 ;
    wire signal_4514 ;
    wire signal_4515 ;
    wire signal_4516 ;
    wire signal_4517 ;
    wire signal_4518 ;
    wire signal_4519 ;
    wire signal_4520 ;
    wire signal_4521 ;
    wire signal_4522 ;
    wire signal_4523 ;
    wire signal_4524 ;
    wire signal_4525 ;
    wire signal_4526 ;
    wire signal_4527 ;
    wire signal_4528 ;
    wire signal_4529 ;
    wire signal_4530 ;
    wire signal_4531 ;
    wire signal_4532 ;
    wire signal_4533 ;
    wire signal_4534 ;
    wire signal_4535 ;
    wire signal_4536 ;
    wire signal_4537 ;
    wire signal_4538 ;
    wire signal_4539 ;
    wire signal_4540 ;
    wire signal_4541 ;
    wire signal_4542 ;
    wire signal_4543 ;
    wire signal_4544 ;
    wire signal_4545 ;
    wire signal_4546 ;
    wire signal_4547 ;
    wire signal_4548 ;
    wire signal_4549 ;
    wire signal_4550 ;
    wire signal_4551 ;
    wire signal_4552 ;
    wire signal_4553 ;
    wire signal_4554 ;
    wire signal_4555 ;
    wire signal_4556 ;
    wire signal_4557 ;
    wire signal_4558 ;
    wire signal_4559 ;
    wire signal_4560 ;
    wire signal_4561 ;
    wire signal_4562 ;
    wire signal_4563 ;
    wire signal_4564 ;
    wire signal_4565 ;
    wire signal_4566 ;
    wire signal_4567 ;
    wire signal_4568 ;
    wire signal_4569 ;
    wire signal_4570 ;
    wire signal_4571 ;
    wire signal_4572 ;
    wire signal_4573 ;
    wire signal_4574 ;
    wire signal_4575 ;
    wire signal_4576 ;
    wire signal_4577 ;
    wire signal_4578 ;
    wire signal_4579 ;
    wire signal_4580 ;
    wire signal_4581 ;
    wire signal_4582 ;
    wire signal_4583 ;
    wire signal_4584 ;
    wire signal_4585 ;
    wire signal_4586 ;
    wire signal_4587 ;
    wire signal_4588 ;
    wire signal_4589 ;
    wire signal_4590 ;
    wire signal_4591 ;
    wire signal_4592 ;
    wire signal_4593 ;
    wire signal_4594 ;
    wire signal_4595 ;
    wire signal_4596 ;
    wire signal_4597 ;
    wire signal_4598 ;
    wire signal_4599 ;
    wire signal_4600 ;
    wire signal_4601 ;
    wire signal_4602 ;
    wire signal_4603 ;
    wire signal_4604 ;
    wire signal_4605 ;
    wire signal_4606 ;
    wire signal_4607 ;
    wire signal_4608 ;
    wire signal_4609 ;
    wire signal_4610 ;
    wire signal_4611 ;
    wire signal_4612 ;
    wire signal_4613 ;
    wire signal_4614 ;
    wire signal_4615 ;
    wire signal_4616 ;
    wire signal_4617 ;
    wire signal_4618 ;
    wire signal_4619 ;
    wire signal_4620 ;
    wire signal_4621 ;
    wire signal_4622 ;
    wire signal_4623 ;
    wire signal_4624 ;
    wire signal_4625 ;
    wire signal_4626 ;
    wire signal_4627 ;
    wire signal_4628 ;
    wire signal_4629 ;
    wire signal_4630 ;
    wire signal_4631 ;
    wire signal_4632 ;
    wire signal_4633 ;
    wire signal_4634 ;
    wire signal_4635 ;
    wire signal_4636 ;
    wire signal_4637 ;
    wire signal_4638 ;
    wire signal_4639 ;
    wire signal_4640 ;
    wire signal_4641 ;
    wire signal_4642 ;
    wire signal_4643 ;
    wire signal_4644 ;
    wire signal_4645 ;
    wire signal_4646 ;
    wire signal_4647 ;
    wire signal_4648 ;
    wire signal_4649 ;
    wire signal_4650 ;
    wire signal_4651 ;
    wire signal_4652 ;
    wire signal_4653 ;
    wire signal_4654 ;
    wire signal_4655 ;
    wire signal_4656 ;
    wire signal_4657 ;
    wire signal_4658 ;
    wire signal_4659 ;
    wire signal_4660 ;
    wire signal_4661 ;
    wire signal_4662 ;
    wire signal_4663 ;
    wire signal_4664 ;
    wire signal_4665 ;
    wire signal_4666 ;
    wire signal_4667 ;
    wire signal_4668 ;
    wire signal_4669 ;
    wire signal_4670 ;
    wire signal_4671 ;
    wire signal_4672 ;
    wire signal_4673 ;
    wire signal_4674 ;
    wire signal_4675 ;
    wire signal_4676 ;
    wire signal_4677 ;
    wire signal_4678 ;
    wire signal_4679 ;
    wire signal_4680 ;
    wire signal_4681 ;
    wire signal_4682 ;
    wire signal_4683 ;
    wire signal_4684 ;
    wire signal_4685 ;
    wire signal_4686 ;
    wire signal_4687 ;
    wire signal_4688 ;
    wire signal_4689 ;
    wire signal_4690 ;
    wire signal_4691 ;
    wire signal_4692 ;
    wire signal_4693 ;
    wire signal_4694 ;
    wire signal_4695 ;
    wire signal_4696 ;
    wire signal_4697 ;
    wire signal_4698 ;
    wire signal_4699 ;
    wire signal_4700 ;
    wire signal_4701 ;
    wire signal_4702 ;
    wire signal_4703 ;
    wire signal_4704 ;
    wire signal_4705 ;
    wire signal_4706 ;
    wire signal_4707 ;
    wire signal_4708 ;
    wire signal_4709 ;
    wire signal_4710 ;
    wire signal_4711 ;
    wire signal_4712 ;
    wire signal_4713 ;
    wire signal_4714 ;
    wire signal_4715 ;
    wire signal_4716 ;
    wire signal_4717 ;
    wire signal_4718 ;
    wire signal_4719 ;
    wire signal_4720 ;
    wire signal_4721 ;
    wire signal_4722 ;
    wire signal_4723 ;
    wire signal_4724 ;
    wire signal_4725 ;
    wire signal_4726 ;
    wire signal_4727 ;
    wire signal_4728 ;
    wire signal_4729 ;
    wire signal_4730 ;
    wire signal_4731 ;

    /* cells in depth 0 */
    NOR2_X1 cell_0 ( .A1 (signal_875), .A2 (signal_878), .ZN (signal_266) ) ;
    NAND2_X1 cell_1 ( .A1 (signal_879), .A2 (signal_266), .ZN (signal_267) ) ;
    NOR2_X1 cell_2 ( .A1 (signal_874), .A2 (signal_267), .ZN (signal_268) ) ;
    NAND2_X1 cell_3 ( .A1 (signal_876), .A2 (signal_268), .ZN (signal_269) ) ;
    NOR2_X1 cell_4 ( .A1 (signal_877), .A2 (signal_269), .ZN (signal_270) ) ;
    NOR2_X1 cell_5 ( .A1 (OUT_done), .A2 (signal_270), .ZN (signal_271) ) ;
    NOR2_X1 cell_6 ( .A1 (IN_reset), .A2 (signal_271), .ZN (signal_265) ) ;
    NAND2_X1 cell_7 ( .A1 (signal_273), .A2 (signal_274), .ZN (signal_272) ) ;
    XNOR2_X1 cell_8 ( .A (signal_304), .B (signal_275), .ZN (signal_274) ) ;
    XOR2_X1 cell_9 ( .A (signal_309), .B (signal_307), .Z (signal_275) ) ;
    NAND2_X1 cell_10 ( .A1 (signal_276), .A2 (signal_277), .ZN (signal_273) ) ;
    NAND2_X1 cell_11 ( .A1 (signal_278), .A2 (signal_279), .ZN (signal_277) ) ;
    NOR2_X1 cell_12 ( .A1 (signal_302), .A2 (signal_289), .ZN (signal_279) ) ;
    NOR2_X1 cell_13 ( .A1 (signal_306), .A2 (signal_309), .ZN (signal_278) ) ;
    NAND2_X1 cell_14 ( .A1 (signal_289), .A2 (signal_280), .ZN (signal_276) ) ;
    AND2_X1 cell_15 ( .A1 (signal_306), .A2 (signal_309), .ZN (signal_280) ) ;
    NAND2_X1 cell_16 ( .A1 (signal_298), .A2 (signal_283), .ZN (signal_282) ) ;
    NOR2_X1 cell_17 ( .A1 (signal_300), .A2 (signal_284), .ZN (signal_283) ) ;
    NAND2_X1 cell_18 ( .A1 (signal_296), .A2 (signal_876), .ZN (signal_284) ) ;
    NAND2_X1 cell_19 ( .A1 (signal_292), .A2 (signal_290), .ZN (signal_281) ) ;
    NOR2_X1 cell_20 ( .A1 (signal_292), .A2 (IN_reset), .ZN (signal_291) ) ;
    NOR2_X1 cell_21 ( .A1 (IN_reset), .A2 (signal_294), .ZN (signal_293) ) ;
    NOR2_X1 cell_22 ( .A1 (IN_reset), .A2 (signal_296), .ZN (signal_295) ) ;
    NOR2_X1 cell_23 ( .A1 (IN_reset), .A2 (signal_298), .ZN (signal_297) ) ;
    NOR2_X1 cell_24 ( .A1 (IN_reset), .A2 (signal_300), .ZN (signal_299) ) ;
    NOR2_X1 cell_25 ( .A1 (signal_289), .A2 (IN_reset), .ZN (signal_303) ) ;
    NOR2_X1 cell_26 ( .A1 (signal_306), .A2 (IN_reset), .ZN (signal_305) ) ;
    NOR2_X1 cell_27 ( .A1 (signal_309), .A2 (IN_reset), .ZN (signal_308) ) ;
    NOR2_X1 cell_28 ( .A1 (signal_288), .A2 (IN_reset), .ZN (signal_310) ) ;
    OR2_X1 cell_29 ( .A1 (signal_288), .A2 (signal_276), .ZN (signal_286) ) ;
    NAND2_X1 cell_30 ( .A1 (signal_272), .A2 (signal_286), .ZN (signal_311) ) ;
    NOR2_X1 cell_31 ( .A1 (signal_281), .A2 (signal_282), .ZN (signal_340) ) ;
    INV_X1 cell_32 ( .A (signal_286), .ZN (signal_285) ) ;
    OR2_X1 cell_33 ( .A1 (IN_reset), .A2 (signal_287), .ZN (signal_301) ) ;
    XNOR2_X1 cell_34 ( .A (signal_292), .B (signal_290), .ZN (signal_287) ) ;
    INV_X1 cell_35 ( .A (signal_340), .ZN (signal_341) ) ;
    INV_X1 cell_36 ( .A (signal_341), .ZN (signal_344) ) ;
    INV_X1 cell_37 ( .A (signal_341), .ZN (signal_342) ) ;
    INV_X1 cell_38 ( .A (signal_341), .ZN (signal_343) ) ;
    INV_X1 cell_167 ( .A (signal_345), .ZN (signal_346) ) ;
    INV_X1 cell_168 ( .A (signal_285), .ZN (signal_345) ) ;
    INV_X1 cell_169 ( .A (signal_345), .ZN (signal_348) ) ;
    INV_X1 cell_170 ( .A (signal_345), .ZN (signal_347) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_171 ( .s (signal_285), .b ({IN_key_s1[64], IN_key_s0[64]}), .a ({IN_key_s1[0], IN_key_s0[0]}), .c ({signal_1658, signal_1135}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_172 ( .s (signal_346), .b ({IN_key_s1[65], IN_key_s0[65]}), .a ({IN_key_s1[1], IN_key_s0[1]}), .c ({signal_1723, signal_1134}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_173 ( .s (signal_346), .b ({IN_key_s1[66], IN_key_s0[66]}), .a ({IN_key_s1[2], IN_key_s0[2]}), .c ({signal_1726, signal_1133}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_174 ( .s (signal_285), .b ({IN_key_s1[67], IN_key_s0[67]}), .a ({IN_key_s1[3], IN_key_s0[3]}), .c ({signal_1661, signal_1132}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_175 ( .s (signal_346), .b ({IN_key_s1[68], IN_key_s0[68]}), .a ({IN_key_s1[4], IN_key_s0[4]}), .c ({signal_1729, signal_1131}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_176 ( .s (signal_346), .b ({IN_key_s1[69], IN_key_s0[69]}), .a ({IN_key_s1[5], IN_key_s0[5]}), .c ({signal_1732, signal_1130}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_177 ( .s (signal_346), .b ({IN_key_s1[70], IN_key_s0[70]}), .a ({IN_key_s1[6], IN_key_s0[6]}), .c ({signal_1735, signal_1129}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_178 ( .s (signal_346), .b ({IN_key_s1[71], IN_key_s0[71]}), .a ({IN_key_s1[7], IN_key_s0[7]}), .c ({signal_1738, signal_1128}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_179 ( .s (signal_346), .b ({IN_key_s1[72], IN_key_s0[72]}), .a ({IN_key_s1[8], IN_key_s0[8]}), .c ({signal_1741, signal_1127}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_180 ( .s (signal_346), .b ({IN_key_s1[73], IN_key_s0[73]}), .a ({IN_key_s1[9], IN_key_s0[9]}), .c ({signal_1744, signal_1126}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_181 ( .s (signal_346), .b ({IN_key_s1[74], IN_key_s0[74]}), .a ({IN_key_s1[10], IN_key_s0[10]}), .c ({signal_1747, signal_1125}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_182 ( .s (signal_346), .b ({IN_key_s1[75], IN_key_s0[75]}), .a ({IN_key_s1[11], IN_key_s0[11]}), .c ({signal_1750, signal_1124}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_183 ( .s (signal_346), .b ({IN_key_s1[76], IN_key_s0[76]}), .a ({IN_key_s1[12], IN_key_s0[12]}), .c ({signal_1753, signal_1123}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_184 ( .s (signal_346), .b ({IN_key_s1[77], IN_key_s0[77]}), .a ({IN_key_s1[13], IN_key_s0[13]}), .c ({signal_1756, signal_1122}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_185 ( .s (signal_346), .b ({IN_key_s1[78], IN_key_s0[78]}), .a ({IN_key_s1[14], IN_key_s0[14]}), .c ({signal_1759, signal_1121}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_186 ( .s (signal_346), .b ({IN_key_s1[79], IN_key_s0[79]}), .a ({IN_key_s1[15], IN_key_s0[15]}), .c ({signal_1762, signal_1120}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_187 ( .s (signal_285), .b ({IN_key_s1[80], IN_key_s0[80]}), .a ({IN_key_s1[16], IN_key_s0[16]}), .c ({signal_1664, signal_1119}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_188 ( .s (signal_347), .b ({IN_key_s1[81], IN_key_s0[81]}), .a ({IN_key_s1[17], IN_key_s0[17]}), .c ({signal_1765, signal_1118}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_189 ( .s (signal_348), .b ({IN_key_s1[82], IN_key_s0[82]}), .a ({IN_key_s1[18], IN_key_s0[18]}), .c ({signal_1768, signal_1117}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_190 ( .s (signal_285), .b ({IN_key_s1[83], IN_key_s0[83]}), .a ({IN_key_s1[19], IN_key_s0[19]}), .c ({signal_1667, signal_1116}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_191 ( .s (signal_346), .b ({IN_key_s1[84], IN_key_s0[84]}), .a ({IN_key_s1[20], IN_key_s0[20]}), .c ({signal_1771, signal_1115}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_192 ( .s (signal_348), .b ({IN_key_s1[85], IN_key_s0[85]}), .a ({IN_key_s1[21], IN_key_s0[21]}), .c ({signal_1774, signal_1114}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_193 ( .s (signal_285), .b ({IN_key_s1[86], IN_key_s0[86]}), .a ({IN_key_s1[22], IN_key_s0[22]}), .c ({signal_1670, signal_1113}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_194 ( .s (signal_348), .b ({IN_key_s1[87], IN_key_s0[87]}), .a ({IN_key_s1[23], IN_key_s0[23]}), .c ({signal_1777, signal_1112}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_195 ( .s (signal_285), .b ({IN_key_s1[88], IN_key_s0[88]}), .a ({IN_key_s1[24], IN_key_s0[24]}), .c ({signal_1673, signal_1111}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_196 ( .s (signal_348), .b ({IN_key_s1[89], IN_key_s0[89]}), .a ({IN_key_s1[25], IN_key_s0[25]}), .c ({signal_1780, signal_1110}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_197 ( .s (signal_285), .b ({IN_key_s1[90], IN_key_s0[90]}), .a ({IN_key_s1[26], IN_key_s0[26]}), .c ({signal_1676, signal_1109}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_198 ( .s (signal_348), .b ({IN_key_s1[91], IN_key_s0[91]}), .a ({IN_key_s1[27], IN_key_s0[27]}), .c ({signal_1783, signal_1108}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_199 ( .s (signal_285), .b ({IN_key_s1[92], IN_key_s0[92]}), .a ({IN_key_s1[28], IN_key_s0[28]}), .c ({signal_1679, signal_1107}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_200 ( .s (signal_347), .b ({IN_key_s1[93], IN_key_s0[93]}), .a ({IN_key_s1[29], IN_key_s0[29]}), .c ({signal_1786, signal_1106}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_201 ( .s (signal_347), .b ({IN_key_s1[94], IN_key_s0[94]}), .a ({IN_key_s1[30], IN_key_s0[30]}), .c ({signal_1789, signal_1105}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_202 ( .s (signal_347), .b ({IN_key_s1[95], IN_key_s0[95]}), .a ({IN_key_s1[31], IN_key_s0[31]}), .c ({signal_1792, signal_1104}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_203 ( .s (signal_285), .b ({IN_key_s1[96], IN_key_s0[96]}), .a ({IN_key_s1[32], IN_key_s0[32]}), .c ({signal_1682, signal_1103}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_204 ( .s (signal_348), .b ({IN_key_s1[97], IN_key_s0[97]}), .a ({IN_key_s1[33], IN_key_s0[33]}), .c ({signal_1795, signal_1102}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_205 ( .s (signal_285), .b ({IN_key_s1[98], IN_key_s0[98]}), .a ({IN_key_s1[34], IN_key_s0[34]}), .c ({signal_1685, signal_1101}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_206 ( .s (signal_285), .b ({IN_key_s1[99], IN_key_s0[99]}), .a ({IN_key_s1[35], IN_key_s0[35]}), .c ({signal_1688, signal_1100}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_207 ( .s (signal_285), .b ({IN_key_s1[100], IN_key_s0[100]}), .a ({IN_key_s1[36], IN_key_s0[36]}), .c ({signal_1691, signal_1099}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_208 ( .s (signal_347), .b ({IN_key_s1[101], IN_key_s0[101]}), .a ({IN_key_s1[37], IN_key_s0[37]}), .c ({signal_1798, signal_1098}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_209 ( .s (signal_347), .b ({IN_key_s1[102], IN_key_s0[102]}), .a ({IN_key_s1[38], IN_key_s0[38]}), .c ({signal_1801, signal_1097}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_210 ( .s (signal_285), .b ({IN_key_s1[103], IN_key_s0[103]}), .a ({IN_key_s1[39], IN_key_s0[39]}), .c ({signal_1694, signal_1096}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_211 ( .s (signal_347), .b ({IN_key_s1[104], IN_key_s0[104]}), .a ({IN_key_s1[40], IN_key_s0[40]}), .c ({signal_1804, signal_1095}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_212 ( .s (signal_347), .b ({IN_key_s1[105], IN_key_s0[105]}), .a ({IN_key_s1[41], IN_key_s0[41]}), .c ({signal_1807, signal_1094}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_213 ( .s (signal_347), .b ({IN_key_s1[106], IN_key_s0[106]}), .a ({IN_key_s1[42], IN_key_s0[42]}), .c ({signal_1810, signal_1093}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_214 ( .s (signal_347), .b ({IN_key_s1[107], IN_key_s0[107]}), .a ({IN_key_s1[43], IN_key_s0[43]}), .c ({signal_1813, signal_1092}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_215 ( .s (signal_347), .b ({IN_key_s1[108], IN_key_s0[108]}), .a ({IN_key_s1[44], IN_key_s0[44]}), .c ({signal_1816, signal_1091}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_216 ( .s (signal_347), .b ({IN_key_s1[109], IN_key_s0[109]}), .a ({IN_key_s1[45], IN_key_s0[45]}), .c ({signal_1819, signal_1090}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_217 ( .s (signal_347), .b ({IN_key_s1[110], IN_key_s0[110]}), .a ({IN_key_s1[46], IN_key_s0[46]}), .c ({signal_1822, signal_1089}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_218 ( .s (signal_347), .b ({IN_key_s1[111], IN_key_s0[111]}), .a ({IN_key_s1[47], IN_key_s0[47]}), .c ({signal_1825, signal_1088}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_219 ( .s (signal_347), .b ({IN_key_s1[112], IN_key_s0[112]}), .a ({IN_key_s1[48], IN_key_s0[48]}), .c ({signal_1828, signal_1087}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_220 ( .s (signal_347), .b ({IN_key_s1[113], IN_key_s0[113]}), .a ({IN_key_s1[49], IN_key_s0[49]}), .c ({signal_1831, signal_1086}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_221 ( .s (signal_347), .b ({IN_key_s1[114], IN_key_s0[114]}), .a ({IN_key_s1[50], IN_key_s0[50]}), .c ({signal_1834, signal_1085}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_222 ( .s (signal_347), .b ({IN_key_s1[115], IN_key_s0[115]}), .a ({IN_key_s1[51], IN_key_s0[51]}), .c ({signal_1837, signal_1084}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_223 ( .s (signal_348), .b ({IN_key_s1[116], IN_key_s0[116]}), .a ({IN_key_s1[52], IN_key_s0[52]}), .c ({signal_1840, signal_1083}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_224 ( .s (signal_348), .b ({IN_key_s1[117], IN_key_s0[117]}), .a ({IN_key_s1[53], IN_key_s0[53]}), .c ({signal_1843, signal_1082}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_225 ( .s (signal_348), .b ({IN_key_s1[118], IN_key_s0[118]}), .a ({IN_key_s1[54], IN_key_s0[54]}), .c ({signal_1846, signal_1081}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_226 ( .s (signal_348), .b ({IN_key_s1[119], IN_key_s0[119]}), .a ({IN_key_s1[55], IN_key_s0[55]}), .c ({signal_1849, signal_1080}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_227 ( .s (signal_348), .b ({IN_key_s1[120], IN_key_s0[120]}), .a ({IN_key_s1[56], IN_key_s0[56]}), .c ({signal_1852, signal_1079}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_228 ( .s (signal_348), .b ({IN_key_s1[121], IN_key_s0[121]}), .a ({IN_key_s1[57], IN_key_s0[57]}), .c ({signal_1855, signal_1078}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_229 ( .s (signal_348), .b ({IN_key_s1[122], IN_key_s0[122]}), .a ({IN_key_s1[58], IN_key_s0[58]}), .c ({signal_1858, signal_1077}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_230 ( .s (signal_348), .b ({IN_key_s1[123], IN_key_s0[123]}), .a ({IN_key_s1[59], IN_key_s0[59]}), .c ({signal_1861, signal_1076}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_231 ( .s (signal_348), .b ({IN_key_s1[124], IN_key_s0[124]}), .a ({IN_key_s1[60], IN_key_s0[60]}), .c ({signal_1864, signal_1075}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_232 ( .s (signal_348), .b ({IN_key_s1[125], IN_key_s0[125]}), .a ({IN_key_s1[61], IN_key_s0[61]}), .c ({signal_1867, signal_1074}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_233 ( .s (signal_348), .b ({IN_key_s1[126], IN_key_s0[126]}), .a ({IN_key_s1[62], IN_key_s0[62]}), .c ({signal_1870, signal_1073}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_234 ( .s (signal_348), .b ({IN_key_s1[127], IN_key_s0[127]}), .a ({IN_key_s1[63], IN_key_s0[63]}), .c ({signal_1873, signal_1072}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_235 ( .a ({OUT_ciphertext_s1[9], OUT_ciphertext_s0[9]}), .b ({signal_1744, signal_1126}), .c ({signal_1882, signal_1062}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_236 ( .a ({OUT_ciphertext_s1[8], OUT_ciphertext_s0[8]}), .b ({signal_1741, signal_1127}), .c ({signal_1884, signal_1063}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_237 ( .a ({OUT_ciphertext_s1[7], OUT_ciphertext_s0[7]}), .b ({signal_1738, signal_1128}), .c ({signal_1886, signal_1064}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_238 ( .a ({OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}), .b ({signal_1735, signal_1129}), .c ({signal_1888, signal_1065}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_239 ( .a ({OUT_ciphertext_s1[63], OUT_ciphertext_s0[63]}), .b ({signal_1873, signal_1072}), .c ({signal_1890, signal_1008}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_240 ( .a ({OUT_ciphertext_s1[62], OUT_ciphertext_s0[62]}), .b ({signal_1870, signal_1073}), .c ({signal_1892, signal_1009}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_241 ( .a ({OUT_ciphertext_s1[61], OUT_ciphertext_s0[61]}), .b ({signal_1867, signal_1074}), .c ({signal_1894, signal_1010}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_242 ( .a ({OUT_ciphertext_s1[60], OUT_ciphertext_s0[60]}), .b ({signal_1864, signal_1075}), .c ({signal_1896, signal_1011}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_243 ( .a ({OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}), .b ({signal_1732, signal_1130}), .c ({signal_1898, signal_1066}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_244 ( .a ({OUT_ciphertext_s1[59], OUT_ciphertext_s0[59]}), .b ({signal_1861, signal_1076}), .c ({signal_1900, signal_1012}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_245 ( .a ({OUT_ciphertext_s1[58], OUT_ciphertext_s0[58]}), .b ({signal_1858, signal_1077}), .c ({signal_1902, signal_1013}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_246 ( .a ({OUT_ciphertext_s1[57], OUT_ciphertext_s0[57]}), .b ({signal_1855, signal_1078}), .c ({signal_1904, signal_1014}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_247 ( .a ({OUT_ciphertext_s1[56], OUT_ciphertext_s0[56]}), .b ({signal_1852, signal_1079}), .c ({signal_1906, signal_1015}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_248 ( .a ({OUT_ciphertext_s1[55], OUT_ciphertext_s0[55]}), .b ({signal_1849, signal_1080}), .c ({signal_1908, signal_1016}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_249 ( .a ({OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}), .b ({signal_1846, signal_1081}), .c ({signal_1910, signal_1017}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_250 ( .a ({OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}), .b ({signal_1843, signal_1082}), .c ({signal_1912, signal_1018}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_251 ( .a ({OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}), .b ({signal_1840, signal_1083}), .c ({signal_1914, signal_1019}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_252 ( .a ({OUT_ciphertext_s1[51], OUT_ciphertext_s0[51]}), .b ({signal_1837, signal_1084}), .c ({signal_1916, signal_1020}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_253 ( .a ({OUT_ciphertext_s1[50], OUT_ciphertext_s0[50]}), .b ({signal_1834, signal_1085}), .c ({signal_1918, signal_1021}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_254 ( .a ({OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}), .b ({signal_1729, signal_1131}), .c ({signal_1920, signal_1067}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_255 ( .a ({OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}), .b ({signal_1831, signal_1086}), .c ({signal_1922, signal_1022}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_256 ( .a ({OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}), .b ({signal_1828, signal_1087}), .c ({signal_1924, signal_1023}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_257 ( .a ({OUT_ciphertext_s1[47], OUT_ciphertext_s0[47]}), .b ({signal_1825, signal_1088}), .c ({signal_1926, signal_1024}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_258 ( .a ({OUT_ciphertext_s1[46], OUT_ciphertext_s0[46]}), .b ({signal_1822, signal_1089}), .c ({signal_1928, signal_1025}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_259 ( .a ({OUT_ciphertext_s1[45], OUT_ciphertext_s0[45]}), .b ({signal_1819, signal_1090}), .c ({signal_1930, signal_1026}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_260 ( .a ({OUT_ciphertext_s1[44], OUT_ciphertext_s0[44]}), .b ({signal_1816, signal_1091}), .c ({signal_1932, signal_1027}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_261 ( .a ({OUT_ciphertext_s1[43], OUT_ciphertext_s0[43]}), .b ({signal_1813, signal_1092}), .c ({signal_1934, signal_1028}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_262 ( .a ({OUT_ciphertext_s1[42], OUT_ciphertext_s0[42]}), .b ({signal_1810, signal_1093}), .c ({signal_1936, signal_1029}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_263 ( .a ({OUT_ciphertext_s1[41], OUT_ciphertext_s0[41]}), .b ({signal_1807, signal_1094}), .c ({signal_1938, signal_1030}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_264 ( .a ({OUT_ciphertext_s1[40], OUT_ciphertext_s0[40]}), .b ({signal_1804, signal_1095}), .c ({signal_1940, signal_1031}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_265 ( .a ({OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}), .b ({signal_1661, signal_1132}), .c ({signal_1696, signal_1068}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_266 ( .a ({OUT_ciphertext_s1[39], OUT_ciphertext_s0[39]}), .b ({signal_1694, signal_1096}), .c ({signal_1698, signal_1032}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_267 ( .a ({OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}), .b ({signal_1801, signal_1097}), .c ({signal_1942, signal_1033}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_268 ( .a ({OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}), .b ({signal_1798, signal_1098}), .c ({signal_1944, signal_1034}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_269 ( .a ({OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}), .b ({signal_1691, signal_1099}), .c ({signal_1700, signal_1035}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_270 ( .a ({OUT_ciphertext_s1[35], OUT_ciphertext_s0[35]}), .b ({signal_1688, signal_1100}), .c ({signal_1702, signal_1036}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_271 ( .a ({OUT_ciphertext_s1[34], OUT_ciphertext_s0[34]}), .b ({signal_1685, signal_1101}), .c ({signal_1704, signal_1037}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_272 ( .a ({OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}), .b ({signal_1795, signal_1102}), .c ({signal_1946, signal_1038}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_273 ( .a ({OUT_ciphertext_s1[32], OUT_ciphertext_s0[32]}), .b ({signal_1682, signal_1103}), .c ({signal_1706, signal_1039}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_274 ( .a ({OUT_ciphertext_s1[31], OUT_ciphertext_s0[31]}), .b ({signal_1792, signal_1104}), .c ({signal_1948, signal_1040}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_275 ( .a ({OUT_ciphertext_s1[30], OUT_ciphertext_s0[30]}), .b ({signal_1789, signal_1105}), .c ({signal_1950, signal_1041}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_276 ( .a ({OUT_ciphertext_s1[2], OUT_ciphertext_s0[2]}), .b ({signal_1726, signal_1133}), .c ({signal_1952, signal_1069}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_277 ( .a ({OUT_ciphertext_s1[29], OUT_ciphertext_s0[29]}), .b ({signal_1786, signal_1106}), .c ({signal_1954, signal_1042}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_278 ( .a ({OUT_ciphertext_s1[28], OUT_ciphertext_s0[28]}), .b ({signal_1679, signal_1107}), .c ({signal_1708, signal_1043}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_279 ( .a ({OUT_ciphertext_s1[27], OUT_ciphertext_s0[27]}), .b ({signal_1783, signal_1108}), .c ({signal_1956, signal_1044}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_280 ( .a ({OUT_ciphertext_s1[26], OUT_ciphertext_s0[26]}), .b ({signal_1676, signal_1109}), .c ({signal_1710, signal_1045}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_281 ( .a ({OUT_ciphertext_s1[25], OUT_ciphertext_s0[25]}), .b ({signal_1780, signal_1110}), .c ({signal_1958, signal_1046}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_282 ( .a ({OUT_ciphertext_s1[24], OUT_ciphertext_s0[24]}), .b ({signal_1673, signal_1111}), .c ({signal_1712, signal_1047}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_283 ( .a ({OUT_ciphertext_s1[23], OUT_ciphertext_s0[23]}), .b ({signal_1777, signal_1112}), .c ({signal_1960, signal_1048}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_284 ( .a ({OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}), .b ({signal_1670, signal_1113}), .c ({signal_1714, signal_1049}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_285 ( .a ({OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}), .b ({signal_1774, signal_1114}), .c ({signal_1962, signal_1050}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_286 ( .a ({OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}), .b ({signal_1771, signal_1115}), .c ({signal_1964, signal_1051}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_287 ( .a ({OUT_ciphertext_s1[1], OUT_ciphertext_s0[1]}), .b ({signal_1723, signal_1134}), .c ({signal_1966, signal_1070}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_288 ( .a ({OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}), .b ({signal_1667, signal_1116}), .c ({signal_1716, signal_1052}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_289 ( .a ({OUT_ciphertext_s1[18], OUT_ciphertext_s0[18]}), .b ({signal_1768, signal_1117}), .c ({signal_1968, signal_1053}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_290 ( .a ({OUT_ciphertext_s1[17], OUT_ciphertext_s0[17]}), .b ({signal_1765, signal_1118}), .c ({signal_1970, signal_1054}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_291 ( .a ({OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}), .b ({signal_1664, signal_1119}), .c ({signal_1718, signal_1055}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_292 ( .a ({OUT_ciphertext_s1[15], OUT_ciphertext_s0[15]}), .b ({signal_1762, signal_1120}), .c ({signal_1972, signal_1056}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_293 ( .a ({OUT_ciphertext_s1[14], OUT_ciphertext_s0[14]}), .b ({signal_1759, signal_1121}), .c ({signal_1974, signal_1057}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_294 ( .a ({OUT_ciphertext_s1[13], OUT_ciphertext_s0[13]}), .b ({signal_1756, signal_1122}), .c ({signal_1976, signal_1058}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_295 ( .a ({OUT_ciphertext_s1[12], OUT_ciphertext_s0[12]}), .b ({signal_1753, signal_1123}), .c ({signal_1978, signal_1059}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_296 ( .a ({OUT_ciphertext_s1[11], OUT_ciphertext_s0[11]}), .b ({signal_1750, signal_1124}), .c ({signal_1980, signal_1060}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_297 ( .a ({OUT_ciphertext_s1[10], OUT_ciphertext_s0[10]}), .b ({signal_1747, signal_1125}), .c ({signal_1982, signal_1061}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_298 ( .a ({OUT_ciphertext_s1[0], OUT_ciphertext_s0[0]}), .b ({signal_1658, signal_1135}), .c ({signal_1720, signal_1071}) ) ;
    INV_X1 cell_299 ( .A (signal_349), .ZN (signal_351) ) ;
    INV_X1 cell_300 ( .A (signal_311), .ZN (signal_349) ) ;
    INV_X1 cell_301 ( .A (signal_349), .ZN (signal_350) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_302 ( .s (signal_311), .b ({OUT_ciphertext_s1[0], OUT_ciphertext_s0[0]}), .a ({signal_1720, signal_1071}), .c ({signal_1874, signal_312}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_303 ( .s (signal_311), .b ({OUT_ciphertext_s1[1], OUT_ciphertext_s0[1]}), .a ({signal_1966, signal_1070}), .c ({signal_1994, signal_313}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_304 ( .s (signal_311), .b ({OUT_ciphertext_s1[2], OUT_ciphertext_s0[2]}), .a ({signal_1952, signal_1069}), .c ({signal_1995, signal_314}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_305 ( .s (signal_311), .b ({OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}), .a ({signal_1696, signal_1068}), .c ({signal_1875, signal_315}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_306 ( .s (signal_350), .b ({OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}), .a ({signal_1920, signal_1067}), .c ({signal_1996, signal_316}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_307 ( .s (signal_350), .b ({OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}), .a ({signal_1898, signal_1066}), .c ({signal_1997, signal_317}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_308 ( .s (signal_350), .b ({OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}), .a ({signal_1888, signal_1065}), .c ({signal_1998, signal_318}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_309 ( .s (signal_350), .b ({OUT_ciphertext_s1[7], OUT_ciphertext_s0[7]}), .a ({signal_1886, signal_1064}), .c ({signal_1999, signal_1000}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_310 ( .s (signal_350), .b ({OUT_ciphertext_s1[8], OUT_ciphertext_s0[8]}), .a ({signal_1884, signal_1063}), .c ({signal_2000, signal_999}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_311 ( .s (signal_350), .b ({OUT_ciphertext_s1[9], OUT_ciphertext_s0[9]}), .a ({signal_1882, signal_1062}), .c ({signal_2001, signal_998}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_312 ( .s (signal_350), .b ({OUT_ciphertext_s1[10], OUT_ciphertext_s0[10]}), .a ({signal_1982, signal_1061}), .c ({signal_2002, signal_997}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_313 ( .s (signal_350), .b ({OUT_ciphertext_s1[11], OUT_ciphertext_s0[11]}), .a ({signal_1980, signal_1060}), .c ({signal_2003, signal_996}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_314 ( .s (signal_350), .b ({OUT_ciphertext_s1[12], OUT_ciphertext_s0[12]}), .a ({signal_1978, signal_1059}), .c ({signal_2004, signal_995}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_315 ( .s (signal_350), .b ({OUT_ciphertext_s1[13], OUT_ciphertext_s0[13]}), .a ({signal_1976, signal_1058}), .c ({signal_2005, signal_994}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_316 ( .s (signal_350), .b ({OUT_ciphertext_s1[14], OUT_ciphertext_s0[14]}), .a ({signal_1974, signal_1057}), .c ({signal_2006, signal_993}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_317 ( .s (signal_350), .b ({OUT_ciphertext_s1[15], OUT_ciphertext_s0[15]}), .a ({signal_1972, signal_1056}), .c ({signal_2007, signal_992}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_318 ( .s (signal_311), .b ({OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}), .a ({signal_1718, signal_1055}), .c ({signal_1876, signal_319}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_319 ( .s (signal_311), .b ({OUT_ciphertext_s1[17], OUT_ciphertext_s0[17]}), .a ({signal_1970, signal_1054}), .c ({signal_2008, signal_320}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_320 ( .s (signal_311), .b ({OUT_ciphertext_s1[18], OUT_ciphertext_s0[18]}), .a ({signal_1968, signal_1053}), .c ({signal_2009, signal_321}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_321 ( .s (signal_311), .b ({OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}), .a ({signal_1716, signal_1052}), .c ({signal_1877, signal_322}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_322 ( .s (signal_350), .b ({OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}), .a ({signal_1964, signal_1051}), .c ({signal_2010, signal_323}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_323 ( .s (signal_311), .b ({OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}), .a ({signal_1962, signal_1050}), .c ({signal_2011, signal_324}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_324 ( .s (signal_311), .b ({OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}), .a ({signal_1714, signal_1049}), .c ({signal_1878, signal_325}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_325 ( .s (signal_311), .b ({OUT_ciphertext_s1[23], OUT_ciphertext_s0[23]}), .a ({signal_1960, signal_1048}), .c ({signal_2012, signal_984}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_326 ( .s (signal_311), .b ({OUT_ciphertext_s1[24], OUT_ciphertext_s0[24]}), .a ({signal_1712, signal_1047}), .c ({signal_1879, signal_983}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_327 ( .s (signal_311), .b ({OUT_ciphertext_s1[25], OUT_ciphertext_s0[25]}), .a ({signal_1958, signal_1046}), .c ({signal_2013, signal_982}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_328 ( .s (signal_311), .b ({OUT_ciphertext_s1[26], OUT_ciphertext_s0[26]}), .a ({signal_1710, signal_1045}), .c ({signal_1880, signal_981}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_329 ( .s (signal_311), .b ({OUT_ciphertext_s1[27], OUT_ciphertext_s0[27]}), .a ({signal_1956, signal_1044}), .c ({signal_2014, signal_980}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_330 ( .s (signal_351), .b ({OUT_ciphertext_s1[28], OUT_ciphertext_s0[28]}), .a ({signal_1708, signal_1043}), .c ({signal_1983, signal_979}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_331 ( .s (signal_351), .b ({OUT_ciphertext_s1[29], OUT_ciphertext_s0[29]}), .a ({signal_1954, signal_1042}), .c ({signal_2015, signal_978}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_332 ( .s (signal_351), .b ({OUT_ciphertext_s1[30], OUT_ciphertext_s0[30]}), .a ({signal_1950, signal_1041}), .c ({signal_2016, signal_977}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_333 ( .s (signal_351), .b ({OUT_ciphertext_s1[31], OUT_ciphertext_s0[31]}), .a ({signal_1948, signal_1040}), .c ({signal_2017, signal_976}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_334 ( .s (signal_351), .b ({OUT_ciphertext_s1[32], OUT_ciphertext_s0[32]}), .a ({signal_1706, signal_1039}), .c ({signal_1984, signal_326}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_335 ( .s (signal_351), .b ({OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}), .a ({signal_1946, signal_1038}), .c ({signal_2018, signal_327}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_336 ( .s (signal_351), .b ({OUT_ciphertext_s1[34], OUT_ciphertext_s0[34]}), .a ({signal_1704, signal_1037}), .c ({signal_1985, signal_328}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_337 ( .s (signal_351), .b ({OUT_ciphertext_s1[35], OUT_ciphertext_s0[35]}), .a ({signal_1702, signal_1036}), .c ({signal_1986, signal_329}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_338 ( .s (signal_351), .b ({OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}), .a ({signal_1700, signal_1035}), .c ({signal_1987, signal_330}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_339 ( .s (signal_311), .b ({OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}), .a ({signal_1944, signal_1034}), .c ({signal_2019, signal_331}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_340 ( .s (signal_351), .b ({OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}), .a ({signal_1942, signal_1033}), .c ({signal_2020, signal_332}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_341 ( .s (signal_351), .b ({OUT_ciphertext_s1[39], OUT_ciphertext_s0[39]}), .a ({signal_1698, signal_1032}), .c ({signal_1988, signal_968}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_342 ( .s (signal_351), .b ({OUT_ciphertext_s1[40], OUT_ciphertext_s0[40]}), .a ({signal_1940, signal_1031}), .c ({signal_2021, signal_967}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_343 ( .s (signal_351), .b ({OUT_ciphertext_s1[41], OUT_ciphertext_s0[41]}), .a ({signal_1938, signal_1030}), .c ({signal_2022, signal_966}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_344 ( .s (signal_351), .b ({OUT_ciphertext_s1[42], OUT_ciphertext_s0[42]}), .a ({signal_1936, signal_1029}), .c ({signal_2023, signal_965}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_345 ( .s (signal_351), .b ({OUT_ciphertext_s1[43], OUT_ciphertext_s0[43]}), .a ({signal_1934, signal_1028}), .c ({signal_2024, signal_964}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_346 ( .s (signal_351), .b ({OUT_ciphertext_s1[44], OUT_ciphertext_s0[44]}), .a ({signal_1932, signal_1027}), .c ({signal_2025, signal_963}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_347 ( .s (signal_351), .b ({OUT_ciphertext_s1[45], OUT_ciphertext_s0[45]}), .a ({signal_1930, signal_1026}), .c ({signal_2026, signal_962}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_348 ( .s (signal_351), .b ({OUT_ciphertext_s1[46], OUT_ciphertext_s0[46]}), .a ({signal_1928, signal_1025}), .c ({signal_2027, signal_961}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_349 ( .s (signal_351), .b ({OUT_ciphertext_s1[47], OUT_ciphertext_s0[47]}), .a ({signal_1926, signal_1024}), .c ({signal_2028, signal_960}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_350 ( .s (signal_351), .b ({OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}), .a ({signal_1924, signal_1023}), .c ({signal_2029, signal_333}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_351 ( .s (signal_351), .b ({OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}), .a ({signal_1922, signal_1022}), .c ({signal_2030, signal_334}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_352 ( .s (signal_311), .b ({OUT_ciphertext_s1[50], OUT_ciphertext_s0[50]}), .a ({signal_1918, signal_1021}), .c ({signal_2031, signal_335}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_353 ( .s (signal_351), .b ({OUT_ciphertext_s1[51], OUT_ciphertext_s0[51]}), .a ({signal_1916, signal_1020}), .c ({signal_2032, signal_336}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_354 ( .s (signal_351), .b ({OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}), .a ({signal_1914, signal_1019}), .c ({signal_2033, signal_337}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_355 ( .s (signal_351), .b ({OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}), .a ({signal_1912, signal_1018}), .c ({signal_2034, signal_338}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_356 ( .s (signal_351), .b ({OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}), .a ({signal_1910, signal_1017}), .c ({signal_2035, signal_339}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_357 ( .s (signal_351), .b ({OUT_ciphertext_s1[55], OUT_ciphertext_s0[55]}), .a ({signal_1908, signal_1016}), .c ({signal_2036, signal_952}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_358 ( .s (signal_351), .b ({OUT_ciphertext_s1[56], OUT_ciphertext_s0[56]}), .a ({signal_1906, signal_1015}), .c ({signal_2037, signal_951}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_359 ( .s (signal_351), .b ({OUT_ciphertext_s1[57], OUT_ciphertext_s0[57]}), .a ({signal_1904, signal_1014}), .c ({signal_2038, signal_950}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_360 ( .s (signal_351), .b ({OUT_ciphertext_s1[58], OUT_ciphertext_s0[58]}), .a ({signal_1902, signal_1013}), .c ({signal_2039, signal_949}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_361 ( .s (signal_351), .b ({OUT_ciphertext_s1[59], OUT_ciphertext_s0[59]}), .a ({signal_1900, signal_1012}), .c ({signal_2040, signal_948}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_362 ( .s (signal_351), .b ({OUT_ciphertext_s1[60], OUT_ciphertext_s0[60]}), .a ({signal_1896, signal_1011}), .c ({signal_2041, signal_947}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_363 ( .s (signal_351), .b ({OUT_ciphertext_s1[61], OUT_ciphertext_s0[61]}), .a ({signal_1894, signal_1010}), .c ({signal_2042, signal_946}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_364 ( .s (signal_351), .b ({OUT_ciphertext_s1[62], OUT_ciphertext_s0[62]}), .a ({signal_1892, signal_1009}), .c ({signal_2043, signal_945}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_365 ( .s (signal_351), .b ({OUT_ciphertext_s1[63], OUT_ciphertext_s0[63]}), .a ({signal_1890, signal_1008}), .c ({signal_2044, signal_944}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_366 ( .a ({1'b0, signal_874}), .b ({signal_1998, signal_318}), .c ({signal_2054, signal_1001}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_367 ( .a ({1'b0, signal_875}), .b ({signal_1997, signal_317}), .c ({signal_2055, signal_1002}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_368 ( .a ({1'b0, signal_877}), .b ({signal_2035, signal_339}), .c ({signal_2056, signal_953}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_369 ( .a ({1'b0, signal_878}), .b ({signal_2034, signal_338}), .c ({signal_2057, signal_954}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_370 ( .a ({1'b0, signal_879}), .b ({signal_2033, signal_337}), .c ({signal_2058, signal_955}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_371 ( .a ({1'b0, 1'b0}), .b ({signal_2032, signal_336}), .c ({signal_2059, signal_956}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_372 ( .a ({1'b0, 1'b0}), .b ({signal_2031, signal_335}), .c ({signal_2060, signal_957}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_373 ( .a ({1'b0, signal_876}), .b ({signal_1996, signal_316}), .c ({signal_2061, signal_1003}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_374 ( .a ({1'b0, 1'b0}), .b ({signal_2030, signal_334}), .c ({signal_2062, signal_958}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_375 ( .a ({1'b0, 1'b0}), .b ({signal_2029, signal_333}), .c ({signal_2063, signal_959}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_376 ( .a ({1'b0, 1'b1}), .b ({signal_1875, signal_315}), .c ({signal_1989, signal_1004}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_377 ( .a ({1'b0, signal_874}), .b ({signal_2020, signal_332}), .c ({signal_2064, signal_969}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_378 ( .a ({1'b0, signal_875}), .b ({signal_2019, signal_331}), .c ({signal_2065, signal_970}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_379 ( .a ({1'b0, signal_876}), .b ({signal_1987, signal_330}), .c ({signal_2045, signal_971}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_380 ( .a ({1'b0, 1'b0}), .b ({signal_1986, signal_329}), .c ({signal_2046, signal_972}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_381 ( .a ({1'b0, 1'b0}), .b ({signal_1985, signal_328}), .c ({signal_2047, signal_973}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_382 ( .a ({1'b0, 1'b0}), .b ({signal_2018, signal_327}), .c ({signal_2066, signal_974}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_383 ( .a ({1'b0, 1'b0}), .b ({signal_1984, signal_326}), .c ({signal_2048, signal_975}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_384 ( .a ({1'b0, 1'b0}), .b ({signal_1995, signal_314}), .c ({signal_2067, signal_1005}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_385 ( .a ({1'b0, signal_877}), .b ({signal_1878, signal_325}), .c ({signal_1990, signal_985}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_386 ( .a ({1'b0, signal_878}), .b ({signal_2011, signal_324}), .c ({signal_2068, signal_986}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_387 ( .a ({1'b0, signal_879}), .b ({signal_2010, signal_323}), .c ({signal_2069, signal_987}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_388 ( .a ({1'b0, 1'b0}), .b ({signal_1994, signal_313}), .c ({signal_2070, signal_1006}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_389 ( .a ({1'b0, 1'b1}), .b ({signal_1877, signal_322}), .c ({signal_1991, signal_988}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_390 ( .a ({1'b0, 1'b0}), .b ({signal_2009, signal_321}), .c ({signal_2071, signal_989}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_391 ( .a ({1'b0, 1'b0}), .b ({signal_2008, signal_320}), .c ({signal_2072, signal_990}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_392 ( .a ({1'b0, 1'b0}), .b ({signal_1876, signal_319}), .c ({signal_1992, signal_991}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_393 ( .a ({1'b0, 1'b0}), .b ({signal_1874, signal_312}), .c ({signal_1993, signal_1007}) ) ;
    INV_X1 cell_978 ( .A (signal_808), .ZN (signal_309) ) ;
    INV_X1 cell_980 ( .A (signal_307), .ZN (signal_306) ) ;
    INV_X1 cell_982 ( .A (signal_304), .ZN (signal_289) ) ;
    INV_X1 cell_984 ( .A (signal_288), .ZN (signal_302) ) ;
    INV_X1 cell_986 ( .A (signal_879), .ZN (signal_300) ) ;
    INV_X1 cell_988 ( .A (signal_878), .ZN (signal_298) ) ;
    INV_X1 cell_990 ( .A (signal_877), .ZN (signal_296) ) ;
    INV_X1 cell_992 ( .A (signal_876), .ZN (signal_294) ) ;
    INV_X1 cell_994 ( .A (signal_875), .ZN (signal_292) ) ;
    INV_X1 cell_996 ( .A (signal_874), .ZN (signal_290) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1128 ( .a ({signal_1988, signal_968}), .b ({signal_2049, signal_1328}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1129 ( .a ({signal_1989, signal_1004}), .b ({signal_2050, signal_1329}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1130 ( .a ({signal_1991, signal_988}), .b ({signal_2051, signal_1330}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1131 ( .a ({signal_1999, signal_1000}), .b ({signal_2073, signal_1331}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1132 ( .a ({signal_2001, signal_998}), .b ({signal_2074, signal_1332}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1133 ( .a ({signal_2003, signal_996}), .b ({signal_2075, signal_1333}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1134 ( .a ({signal_2005, signal_994}), .b ({signal_2076, signal_1334}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1135 ( .a ({signal_2007, signal_992}), .b ({signal_2077, signal_1335}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1136 ( .a ({signal_2012, signal_984}), .b ({signal_2078, signal_1336}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1137 ( .a ({signal_2013, signal_982}), .b ({signal_2079, signal_1337}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1138 ( .a ({signal_2014, signal_980}), .b ({signal_2080, signal_1338}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1139 ( .a ({signal_2015, signal_978}), .b ({signal_2081, signal_1339}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1140 ( .a ({signal_2017, signal_976}), .b ({signal_2082, signal_1340}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1141 ( .a ({signal_2022, signal_966}), .b ({signal_2083, signal_1341}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1142 ( .a ({signal_2024, signal_964}), .b ({signal_2084, signal_1342}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1143 ( .a ({signal_2026, signal_962}), .b ({signal_2085, signal_1343}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1144 ( .a ({signal_2028, signal_960}), .b ({signal_2086, signal_1344}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1145 ( .a ({signal_2036, signal_952}), .b ({signal_2087, signal_1345}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1146 ( .a ({signal_2038, signal_950}), .b ({signal_2088, signal_1346}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1147 ( .a ({signal_2040, signal_948}), .b ({signal_2089, signal_1347}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1148 ( .a ({signal_2042, signal_946}), .b ({signal_2090, signal_1348}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1149 ( .a ({signal_2044, signal_944}), .b ({signal_2091, signal_1349}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1150 ( .a ({signal_2046, signal_972}), .b ({signal_2092, signal_1350}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1151 ( .a ({signal_2055, signal_1002}), .b ({signal_2127, signal_1351}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1152 ( .a ({signal_2057, signal_954}), .b ({signal_2128, signal_1352}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1153 ( .a ({signal_2059, signal_956}), .b ({signal_2129, signal_1353}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1154 ( .a ({signal_2062, signal_958}), .b ({signal_2130, signal_1354}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1155 ( .a ({signal_2065, signal_970}), .b ({signal_2131, signal_1355}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1156 ( .a ({signal_2066, signal_974}), .b ({signal_2132, signal_1356}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1157 ( .a ({signal_2068, signal_986}), .b ({signal_2133, signal_1357}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1158 ( .a ({signal_2070, signal_1006}), .b ({signal_2134, signal_1358}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1159 ( .a ({signal_2072, signal_990}), .b ({signal_2135, signal_1359}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1160 ( .a ({signal_2067, signal_1005}), .b ({signal_2070, signal_1006}), .c ({signal_2136, signal_1360}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1161 ( .a ({signal_1993, signal_1007}), .b ({signal_2070, signal_1006}), .c ({signal_2137, signal_1361}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1162 ( .a ({signal_1989, signal_1004}), .b ({signal_1993, signal_1007}), .c ({signal_2052, signal_1362}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1163 ( .a ({signal_1989, signal_1004}), .b ({signal_2070, signal_1006}), .c ({signal_2138, signal_1363}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1164 ( .a ({signal_2054, signal_1001}), .b ({signal_2055, signal_1002}), .c ({signal_2139, signal_1364}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1165 ( .a ({signal_2055, signal_1002}), .b ({signal_2061, signal_1003}), .c ({signal_2140, signal_1365}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1166 ( .a ({signal_1999, signal_1000}), .b ({signal_2061, signal_1003}), .c ({signal_2141, signal_1366}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1167 ( .a ({signal_1999, signal_1000}), .b ({signal_2055, signal_1002}), .c ({signal_2142, signal_1367}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1168 ( .a ({signal_2001, signal_998}), .b ({signal_2002, signal_997}), .c ({signal_2093, signal_1368}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1169 ( .a ({signal_2000, signal_999}), .b ({signal_2001, signal_998}), .c ({signal_2094, signal_1369}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1170 ( .a ({signal_2000, signal_999}), .b ({signal_2003, signal_996}), .c ({signal_2095, signal_1370}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1171 ( .a ({signal_2001, signal_998}), .b ({signal_2003, signal_996}), .c ({signal_2096, signal_1371}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1172 ( .a ({signal_2005, signal_994}), .b ({signal_2006, signal_993}), .c ({signal_2097, signal_1372}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1173 ( .a ({signal_2004, signal_995}), .b ({signal_2005, signal_994}), .c ({signal_2098, signal_1373}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1174 ( .a ({signal_2004, signal_995}), .b ({signal_2007, signal_992}), .c ({signal_2099, signal_1374}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1175 ( .a ({signal_2005, signal_994}), .b ({signal_2007, signal_992}), .c ({signal_2100, signal_1375}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1176 ( .a ({signal_2071, signal_989}), .b ({signal_2072, signal_990}), .c ({signal_2143, signal_1376}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1177 ( .a ({signal_1992, signal_991}), .b ({signal_2072, signal_990}), .c ({signal_2144, signal_1377}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1178 ( .a ({signal_1991, signal_988}), .b ({signal_1992, signal_991}), .c ({signal_2053, signal_1378}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1179 ( .a ({signal_1991, signal_988}), .b ({signal_2072, signal_990}), .c ({signal_2145, signal_1379}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1180 ( .a ({signal_1990, signal_985}), .b ({signal_2068, signal_986}), .c ({signal_2146, signal_1380}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1181 ( .a ({signal_2068, signal_986}), .b ({signal_2069, signal_987}), .c ({signal_2147, signal_1381}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1182 ( .a ({signal_2012, signal_984}), .b ({signal_2069, signal_987}), .c ({signal_2148, signal_1382}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1183 ( .a ({signal_2012, signal_984}), .b ({signal_2068, signal_986}), .c ({signal_2149, signal_1383}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1184 ( .a ({signal_1880, signal_981}), .b ({signal_2013, signal_982}), .c ({signal_2101, signal_1384}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1185 ( .a ({signal_1879, signal_983}), .b ({signal_2013, signal_982}), .c ({signal_2102, signal_1385}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1186 ( .a ({signal_1879, signal_983}), .b ({signal_2014, signal_980}), .c ({signal_2103, signal_1386}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1187 ( .a ({signal_2013, signal_982}), .b ({signal_2014, signal_980}), .c ({signal_2104, signal_1387}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1188 ( .a ({signal_2015, signal_978}), .b ({signal_2016, signal_977}), .c ({signal_2105, signal_1388}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1189 ( .a ({signal_1983, signal_979}), .b ({signal_2015, signal_978}), .c ({signal_2106, signal_1389}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1190 ( .a ({signal_1983, signal_979}), .b ({signal_2017, signal_976}), .c ({signal_2107, signal_1390}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1191 ( .a ({signal_2015, signal_978}), .b ({signal_2017, signal_976}), .c ({signal_2108, signal_1391}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1192 ( .a ({signal_2047, signal_973}), .b ({signal_2066, signal_974}), .c ({signal_2150, signal_1392}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1193 ( .a ({signal_2048, signal_975}), .b ({signal_2066, signal_974}), .c ({signal_2151, signal_1393}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1194 ( .a ({signal_2046, signal_972}), .b ({signal_2048, signal_975}), .c ({signal_2109, signal_1394}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1195 ( .a ({signal_2046, signal_972}), .b ({signal_2066, signal_974}), .c ({signal_2152, signal_1395}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1196 ( .a ({signal_2064, signal_969}), .b ({signal_2065, signal_970}), .c ({signal_2153, signal_1396}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1197 ( .a ({signal_2045, signal_971}), .b ({signal_2065, signal_970}), .c ({signal_2154, signal_1397}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1198 ( .a ({signal_1988, signal_968}), .b ({signal_2045, signal_971}), .c ({signal_2110, signal_1398}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1199 ( .a ({signal_1988, signal_968}), .b ({signal_2065, signal_970}), .c ({signal_2155, signal_1399}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1200 ( .a ({signal_2022, signal_966}), .b ({signal_2023, signal_965}), .c ({signal_2111, signal_1400}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1201 ( .a ({signal_2021, signal_967}), .b ({signal_2022, signal_966}), .c ({signal_2112, signal_1401}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1202 ( .a ({signal_2021, signal_967}), .b ({signal_2024, signal_964}), .c ({signal_2113, signal_1402}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1203 ( .a ({signal_2022, signal_966}), .b ({signal_2024, signal_964}), .c ({signal_2114, signal_1403}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1204 ( .a ({signal_2026, signal_962}), .b ({signal_2027, signal_961}), .c ({signal_2115, signal_1404}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1205 ( .a ({signal_2025, signal_963}), .b ({signal_2026, signal_962}), .c ({signal_2116, signal_1405}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1206 ( .a ({signal_2025, signal_963}), .b ({signal_2028, signal_960}), .c ({signal_2117, signal_1406}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1207 ( .a ({signal_2026, signal_962}), .b ({signal_2028, signal_960}), .c ({signal_2118, signal_1407}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1208 ( .a ({signal_2060, signal_957}), .b ({signal_2062, signal_958}), .c ({signal_2156, signal_1408}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1209 ( .a ({signal_2062, signal_958}), .b ({signal_2063, signal_959}), .c ({signal_2157, signal_1409}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1210 ( .a ({signal_2059, signal_956}), .b ({signal_2063, signal_959}), .c ({signal_2158, signal_1410}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1211 ( .a ({signal_2059, signal_956}), .b ({signal_2062, signal_958}), .c ({signal_2159, signal_1411}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1212 ( .a ({signal_2056, signal_953}), .b ({signal_2057, signal_954}), .c ({signal_2160, signal_1412}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1213 ( .a ({signal_2057, signal_954}), .b ({signal_2058, signal_955}), .c ({signal_2161, signal_1413}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1214 ( .a ({signal_2036, signal_952}), .b ({signal_2058, signal_955}), .c ({signal_2162, signal_1414}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1215 ( .a ({signal_2036, signal_952}), .b ({signal_2057, signal_954}), .c ({signal_2163, signal_1415}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1216 ( .a ({signal_2038, signal_950}), .b ({signal_2039, signal_949}), .c ({signal_2119, signal_1416}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1217 ( .a ({signal_2037, signal_951}), .b ({signal_2038, signal_950}), .c ({signal_2120, signal_1417}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1218 ( .a ({signal_2037, signal_951}), .b ({signal_2040, signal_948}), .c ({signal_2121, signal_1418}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1219 ( .a ({signal_2038, signal_950}), .b ({signal_2040, signal_948}), .c ({signal_2122, signal_1419}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1220 ( .a ({signal_2042, signal_946}), .b ({signal_2043, signal_945}), .c ({signal_2123, signal_1420}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1221 ( .a ({signal_2041, signal_947}), .b ({signal_2042, signal_946}), .c ({signal_2124, signal_1421}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1222 ( .a ({signal_2041, signal_947}), .b ({signal_2044, signal_944}), .c ({signal_2125, signal_1422}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1223 ( .a ({signal_2042, signal_946}), .b ({signal_2044, signal_944}), .c ({signal_2126, signal_1423}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1224 ( .a ({signal_2136, signal_1360}), .b ({signal_2204, signal_1424}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1225 ( .a ({signal_2139, signal_1364}), .b ({signal_2205, signal_1425}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1226 ( .a ({signal_2093, signal_1368}), .b ({signal_2164, signal_1426}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1227 ( .a ({signal_2097, signal_1372}), .b ({signal_2165, signal_1427}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1228 ( .a ({signal_2143, signal_1376}), .b ({signal_2206, signal_1428}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1229 ( .a ({signal_2146, signal_1380}), .b ({signal_2207, signal_1429}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1230 ( .a ({signal_2101, signal_1384}), .b ({signal_2166, signal_1430}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1231 ( .a ({signal_2105, signal_1388}), .b ({signal_2167, signal_1431}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1232 ( .a ({signal_2150, signal_1392}), .b ({signal_2208, signal_1432}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1233 ( .a ({signal_2153, signal_1396}), .b ({signal_2209, signal_1433}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1234 ( .a ({signal_2111, signal_1400}), .b ({signal_2168, signal_1434}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1235 ( .a ({signal_2115, signal_1404}), .b ({signal_2169, signal_1435}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1236 ( .a ({signal_2156, signal_1408}), .b ({signal_2210, signal_1436}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1237 ( .a ({signal_2160, signal_1412}), .b ({signal_2211, signal_1437}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1238 ( .a ({signal_2119, signal_1416}), .b ({signal_2170, signal_1438}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1239 ( .a ({signal_2123, signal_1420}), .b ({signal_2171, signal_1439}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1256 ( .a ({signal_1989, signal_1004}), .b ({signal_2137, signal_1361}), .c ({signal_2220, signal_1456}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1257 ( .a ({signal_2136, signal_1360}), .b ({signal_2052, signal_1362}), .c ({signal_2221, signal_1457}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1258 ( .a ({signal_2067, signal_1005}), .b ({signal_2137, signal_1361}), .c ({signal_2222, signal_1458}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1259 ( .a ({signal_1999, signal_1000}), .b ({signal_2140, signal_1365}), .c ({signal_2223, signal_1459}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1260 ( .a ({signal_2139, signal_1364}), .b ({signal_2141, signal_1366}), .c ({signal_2224, signal_1460}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1261 ( .a ({signal_2054, signal_1001}), .b ({signal_2140, signal_1365}), .c ({signal_2225, signal_1461}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1262 ( .a ({signal_2003, signal_996}), .b ({signal_2094, signal_1369}), .c ({signal_2180, signal_1462}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1263 ( .a ({signal_2093, signal_1368}), .b ({signal_2095, signal_1370}), .c ({signal_2181, signal_1463}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1264 ( .a ({signal_2002, signal_997}), .b ({signal_2094, signal_1369}), .c ({signal_2182, signal_1464}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1265 ( .a ({signal_2007, signal_992}), .b ({signal_2098, signal_1373}), .c ({signal_2183, signal_1465}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1266 ( .a ({signal_2097, signal_1372}), .b ({signal_2099, signal_1374}), .c ({signal_2184, signal_1466}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1267 ( .a ({signal_2006, signal_993}), .b ({signal_2098, signal_1373}), .c ({signal_2185, signal_1467}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1268 ( .a ({signal_1991, signal_988}), .b ({signal_2144, signal_1377}), .c ({signal_2226, signal_1468}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1269 ( .a ({signal_2143, signal_1376}), .b ({signal_2053, signal_1378}), .c ({signal_2227, signal_1469}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1270 ( .a ({signal_2071, signal_989}), .b ({signal_2144, signal_1377}), .c ({signal_2228, signal_1470}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1271 ( .a ({signal_2012, signal_984}), .b ({signal_2147, signal_1381}), .c ({signal_2229, signal_1471}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1272 ( .a ({signal_2146, signal_1380}), .b ({signal_2148, signal_1382}), .c ({signal_2230, signal_1472}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1273 ( .a ({signal_1990, signal_985}), .b ({signal_2147, signal_1381}), .c ({signal_2231, signal_1473}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1274 ( .a ({signal_2014, signal_980}), .b ({signal_2102, signal_1385}), .c ({signal_2186, signal_1474}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1275 ( .a ({signal_2101, signal_1384}), .b ({signal_2103, signal_1386}), .c ({signal_2187, signal_1475}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1276 ( .a ({signal_1880, signal_981}), .b ({signal_2102, signal_1385}), .c ({signal_2188, signal_1476}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1277 ( .a ({signal_2017, signal_976}), .b ({signal_2106, signal_1389}), .c ({signal_2189, signal_1477}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1278 ( .a ({signal_2105, signal_1388}), .b ({signal_2107, signal_1390}), .c ({signal_2190, signal_1478}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1279 ( .a ({signal_2016, signal_977}), .b ({signal_2106, signal_1389}), .c ({signal_2191, signal_1479}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1280 ( .a ({signal_2046, signal_972}), .b ({signal_2151, signal_1393}), .c ({signal_2232, signal_1480}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1281 ( .a ({signal_2150, signal_1392}), .b ({signal_2109, signal_1394}), .c ({signal_2233, signal_1481}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1282 ( .a ({signal_2047, signal_973}), .b ({signal_2151, signal_1393}), .c ({signal_2234, signal_1482}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1283 ( .a ({signal_1988, signal_968}), .b ({signal_2154, signal_1397}), .c ({signal_2235, signal_1483}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1284 ( .a ({signal_2153, signal_1396}), .b ({signal_2110, signal_1398}), .c ({signal_2236, signal_1484}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1285 ( .a ({signal_2064, signal_969}), .b ({signal_2154, signal_1397}), .c ({signal_2237, signal_1485}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1286 ( .a ({signal_2024, signal_964}), .b ({signal_2112, signal_1401}), .c ({signal_2192, signal_1486}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1287 ( .a ({signal_2111, signal_1400}), .b ({signal_2113, signal_1402}), .c ({signal_2193, signal_1487}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1288 ( .a ({signal_2023, signal_965}), .b ({signal_2112, signal_1401}), .c ({signal_2194, signal_1488}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1289 ( .a ({signal_2028, signal_960}), .b ({signal_2116, signal_1405}), .c ({signal_2195, signal_1489}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1290 ( .a ({signal_2115, signal_1404}), .b ({signal_2117, signal_1406}), .c ({signal_2196, signal_1490}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1291 ( .a ({signal_2027, signal_961}), .b ({signal_2116, signal_1405}), .c ({signal_2197, signal_1491}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1292 ( .a ({signal_2059, signal_956}), .b ({signal_2157, signal_1409}), .c ({signal_2238, signal_1492}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1293 ( .a ({signal_2156, signal_1408}), .b ({signal_2158, signal_1410}), .c ({signal_2239, signal_1493}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1294 ( .a ({signal_2060, signal_957}), .b ({signal_2157, signal_1409}), .c ({signal_2240, signal_1494}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1295 ( .a ({signal_2036, signal_952}), .b ({signal_2161, signal_1413}), .c ({signal_2241, signal_1495}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1296 ( .a ({signal_2160, signal_1412}), .b ({signal_2162, signal_1414}), .c ({signal_2242, signal_1496}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1297 ( .a ({signal_2056, signal_953}), .b ({signal_2161, signal_1413}), .c ({signal_2243, signal_1497}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1298 ( .a ({signal_2040, signal_948}), .b ({signal_2120, signal_1417}), .c ({signal_2198, signal_1498}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1299 ( .a ({signal_2119, signal_1416}), .b ({signal_2121, signal_1418}), .c ({signal_2199, signal_1499}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1300 ( .a ({signal_2039, signal_949}), .b ({signal_2120, signal_1417}), .c ({signal_2200, signal_1500}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1301 ( .a ({signal_2044, signal_944}), .b ({signal_2124, signal_1421}), .c ({signal_2201, signal_1501}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1302 ( .a ({signal_2123, signal_1420}), .b ({signal_2125, signal_1422}), .c ({signal_2202, signal_1502}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1303 ( .a ({signal_2043, signal_945}), .b ({signal_2124, signal_1421}), .c ({signal_2203, signal_1503}) ) ;

    /* cells in depth 1 */
    buf_clk cell_1528 ( .C (CLK), .D (signal_1362), .Q (signal_2940) ) ;
    buf_clk cell_1530 ( .C (CLK), .D (signal_2052), .Q (signal_2942) ) ;
    buf_clk cell_1532 ( .C (CLK), .D (signal_1366), .Q (signal_2944) ) ;
    buf_clk cell_1534 ( .C (CLK), .D (signal_2141), .Q (signal_2946) ) ;
    buf_clk cell_1536 ( .C (CLK), .D (signal_1370), .Q (signal_2948) ) ;
    buf_clk cell_1538 ( .C (CLK), .D (signal_2095), .Q (signal_2950) ) ;
    buf_clk cell_1540 ( .C (CLK), .D (signal_1374), .Q (signal_2952) ) ;
    buf_clk cell_1542 ( .C (CLK), .D (signal_2099), .Q (signal_2954) ) ;
    buf_clk cell_1544 ( .C (CLK), .D (signal_1378), .Q (signal_2956) ) ;
    buf_clk cell_1546 ( .C (CLK), .D (signal_2053), .Q (signal_2958) ) ;
    buf_clk cell_1548 ( .C (CLK), .D (signal_1382), .Q (signal_2960) ) ;
    buf_clk cell_1550 ( .C (CLK), .D (signal_2148), .Q (signal_2962) ) ;
    buf_clk cell_1552 ( .C (CLK), .D (signal_1386), .Q (signal_2964) ) ;
    buf_clk cell_1554 ( .C (CLK), .D (signal_2103), .Q (signal_2966) ) ;
    buf_clk cell_1556 ( .C (CLK), .D (signal_1390), .Q (signal_2968) ) ;
    buf_clk cell_1558 ( .C (CLK), .D (signal_2107), .Q (signal_2970) ) ;
    buf_clk cell_1560 ( .C (CLK), .D (signal_1394), .Q (signal_2972) ) ;
    buf_clk cell_1562 ( .C (CLK), .D (signal_2109), .Q (signal_2974) ) ;
    buf_clk cell_1564 ( .C (CLK), .D (signal_1398), .Q (signal_2976) ) ;
    buf_clk cell_1566 ( .C (CLK), .D (signal_2110), .Q (signal_2978) ) ;
    buf_clk cell_1568 ( .C (CLK), .D (signal_1402), .Q (signal_2980) ) ;
    buf_clk cell_1570 ( .C (CLK), .D (signal_2113), .Q (signal_2982) ) ;
    buf_clk cell_1572 ( .C (CLK), .D (signal_1406), .Q (signal_2984) ) ;
    buf_clk cell_1574 ( .C (CLK), .D (signal_2117), .Q (signal_2986) ) ;
    buf_clk cell_1576 ( .C (CLK), .D (signal_1410), .Q (signal_2988) ) ;
    buf_clk cell_1578 ( .C (CLK), .D (signal_2158), .Q (signal_2990) ) ;
    buf_clk cell_1580 ( .C (CLK), .D (signal_1414), .Q (signal_2992) ) ;
    buf_clk cell_1582 ( .C (CLK), .D (signal_2162), .Q (signal_2994) ) ;
    buf_clk cell_1584 ( .C (CLK), .D (signal_1418), .Q (signal_2996) ) ;
    buf_clk cell_1586 ( .C (CLK), .D (signal_2121), .Q (signal_2998) ) ;
    buf_clk cell_1588 ( .C (CLK), .D (signal_1422), .Q (signal_3000) ) ;
    buf_clk cell_1590 ( .C (CLK), .D (signal_2125), .Q (signal_3002) ) ;
    buf_clk cell_1592 ( .C (CLK), .D (signal_1456), .Q (signal_3004) ) ;
    buf_clk cell_1594 ( .C (CLK), .D (signal_2220), .Q (signal_3006) ) ;
    buf_clk cell_1596 ( .C (CLK), .D (signal_1459), .Q (signal_3008) ) ;
    buf_clk cell_1598 ( .C (CLK), .D (signal_2223), .Q (signal_3010) ) ;
    buf_clk cell_1600 ( .C (CLK), .D (signal_1462), .Q (signal_3012) ) ;
    buf_clk cell_1602 ( .C (CLK), .D (signal_2180), .Q (signal_3014) ) ;
    buf_clk cell_1604 ( .C (CLK), .D (signal_1465), .Q (signal_3016) ) ;
    buf_clk cell_1606 ( .C (CLK), .D (signal_2183), .Q (signal_3018) ) ;
    buf_clk cell_1608 ( .C (CLK), .D (signal_1468), .Q (signal_3020) ) ;
    buf_clk cell_1610 ( .C (CLK), .D (signal_2226), .Q (signal_3022) ) ;
    buf_clk cell_1612 ( .C (CLK), .D (signal_1471), .Q (signal_3024) ) ;
    buf_clk cell_1614 ( .C (CLK), .D (signal_2229), .Q (signal_3026) ) ;
    buf_clk cell_1616 ( .C (CLK), .D (signal_1474), .Q (signal_3028) ) ;
    buf_clk cell_1618 ( .C (CLK), .D (signal_2186), .Q (signal_3030) ) ;
    buf_clk cell_1620 ( .C (CLK), .D (signal_1477), .Q (signal_3032) ) ;
    buf_clk cell_1622 ( .C (CLK), .D (signal_2189), .Q (signal_3034) ) ;
    buf_clk cell_1624 ( .C (CLK), .D (signal_1480), .Q (signal_3036) ) ;
    buf_clk cell_1626 ( .C (CLK), .D (signal_2232), .Q (signal_3038) ) ;
    buf_clk cell_1628 ( .C (CLK), .D (signal_1483), .Q (signal_3040) ) ;
    buf_clk cell_1630 ( .C (CLK), .D (signal_2235), .Q (signal_3042) ) ;
    buf_clk cell_1632 ( .C (CLK), .D (signal_1486), .Q (signal_3044) ) ;
    buf_clk cell_1634 ( .C (CLK), .D (signal_2192), .Q (signal_3046) ) ;
    buf_clk cell_1636 ( .C (CLK), .D (signal_1489), .Q (signal_3048) ) ;
    buf_clk cell_1638 ( .C (CLK), .D (signal_2195), .Q (signal_3050) ) ;
    buf_clk cell_1640 ( .C (CLK), .D (signal_1492), .Q (signal_3052) ) ;
    buf_clk cell_1642 ( .C (CLK), .D (signal_2238), .Q (signal_3054) ) ;
    buf_clk cell_1644 ( .C (CLK), .D (signal_1495), .Q (signal_3056) ) ;
    buf_clk cell_1646 ( .C (CLK), .D (signal_2241), .Q (signal_3058) ) ;
    buf_clk cell_1648 ( .C (CLK), .D (signal_1498), .Q (signal_3060) ) ;
    buf_clk cell_1650 ( .C (CLK), .D (signal_2198), .Q (signal_3062) ) ;
    buf_clk cell_1652 ( .C (CLK), .D (signal_1501), .Q (signal_3064) ) ;
    buf_clk cell_1654 ( .C (CLK), .D (signal_2201), .Q (signal_3066) ) ;
    buf_clk cell_1656 ( .C (CLK), .D (signal_1363), .Q (signal_3068) ) ;
    buf_clk cell_1658 ( .C (CLK), .D (signal_2138), .Q (signal_3070) ) ;
    buf_clk cell_1660 ( .C (CLK), .D (signal_1367), .Q (signal_3072) ) ;
    buf_clk cell_1662 ( .C (CLK), .D (signal_2142), .Q (signal_3074) ) ;
    buf_clk cell_1664 ( .C (CLK), .D (signal_1371), .Q (signal_3076) ) ;
    buf_clk cell_1666 ( .C (CLK), .D (signal_2096), .Q (signal_3078) ) ;
    buf_clk cell_1668 ( .C (CLK), .D (signal_1375), .Q (signal_3080) ) ;
    buf_clk cell_1670 ( .C (CLK), .D (signal_2100), .Q (signal_3082) ) ;
    buf_clk cell_1672 ( .C (CLK), .D (signal_1379), .Q (signal_3084) ) ;
    buf_clk cell_1674 ( .C (CLK), .D (signal_2145), .Q (signal_3086) ) ;
    buf_clk cell_1676 ( .C (CLK), .D (signal_1383), .Q (signal_3088) ) ;
    buf_clk cell_1678 ( .C (CLK), .D (signal_2149), .Q (signal_3090) ) ;
    buf_clk cell_1680 ( .C (CLK), .D (signal_1387), .Q (signal_3092) ) ;
    buf_clk cell_1682 ( .C (CLK), .D (signal_2104), .Q (signal_3094) ) ;
    buf_clk cell_1684 ( .C (CLK), .D (signal_1391), .Q (signal_3096) ) ;
    buf_clk cell_1686 ( .C (CLK), .D (signal_2108), .Q (signal_3098) ) ;
    buf_clk cell_1688 ( .C (CLK), .D (signal_1395), .Q (signal_3100) ) ;
    buf_clk cell_1690 ( .C (CLK), .D (signal_2152), .Q (signal_3102) ) ;
    buf_clk cell_1692 ( .C (CLK), .D (signal_1399), .Q (signal_3104) ) ;
    buf_clk cell_1694 ( .C (CLK), .D (signal_2155), .Q (signal_3106) ) ;
    buf_clk cell_1696 ( .C (CLK), .D (signal_1403), .Q (signal_3108) ) ;
    buf_clk cell_1698 ( .C (CLK), .D (signal_2114), .Q (signal_3110) ) ;
    buf_clk cell_1700 ( .C (CLK), .D (signal_1407), .Q (signal_3112) ) ;
    buf_clk cell_1702 ( .C (CLK), .D (signal_2118), .Q (signal_3114) ) ;
    buf_clk cell_1704 ( .C (CLK), .D (signal_1411), .Q (signal_3116) ) ;
    buf_clk cell_1706 ( .C (CLK), .D (signal_2159), .Q (signal_3118) ) ;
    buf_clk cell_1708 ( .C (CLK), .D (signal_1415), .Q (signal_3120) ) ;
    buf_clk cell_1710 ( .C (CLK), .D (signal_2163), .Q (signal_3122) ) ;
    buf_clk cell_1712 ( .C (CLK), .D (signal_1419), .Q (signal_3124) ) ;
    buf_clk cell_1714 ( .C (CLK), .D (signal_2122), .Q (signal_3126) ) ;
    buf_clk cell_1716 ( .C (CLK), .D (signal_1423), .Q (signal_3128) ) ;
    buf_clk cell_1718 ( .C (CLK), .D (signal_2126), .Q (signal_3130) ) ;
    buf_clk cell_1720 ( .C (CLK), .D (signal_343), .Q (signal_3132) ) ;
    buf_clk cell_1724 ( .C (CLK), .D (signal_312), .Q (signal_3136) ) ;
    buf_clk cell_1728 ( .C (CLK), .D (signal_1874), .Q (signal_3140) ) ;
    buf_clk cell_1732 ( .C (CLK), .D (signal_313), .Q (signal_3144) ) ;
    buf_clk cell_1736 ( .C (CLK), .D (signal_1994), .Q (signal_3148) ) ;
    buf_clk cell_1740 ( .C (CLK), .D (signal_344), .Q (signal_3152) ) ;
    buf_clk cell_1744 ( .C (CLK), .D (signal_314), .Q (signal_3156) ) ;
    buf_clk cell_1748 ( .C (CLK), .D (signal_1995), .Q (signal_3160) ) ;
    buf_clk cell_1752 ( .C (CLK), .D (signal_342), .Q (signal_3164) ) ;
    buf_clk cell_1756 ( .C (CLK), .D (signal_315), .Q (signal_3168) ) ;
    buf_clk cell_1760 ( .C (CLK), .D (signal_1875), .Q (signal_3172) ) ;
    buf_clk cell_1764 ( .C (CLK), .D (signal_316), .Q (signal_3176) ) ;
    buf_clk cell_1768 ( .C (CLK), .D (signal_1996), .Q (signal_3180) ) ;
    buf_clk cell_1772 ( .C (CLK), .D (signal_317), .Q (signal_3184) ) ;
    buf_clk cell_1776 ( .C (CLK), .D (signal_1997), .Q (signal_3188) ) ;
    buf_clk cell_1780 ( .C (CLK), .D (signal_318), .Q (signal_3192) ) ;
    buf_clk cell_1784 ( .C (CLK), .D (signal_1998), .Q (signal_3196) ) ;
    buf_clk cell_1788 ( .C (CLK), .D (signal_1000), .Q (signal_3200) ) ;
    buf_clk cell_1792 ( .C (CLK), .D (signal_1999), .Q (signal_3204) ) ;
    buf_clk cell_1796 ( .C (CLK), .D (signal_999), .Q (signal_3208) ) ;
    buf_clk cell_1800 ( .C (CLK), .D (signal_2000), .Q (signal_3212) ) ;
    buf_clk cell_1804 ( .C (CLK), .D (signal_998), .Q (signal_3216) ) ;
    buf_clk cell_1808 ( .C (CLK), .D (signal_2001), .Q (signal_3220) ) ;
    buf_clk cell_1812 ( .C (CLK), .D (signal_997), .Q (signal_3224) ) ;
    buf_clk cell_1816 ( .C (CLK), .D (signal_2002), .Q (signal_3228) ) ;
    buf_clk cell_1820 ( .C (CLK), .D (signal_996), .Q (signal_3232) ) ;
    buf_clk cell_1824 ( .C (CLK), .D (signal_2003), .Q (signal_3236) ) ;
    buf_clk cell_1828 ( .C (CLK), .D (signal_995), .Q (signal_3240) ) ;
    buf_clk cell_1832 ( .C (CLK), .D (signal_2004), .Q (signal_3244) ) ;
    buf_clk cell_1836 ( .C (CLK), .D (signal_994), .Q (signal_3248) ) ;
    buf_clk cell_1840 ( .C (CLK), .D (signal_2005), .Q (signal_3252) ) ;
    buf_clk cell_1844 ( .C (CLK), .D (signal_993), .Q (signal_3256) ) ;
    buf_clk cell_1848 ( .C (CLK), .D (signal_2006), .Q (signal_3260) ) ;
    buf_clk cell_1852 ( .C (CLK), .D (signal_992), .Q (signal_3264) ) ;
    buf_clk cell_1856 ( .C (CLK), .D (signal_2007), .Q (signal_3268) ) ;
    buf_clk cell_1860 ( .C (CLK), .D (signal_319), .Q (signal_3272) ) ;
    buf_clk cell_1864 ( .C (CLK), .D (signal_1876), .Q (signal_3276) ) ;
    buf_clk cell_1868 ( .C (CLK), .D (signal_320), .Q (signal_3280) ) ;
    buf_clk cell_1872 ( .C (CLK), .D (signal_2008), .Q (signal_3284) ) ;
    buf_clk cell_1876 ( .C (CLK), .D (signal_321), .Q (signal_3288) ) ;
    buf_clk cell_1880 ( .C (CLK), .D (signal_2009), .Q (signal_3292) ) ;
    buf_clk cell_1884 ( .C (CLK), .D (signal_322), .Q (signal_3296) ) ;
    buf_clk cell_1888 ( .C (CLK), .D (signal_1877), .Q (signal_3300) ) ;
    buf_clk cell_1892 ( .C (CLK), .D (signal_323), .Q (signal_3304) ) ;
    buf_clk cell_1896 ( .C (CLK), .D (signal_2010), .Q (signal_3308) ) ;
    buf_clk cell_1900 ( .C (CLK), .D (signal_324), .Q (signal_3312) ) ;
    buf_clk cell_1904 ( .C (CLK), .D (signal_2011), .Q (signal_3316) ) ;
    buf_clk cell_1908 ( .C (CLK), .D (signal_325), .Q (signal_3320) ) ;
    buf_clk cell_1912 ( .C (CLK), .D (signal_1878), .Q (signal_3324) ) ;
    buf_clk cell_1916 ( .C (CLK), .D (signal_984), .Q (signal_3328) ) ;
    buf_clk cell_1920 ( .C (CLK), .D (signal_2012), .Q (signal_3332) ) ;
    buf_clk cell_1924 ( .C (CLK), .D (signal_983), .Q (signal_3336) ) ;
    buf_clk cell_1928 ( .C (CLK), .D (signal_1879), .Q (signal_3340) ) ;
    buf_clk cell_1932 ( .C (CLK), .D (signal_982), .Q (signal_3344) ) ;
    buf_clk cell_1936 ( .C (CLK), .D (signal_2013), .Q (signal_3348) ) ;
    buf_clk cell_1940 ( .C (CLK), .D (signal_981), .Q (signal_3352) ) ;
    buf_clk cell_1944 ( .C (CLK), .D (signal_1880), .Q (signal_3356) ) ;
    buf_clk cell_1948 ( .C (CLK), .D (signal_980), .Q (signal_3360) ) ;
    buf_clk cell_1952 ( .C (CLK), .D (signal_2014), .Q (signal_3364) ) ;
    buf_clk cell_1956 ( .C (CLK), .D (signal_979), .Q (signal_3368) ) ;
    buf_clk cell_1960 ( .C (CLK), .D (signal_1983), .Q (signal_3372) ) ;
    buf_clk cell_1964 ( .C (CLK), .D (signal_978), .Q (signal_3376) ) ;
    buf_clk cell_1968 ( .C (CLK), .D (signal_2015), .Q (signal_3380) ) ;
    buf_clk cell_1972 ( .C (CLK), .D (signal_977), .Q (signal_3384) ) ;
    buf_clk cell_1976 ( .C (CLK), .D (signal_2016), .Q (signal_3388) ) ;
    buf_clk cell_1980 ( .C (CLK), .D (signal_976), .Q (signal_3392) ) ;
    buf_clk cell_1984 ( .C (CLK), .D (signal_2017), .Q (signal_3396) ) ;
    buf_clk cell_1988 ( .C (CLK), .D (signal_326), .Q (signal_3400) ) ;
    buf_clk cell_1992 ( .C (CLK), .D (signal_1984), .Q (signal_3404) ) ;
    buf_clk cell_1996 ( .C (CLK), .D (signal_327), .Q (signal_3408) ) ;
    buf_clk cell_2000 ( .C (CLK), .D (signal_2018), .Q (signal_3412) ) ;
    buf_clk cell_2004 ( .C (CLK), .D (signal_328), .Q (signal_3416) ) ;
    buf_clk cell_2008 ( .C (CLK), .D (signal_1985), .Q (signal_3420) ) ;
    buf_clk cell_2012 ( .C (CLK), .D (signal_329), .Q (signal_3424) ) ;
    buf_clk cell_2016 ( .C (CLK), .D (signal_1986), .Q (signal_3428) ) ;
    buf_clk cell_2020 ( .C (CLK), .D (signal_330), .Q (signal_3432) ) ;
    buf_clk cell_2024 ( .C (CLK), .D (signal_1987), .Q (signal_3436) ) ;
    buf_clk cell_2028 ( .C (CLK), .D (signal_331), .Q (signal_3440) ) ;
    buf_clk cell_2032 ( .C (CLK), .D (signal_2019), .Q (signal_3444) ) ;
    buf_clk cell_2036 ( .C (CLK), .D (signal_332), .Q (signal_3448) ) ;
    buf_clk cell_2040 ( .C (CLK), .D (signal_2020), .Q (signal_3452) ) ;
    buf_clk cell_2044 ( .C (CLK), .D (signal_968), .Q (signal_3456) ) ;
    buf_clk cell_2048 ( .C (CLK), .D (signal_1988), .Q (signal_3460) ) ;
    buf_clk cell_2052 ( .C (CLK), .D (signal_967), .Q (signal_3464) ) ;
    buf_clk cell_2056 ( .C (CLK), .D (signal_2021), .Q (signal_3468) ) ;
    buf_clk cell_2060 ( .C (CLK), .D (signal_966), .Q (signal_3472) ) ;
    buf_clk cell_2064 ( .C (CLK), .D (signal_2022), .Q (signal_3476) ) ;
    buf_clk cell_2068 ( .C (CLK), .D (signal_965), .Q (signal_3480) ) ;
    buf_clk cell_2072 ( .C (CLK), .D (signal_2023), .Q (signal_3484) ) ;
    buf_clk cell_2076 ( .C (CLK), .D (signal_340), .Q (signal_3488) ) ;
    buf_clk cell_2080 ( .C (CLK), .D (signal_964), .Q (signal_3492) ) ;
    buf_clk cell_2084 ( .C (CLK), .D (signal_2024), .Q (signal_3496) ) ;
    buf_clk cell_2088 ( .C (CLK), .D (signal_963), .Q (signal_3500) ) ;
    buf_clk cell_2092 ( .C (CLK), .D (signal_2025), .Q (signal_3504) ) ;
    buf_clk cell_2096 ( .C (CLK), .D (signal_962), .Q (signal_3508) ) ;
    buf_clk cell_2100 ( .C (CLK), .D (signal_2026), .Q (signal_3512) ) ;
    buf_clk cell_2104 ( .C (CLK), .D (signal_961), .Q (signal_3516) ) ;
    buf_clk cell_2108 ( .C (CLK), .D (signal_2027), .Q (signal_3520) ) ;
    buf_clk cell_2112 ( .C (CLK), .D (signal_960), .Q (signal_3524) ) ;
    buf_clk cell_2116 ( .C (CLK), .D (signal_2028), .Q (signal_3528) ) ;
    buf_clk cell_2120 ( .C (CLK), .D (signal_333), .Q (signal_3532) ) ;
    buf_clk cell_2124 ( .C (CLK), .D (signal_2029), .Q (signal_3536) ) ;
    buf_clk cell_2128 ( .C (CLK), .D (signal_334), .Q (signal_3540) ) ;
    buf_clk cell_2132 ( .C (CLK), .D (signal_2030), .Q (signal_3544) ) ;
    buf_clk cell_2136 ( .C (CLK), .D (signal_335), .Q (signal_3548) ) ;
    buf_clk cell_2140 ( .C (CLK), .D (signal_2031), .Q (signal_3552) ) ;
    buf_clk cell_2144 ( .C (CLK), .D (signal_336), .Q (signal_3556) ) ;
    buf_clk cell_2148 ( .C (CLK), .D (signal_2032), .Q (signal_3560) ) ;
    buf_clk cell_2152 ( .C (CLK), .D (signal_337), .Q (signal_3564) ) ;
    buf_clk cell_2156 ( .C (CLK), .D (signal_2033), .Q (signal_3568) ) ;
    buf_clk cell_2160 ( .C (CLK), .D (signal_338), .Q (signal_3572) ) ;
    buf_clk cell_2164 ( .C (CLK), .D (signal_2034), .Q (signal_3576) ) ;
    buf_clk cell_2168 ( .C (CLK), .D (signal_339), .Q (signal_3580) ) ;
    buf_clk cell_2172 ( .C (CLK), .D (signal_2035), .Q (signal_3584) ) ;
    buf_clk cell_2176 ( .C (CLK), .D (signal_952), .Q (signal_3588) ) ;
    buf_clk cell_2180 ( .C (CLK), .D (signal_2036), .Q (signal_3592) ) ;
    buf_clk cell_2184 ( .C (CLK), .D (signal_951), .Q (signal_3596) ) ;
    buf_clk cell_2188 ( .C (CLK), .D (signal_2037), .Q (signal_3600) ) ;
    buf_clk cell_2192 ( .C (CLK), .D (signal_950), .Q (signal_3604) ) ;
    buf_clk cell_2196 ( .C (CLK), .D (signal_2038), .Q (signal_3608) ) ;
    buf_clk cell_2200 ( .C (CLK), .D (signal_949), .Q (signal_3612) ) ;
    buf_clk cell_2204 ( .C (CLK), .D (signal_2039), .Q (signal_3616) ) ;
    buf_clk cell_2208 ( .C (CLK), .D (signal_948), .Q (signal_3620) ) ;
    buf_clk cell_2212 ( .C (CLK), .D (signal_2040), .Q (signal_3624) ) ;
    buf_clk cell_2216 ( .C (CLK), .D (signal_947), .Q (signal_3628) ) ;
    buf_clk cell_2220 ( .C (CLK), .D (signal_2041), .Q (signal_3632) ) ;
    buf_clk cell_2224 ( .C (CLK), .D (signal_946), .Q (signal_3636) ) ;
    buf_clk cell_2228 ( .C (CLK), .D (signal_2042), .Q (signal_3640) ) ;
    buf_clk cell_2232 ( .C (CLK), .D (signal_945), .Q (signal_3644) ) ;
    buf_clk cell_2236 ( .C (CLK), .D (signal_2043), .Q (signal_3648) ) ;
    buf_clk cell_2240 ( .C (CLK), .D (signal_944), .Q (signal_3652) ) ;
    buf_clk cell_2244 ( .C (CLK), .D (signal_2044), .Q (signal_3656) ) ;
    buf_clk cell_2248 ( .C (CLK), .D (IN_reset), .Q (signal_3660) ) ;
    buf_clk cell_2252 ( .C (CLK), .D (IN_plaintext_s0[0]), .Q (signal_3664) ) ;
    buf_clk cell_2256 ( .C (CLK), .D (IN_plaintext_s1[0]), .Q (signal_3668) ) ;
    buf_clk cell_2260 ( .C (CLK), .D (IN_plaintext_s0[1]), .Q (signal_3672) ) ;
    buf_clk cell_2264 ( .C (CLK), .D (IN_plaintext_s1[1]), .Q (signal_3676) ) ;
    buf_clk cell_2268 ( .C (CLK), .D (IN_plaintext_s0[2]), .Q (signal_3680) ) ;
    buf_clk cell_2272 ( .C (CLK), .D (IN_plaintext_s1[2]), .Q (signal_3684) ) ;
    buf_clk cell_2276 ( .C (CLK), .D (IN_plaintext_s0[3]), .Q (signal_3688) ) ;
    buf_clk cell_2280 ( .C (CLK), .D (IN_plaintext_s1[3]), .Q (signal_3692) ) ;
    buf_clk cell_2284 ( .C (CLK), .D (IN_plaintext_s0[4]), .Q (signal_3696) ) ;
    buf_clk cell_2288 ( .C (CLK), .D (IN_plaintext_s1[4]), .Q (signal_3700) ) ;
    buf_clk cell_2292 ( .C (CLK), .D (IN_plaintext_s0[5]), .Q (signal_3704) ) ;
    buf_clk cell_2296 ( .C (CLK), .D (IN_plaintext_s1[5]), .Q (signal_3708) ) ;
    buf_clk cell_2300 ( .C (CLK), .D (IN_plaintext_s0[6]), .Q (signal_3712) ) ;
    buf_clk cell_2304 ( .C (CLK), .D (IN_plaintext_s1[6]), .Q (signal_3716) ) ;
    buf_clk cell_2308 ( .C (CLK), .D (IN_plaintext_s0[7]), .Q (signal_3720) ) ;
    buf_clk cell_2312 ( .C (CLK), .D (IN_plaintext_s1[7]), .Q (signal_3724) ) ;
    buf_clk cell_2316 ( .C (CLK), .D (IN_plaintext_s0[8]), .Q (signal_3728) ) ;
    buf_clk cell_2320 ( .C (CLK), .D (IN_plaintext_s1[8]), .Q (signal_3732) ) ;
    buf_clk cell_2324 ( .C (CLK), .D (IN_plaintext_s0[9]), .Q (signal_3736) ) ;
    buf_clk cell_2328 ( .C (CLK), .D (IN_plaintext_s1[9]), .Q (signal_3740) ) ;
    buf_clk cell_2332 ( .C (CLK), .D (IN_plaintext_s0[10]), .Q (signal_3744) ) ;
    buf_clk cell_2336 ( .C (CLK), .D (IN_plaintext_s1[10]), .Q (signal_3748) ) ;
    buf_clk cell_2340 ( .C (CLK), .D (IN_plaintext_s0[11]), .Q (signal_3752) ) ;
    buf_clk cell_2344 ( .C (CLK), .D (IN_plaintext_s1[11]), .Q (signal_3756) ) ;
    buf_clk cell_2348 ( .C (CLK), .D (IN_plaintext_s0[12]), .Q (signal_3760) ) ;
    buf_clk cell_2352 ( .C (CLK), .D (IN_plaintext_s1[12]), .Q (signal_3764) ) ;
    buf_clk cell_2356 ( .C (CLK), .D (IN_plaintext_s0[13]), .Q (signal_3768) ) ;
    buf_clk cell_2360 ( .C (CLK), .D (IN_plaintext_s1[13]), .Q (signal_3772) ) ;
    buf_clk cell_2364 ( .C (CLK), .D (IN_plaintext_s0[14]), .Q (signal_3776) ) ;
    buf_clk cell_2368 ( .C (CLK), .D (IN_plaintext_s1[14]), .Q (signal_3780) ) ;
    buf_clk cell_2372 ( .C (CLK), .D (IN_plaintext_s0[15]), .Q (signal_3784) ) ;
    buf_clk cell_2376 ( .C (CLK), .D (IN_plaintext_s1[15]), .Q (signal_3788) ) ;
    buf_clk cell_2380 ( .C (CLK), .D (IN_plaintext_s0[16]), .Q (signal_3792) ) ;
    buf_clk cell_2384 ( .C (CLK), .D (IN_plaintext_s1[16]), .Q (signal_3796) ) ;
    buf_clk cell_2388 ( .C (CLK), .D (IN_plaintext_s0[17]), .Q (signal_3800) ) ;
    buf_clk cell_2392 ( .C (CLK), .D (IN_plaintext_s1[17]), .Q (signal_3804) ) ;
    buf_clk cell_2396 ( .C (CLK), .D (IN_plaintext_s0[18]), .Q (signal_3808) ) ;
    buf_clk cell_2400 ( .C (CLK), .D (IN_plaintext_s1[18]), .Q (signal_3812) ) ;
    buf_clk cell_2404 ( .C (CLK), .D (IN_plaintext_s0[19]), .Q (signal_3816) ) ;
    buf_clk cell_2408 ( .C (CLK), .D (IN_plaintext_s1[19]), .Q (signal_3820) ) ;
    buf_clk cell_2412 ( .C (CLK), .D (IN_plaintext_s0[20]), .Q (signal_3824) ) ;
    buf_clk cell_2416 ( .C (CLK), .D (IN_plaintext_s1[20]), .Q (signal_3828) ) ;
    buf_clk cell_2420 ( .C (CLK), .D (IN_plaintext_s0[21]), .Q (signal_3832) ) ;
    buf_clk cell_2424 ( .C (CLK), .D (IN_plaintext_s1[21]), .Q (signal_3836) ) ;
    buf_clk cell_2428 ( .C (CLK), .D (IN_plaintext_s0[22]), .Q (signal_3840) ) ;
    buf_clk cell_2432 ( .C (CLK), .D (IN_plaintext_s1[22]), .Q (signal_3844) ) ;
    buf_clk cell_2436 ( .C (CLK), .D (IN_plaintext_s0[23]), .Q (signal_3848) ) ;
    buf_clk cell_2440 ( .C (CLK), .D (IN_plaintext_s1[23]), .Q (signal_3852) ) ;
    buf_clk cell_2444 ( .C (CLK), .D (IN_plaintext_s0[24]), .Q (signal_3856) ) ;
    buf_clk cell_2448 ( .C (CLK), .D (IN_plaintext_s1[24]), .Q (signal_3860) ) ;
    buf_clk cell_2452 ( .C (CLK), .D (IN_plaintext_s0[25]), .Q (signal_3864) ) ;
    buf_clk cell_2456 ( .C (CLK), .D (IN_plaintext_s1[25]), .Q (signal_3868) ) ;
    buf_clk cell_2460 ( .C (CLK), .D (IN_plaintext_s0[26]), .Q (signal_3872) ) ;
    buf_clk cell_2464 ( .C (CLK), .D (IN_plaintext_s1[26]), .Q (signal_3876) ) ;
    buf_clk cell_2468 ( .C (CLK), .D (IN_plaintext_s0[27]), .Q (signal_3880) ) ;
    buf_clk cell_2472 ( .C (CLK), .D (IN_plaintext_s1[27]), .Q (signal_3884) ) ;
    buf_clk cell_2476 ( .C (CLK), .D (IN_plaintext_s0[28]), .Q (signal_3888) ) ;
    buf_clk cell_2480 ( .C (CLK), .D (IN_plaintext_s1[28]), .Q (signal_3892) ) ;
    buf_clk cell_2484 ( .C (CLK), .D (IN_plaintext_s0[29]), .Q (signal_3896) ) ;
    buf_clk cell_2488 ( .C (CLK), .D (IN_plaintext_s1[29]), .Q (signal_3900) ) ;
    buf_clk cell_2492 ( .C (CLK), .D (IN_plaintext_s0[30]), .Q (signal_3904) ) ;
    buf_clk cell_2496 ( .C (CLK), .D (IN_plaintext_s1[30]), .Q (signal_3908) ) ;
    buf_clk cell_2500 ( .C (CLK), .D (IN_plaintext_s0[31]), .Q (signal_3912) ) ;
    buf_clk cell_2504 ( .C (CLK), .D (IN_plaintext_s1[31]), .Q (signal_3916) ) ;
    buf_clk cell_2508 ( .C (CLK), .D (IN_plaintext_s0[32]), .Q (signal_3920) ) ;
    buf_clk cell_2512 ( .C (CLK), .D (IN_plaintext_s1[32]), .Q (signal_3924) ) ;
    buf_clk cell_2516 ( .C (CLK), .D (IN_plaintext_s0[33]), .Q (signal_3928) ) ;
    buf_clk cell_2520 ( .C (CLK), .D (IN_plaintext_s1[33]), .Q (signal_3932) ) ;
    buf_clk cell_2524 ( .C (CLK), .D (IN_plaintext_s0[34]), .Q (signal_3936) ) ;
    buf_clk cell_2528 ( .C (CLK), .D (IN_plaintext_s1[34]), .Q (signal_3940) ) ;
    buf_clk cell_2532 ( .C (CLK), .D (IN_plaintext_s0[35]), .Q (signal_3944) ) ;
    buf_clk cell_2536 ( .C (CLK), .D (IN_plaintext_s1[35]), .Q (signal_3948) ) ;
    buf_clk cell_2540 ( .C (CLK), .D (IN_plaintext_s0[36]), .Q (signal_3952) ) ;
    buf_clk cell_2544 ( .C (CLK), .D (IN_plaintext_s1[36]), .Q (signal_3956) ) ;
    buf_clk cell_2548 ( .C (CLK), .D (IN_plaintext_s0[37]), .Q (signal_3960) ) ;
    buf_clk cell_2552 ( .C (CLK), .D (IN_plaintext_s1[37]), .Q (signal_3964) ) ;
    buf_clk cell_2556 ( .C (CLK), .D (IN_plaintext_s0[38]), .Q (signal_3968) ) ;
    buf_clk cell_2560 ( .C (CLK), .D (IN_plaintext_s1[38]), .Q (signal_3972) ) ;
    buf_clk cell_2564 ( .C (CLK), .D (IN_plaintext_s0[39]), .Q (signal_3976) ) ;
    buf_clk cell_2568 ( .C (CLK), .D (IN_plaintext_s1[39]), .Q (signal_3980) ) ;
    buf_clk cell_2572 ( .C (CLK), .D (IN_plaintext_s0[40]), .Q (signal_3984) ) ;
    buf_clk cell_2576 ( .C (CLK), .D (IN_plaintext_s1[40]), .Q (signal_3988) ) ;
    buf_clk cell_2580 ( .C (CLK), .D (IN_plaintext_s0[41]), .Q (signal_3992) ) ;
    buf_clk cell_2584 ( .C (CLK), .D (IN_plaintext_s1[41]), .Q (signal_3996) ) ;
    buf_clk cell_2588 ( .C (CLK), .D (IN_plaintext_s0[42]), .Q (signal_4000) ) ;
    buf_clk cell_2592 ( .C (CLK), .D (IN_plaintext_s1[42]), .Q (signal_4004) ) ;
    buf_clk cell_2596 ( .C (CLK), .D (IN_plaintext_s0[43]), .Q (signal_4008) ) ;
    buf_clk cell_2600 ( .C (CLK), .D (IN_plaintext_s1[43]), .Q (signal_4012) ) ;
    buf_clk cell_2604 ( .C (CLK), .D (IN_plaintext_s0[44]), .Q (signal_4016) ) ;
    buf_clk cell_2608 ( .C (CLK), .D (IN_plaintext_s1[44]), .Q (signal_4020) ) ;
    buf_clk cell_2612 ( .C (CLK), .D (IN_plaintext_s0[45]), .Q (signal_4024) ) ;
    buf_clk cell_2616 ( .C (CLK), .D (IN_plaintext_s1[45]), .Q (signal_4028) ) ;
    buf_clk cell_2620 ( .C (CLK), .D (IN_plaintext_s0[46]), .Q (signal_4032) ) ;
    buf_clk cell_2624 ( .C (CLK), .D (IN_plaintext_s1[46]), .Q (signal_4036) ) ;
    buf_clk cell_2628 ( .C (CLK), .D (IN_plaintext_s0[47]), .Q (signal_4040) ) ;
    buf_clk cell_2632 ( .C (CLK), .D (IN_plaintext_s1[47]), .Q (signal_4044) ) ;
    buf_clk cell_2636 ( .C (CLK), .D (IN_plaintext_s0[48]), .Q (signal_4048) ) ;
    buf_clk cell_2640 ( .C (CLK), .D (IN_plaintext_s1[48]), .Q (signal_4052) ) ;
    buf_clk cell_2644 ( .C (CLK), .D (IN_plaintext_s0[49]), .Q (signal_4056) ) ;
    buf_clk cell_2648 ( .C (CLK), .D (IN_plaintext_s1[49]), .Q (signal_4060) ) ;
    buf_clk cell_2652 ( .C (CLK), .D (IN_plaintext_s0[50]), .Q (signal_4064) ) ;
    buf_clk cell_2656 ( .C (CLK), .D (IN_plaintext_s1[50]), .Q (signal_4068) ) ;
    buf_clk cell_2660 ( .C (CLK), .D (IN_plaintext_s0[51]), .Q (signal_4072) ) ;
    buf_clk cell_2664 ( .C (CLK), .D (IN_plaintext_s1[51]), .Q (signal_4076) ) ;
    buf_clk cell_2668 ( .C (CLK), .D (IN_plaintext_s0[52]), .Q (signal_4080) ) ;
    buf_clk cell_2672 ( .C (CLK), .D (IN_plaintext_s1[52]), .Q (signal_4084) ) ;
    buf_clk cell_2676 ( .C (CLK), .D (IN_plaintext_s0[53]), .Q (signal_4088) ) ;
    buf_clk cell_2680 ( .C (CLK), .D (IN_plaintext_s1[53]), .Q (signal_4092) ) ;
    buf_clk cell_2684 ( .C (CLK), .D (IN_plaintext_s0[54]), .Q (signal_4096) ) ;
    buf_clk cell_2688 ( .C (CLK), .D (IN_plaintext_s1[54]), .Q (signal_4100) ) ;
    buf_clk cell_2692 ( .C (CLK), .D (IN_plaintext_s0[55]), .Q (signal_4104) ) ;
    buf_clk cell_2696 ( .C (CLK), .D (IN_plaintext_s1[55]), .Q (signal_4108) ) ;
    buf_clk cell_2700 ( .C (CLK), .D (IN_plaintext_s0[56]), .Q (signal_4112) ) ;
    buf_clk cell_2704 ( .C (CLK), .D (IN_plaintext_s1[56]), .Q (signal_4116) ) ;
    buf_clk cell_2708 ( .C (CLK), .D (IN_plaintext_s0[57]), .Q (signal_4120) ) ;
    buf_clk cell_2712 ( .C (CLK), .D (IN_plaintext_s1[57]), .Q (signal_4124) ) ;
    buf_clk cell_2716 ( .C (CLK), .D (IN_plaintext_s0[58]), .Q (signal_4128) ) ;
    buf_clk cell_2720 ( .C (CLK), .D (IN_plaintext_s1[58]), .Q (signal_4132) ) ;
    buf_clk cell_2724 ( .C (CLK), .D (IN_plaintext_s0[59]), .Q (signal_4136) ) ;
    buf_clk cell_2728 ( .C (CLK), .D (IN_plaintext_s1[59]), .Q (signal_4140) ) ;
    buf_clk cell_2732 ( .C (CLK), .D (IN_plaintext_s0[60]), .Q (signal_4144) ) ;
    buf_clk cell_2736 ( .C (CLK), .D (IN_plaintext_s1[60]), .Q (signal_4148) ) ;
    buf_clk cell_2740 ( .C (CLK), .D (IN_plaintext_s0[61]), .Q (signal_4152) ) ;
    buf_clk cell_2744 ( .C (CLK), .D (IN_plaintext_s1[61]), .Q (signal_4156) ) ;
    buf_clk cell_2748 ( .C (CLK), .D (IN_plaintext_s0[62]), .Q (signal_4160) ) ;
    buf_clk cell_2752 ( .C (CLK), .D (IN_plaintext_s1[62]), .Q (signal_4164) ) ;
    buf_clk cell_2756 ( .C (CLK), .D (IN_plaintext_s0[63]), .Q (signal_4168) ) ;
    buf_clk cell_2760 ( .C (CLK), .D (IN_plaintext_s1[63]), .Q (signal_4172) ) ;
    buf_clk cell_2764 ( .C (CLK), .D (signal_1007), .Q (signal_4176) ) ;
    buf_clk cell_2768 ( .C (CLK), .D (signal_1993), .Q (signal_4180) ) ;
    buf_clk cell_2772 ( .C (CLK), .D (signal_1003), .Q (signal_4184) ) ;
    buf_clk cell_2776 ( .C (CLK), .D (signal_2061), .Q (signal_4188) ) ;
    buf_clk cell_2780 ( .C (CLK), .D (signal_991), .Q (signal_4192) ) ;
    buf_clk cell_2784 ( .C (CLK), .D (signal_1992), .Q (signal_4196) ) ;
    buf_clk cell_2788 ( .C (CLK), .D (signal_987), .Q (signal_4200) ) ;
    buf_clk cell_2792 ( .C (CLK), .D (signal_2069), .Q (signal_4204) ) ;
    buf_clk cell_2796 ( .C (CLK), .D (signal_975), .Q (signal_4208) ) ;
    buf_clk cell_2800 ( .C (CLK), .D (signal_2048), .Q (signal_4212) ) ;
    buf_clk cell_2804 ( .C (CLK), .D (signal_971), .Q (signal_4216) ) ;
    buf_clk cell_2808 ( .C (CLK), .D (signal_2045), .Q (signal_4220) ) ;
    buf_clk cell_2812 ( .C (CLK), .D (signal_959), .Q (signal_4224) ) ;
    buf_clk cell_2816 ( .C (CLK), .D (signal_2063), .Q (signal_4228) ) ;
    buf_clk cell_2820 ( .C (CLK), .D (signal_955), .Q (signal_4232) ) ;
    buf_clk cell_2824 ( .C (CLK), .D (signal_2058), .Q (signal_4236) ) ;
    buf_clk cell_2876 ( .C (CLK), .D (signal_1457), .Q (signal_4288) ) ;
    buf_clk cell_2878 ( .C (CLK), .D (signal_2221), .Q (signal_4290) ) ;
    buf_clk cell_2880 ( .C (CLK), .D (signal_1460), .Q (signal_4292) ) ;
    buf_clk cell_2882 ( .C (CLK), .D (signal_2224), .Q (signal_4294) ) ;
    buf_clk cell_2884 ( .C (CLK), .D (signal_1463), .Q (signal_4296) ) ;
    buf_clk cell_2886 ( .C (CLK), .D (signal_2181), .Q (signal_4298) ) ;
    buf_clk cell_2888 ( .C (CLK), .D (signal_1466), .Q (signal_4300) ) ;
    buf_clk cell_2890 ( .C (CLK), .D (signal_2184), .Q (signal_4302) ) ;
    buf_clk cell_2892 ( .C (CLK), .D (signal_1469), .Q (signal_4304) ) ;
    buf_clk cell_2894 ( .C (CLK), .D (signal_2227), .Q (signal_4306) ) ;
    buf_clk cell_2896 ( .C (CLK), .D (signal_1472), .Q (signal_4308) ) ;
    buf_clk cell_2898 ( .C (CLK), .D (signal_2230), .Q (signal_4310) ) ;
    buf_clk cell_2900 ( .C (CLK), .D (signal_1475), .Q (signal_4312) ) ;
    buf_clk cell_2902 ( .C (CLK), .D (signal_2187), .Q (signal_4314) ) ;
    buf_clk cell_2904 ( .C (CLK), .D (signal_1478), .Q (signal_4316) ) ;
    buf_clk cell_2906 ( .C (CLK), .D (signal_2190), .Q (signal_4318) ) ;
    buf_clk cell_2908 ( .C (CLK), .D (signal_1481), .Q (signal_4320) ) ;
    buf_clk cell_2910 ( .C (CLK), .D (signal_2233), .Q (signal_4322) ) ;
    buf_clk cell_2912 ( .C (CLK), .D (signal_1484), .Q (signal_4324) ) ;
    buf_clk cell_2914 ( .C (CLK), .D (signal_2236), .Q (signal_4326) ) ;
    buf_clk cell_2916 ( .C (CLK), .D (signal_1487), .Q (signal_4328) ) ;
    buf_clk cell_2918 ( .C (CLK), .D (signal_2193), .Q (signal_4330) ) ;
    buf_clk cell_2920 ( .C (CLK), .D (signal_1490), .Q (signal_4332) ) ;
    buf_clk cell_2922 ( .C (CLK), .D (signal_2196), .Q (signal_4334) ) ;
    buf_clk cell_2924 ( .C (CLK), .D (signal_1493), .Q (signal_4336) ) ;
    buf_clk cell_2926 ( .C (CLK), .D (signal_2239), .Q (signal_4338) ) ;
    buf_clk cell_2928 ( .C (CLK), .D (signal_1496), .Q (signal_4340) ) ;
    buf_clk cell_2930 ( .C (CLK), .D (signal_2242), .Q (signal_4342) ) ;
    buf_clk cell_2932 ( .C (CLK), .D (signal_1499), .Q (signal_4344) ) ;
    buf_clk cell_2934 ( .C (CLK), .D (signal_2199), .Q (signal_4346) ) ;
    buf_clk cell_2936 ( .C (CLK), .D (signal_1502), .Q (signal_4348) ) ;
    buf_clk cell_2938 ( .C (CLK), .D (signal_2202), .Q (signal_4350) ) ;
    buf_clk cell_2940 ( .C (CLK), .D (signal_1458), .Q (signal_4352) ) ;
    buf_clk cell_2942 ( .C (CLK), .D (signal_2222), .Q (signal_4354) ) ;
    buf_clk cell_2944 ( .C (CLK), .D (signal_1461), .Q (signal_4356) ) ;
    buf_clk cell_2946 ( .C (CLK), .D (signal_2225), .Q (signal_4358) ) ;
    buf_clk cell_2948 ( .C (CLK), .D (signal_1464), .Q (signal_4360) ) ;
    buf_clk cell_2950 ( .C (CLK), .D (signal_2182), .Q (signal_4362) ) ;
    buf_clk cell_2952 ( .C (CLK), .D (signal_1467), .Q (signal_4364) ) ;
    buf_clk cell_2954 ( .C (CLK), .D (signal_2185), .Q (signal_4366) ) ;
    buf_clk cell_2956 ( .C (CLK), .D (signal_1470), .Q (signal_4368) ) ;
    buf_clk cell_2958 ( .C (CLK), .D (signal_2228), .Q (signal_4370) ) ;
    buf_clk cell_2960 ( .C (CLK), .D (signal_1473), .Q (signal_4372) ) ;
    buf_clk cell_2962 ( .C (CLK), .D (signal_2231), .Q (signal_4374) ) ;
    buf_clk cell_2964 ( .C (CLK), .D (signal_1476), .Q (signal_4376) ) ;
    buf_clk cell_2966 ( .C (CLK), .D (signal_2188), .Q (signal_4378) ) ;
    buf_clk cell_2968 ( .C (CLK), .D (signal_1479), .Q (signal_4380) ) ;
    buf_clk cell_2970 ( .C (CLK), .D (signal_2191), .Q (signal_4382) ) ;
    buf_clk cell_2972 ( .C (CLK), .D (signal_1482), .Q (signal_4384) ) ;
    buf_clk cell_2974 ( .C (CLK), .D (signal_2234), .Q (signal_4386) ) ;
    buf_clk cell_2976 ( .C (CLK), .D (signal_1485), .Q (signal_4388) ) ;
    buf_clk cell_2978 ( .C (CLK), .D (signal_2237), .Q (signal_4390) ) ;
    buf_clk cell_2980 ( .C (CLK), .D (signal_1488), .Q (signal_4392) ) ;
    buf_clk cell_2982 ( .C (CLK), .D (signal_2194), .Q (signal_4394) ) ;
    buf_clk cell_2984 ( .C (CLK), .D (signal_1491), .Q (signal_4396) ) ;
    buf_clk cell_2986 ( .C (CLK), .D (signal_2197), .Q (signal_4398) ) ;
    buf_clk cell_2988 ( .C (CLK), .D (signal_1494), .Q (signal_4400) ) ;
    buf_clk cell_2990 ( .C (CLK), .D (signal_2240), .Q (signal_4402) ) ;
    buf_clk cell_2992 ( .C (CLK), .D (signal_1497), .Q (signal_4404) ) ;
    buf_clk cell_2994 ( .C (CLK), .D (signal_2243), .Q (signal_4406) ) ;
    buf_clk cell_2996 ( .C (CLK), .D (signal_1500), .Q (signal_4408) ) ;
    buf_clk cell_2998 ( .C (CLK), .D (signal_2200), .Q (signal_4410) ) ;
    buf_clk cell_3000 ( .C (CLK), .D (signal_1503), .Q (signal_4412) ) ;
    buf_clk cell_3002 ( .C (CLK), .D (signal_2203), .Q (signal_4414) ) ;
    buf_clk cell_3068 ( .C (CLK), .D (signal_1361), .Q (signal_4480) ) ;
    buf_clk cell_3072 ( .C (CLK), .D (signal_2137), .Q (signal_4484) ) ;
    buf_clk cell_3080 ( .C (CLK), .D (signal_1365), .Q (signal_4492) ) ;
    buf_clk cell_3084 ( .C (CLK), .D (signal_2140), .Q (signal_4496) ) ;
    buf_clk cell_3092 ( .C (CLK), .D (signal_1369), .Q (signal_4504) ) ;
    buf_clk cell_3096 ( .C (CLK), .D (signal_2094), .Q (signal_4508) ) ;
    buf_clk cell_3104 ( .C (CLK), .D (signal_1373), .Q (signal_4516) ) ;
    buf_clk cell_3108 ( .C (CLK), .D (signal_2098), .Q (signal_4520) ) ;
    buf_clk cell_3116 ( .C (CLK), .D (signal_1377), .Q (signal_4528) ) ;
    buf_clk cell_3120 ( .C (CLK), .D (signal_2144), .Q (signal_4532) ) ;
    buf_clk cell_3128 ( .C (CLK), .D (signal_1381), .Q (signal_4540) ) ;
    buf_clk cell_3132 ( .C (CLK), .D (signal_2147), .Q (signal_4544) ) ;
    buf_clk cell_3140 ( .C (CLK), .D (signal_1385), .Q (signal_4552) ) ;
    buf_clk cell_3144 ( .C (CLK), .D (signal_2102), .Q (signal_4556) ) ;
    buf_clk cell_3152 ( .C (CLK), .D (signal_1389), .Q (signal_4564) ) ;
    buf_clk cell_3156 ( .C (CLK), .D (signal_2106), .Q (signal_4568) ) ;
    buf_clk cell_3164 ( .C (CLK), .D (signal_1393), .Q (signal_4576) ) ;
    buf_clk cell_3168 ( .C (CLK), .D (signal_2151), .Q (signal_4580) ) ;
    buf_clk cell_3176 ( .C (CLK), .D (signal_1397), .Q (signal_4588) ) ;
    buf_clk cell_3180 ( .C (CLK), .D (signal_2154), .Q (signal_4592) ) ;
    buf_clk cell_3188 ( .C (CLK), .D (signal_1401), .Q (signal_4600) ) ;
    buf_clk cell_3192 ( .C (CLK), .D (signal_2112), .Q (signal_4604) ) ;
    buf_clk cell_3200 ( .C (CLK), .D (signal_1405), .Q (signal_4612) ) ;
    buf_clk cell_3204 ( .C (CLK), .D (signal_2116), .Q (signal_4616) ) ;
    buf_clk cell_3212 ( .C (CLK), .D (signal_1409), .Q (signal_4624) ) ;
    buf_clk cell_3216 ( .C (CLK), .D (signal_2157), .Q (signal_4628) ) ;
    buf_clk cell_3224 ( .C (CLK), .D (signal_1413), .Q (signal_4636) ) ;
    buf_clk cell_3228 ( .C (CLK), .D (signal_2161), .Q (signal_4640) ) ;
    buf_clk cell_3236 ( .C (CLK), .D (signal_1417), .Q (signal_4648) ) ;
    buf_clk cell_3240 ( .C (CLK), .D (signal_2120), .Q (signal_4652) ) ;
    buf_clk cell_3248 ( .C (CLK), .D (signal_1421), .Q (signal_4660) ) ;
    buf_clk cell_3252 ( .C (CLK), .D (signal_2124), .Q (signal_4664) ) ;
    buf_clk cell_3276 ( .C (CLK), .D (signal_310), .Q (signal_4688) ) ;
    buf_clk cell_3280 ( .C (CLK), .D (signal_308), .Q (signal_4692) ) ;
    buf_clk cell_3284 ( .C (CLK), .D (signal_305), .Q (signal_4696) ) ;
    buf_clk cell_3288 ( .C (CLK), .D (signal_303), .Q (signal_4700) ) ;
    buf_clk cell_3292 ( .C (CLK), .D (signal_301), .Q (signal_4704) ) ;
    buf_clk cell_3296 ( .C (CLK), .D (signal_299), .Q (signal_4708) ) ;
    buf_clk cell_3300 ( .C (CLK), .D (signal_297), .Q (signal_4712) ) ;
    buf_clk cell_3304 ( .C (CLK), .D (signal_295), .Q (signal_4716) ) ;
    buf_clk cell_3308 ( .C (CLK), .D (signal_293), .Q (signal_4720) ) ;
    buf_clk cell_3312 ( .C (CLK), .D (signal_291), .Q (signal_4724) ) ;
    buf_clk cell_3316 ( .C (CLK), .D (signal_265), .Q (signal_4728) ) ;

    /* cells in depth 2 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1240 ( .a ({signal_2067, signal_1005}), .b ({signal_2134, signal_1358}), .clk (CLK), .r (Fresh[0]), .c ({signal_2212, signal_1440}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1241 ( .a ({signal_2054, signal_1001}), .b ({signal_2127, signal_1351}), .clk (CLK), .r (Fresh[1]), .c ({signal_2213, signal_1441}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1242 ( .a ({signal_2074, signal_1332}), .b ({signal_2002, signal_997}), .clk (CLK), .r (Fresh[2]), .c ({signal_2172, signal_1442}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1243 ( .a ({signal_2076, signal_1334}), .b ({signal_2006, signal_993}), .clk (CLK), .r (Fresh[3]), .c ({signal_2173, signal_1443}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1244 ( .a ({signal_2071, signal_989}), .b ({signal_2135, signal_1359}), .clk (CLK), .r (Fresh[4]), .c ({signal_2214, signal_1444}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1245 ( .a ({signal_1990, signal_985}), .b ({signal_2133, signal_1357}), .clk (CLK), .r (Fresh[5]), .c ({signal_2215, signal_1445}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1246 ( .a ({signal_1880, signal_981}), .b ({signal_2079, signal_1337}), .clk (CLK), .r (Fresh[6]), .c ({signal_2174, signal_1446}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1247 ( .a ({signal_2081, signal_1339}), .b ({signal_2016, signal_977}), .clk (CLK), .r (Fresh[7]), .c ({signal_2175, signal_1447}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1248 ( .a ({signal_2047, signal_973}), .b ({signal_2132, signal_1356}), .clk (CLK), .r (Fresh[8]), .c ({signal_2216, signal_1448}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1249 ( .a ({signal_2064, signal_969}), .b ({signal_2131, signal_1355}), .clk (CLK), .r (Fresh[9]), .c ({signal_2217, signal_1449}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1250 ( .a ({signal_2083, signal_1341}), .b ({signal_2023, signal_965}), .clk (CLK), .r (Fresh[10]), .c ({signal_2176, signal_1450}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1251 ( .a ({signal_2085, signal_1343}), .b ({signal_2027, signal_961}), .clk (CLK), .r (Fresh[11]), .c ({signal_2177, signal_1451}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1252 ( .a ({signal_2060, signal_957}), .b ({signal_2130, signal_1354}), .clk (CLK), .r (Fresh[12]), .c ({signal_2218, signal_1452}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1253 ( .a ({signal_2056, signal_953}), .b ({signal_2128, signal_1352}), .clk (CLK), .r (Fresh[13]), .c ({signal_2219, signal_1453}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1254 ( .a ({signal_2088, signal_1346}), .b ({signal_2039, signal_949}), .clk (CLK), .r (Fresh[14]), .c ({signal_2178, signal_1454}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1255 ( .a ({signal_2090, signal_1348}), .b ({signal_2043, signal_945}), .clk (CLK), .r (Fresh[15]), .c ({signal_2179, signal_1455}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1304 ( .a ({signal_2050, signal_1329}), .b ({signal_2204, signal_1424}), .clk (CLK), .r (Fresh[16]), .c ({signal_2260, signal_1504}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1305 ( .a ({signal_2073, signal_1331}), .b ({signal_2205, signal_1425}), .clk (CLK), .r (Fresh[17]), .c ({signal_2261, signal_1505}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1306 ( .a ({signal_2075, signal_1333}), .b ({signal_2164, signal_1426}), .clk (CLK), .r (Fresh[18]), .c ({signal_2244, signal_1506}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1307 ( .a ({signal_2077, signal_1335}), .b ({signal_2165, signal_1427}), .clk (CLK), .r (Fresh[19]), .c ({signal_2245, signal_1507}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1308 ( .a ({signal_2051, signal_1330}), .b ({signal_2206, signal_1428}), .clk (CLK), .r (Fresh[20]), .c ({signal_2262, signal_1508}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1309 ( .a ({signal_2078, signal_1336}), .b ({signal_2207, signal_1429}), .clk (CLK), .r (Fresh[21]), .c ({signal_2263, signal_1509}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1310 ( .a ({signal_2080, signal_1338}), .b ({signal_2166, signal_1430}), .clk (CLK), .r (Fresh[22]), .c ({signal_2246, signal_1510}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1311 ( .a ({signal_2082, signal_1340}), .b ({signal_2167, signal_1431}), .clk (CLK), .r (Fresh[23]), .c ({signal_2247, signal_1511}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1312 ( .a ({signal_2092, signal_1350}), .b ({signal_2208, signal_1432}), .clk (CLK), .r (Fresh[24]), .c ({signal_2264, signal_1512}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1313 ( .a ({signal_2049, signal_1328}), .b ({signal_2209, signal_1433}), .clk (CLK), .r (Fresh[25]), .c ({signal_2265, signal_1513}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1314 ( .a ({signal_2084, signal_1342}), .b ({signal_2168, signal_1434}), .clk (CLK), .r (Fresh[26]), .c ({signal_2248, signal_1514}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1315 ( .a ({signal_2086, signal_1344}), .b ({signal_2169, signal_1435}), .clk (CLK), .r (Fresh[27]), .c ({signal_2249, signal_1515}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1316 ( .a ({signal_2129, signal_1353}), .b ({signal_2210, signal_1436}), .clk (CLK), .r (Fresh[28]), .c ({signal_2266, signal_1516}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1317 ( .a ({signal_2087, signal_1345}), .b ({signal_2211, signal_1437}), .clk (CLK), .r (Fresh[29]), .c ({signal_2267, signal_1517}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1318 ( .a ({signal_2089, signal_1347}), .b ({signal_2170, signal_1438}), .clk (CLK), .r (Fresh[30]), .c ({signal_2250, signal_1518}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1319 ( .a ({signal_2091, signal_1349}), .b ({signal_2171, signal_1439}), .clk (CLK), .r (Fresh[31]), .c ({signal_2251, signal_1519}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1320 ( .a ({signal_2943, signal_2941}), .b ({signal_2212, signal_1440}), .c ({signal_2268, signal_1520}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1321 ( .a ({signal_2947, signal_2945}), .b ({signal_2213, signal_1441}), .c ({signal_2269, signal_1521}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1322 ( .a ({signal_2951, signal_2949}), .b ({signal_2172, signal_1442}), .c ({signal_2252, signal_1522}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1323 ( .a ({signal_2955, signal_2953}), .b ({signal_2173, signal_1443}), .c ({signal_2253, signal_1523}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1324 ( .a ({signal_2959, signal_2957}), .b ({signal_2214, signal_1444}), .c ({signal_2270, signal_927}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1325 ( .a ({signal_2963, signal_2961}), .b ({signal_2215, signal_1445}), .c ({signal_2271, signal_923}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1326 ( .a ({signal_2967, signal_2965}), .b ({signal_2174, signal_1446}), .c ({signal_2254, signal_919}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1327 ( .a ({signal_2971, signal_2969}), .b ({signal_2175, signal_1447}), .c ({signal_2255, signal_915}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1328 ( .a ({signal_2975, signal_2973}), .b ({signal_2216, signal_1448}), .c ({signal_2272, signal_911}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1329 ( .a ({signal_2979, signal_2977}), .b ({signal_2217, signal_1449}), .c ({signal_2273, signal_907}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1330 ( .a ({signal_2983, signal_2981}), .b ({signal_2176, signal_1450}), .c ({signal_2256, signal_903}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1331 ( .a ({signal_2987, signal_2985}), .b ({signal_2177, signal_1451}), .c ({signal_2257, signal_899}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1332 ( .a ({signal_2991, signal_2989}), .b ({signal_2218, signal_1452}), .c ({signal_2274, signal_895}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1333 ( .a ({signal_2995, signal_2993}), .b ({signal_2219, signal_1453}), .c ({signal_2275, signal_891}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1334 ( .a ({signal_2999, signal_2997}), .b ({signal_2178, signal_1454}), .c ({signal_2258, signal_887}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1335 ( .a ({signal_3003, signal_3001}), .b ({signal_2179, signal_1455}), .c ({signal_2259, signal_883}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1336 ( .a ({signal_3007, signal_3005}), .b ({signal_2260, signal_1504}), .c ({signal_2292, signal_1524}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1337 ( .a ({signal_2212, signal_1440}), .b ({signal_2260, signal_1504}), .c ({signal_2293, signal_1525}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1338 ( .a ({signal_3011, signal_3009}), .b ({signal_2261, signal_1505}), .c ({signal_2294, signal_1526}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1339 ( .a ({signal_2213, signal_1441}), .b ({signal_2261, signal_1505}), .c ({signal_2295, signal_1527}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1340 ( .a ({signal_3015, signal_3013}), .b ({signal_2244, signal_1506}), .c ({signal_2276, signal_1528}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1341 ( .a ({signal_2172, signal_1442}), .b ({signal_2244, signal_1506}), .c ({signal_2277, signal_1529}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1342 ( .a ({signal_3019, signal_3017}), .b ({signal_2245, signal_1507}), .c ({signal_2278, signal_1530}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1343 ( .a ({signal_2173, signal_1443}), .b ({signal_2245, signal_1507}), .c ({signal_2279, signal_1531}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1344 ( .a ({signal_3023, signal_3021}), .b ({signal_2262, signal_1508}), .c ({signal_2296, signal_1532}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1345 ( .a ({signal_2214, signal_1444}), .b ({signal_2262, signal_1508}), .c ({signal_2297, signal_1533}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1346 ( .a ({signal_3027, signal_3025}), .b ({signal_2263, signal_1509}), .c ({signal_2298, signal_1534}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1347 ( .a ({signal_2215, signal_1445}), .b ({signal_2263, signal_1509}), .c ({signal_2299, signal_1535}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1348 ( .a ({signal_3031, signal_3029}), .b ({signal_2246, signal_1510}), .c ({signal_2280, signal_1536}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1349 ( .a ({signal_2174, signal_1446}), .b ({signal_2246, signal_1510}), .c ({signal_2281, signal_1537}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1350 ( .a ({signal_3035, signal_3033}), .b ({signal_2247, signal_1511}), .c ({signal_2282, signal_1538}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1351 ( .a ({signal_2175, signal_1447}), .b ({signal_2247, signal_1511}), .c ({signal_2283, signal_1539}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1352 ( .a ({signal_3039, signal_3037}), .b ({signal_2264, signal_1512}), .c ({signal_2300, signal_1540}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1353 ( .a ({signal_2216, signal_1448}), .b ({signal_2264, signal_1512}), .c ({signal_2301, signal_1541}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1354 ( .a ({signal_3043, signal_3041}), .b ({signal_2265, signal_1513}), .c ({signal_2302, signal_1542}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1355 ( .a ({signal_2217, signal_1449}), .b ({signal_2265, signal_1513}), .c ({signal_2303, signal_1543}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1356 ( .a ({signal_3047, signal_3045}), .b ({signal_2248, signal_1514}), .c ({signal_2284, signal_1544}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1357 ( .a ({signal_2176, signal_1450}), .b ({signal_2248, signal_1514}), .c ({signal_2285, signal_1545}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1358 ( .a ({signal_3051, signal_3049}), .b ({signal_2249, signal_1515}), .c ({signal_2286, signal_1546}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1359 ( .a ({signal_2177, signal_1451}), .b ({signal_2249, signal_1515}), .c ({signal_2287, signal_1547}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1360 ( .a ({signal_3055, signal_3053}), .b ({signal_2266, signal_1516}), .c ({signal_2304, signal_1548}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1361 ( .a ({signal_2218, signal_1452}), .b ({signal_2266, signal_1516}), .c ({signal_2305, signal_1549}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1362 ( .a ({signal_3059, signal_3057}), .b ({signal_2267, signal_1517}), .c ({signal_2306, signal_1550}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1363 ( .a ({signal_2219, signal_1453}), .b ({signal_2267, signal_1517}), .c ({signal_2307, signal_1551}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1364 ( .a ({signal_3063, signal_3061}), .b ({signal_2250, signal_1518}), .c ({signal_2288, signal_1552}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1365 ( .a ({signal_2178, signal_1454}), .b ({signal_2250, signal_1518}), .c ({signal_2289, signal_1553}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1366 ( .a ({signal_3067, signal_3065}), .b ({signal_2251, signal_1519}), .c ({signal_2290, signal_1554}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1367 ( .a ({signal_2179, signal_1455}), .b ({signal_2251, signal_1519}), .c ({signal_2291, signal_1555}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1368 ( .a ({signal_2292, signal_1524}), .b ({signal_2324, signal_1556}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1369 ( .a ({signal_2294, signal_1526}), .b ({signal_2325, signal_1557}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1370 ( .a ({signal_2276, signal_1528}), .b ({signal_2308, signal_1558}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1371 ( .a ({signal_2278, signal_1530}), .b ({signal_2309, signal_1559}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1372 ( .a ({signal_2296, signal_1532}), .b ({signal_2326, signal_1560}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1373 ( .a ({signal_2298, signal_1534}), .b ({signal_2327, signal_1561}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1374 ( .a ({signal_2280, signal_1536}), .b ({signal_2310, signal_1562}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1375 ( .a ({signal_2282, signal_1538}), .b ({signal_2311, signal_1563}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1376 ( .a ({signal_2300, signal_1540}), .b ({signal_2328, signal_1564}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1377 ( .a ({signal_2302, signal_1542}), .b ({signal_2329, signal_1565}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1378 ( .a ({signal_2284, signal_1544}), .b ({signal_2312, signal_1566}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1379 ( .a ({signal_2286, signal_1546}), .b ({signal_2313, signal_1567}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1380 ( .a ({signal_2304, signal_1548}), .b ({signal_2330, signal_1568}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1381 ( .a ({signal_2306, signal_1550}), .b ({signal_2331, signal_1569}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1382 ( .a ({signal_2288, signal_1552}), .b ({signal_2314, signal_1570}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1383 ( .a ({signal_2290, signal_1554}), .b ({signal_2315, signal_1571}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1384 ( .a ({signal_3071, signal_3069}), .b ({signal_2293, signal_1525}), .c ({signal_2332, signal_1572}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1385 ( .a ({signal_3075, signal_3073}), .b ({signal_2295, signal_1527}), .c ({signal_2333, signal_1573}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1386 ( .a ({signal_3079, signal_3077}), .b ({signal_2277, signal_1529}), .c ({signal_2316, signal_1574}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1387 ( .a ({signal_3083, signal_3081}), .b ({signal_2279, signal_1531}), .c ({signal_2317, signal_1575}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1388 ( .a ({signal_3087, signal_3085}), .b ({signal_2297, signal_1533}), .c ({signal_2334, signal_1576}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1389 ( .a ({signal_3091, signal_3089}), .b ({signal_2299, signal_1535}), .c ({signal_2335, signal_1577}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1390 ( .a ({signal_3095, signal_3093}), .b ({signal_2281, signal_1537}), .c ({signal_2318, signal_1578}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1391 ( .a ({signal_3099, signal_3097}), .b ({signal_2283, signal_1539}), .c ({signal_2319, signal_1579}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1392 ( .a ({signal_3103, signal_3101}), .b ({signal_2301, signal_1541}), .c ({signal_2336, signal_1580}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1393 ( .a ({signal_3107, signal_3105}), .b ({signal_2303, signal_1543}), .c ({signal_2337, signal_1581}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1394 ( .a ({signal_3111, signal_3109}), .b ({signal_2285, signal_1545}), .c ({signal_2320, signal_1582}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1395 ( .a ({signal_3115, signal_3113}), .b ({signal_2287, signal_1547}), .c ({signal_2321, signal_1583}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1396 ( .a ({signal_3119, signal_3117}), .b ({signal_2305, signal_1549}), .c ({signal_2338, signal_1584}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1397 ( .a ({signal_3123, signal_3121}), .b ({signal_2307, signal_1551}), .c ({signal_2339, signal_1585}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1398 ( .a ({signal_3127, signal_3125}), .b ({signal_2289, signal_1553}), .c ({signal_2322, signal_1586}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1399 ( .a ({signal_3131, signal_3129}), .b ({signal_2291, signal_1555}), .c ({signal_2323, signal_1587}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1400 ( .a ({signal_2332, signal_1572}), .b ({signal_2356, signal_1588}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1401 ( .a ({signal_2333, signal_1573}), .b ({signal_2357, signal_1589}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1402 ( .a ({signal_2316, signal_1574}), .b ({signal_2340, signal_1590}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1403 ( .a ({signal_2317, signal_1575}), .b ({signal_2341, signal_1591}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1404 ( .a ({signal_2334, signal_1576}), .b ({signal_2358, signal_1592}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1405 ( .a ({signal_2335, signal_1577}), .b ({signal_2359, signal_1593}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1406 ( .a ({signal_2318, signal_1578}), .b ({signal_2342, signal_1594}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1407 ( .a ({signal_2319, signal_1579}), .b ({signal_2343, signal_1595}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1408 ( .a ({signal_2336, signal_1580}), .b ({signal_2360, signal_1596}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1409 ( .a ({signal_2337, signal_1581}), .b ({signal_2361, signal_1597}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1410 ( .a ({signal_2320, signal_1582}), .b ({signal_2344, signal_1598}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1411 ( .a ({signal_2321, signal_1583}), .b ({signal_2345, signal_1599}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1412 ( .a ({signal_2338, signal_1584}), .b ({signal_2362, signal_1600}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1413 ( .a ({signal_2339, signal_1585}), .b ({signal_2363, signal_1601}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1414 ( .a ({signal_2322, signal_1586}), .b ({signal_2346, signal_1602}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1415 ( .a ({signal_2323, signal_1587}), .b ({signal_2347, signal_1603}) ) ;
    buf_clk cell_1529 ( .C (CLK), .D (signal_2940), .Q (signal_2941) ) ;
    buf_clk cell_1531 ( .C (CLK), .D (signal_2942), .Q (signal_2943) ) ;
    buf_clk cell_1533 ( .C (CLK), .D (signal_2944), .Q (signal_2945) ) ;
    buf_clk cell_1535 ( .C (CLK), .D (signal_2946), .Q (signal_2947) ) ;
    buf_clk cell_1537 ( .C (CLK), .D (signal_2948), .Q (signal_2949) ) ;
    buf_clk cell_1539 ( .C (CLK), .D (signal_2950), .Q (signal_2951) ) ;
    buf_clk cell_1541 ( .C (CLK), .D (signal_2952), .Q (signal_2953) ) ;
    buf_clk cell_1543 ( .C (CLK), .D (signal_2954), .Q (signal_2955) ) ;
    buf_clk cell_1545 ( .C (CLK), .D (signal_2956), .Q (signal_2957) ) ;
    buf_clk cell_1547 ( .C (CLK), .D (signal_2958), .Q (signal_2959) ) ;
    buf_clk cell_1549 ( .C (CLK), .D (signal_2960), .Q (signal_2961) ) ;
    buf_clk cell_1551 ( .C (CLK), .D (signal_2962), .Q (signal_2963) ) ;
    buf_clk cell_1553 ( .C (CLK), .D (signal_2964), .Q (signal_2965) ) ;
    buf_clk cell_1555 ( .C (CLK), .D (signal_2966), .Q (signal_2967) ) ;
    buf_clk cell_1557 ( .C (CLK), .D (signal_2968), .Q (signal_2969) ) ;
    buf_clk cell_1559 ( .C (CLK), .D (signal_2970), .Q (signal_2971) ) ;
    buf_clk cell_1561 ( .C (CLK), .D (signal_2972), .Q (signal_2973) ) ;
    buf_clk cell_1563 ( .C (CLK), .D (signal_2974), .Q (signal_2975) ) ;
    buf_clk cell_1565 ( .C (CLK), .D (signal_2976), .Q (signal_2977) ) ;
    buf_clk cell_1567 ( .C (CLK), .D (signal_2978), .Q (signal_2979) ) ;
    buf_clk cell_1569 ( .C (CLK), .D (signal_2980), .Q (signal_2981) ) ;
    buf_clk cell_1571 ( .C (CLK), .D (signal_2982), .Q (signal_2983) ) ;
    buf_clk cell_1573 ( .C (CLK), .D (signal_2984), .Q (signal_2985) ) ;
    buf_clk cell_1575 ( .C (CLK), .D (signal_2986), .Q (signal_2987) ) ;
    buf_clk cell_1577 ( .C (CLK), .D (signal_2988), .Q (signal_2989) ) ;
    buf_clk cell_1579 ( .C (CLK), .D (signal_2990), .Q (signal_2991) ) ;
    buf_clk cell_1581 ( .C (CLK), .D (signal_2992), .Q (signal_2993) ) ;
    buf_clk cell_1583 ( .C (CLK), .D (signal_2994), .Q (signal_2995) ) ;
    buf_clk cell_1585 ( .C (CLK), .D (signal_2996), .Q (signal_2997) ) ;
    buf_clk cell_1587 ( .C (CLK), .D (signal_2998), .Q (signal_2999) ) ;
    buf_clk cell_1589 ( .C (CLK), .D (signal_3000), .Q (signal_3001) ) ;
    buf_clk cell_1591 ( .C (CLK), .D (signal_3002), .Q (signal_3003) ) ;
    buf_clk cell_1593 ( .C (CLK), .D (signal_3004), .Q (signal_3005) ) ;
    buf_clk cell_1595 ( .C (CLK), .D (signal_3006), .Q (signal_3007) ) ;
    buf_clk cell_1597 ( .C (CLK), .D (signal_3008), .Q (signal_3009) ) ;
    buf_clk cell_1599 ( .C (CLK), .D (signal_3010), .Q (signal_3011) ) ;
    buf_clk cell_1601 ( .C (CLK), .D (signal_3012), .Q (signal_3013) ) ;
    buf_clk cell_1603 ( .C (CLK), .D (signal_3014), .Q (signal_3015) ) ;
    buf_clk cell_1605 ( .C (CLK), .D (signal_3016), .Q (signal_3017) ) ;
    buf_clk cell_1607 ( .C (CLK), .D (signal_3018), .Q (signal_3019) ) ;
    buf_clk cell_1609 ( .C (CLK), .D (signal_3020), .Q (signal_3021) ) ;
    buf_clk cell_1611 ( .C (CLK), .D (signal_3022), .Q (signal_3023) ) ;
    buf_clk cell_1613 ( .C (CLK), .D (signal_3024), .Q (signal_3025) ) ;
    buf_clk cell_1615 ( .C (CLK), .D (signal_3026), .Q (signal_3027) ) ;
    buf_clk cell_1617 ( .C (CLK), .D (signal_3028), .Q (signal_3029) ) ;
    buf_clk cell_1619 ( .C (CLK), .D (signal_3030), .Q (signal_3031) ) ;
    buf_clk cell_1621 ( .C (CLK), .D (signal_3032), .Q (signal_3033) ) ;
    buf_clk cell_1623 ( .C (CLK), .D (signal_3034), .Q (signal_3035) ) ;
    buf_clk cell_1625 ( .C (CLK), .D (signal_3036), .Q (signal_3037) ) ;
    buf_clk cell_1627 ( .C (CLK), .D (signal_3038), .Q (signal_3039) ) ;
    buf_clk cell_1629 ( .C (CLK), .D (signal_3040), .Q (signal_3041) ) ;
    buf_clk cell_1631 ( .C (CLK), .D (signal_3042), .Q (signal_3043) ) ;
    buf_clk cell_1633 ( .C (CLK), .D (signal_3044), .Q (signal_3045) ) ;
    buf_clk cell_1635 ( .C (CLK), .D (signal_3046), .Q (signal_3047) ) ;
    buf_clk cell_1637 ( .C (CLK), .D (signal_3048), .Q (signal_3049) ) ;
    buf_clk cell_1639 ( .C (CLK), .D (signal_3050), .Q (signal_3051) ) ;
    buf_clk cell_1641 ( .C (CLK), .D (signal_3052), .Q (signal_3053) ) ;
    buf_clk cell_1643 ( .C (CLK), .D (signal_3054), .Q (signal_3055) ) ;
    buf_clk cell_1645 ( .C (CLK), .D (signal_3056), .Q (signal_3057) ) ;
    buf_clk cell_1647 ( .C (CLK), .D (signal_3058), .Q (signal_3059) ) ;
    buf_clk cell_1649 ( .C (CLK), .D (signal_3060), .Q (signal_3061) ) ;
    buf_clk cell_1651 ( .C (CLK), .D (signal_3062), .Q (signal_3063) ) ;
    buf_clk cell_1653 ( .C (CLK), .D (signal_3064), .Q (signal_3065) ) ;
    buf_clk cell_1655 ( .C (CLK), .D (signal_3066), .Q (signal_3067) ) ;
    buf_clk cell_1657 ( .C (CLK), .D (signal_3068), .Q (signal_3069) ) ;
    buf_clk cell_1659 ( .C (CLK), .D (signal_3070), .Q (signal_3071) ) ;
    buf_clk cell_1661 ( .C (CLK), .D (signal_3072), .Q (signal_3073) ) ;
    buf_clk cell_1663 ( .C (CLK), .D (signal_3074), .Q (signal_3075) ) ;
    buf_clk cell_1665 ( .C (CLK), .D (signal_3076), .Q (signal_3077) ) ;
    buf_clk cell_1667 ( .C (CLK), .D (signal_3078), .Q (signal_3079) ) ;
    buf_clk cell_1669 ( .C (CLK), .D (signal_3080), .Q (signal_3081) ) ;
    buf_clk cell_1671 ( .C (CLK), .D (signal_3082), .Q (signal_3083) ) ;
    buf_clk cell_1673 ( .C (CLK), .D (signal_3084), .Q (signal_3085) ) ;
    buf_clk cell_1675 ( .C (CLK), .D (signal_3086), .Q (signal_3087) ) ;
    buf_clk cell_1677 ( .C (CLK), .D (signal_3088), .Q (signal_3089) ) ;
    buf_clk cell_1679 ( .C (CLK), .D (signal_3090), .Q (signal_3091) ) ;
    buf_clk cell_1681 ( .C (CLK), .D (signal_3092), .Q (signal_3093) ) ;
    buf_clk cell_1683 ( .C (CLK), .D (signal_3094), .Q (signal_3095) ) ;
    buf_clk cell_1685 ( .C (CLK), .D (signal_3096), .Q (signal_3097) ) ;
    buf_clk cell_1687 ( .C (CLK), .D (signal_3098), .Q (signal_3099) ) ;
    buf_clk cell_1689 ( .C (CLK), .D (signal_3100), .Q (signal_3101) ) ;
    buf_clk cell_1691 ( .C (CLK), .D (signal_3102), .Q (signal_3103) ) ;
    buf_clk cell_1693 ( .C (CLK), .D (signal_3104), .Q (signal_3105) ) ;
    buf_clk cell_1695 ( .C (CLK), .D (signal_3106), .Q (signal_3107) ) ;
    buf_clk cell_1697 ( .C (CLK), .D (signal_3108), .Q (signal_3109) ) ;
    buf_clk cell_1699 ( .C (CLK), .D (signal_3110), .Q (signal_3111) ) ;
    buf_clk cell_1701 ( .C (CLK), .D (signal_3112), .Q (signal_3113) ) ;
    buf_clk cell_1703 ( .C (CLK), .D (signal_3114), .Q (signal_3115) ) ;
    buf_clk cell_1705 ( .C (CLK), .D (signal_3116), .Q (signal_3117) ) ;
    buf_clk cell_1707 ( .C (CLK), .D (signal_3118), .Q (signal_3119) ) ;
    buf_clk cell_1709 ( .C (CLK), .D (signal_3120), .Q (signal_3121) ) ;
    buf_clk cell_1711 ( .C (CLK), .D (signal_3122), .Q (signal_3123) ) ;
    buf_clk cell_1713 ( .C (CLK), .D (signal_3124), .Q (signal_3125) ) ;
    buf_clk cell_1715 ( .C (CLK), .D (signal_3126), .Q (signal_3127) ) ;
    buf_clk cell_1717 ( .C (CLK), .D (signal_3128), .Q (signal_3129) ) ;
    buf_clk cell_1719 ( .C (CLK), .D (signal_3130), .Q (signal_3131) ) ;
    buf_clk cell_1721 ( .C (CLK), .D (signal_3132), .Q (signal_3133) ) ;
    buf_clk cell_1725 ( .C (CLK), .D (signal_3136), .Q (signal_3137) ) ;
    buf_clk cell_1729 ( .C (CLK), .D (signal_3140), .Q (signal_3141) ) ;
    buf_clk cell_1733 ( .C (CLK), .D (signal_3144), .Q (signal_3145) ) ;
    buf_clk cell_1737 ( .C (CLK), .D (signal_3148), .Q (signal_3149) ) ;
    buf_clk cell_1741 ( .C (CLK), .D (signal_3152), .Q (signal_3153) ) ;
    buf_clk cell_1745 ( .C (CLK), .D (signal_3156), .Q (signal_3157) ) ;
    buf_clk cell_1749 ( .C (CLK), .D (signal_3160), .Q (signal_3161) ) ;
    buf_clk cell_1753 ( .C (CLK), .D (signal_3164), .Q (signal_3165) ) ;
    buf_clk cell_1757 ( .C (CLK), .D (signal_3168), .Q (signal_3169) ) ;
    buf_clk cell_1761 ( .C (CLK), .D (signal_3172), .Q (signal_3173) ) ;
    buf_clk cell_1765 ( .C (CLK), .D (signal_3176), .Q (signal_3177) ) ;
    buf_clk cell_1769 ( .C (CLK), .D (signal_3180), .Q (signal_3181) ) ;
    buf_clk cell_1773 ( .C (CLK), .D (signal_3184), .Q (signal_3185) ) ;
    buf_clk cell_1777 ( .C (CLK), .D (signal_3188), .Q (signal_3189) ) ;
    buf_clk cell_1781 ( .C (CLK), .D (signal_3192), .Q (signal_3193) ) ;
    buf_clk cell_1785 ( .C (CLK), .D (signal_3196), .Q (signal_3197) ) ;
    buf_clk cell_1789 ( .C (CLK), .D (signal_3200), .Q (signal_3201) ) ;
    buf_clk cell_1793 ( .C (CLK), .D (signal_3204), .Q (signal_3205) ) ;
    buf_clk cell_1797 ( .C (CLK), .D (signal_3208), .Q (signal_3209) ) ;
    buf_clk cell_1801 ( .C (CLK), .D (signal_3212), .Q (signal_3213) ) ;
    buf_clk cell_1805 ( .C (CLK), .D (signal_3216), .Q (signal_3217) ) ;
    buf_clk cell_1809 ( .C (CLK), .D (signal_3220), .Q (signal_3221) ) ;
    buf_clk cell_1813 ( .C (CLK), .D (signal_3224), .Q (signal_3225) ) ;
    buf_clk cell_1817 ( .C (CLK), .D (signal_3228), .Q (signal_3229) ) ;
    buf_clk cell_1821 ( .C (CLK), .D (signal_3232), .Q (signal_3233) ) ;
    buf_clk cell_1825 ( .C (CLK), .D (signal_3236), .Q (signal_3237) ) ;
    buf_clk cell_1829 ( .C (CLK), .D (signal_3240), .Q (signal_3241) ) ;
    buf_clk cell_1833 ( .C (CLK), .D (signal_3244), .Q (signal_3245) ) ;
    buf_clk cell_1837 ( .C (CLK), .D (signal_3248), .Q (signal_3249) ) ;
    buf_clk cell_1841 ( .C (CLK), .D (signal_3252), .Q (signal_3253) ) ;
    buf_clk cell_1845 ( .C (CLK), .D (signal_3256), .Q (signal_3257) ) ;
    buf_clk cell_1849 ( .C (CLK), .D (signal_3260), .Q (signal_3261) ) ;
    buf_clk cell_1853 ( .C (CLK), .D (signal_3264), .Q (signal_3265) ) ;
    buf_clk cell_1857 ( .C (CLK), .D (signal_3268), .Q (signal_3269) ) ;
    buf_clk cell_1861 ( .C (CLK), .D (signal_3272), .Q (signal_3273) ) ;
    buf_clk cell_1865 ( .C (CLK), .D (signal_3276), .Q (signal_3277) ) ;
    buf_clk cell_1869 ( .C (CLK), .D (signal_3280), .Q (signal_3281) ) ;
    buf_clk cell_1873 ( .C (CLK), .D (signal_3284), .Q (signal_3285) ) ;
    buf_clk cell_1877 ( .C (CLK), .D (signal_3288), .Q (signal_3289) ) ;
    buf_clk cell_1881 ( .C (CLK), .D (signal_3292), .Q (signal_3293) ) ;
    buf_clk cell_1885 ( .C (CLK), .D (signal_3296), .Q (signal_3297) ) ;
    buf_clk cell_1889 ( .C (CLK), .D (signal_3300), .Q (signal_3301) ) ;
    buf_clk cell_1893 ( .C (CLK), .D (signal_3304), .Q (signal_3305) ) ;
    buf_clk cell_1897 ( .C (CLK), .D (signal_3308), .Q (signal_3309) ) ;
    buf_clk cell_1901 ( .C (CLK), .D (signal_3312), .Q (signal_3313) ) ;
    buf_clk cell_1905 ( .C (CLK), .D (signal_3316), .Q (signal_3317) ) ;
    buf_clk cell_1909 ( .C (CLK), .D (signal_3320), .Q (signal_3321) ) ;
    buf_clk cell_1913 ( .C (CLK), .D (signal_3324), .Q (signal_3325) ) ;
    buf_clk cell_1917 ( .C (CLK), .D (signal_3328), .Q (signal_3329) ) ;
    buf_clk cell_1921 ( .C (CLK), .D (signal_3332), .Q (signal_3333) ) ;
    buf_clk cell_1925 ( .C (CLK), .D (signal_3336), .Q (signal_3337) ) ;
    buf_clk cell_1929 ( .C (CLK), .D (signal_3340), .Q (signal_3341) ) ;
    buf_clk cell_1933 ( .C (CLK), .D (signal_3344), .Q (signal_3345) ) ;
    buf_clk cell_1937 ( .C (CLK), .D (signal_3348), .Q (signal_3349) ) ;
    buf_clk cell_1941 ( .C (CLK), .D (signal_3352), .Q (signal_3353) ) ;
    buf_clk cell_1945 ( .C (CLK), .D (signal_3356), .Q (signal_3357) ) ;
    buf_clk cell_1949 ( .C (CLK), .D (signal_3360), .Q (signal_3361) ) ;
    buf_clk cell_1953 ( .C (CLK), .D (signal_3364), .Q (signal_3365) ) ;
    buf_clk cell_1957 ( .C (CLK), .D (signal_3368), .Q (signal_3369) ) ;
    buf_clk cell_1961 ( .C (CLK), .D (signal_3372), .Q (signal_3373) ) ;
    buf_clk cell_1965 ( .C (CLK), .D (signal_3376), .Q (signal_3377) ) ;
    buf_clk cell_1969 ( .C (CLK), .D (signal_3380), .Q (signal_3381) ) ;
    buf_clk cell_1973 ( .C (CLK), .D (signal_3384), .Q (signal_3385) ) ;
    buf_clk cell_1977 ( .C (CLK), .D (signal_3388), .Q (signal_3389) ) ;
    buf_clk cell_1981 ( .C (CLK), .D (signal_3392), .Q (signal_3393) ) ;
    buf_clk cell_1985 ( .C (CLK), .D (signal_3396), .Q (signal_3397) ) ;
    buf_clk cell_1989 ( .C (CLK), .D (signal_3400), .Q (signal_3401) ) ;
    buf_clk cell_1993 ( .C (CLK), .D (signal_3404), .Q (signal_3405) ) ;
    buf_clk cell_1997 ( .C (CLK), .D (signal_3408), .Q (signal_3409) ) ;
    buf_clk cell_2001 ( .C (CLK), .D (signal_3412), .Q (signal_3413) ) ;
    buf_clk cell_2005 ( .C (CLK), .D (signal_3416), .Q (signal_3417) ) ;
    buf_clk cell_2009 ( .C (CLK), .D (signal_3420), .Q (signal_3421) ) ;
    buf_clk cell_2013 ( .C (CLK), .D (signal_3424), .Q (signal_3425) ) ;
    buf_clk cell_2017 ( .C (CLK), .D (signal_3428), .Q (signal_3429) ) ;
    buf_clk cell_2021 ( .C (CLK), .D (signal_3432), .Q (signal_3433) ) ;
    buf_clk cell_2025 ( .C (CLK), .D (signal_3436), .Q (signal_3437) ) ;
    buf_clk cell_2029 ( .C (CLK), .D (signal_3440), .Q (signal_3441) ) ;
    buf_clk cell_2033 ( .C (CLK), .D (signal_3444), .Q (signal_3445) ) ;
    buf_clk cell_2037 ( .C (CLK), .D (signal_3448), .Q (signal_3449) ) ;
    buf_clk cell_2041 ( .C (CLK), .D (signal_3452), .Q (signal_3453) ) ;
    buf_clk cell_2045 ( .C (CLK), .D (signal_3456), .Q (signal_3457) ) ;
    buf_clk cell_2049 ( .C (CLK), .D (signal_3460), .Q (signal_3461) ) ;
    buf_clk cell_2053 ( .C (CLK), .D (signal_3464), .Q (signal_3465) ) ;
    buf_clk cell_2057 ( .C (CLK), .D (signal_3468), .Q (signal_3469) ) ;
    buf_clk cell_2061 ( .C (CLK), .D (signal_3472), .Q (signal_3473) ) ;
    buf_clk cell_2065 ( .C (CLK), .D (signal_3476), .Q (signal_3477) ) ;
    buf_clk cell_2069 ( .C (CLK), .D (signal_3480), .Q (signal_3481) ) ;
    buf_clk cell_2073 ( .C (CLK), .D (signal_3484), .Q (signal_3485) ) ;
    buf_clk cell_2077 ( .C (CLK), .D (signal_3488), .Q (signal_3489) ) ;
    buf_clk cell_2081 ( .C (CLK), .D (signal_3492), .Q (signal_3493) ) ;
    buf_clk cell_2085 ( .C (CLK), .D (signal_3496), .Q (signal_3497) ) ;
    buf_clk cell_2089 ( .C (CLK), .D (signal_3500), .Q (signal_3501) ) ;
    buf_clk cell_2093 ( .C (CLK), .D (signal_3504), .Q (signal_3505) ) ;
    buf_clk cell_2097 ( .C (CLK), .D (signal_3508), .Q (signal_3509) ) ;
    buf_clk cell_2101 ( .C (CLK), .D (signal_3512), .Q (signal_3513) ) ;
    buf_clk cell_2105 ( .C (CLK), .D (signal_3516), .Q (signal_3517) ) ;
    buf_clk cell_2109 ( .C (CLK), .D (signal_3520), .Q (signal_3521) ) ;
    buf_clk cell_2113 ( .C (CLK), .D (signal_3524), .Q (signal_3525) ) ;
    buf_clk cell_2117 ( .C (CLK), .D (signal_3528), .Q (signal_3529) ) ;
    buf_clk cell_2121 ( .C (CLK), .D (signal_3532), .Q (signal_3533) ) ;
    buf_clk cell_2125 ( .C (CLK), .D (signal_3536), .Q (signal_3537) ) ;
    buf_clk cell_2129 ( .C (CLK), .D (signal_3540), .Q (signal_3541) ) ;
    buf_clk cell_2133 ( .C (CLK), .D (signal_3544), .Q (signal_3545) ) ;
    buf_clk cell_2137 ( .C (CLK), .D (signal_3548), .Q (signal_3549) ) ;
    buf_clk cell_2141 ( .C (CLK), .D (signal_3552), .Q (signal_3553) ) ;
    buf_clk cell_2145 ( .C (CLK), .D (signal_3556), .Q (signal_3557) ) ;
    buf_clk cell_2149 ( .C (CLK), .D (signal_3560), .Q (signal_3561) ) ;
    buf_clk cell_2153 ( .C (CLK), .D (signal_3564), .Q (signal_3565) ) ;
    buf_clk cell_2157 ( .C (CLK), .D (signal_3568), .Q (signal_3569) ) ;
    buf_clk cell_2161 ( .C (CLK), .D (signal_3572), .Q (signal_3573) ) ;
    buf_clk cell_2165 ( .C (CLK), .D (signal_3576), .Q (signal_3577) ) ;
    buf_clk cell_2169 ( .C (CLK), .D (signal_3580), .Q (signal_3581) ) ;
    buf_clk cell_2173 ( .C (CLK), .D (signal_3584), .Q (signal_3585) ) ;
    buf_clk cell_2177 ( .C (CLK), .D (signal_3588), .Q (signal_3589) ) ;
    buf_clk cell_2181 ( .C (CLK), .D (signal_3592), .Q (signal_3593) ) ;
    buf_clk cell_2185 ( .C (CLK), .D (signal_3596), .Q (signal_3597) ) ;
    buf_clk cell_2189 ( .C (CLK), .D (signal_3600), .Q (signal_3601) ) ;
    buf_clk cell_2193 ( .C (CLK), .D (signal_3604), .Q (signal_3605) ) ;
    buf_clk cell_2197 ( .C (CLK), .D (signal_3608), .Q (signal_3609) ) ;
    buf_clk cell_2201 ( .C (CLK), .D (signal_3612), .Q (signal_3613) ) ;
    buf_clk cell_2205 ( .C (CLK), .D (signal_3616), .Q (signal_3617) ) ;
    buf_clk cell_2209 ( .C (CLK), .D (signal_3620), .Q (signal_3621) ) ;
    buf_clk cell_2213 ( .C (CLK), .D (signal_3624), .Q (signal_3625) ) ;
    buf_clk cell_2217 ( .C (CLK), .D (signal_3628), .Q (signal_3629) ) ;
    buf_clk cell_2221 ( .C (CLK), .D (signal_3632), .Q (signal_3633) ) ;
    buf_clk cell_2225 ( .C (CLK), .D (signal_3636), .Q (signal_3637) ) ;
    buf_clk cell_2229 ( .C (CLK), .D (signal_3640), .Q (signal_3641) ) ;
    buf_clk cell_2233 ( .C (CLK), .D (signal_3644), .Q (signal_3645) ) ;
    buf_clk cell_2237 ( .C (CLK), .D (signal_3648), .Q (signal_3649) ) ;
    buf_clk cell_2241 ( .C (CLK), .D (signal_3652), .Q (signal_3653) ) ;
    buf_clk cell_2245 ( .C (CLK), .D (signal_3656), .Q (signal_3657) ) ;
    buf_clk cell_2249 ( .C (CLK), .D (signal_3660), .Q (signal_3661) ) ;
    buf_clk cell_2253 ( .C (CLK), .D (signal_3664), .Q (signal_3665) ) ;
    buf_clk cell_2257 ( .C (CLK), .D (signal_3668), .Q (signal_3669) ) ;
    buf_clk cell_2261 ( .C (CLK), .D (signal_3672), .Q (signal_3673) ) ;
    buf_clk cell_2265 ( .C (CLK), .D (signal_3676), .Q (signal_3677) ) ;
    buf_clk cell_2269 ( .C (CLK), .D (signal_3680), .Q (signal_3681) ) ;
    buf_clk cell_2273 ( .C (CLK), .D (signal_3684), .Q (signal_3685) ) ;
    buf_clk cell_2277 ( .C (CLK), .D (signal_3688), .Q (signal_3689) ) ;
    buf_clk cell_2281 ( .C (CLK), .D (signal_3692), .Q (signal_3693) ) ;
    buf_clk cell_2285 ( .C (CLK), .D (signal_3696), .Q (signal_3697) ) ;
    buf_clk cell_2289 ( .C (CLK), .D (signal_3700), .Q (signal_3701) ) ;
    buf_clk cell_2293 ( .C (CLK), .D (signal_3704), .Q (signal_3705) ) ;
    buf_clk cell_2297 ( .C (CLK), .D (signal_3708), .Q (signal_3709) ) ;
    buf_clk cell_2301 ( .C (CLK), .D (signal_3712), .Q (signal_3713) ) ;
    buf_clk cell_2305 ( .C (CLK), .D (signal_3716), .Q (signal_3717) ) ;
    buf_clk cell_2309 ( .C (CLK), .D (signal_3720), .Q (signal_3721) ) ;
    buf_clk cell_2313 ( .C (CLK), .D (signal_3724), .Q (signal_3725) ) ;
    buf_clk cell_2317 ( .C (CLK), .D (signal_3728), .Q (signal_3729) ) ;
    buf_clk cell_2321 ( .C (CLK), .D (signal_3732), .Q (signal_3733) ) ;
    buf_clk cell_2325 ( .C (CLK), .D (signal_3736), .Q (signal_3737) ) ;
    buf_clk cell_2329 ( .C (CLK), .D (signal_3740), .Q (signal_3741) ) ;
    buf_clk cell_2333 ( .C (CLK), .D (signal_3744), .Q (signal_3745) ) ;
    buf_clk cell_2337 ( .C (CLK), .D (signal_3748), .Q (signal_3749) ) ;
    buf_clk cell_2341 ( .C (CLK), .D (signal_3752), .Q (signal_3753) ) ;
    buf_clk cell_2345 ( .C (CLK), .D (signal_3756), .Q (signal_3757) ) ;
    buf_clk cell_2349 ( .C (CLK), .D (signal_3760), .Q (signal_3761) ) ;
    buf_clk cell_2353 ( .C (CLK), .D (signal_3764), .Q (signal_3765) ) ;
    buf_clk cell_2357 ( .C (CLK), .D (signal_3768), .Q (signal_3769) ) ;
    buf_clk cell_2361 ( .C (CLK), .D (signal_3772), .Q (signal_3773) ) ;
    buf_clk cell_2365 ( .C (CLK), .D (signal_3776), .Q (signal_3777) ) ;
    buf_clk cell_2369 ( .C (CLK), .D (signal_3780), .Q (signal_3781) ) ;
    buf_clk cell_2373 ( .C (CLK), .D (signal_3784), .Q (signal_3785) ) ;
    buf_clk cell_2377 ( .C (CLK), .D (signal_3788), .Q (signal_3789) ) ;
    buf_clk cell_2381 ( .C (CLK), .D (signal_3792), .Q (signal_3793) ) ;
    buf_clk cell_2385 ( .C (CLK), .D (signal_3796), .Q (signal_3797) ) ;
    buf_clk cell_2389 ( .C (CLK), .D (signal_3800), .Q (signal_3801) ) ;
    buf_clk cell_2393 ( .C (CLK), .D (signal_3804), .Q (signal_3805) ) ;
    buf_clk cell_2397 ( .C (CLK), .D (signal_3808), .Q (signal_3809) ) ;
    buf_clk cell_2401 ( .C (CLK), .D (signal_3812), .Q (signal_3813) ) ;
    buf_clk cell_2405 ( .C (CLK), .D (signal_3816), .Q (signal_3817) ) ;
    buf_clk cell_2409 ( .C (CLK), .D (signal_3820), .Q (signal_3821) ) ;
    buf_clk cell_2413 ( .C (CLK), .D (signal_3824), .Q (signal_3825) ) ;
    buf_clk cell_2417 ( .C (CLK), .D (signal_3828), .Q (signal_3829) ) ;
    buf_clk cell_2421 ( .C (CLK), .D (signal_3832), .Q (signal_3833) ) ;
    buf_clk cell_2425 ( .C (CLK), .D (signal_3836), .Q (signal_3837) ) ;
    buf_clk cell_2429 ( .C (CLK), .D (signal_3840), .Q (signal_3841) ) ;
    buf_clk cell_2433 ( .C (CLK), .D (signal_3844), .Q (signal_3845) ) ;
    buf_clk cell_2437 ( .C (CLK), .D (signal_3848), .Q (signal_3849) ) ;
    buf_clk cell_2441 ( .C (CLK), .D (signal_3852), .Q (signal_3853) ) ;
    buf_clk cell_2445 ( .C (CLK), .D (signal_3856), .Q (signal_3857) ) ;
    buf_clk cell_2449 ( .C (CLK), .D (signal_3860), .Q (signal_3861) ) ;
    buf_clk cell_2453 ( .C (CLK), .D (signal_3864), .Q (signal_3865) ) ;
    buf_clk cell_2457 ( .C (CLK), .D (signal_3868), .Q (signal_3869) ) ;
    buf_clk cell_2461 ( .C (CLK), .D (signal_3872), .Q (signal_3873) ) ;
    buf_clk cell_2465 ( .C (CLK), .D (signal_3876), .Q (signal_3877) ) ;
    buf_clk cell_2469 ( .C (CLK), .D (signal_3880), .Q (signal_3881) ) ;
    buf_clk cell_2473 ( .C (CLK), .D (signal_3884), .Q (signal_3885) ) ;
    buf_clk cell_2477 ( .C (CLK), .D (signal_3888), .Q (signal_3889) ) ;
    buf_clk cell_2481 ( .C (CLK), .D (signal_3892), .Q (signal_3893) ) ;
    buf_clk cell_2485 ( .C (CLK), .D (signal_3896), .Q (signal_3897) ) ;
    buf_clk cell_2489 ( .C (CLK), .D (signal_3900), .Q (signal_3901) ) ;
    buf_clk cell_2493 ( .C (CLK), .D (signal_3904), .Q (signal_3905) ) ;
    buf_clk cell_2497 ( .C (CLK), .D (signal_3908), .Q (signal_3909) ) ;
    buf_clk cell_2501 ( .C (CLK), .D (signal_3912), .Q (signal_3913) ) ;
    buf_clk cell_2505 ( .C (CLK), .D (signal_3916), .Q (signal_3917) ) ;
    buf_clk cell_2509 ( .C (CLK), .D (signal_3920), .Q (signal_3921) ) ;
    buf_clk cell_2513 ( .C (CLK), .D (signal_3924), .Q (signal_3925) ) ;
    buf_clk cell_2517 ( .C (CLK), .D (signal_3928), .Q (signal_3929) ) ;
    buf_clk cell_2521 ( .C (CLK), .D (signal_3932), .Q (signal_3933) ) ;
    buf_clk cell_2525 ( .C (CLK), .D (signal_3936), .Q (signal_3937) ) ;
    buf_clk cell_2529 ( .C (CLK), .D (signal_3940), .Q (signal_3941) ) ;
    buf_clk cell_2533 ( .C (CLK), .D (signal_3944), .Q (signal_3945) ) ;
    buf_clk cell_2537 ( .C (CLK), .D (signal_3948), .Q (signal_3949) ) ;
    buf_clk cell_2541 ( .C (CLK), .D (signal_3952), .Q (signal_3953) ) ;
    buf_clk cell_2545 ( .C (CLK), .D (signal_3956), .Q (signal_3957) ) ;
    buf_clk cell_2549 ( .C (CLK), .D (signal_3960), .Q (signal_3961) ) ;
    buf_clk cell_2553 ( .C (CLK), .D (signal_3964), .Q (signal_3965) ) ;
    buf_clk cell_2557 ( .C (CLK), .D (signal_3968), .Q (signal_3969) ) ;
    buf_clk cell_2561 ( .C (CLK), .D (signal_3972), .Q (signal_3973) ) ;
    buf_clk cell_2565 ( .C (CLK), .D (signal_3976), .Q (signal_3977) ) ;
    buf_clk cell_2569 ( .C (CLK), .D (signal_3980), .Q (signal_3981) ) ;
    buf_clk cell_2573 ( .C (CLK), .D (signal_3984), .Q (signal_3985) ) ;
    buf_clk cell_2577 ( .C (CLK), .D (signal_3988), .Q (signal_3989) ) ;
    buf_clk cell_2581 ( .C (CLK), .D (signal_3992), .Q (signal_3993) ) ;
    buf_clk cell_2585 ( .C (CLK), .D (signal_3996), .Q (signal_3997) ) ;
    buf_clk cell_2589 ( .C (CLK), .D (signal_4000), .Q (signal_4001) ) ;
    buf_clk cell_2593 ( .C (CLK), .D (signal_4004), .Q (signal_4005) ) ;
    buf_clk cell_2597 ( .C (CLK), .D (signal_4008), .Q (signal_4009) ) ;
    buf_clk cell_2601 ( .C (CLK), .D (signal_4012), .Q (signal_4013) ) ;
    buf_clk cell_2605 ( .C (CLK), .D (signal_4016), .Q (signal_4017) ) ;
    buf_clk cell_2609 ( .C (CLK), .D (signal_4020), .Q (signal_4021) ) ;
    buf_clk cell_2613 ( .C (CLK), .D (signal_4024), .Q (signal_4025) ) ;
    buf_clk cell_2617 ( .C (CLK), .D (signal_4028), .Q (signal_4029) ) ;
    buf_clk cell_2621 ( .C (CLK), .D (signal_4032), .Q (signal_4033) ) ;
    buf_clk cell_2625 ( .C (CLK), .D (signal_4036), .Q (signal_4037) ) ;
    buf_clk cell_2629 ( .C (CLK), .D (signal_4040), .Q (signal_4041) ) ;
    buf_clk cell_2633 ( .C (CLK), .D (signal_4044), .Q (signal_4045) ) ;
    buf_clk cell_2637 ( .C (CLK), .D (signal_4048), .Q (signal_4049) ) ;
    buf_clk cell_2641 ( .C (CLK), .D (signal_4052), .Q (signal_4053) ) ;
    buf_clk cell_2645 ( .C (CLK), .D (signal_4056), .Q (signal_4057) ) ;
    buf_clk cell_2649 ( .C (CLK), .D (signal_4060), .Q (signal_4061) ) ;
    buf_clk cell_2653 ( .C (CLK), .D (signal_4064), .Q (signal_4065) ) ;
    buf_clk cell_2657 ( .C (CLK), .D (signal_4068), .Q (signal_4069) ) ;
    buf_clk cell_2661 ( .C (CLK), .D (signal_4072), .Q (signal_4073) ) ;
    buf_clk cell_2665 ( .C (CLK), .D (signal_4076), .Q (signal_4077) ) ;
    buf_clk cell_2669 ( .C (CLK), .D (signal_4080), .Q (signal_4081) ) ;
    buf_clk cell_2673 ( .C (CLK), .D (signal_4084), .Q (signal_4085) ) ;
    buf_clk cell_2677 ( .C (CLK), .D (signal_4088), .Q (signal_4089) ) ;
    buf_clk cell_2681 ( .C (CLK), .D (signal_4092), .Q (signal_4093) ) ;
    buf_clk cell_2685 ( .C (CLK), .D (signal_4096), .Q (signal_4097) ) ;
    buf_clk cell_2689 ( .C (CLK), .D (signal_4100), .Q (signal_4101) ) ;
    buf_clk cell_2693 ( .C (CLK), .D (signal_4104), .Q (signal_4105) ) ;
    buf_clk cell_2697 ( .C (CLK), .D (signal_4108), .Q (signal_4109) ) ;
    buf_clk cell_2701 ( .C (CLK), .D (signal_4112), .Q (signal_4113) ) ;
    buf_clk cell_2705 ( .C (CLK), .D (signal_4116), .Q (signal_4117) ) ;
    buf_clk cell_2709 ( .C (CLK), .D (signal_4120), .Q (signal_4121) ) ;
    buf_clk cell_2713 ( .C (CLK), .D (signal_4124), .Q (signal_4125) ) ;
    buf_clk cell_2717 ( .C (CLK), .D (signal_4128), .Q (signal_4129) ) ;
    buf_clk cell_2721 ( .C (CLK), .D (signal_4132), .Q (signal_4133) ) ;
    buf_clk cell_2725 ( .C (CLK), .D (signal_4136), .Q (signal_4137) ) ;
    buf_clk cell_2729 ( .C (CLK), .D (signal_4140), .Q (signal_4141) ) ;
    buf_clk cell_2733 ( .C (CLK), .D (signal_4144), .Q (signal_4145) ) ;
    buf_clk cell_2737 ( .C (CLK), .D (signal_4148), .Q (signal_4149) ) ;
    buf_clk cell_2741 ( .C (CLK), .D (signal_4152), .Q (signal_4153) ) ;
    buf_clk cell_2745 ( .C (CLK), .D (signal_4156), .Q (signal_4157) ) ;
    buf_clk cell_2749 ( .C (CLK), .D (signal_4160), .Q (signal_4161) ) ;
    buf_clk cell_2753 ( .C (CLK), .D (signal_4164), .Q (signal_4165) ) ;
    buf_clk cell_2757 ( .C (CLK), .D (signal_4168), .Q (signal_4169) ) ;
    buf_clk cell_2761 ( .C (CLK), .D (signal_4172), .Q (signal_4173) ) ;
    buf_clk cell_2765 ( .C (CLK), .D (signal_4176), .Q (signal_4177) ) ;
    buf_clk cell_2769 ( .C (CLK), .D (signal_4180), .Q (signal_4181) ) ;
    buf_clk cell_2773 ( .C (CLK), .D (signal_4184), .Q (signal_4185) ) ;
    buf_clk cell_2777 ( .C (CLK), .D (signal_4188), .Q (signal_4189) ) ;
    buf_clk cell_2781 ( .C (CLK), .D (signal_4192), .Q (signal_4193) ) ;
    buf_clk cell_2785 ( .C (CLK), .D (signal_4196), .Q (signal_4197) ) ;
    buf_clk cell_2789 ( .C (CLK), .D (signal_4200), .Q (signal_4201) ) ;
    buf_clk cell_2793 ( .C (CLK), .D (signal_4204), .Q (signal_4205) ) ;
    buf_clk cell_2797 ( .C (CLK), .D (signal_4208), .Q (signal_4209) ) ;
    buf_clk cell_2801 ( .C (CLK), .D (signal_4212), .Q (signal_4213) ) ;
    buf_clk cell_2805 ( .C (CLK), .D (signal_4216), .Q (signal_4217) ) ;
    buf_clk cell_2809 ( .C (CLK), .D (signal_4220), .Q (signal_4221) ) ;
    buf_clk cell_2813 ( .C (CLK), .D (signal_4224), .Q (signal_4225) ) ;
    buf_clk cell_2817 ( .C (CLK), .D (signal_4228), .Q (signal_4229) ) ;
    buf_clk cell_2821 ( .C (CLK), .D (signal_4232), .Q (signal_4233) ) ;
    buf_clk cell_2825 ( .C (CLK), .D (signal_4236), .Q (signal_4237) ) ;
    buf_clk cell_2877 ( .C (CLK), .D (signal_4288), .Q (signal_4289) ) ;
    buf_clk cell_2879 ( .C (CLK), .D (signal_4290), .Q (signal_4291) ) ;
    buf_clk cell_2881 ( .C (CLK), .D (signal_4292), .Q (signal_4293) ) ;
    buf_clk cell_2883 ( .C (CLK), .D (signal_4294), .Q (signal_4295) ) ;
    buf_clk cell_2885 ( .C (CLK), .D (signal_4296), .Q (signal_4297) ) ;
    buf_clk cell_2887 ( .C (CLK), .D (signal_4298), .Q (signal_4299) ) ;
    buf_clk cell_2889 ( .C (CLK), .D (signal_4300), .Q (signal_4301) ) ;
    buf_clk cell_2891 ( .C (CLK), .D (signal_4302), .Q (signal_4303) ) ;
    buf_clk cell_2893 ( .C (CLK), .D (signal_4304), .Q (signal_4305) ) ;
    buf_clk cell_2895 ( .C (CLK), .D (signal_4306), .Q (signal_4307) ) ;
    buf_clk cell_2897 ( .C (CLK), .D (signal_4308), .Q (signal_4309) ) ;
    buf_clk cell_2899 ( .C (CLK), .D (signal_4310), .Q (signal_4311) ) ;
    buf_clk cell_2901 ( .C (CLK), .D (signal_4312), .Q (signal_4313) ) ;
    buf_clk cell_2903 ( .C (CLK), .D (signal_4314), .Q (signal_4315) ) ;
    buf_clk cell_2905 ( .C (CLK), .D (signal_4316), .Q (signal_4317) ) ;
    buf_clk cell_2907 ( .C (CLK), .D (signal_4318), .Q (signal_4319) ) ;
    buf_clk cell_2909 ( .C (CLK), .D (signal_4320), .Q (signal_4321) ) ;
    buf_clk cell_2911 ( .C (CLK), .D (signal_4322), .Q (signal_4323) ) ;
    buf_clk cell_2913 ( .C (CLK), .D (signal_4324), .Q (signal_4325) ) ;
    buf_clk cell_2915 ( .C (CLK), .D (signal_4326), .Q (signal_4327) ) ;
    buf_clk cell_2917 ( .C (CLK), .D (signal_4328), .Q (signal_4329) ) ;
    buf_clk cell_2919 ( .C (CLK), .D (signal_4330), .Q (signal_4331) ) ;
    buf_clk cell_2921 ( .C (CLK), .D (signal_4332), .Q (signal_4333) ) ;
    buf_clk cell_2923 ( .C (CLK), .D (signal_4334), .Q (signal_4335) ) ;
    buf_clk cell_2925 ( .C (CLK), .D (signal_4336), .Q (signal_4337) ) ;
    buf_clk cell_2927 ( .C (CLK), .D (signal_4338), .Q (signal_4339) ) ;
    buf_clk cell_2929 ( .C (CLK), .D (signal_4340), .Q (signal_4341) ) ;
    buf_clk cell_2931 ( .C (CLK), .D (signal_4342), .Q (signal_4343) ) ;
    buf_clk cell_2933 ( .C (CLK), .D (signal_4344), .Q (signal_4345) ) ;
    buf_clk cell_2935 ( .C (CLK), .D (signal_4346), .Q (signal_4347) ) ;
    buf_clk cell_2937 ( .C (CLK), .D (signal_4348), .Q (signal_4349) ) ;
    buf_clk cell_2939 ( .C (CLK), .D (signal_4350), .Q (signal_4351) ) ;
    buf_clk cell_2941 ( .C (CLK), .D (signal_4352), .Q (signal_4353) ) ;
    buf_clk cell_2943 ( .C (CLK), .D (signal_4354), .Q (signal_4355) ) ;
    buf_clk cell_2945 ( .C (CLK), .D (signal_4356), .Q (signal_4357) ) ;
    buf_clk cell_2947 ( .C (CLK), .D (signal_4358), .Q (signal_4359) ) ;
    buf_clk cell_2949 ( .C (CLK), .D (signal_4360), .Q (signal_4361) ) ;
    buf_clk cell_2951 ( .C (CLK), .D (signal_4362), .Q (signal_4363) ) ;
    buf_clk cell_2953 ( .C (CLK), .D (signal_4364), .Q (signal_4365) ) ;
    buf_clk cell_2955 ( .C (CLK), .D (signal_4366), .Q (signal_4367) ) ;
    buf_clk cell_2957 ( .C (CLK), .D (signal_4368), .Q (signal_4369) ) ;
    buf_clk cell_2959 ( .C (CLK), .D (signal_4370), .Q (signal_4371) ) ;
    buf_clk cell_2961 ( .C (CLK), .D (signal_4372), .Q (signal_4373) ) ;
    buf_clk cell_2963 ( .C (CLK), .D (signal_4374), .Q (signal_4375) ) ;
    buf_clk cell_2965 ( .C (CLK), .D (signal_4376), .Q (signal_4377) ) ;
    buf_clk cell_2967 ( .C (CLK), .D (signal_4378), .Q (signal_4379) ) ;
    buf_clk cell_2969 ( .C (CLK), .D (signal_4380), .Q (signal_4381) ) ;
    buf_clk cell_2971 ( .C (CLK), .D (signal_4382), .Q (signal_4383) ) ;
    buf_clk cell_2973 ( .C (CLK), .D (signal_4384), .Q (signal_4385) ) ;
    buf_clk cell_2975 ( .C (CLK), .D (signal_4386), .Q (signal_4387) ) ;
    buf_clk cell_2977 ( .C (CLK), .D (signal_4388), .Q (signal_4389) ) ;
    buf_clk cell_2979 ( .C (CLK), .D (signal_4390), .Q (signal_4391) ) ;
    buf_clk cell_2981 ( .C (CLK), .D (signal_4392), .Q (signal_4393) ) ;
    buf_clk cell_2983 ( .C (CLK), .D (signal_4394), .Q (signal_4395) ) ;
    buf_clk cell_2985 ( .C (CLK), .D (signal_4396), .Q (signal_4397) ) ;
    buf_clk cell_2987 ( .C (CLK), .D (signal_4398), .Q (signal_4399) ) ;
    buf_clk cell_2989 ( .C (CLK), .D (signal_4400), .Q (signal_4401) ) ;
    buf_clk cell_2991 ( .C (CLK), .D (signal_4402), .Q (signal_4403) ) ;
    buf_clk cell_2993 ( .C (CLK), .D (signal_4404), .Q (signal_4405) ) ;
    buf_clk cell_2995 ( .C (CLK), .D (signal_4406), .Q (signal_4407) ) ;
    buf_clk cell_2997 ( .C (CLK), .D (signal_4408), .Q (signal_4409) ) ;
    buf_clk cell_2999 ( .C (CLK), .D (signal_4410), .Q (signal_4411) ) ;
    buf_clk cell_3001 ( .C (CLK), .D (signal_4412), .Q (signal_4413) ) ;
    buf_clk cell_3003 ( .C (CLK), .D (signal_4414), .Q (signal_4415) ) ;
    buf_clk cell_3069 ( .C (CLK), .D (signal_4480), .Q (signal_4481) ) ;
    buf_clk cell_3073 ( .C (CLK), .D (signal_4484), .Q (signal_4485) ) ;
    buf_clk cell_3081 ( .C (CLK), .D (signal_4492), .Q (signal_4493) ) ;
    buf_clk cell_3085 ( .C (CLK), .D (signal_4496), .Q (signal_4497) ) ;
    buf_clk cell_3093 ( .C (CLK), .D (signal_4504), .Q (signal_4505) ) ;
    buf_clk cell_3097 ( .C (CLK), .D (signal_4508), .Q (signal_4509) ) ;
    buf_clk cell_3105 ( .C (CLK), .D (signal_4516), .Q (signal_4517) ) ;
    buf_clk cell_3109 ( .C (CLK), .D (signal_4520), .Q (signal_4521) ) ;
    buf_clk cell_3117 ( .C (CLK), .D (signal_4528), .Q (signal_4529) ) ;
    buf_clk cell_3121 ( .C (CLK), .D (signal_4532), .Q (signal_4533) ) ;
    buf_clk cell_3129 ( .C (CLK), .D (signal_4540), .Q (signal_4541) ) ;
    buf_clk cell_3133 ( .C (CLK), .D (signal_4544), .Q (signal_4545) ) ;
    buf_clk cell_3141 ( .C (CLK), .D (signal_4552), .Q (signal_4553) ) ;
    buf_clk cell_3145 ( .C (CLK), .D (signal_4556), .Q (signal_4557) ) ;
    buf_clk cell_3153 ( .C (CLK), .D (signal_4564), .Q (signal_4565) ) ;
    buf_clk cell_3157 ( .C (CLK), .D (signal_4568), .Q (signal_4569) ) ;
    buf_clk cell_3165 ( .C (CLK), .D (signal_4576), .Q (signal_4577) ) ;
    buf_clk cell_3169 ( .C (CLK), .D (signal_4580), .Q (signal_4581) ) ;
    buf_clk cell_3177 ( .C (CLK), .D (signal_4588), .Q (signal_4589) ) ;
    buf_clk cell_3181 ( .C (CLK), .D (signal_4592), .Q (signal_4593) ) ;
    buf_clk cell_3189 ( .C (CLK), .D (signal_4600), .Q (signal_4601) ) ;
    buf_clk cell_3193 ( .C (CLK), .D (signal_4604), .Q (signal_4605) ) ;
    buf_clk cell_3201 ( .C (CLK), .D (signal_4612), .Q (signal_4613) ) ;
    buf_clk cell_3205 ( .C (CLK), .D (signal_4616), .Q (signal_4617) ) ;
    buf_clk cell_3213 ( .C (CLK), .D (signal_4624), .Q (signal_4625) ) ;
    buf_clk cell_3217 ( .C (CLK), .D (signal_4628), .Q (signal_4629) ) ;
    buf_clk cell_3225 ( .C (CLK), .D (signal_4636), .Q (signal_4637) ) ;
    buf_clk cell_3229 ( .C (CLK), .D (signal_4640), .Q (signal_4641) ) ;
    buf_clk cell_3237 ( .C (CLK), .D (signal_4648), .Q (signal_4649) ) ;
    buf_clk cell_3241 ( .C (CLK), .D (signal_4652), .Q (signal_4653) ) ;
    buf_clk cell_3249 ( .C (CLK), .D (signal_4660), .Q (signal_4661) ) ;
    buf_clk cell_3253 ( .C (CLK), .D (signal_4664), .Q (signal_4665) ) ;
    buf_clk cell_3277 ( .C (CLK), .D (signal_4688), .Q (signal_4689) ) ;
    buf_clk cell_3281 ( .C (CLK), .D (signal_4692), .Q (signal_4693) ) ;
    buf_clk cell_3285 ( .C (CLK), .D (signal_4696), .Q (signal_4697) ) ;
    buf_clk cell_3289 ( .C (CLK), .D (signal_4700), .Q (signal_4701) ) ;
    buf_clk cell_3293 ( .C (CLK), .D (signal_4704), .Q (signal_4705) ) ;
    buf_clk cell_3297 ( .C (CLK), .D (signal_4708), .Q (signal_4709) ) ;
    buf_clk cell_3301 ( .C (CLK), .D (signal_4712), .Q (signal_4713) ) ;
    buf_clk cell_3305 ( .C (CLK), .D (signal_4716), .Q (signal_4717) ) ;
    buf_clk cell_3309 ( .C (CLK), .D (signal_4720), .Q (signal_4721) ) ;
    buf_clk cell_3313 ( .C (CLK), .D (signal_4724), .Q (signal_4725) ) ;
    buf_clk cell_3317 ( .C (CLK), .D (signal_4728), .Q (signal_4729) ) ;

    /* cells in depth 3 */
    buf_clk cell_1722 ( .C (CLK), .D (signal_3133), .Q (signal_3134) ) ;
    buf_clk cell_1726 ( .C (CLK), .D (signal_3137), .Q (signal_3138) ) ;
    buf_clk cell_1730 ( .C (CLK), .D (signal_3141), .Q (signal_3142) ) ;
    buf_clk cell_1734 ( .C (CLK), .D (signal_3145), .Q (signal_3146) ) ;
    buf_clk cell_1738 ( .C (CLK), .D (signal_3149), .Q (signal_3150) ) ;
    buf_clk cell_1742 ( .C (CLK), .D (signal_3153), .Q (signal_3154) ) ;
    buf_clk cell_1746 ( .C (CLK), .D (signal_3157), .Q (signal_3158) ) ;
    buf_clk cell_1750 ( .C (CLK), .D (signal_3161), .Q (signal_3162) ) ;
    buf_clk cell_1754 ( .C (CLK), .D (signal_3165), .Q (signal_3166) ) ;
    buf_clk cell_1758 ( .C (CLK), .D (signal_3169), .Q (signal_3170) ) ;
    buf_clk cell_1762 ( .C (CLK), .D (signal_3173), .Q (signal_3174) ) ;
    buf_clk cell_1766 ( .C (CLK), .D (signal_3177), .Q (signal_3178) ) ;
    buf_clk cell_1770 ( .C (CLK), .D (signal_3181), .Q (signal_3182) ) ;
    buf_clk cell_1774 ( .C (CLK), .D (signal_3185), .Q (signal_3186) ) ;
    buf_clk cell_1778 ( .C (CLK), .D (signal_3189), .Q (signal_3190) ) ;
    buf_clk cell_1782 ( .C (CLK), .D (signal_3193), .Q (signal_3194) ) ;
    buf_clk cell_1786 ( .C (CLK), .D (signal_3197), .Q (signal_3198) ) ;
    buf_clk cell_1790 ( .C (CLK), .D (signal_3201), .Q (signal_3202) ) ;
    buf_clk cell_1794 ( .C (CLK), .D (signal_3205), .Q (signal_3206) ) ;
    buf_clk cell_1798 ( .C (CLK), .D (signal_3209), .Q (signal_3210) ) ;
    buf_clk cell_1802 ( .C (CLK), .D (signal_3213), .Q (signal_3214) ) ;
    buf_clk cell_1806 ( .C (CLK), .D (signal_3217), .Q (signal_3218) ) ;
    buf_clk cell_1810 ( .C (CLK), .D (signal_3221), .Q (signal_3222) ) ;
    buf_clk cell_1814 ( .C (CLK), .D (signal_3225), .Q (signal_3226) ) ;
    buf_clk cell_1818 ( .C (CLK), .D (signal_3229), .Q (signal_3230) ) ;
    buf_clk cell_1822 ( .C (CLK), .D (signal_3233), .Q (signal_3234) ) ;
    buf_clk cell_1826 ( .C (CLK), .D (signal_3237), .Q (signal_3238) ) ;
    buf_clk cell_1830 ( .C (CLK), .D (signal_3241), .Q (signal_3242) ) ;
    buf_clk cell_1834 ( .C (CLK), .D (signal_3245), .Q (signal_3246) ) ;
    buf_clk cell_1838 ( .C (CLK), .D (signal_3249), .Q (signal_3250) ) ;
    buf_clk cell_1842 ( .C (CLK), .D (signal_3253), .Q (signal_3254) ) ;
    buf_clk cell_1846 ( .C (CLK), .D (signal_3257), .Q (signal_3258) ) ;
    buf_clk cell_1850 ( .C (CLK), .D (signal_3261), .Q (signal_3262) ) ;
    buf_clk cell_1854 ( .C (CLK), .D (signal_3265), .Q (signal_3266) ) ;
    buf_clk cell_1858 ( .C (CLK), .D (signal_3269), .Q (signal_3270) ) ;
    buf_clk cell_1862 ( .C (CLK), .D (signal_3273), .Q (signal_3274) ) ;
    buf_clk cell_1866 ( .C (CLK), .D (signal_3277), .Q (signal_3278) ) ;
    buf_clk cell_1870 ( .C (CLK), .D (signal_3281), .Q (signal_3282) ) ;
    buf_clk cell_1874 ( .C (CLK), .D (signal_3285), .Q (signal_3286) ) ;
    buf_clk cell_1878 ( .C (CLK), .D (signal_3289), .Q (signal_3290) ) ;
    buf_clk cell_1882 ( .C (CLK), .D (signal_3293), .Q (signal_3294) ) ;
    buf_clk cell_1886 ( .C (CLK), .D (signal_3297), .Q (signal_3298) ) ;
    buf_clk cell_1890 ( .C (CLK), .D (signal_3301), .Q (signal_3302) ) ;
    buf_clk cell_1894 ( .C (CLK), .D (signal_3305), .Q (signal_3306) ) ;
    buf_clk cell_1898 ( .C (CLK), .D (signal_3309), .Q (signal_3310) ) ;
    buf_clk cell_1902 ( .C (CLK), .D (signal_3313), .Q (signal_3314) ) ;
    buf_clk cell_1906 ( .C (CLK), .D (signal_3317), .Q (signal_3318) ) ;
    buf_clk cell_1910 ( .C (CLK), .D (signal_3321), .Q (signal_3322) ) ;
    buf_clk cell_1914 ( .C (CLK), .D (signal_3325), .Q (signal_3326) ) ;
    buf_clk cell_1918 ( .C (CLK), .D (signal_3329), .Q (signal_3330) ) ;
    buf_clk cell_1922 ( .C (CLK), .D (signal_3333), .Q (signal_3334) ) ;
    buf_clk cell_1926 ( .C (CLK), .D (signal_3337), .Q (signal_3338) ) ;
    buf_clk cell_1930 ( .C (CLK), .D (signal_3341), .Q (signal_3342) ) ;
    buf_clk cell_1934 ( .C (CLK), .D (signal_3345), .Q (signal_3346) ) ;
    buf_clk cell_1938 ( .C (CLK), .D (signal_3349), .Q (signal_3350) ) ;
    buf_clk cell_1942 ( .C (CLK), .D (signal_3353), .Q (signal_3354) ) ;
    buf_clk cell_1946 ( .C (CLK), .D (signal_3357), .Q (signal_3358) ) ;
    buf_clk cell_1950 ( .C (CLK), .D (signal_3361), .Q (signal_3362) ) ;
    buf_clk cell_1954 ( .C (CLK), .D (signal_3365), .Q (signal_3366) ) ;
    buf_clk cell_1958 ( .C (CLK), .D (signal_3369), .Q (signal_3370) ) ;
    buf_clk cell_1962 ( .C (CLK), .D (signal_3373), .Q (signal_3374) ) ;
    buf_clk cell_1966 ( .C (CLK), .D (signal_3377), .Q (signal_3378) ) ;
    buf_clk cell_1970 ( .C (CLK), .D (signal_3381), .Q (signal_3382) ) ;
    buf_clk cell_1974 ( .C (CLK), .D (signal_3385), .Q (signal_3386) ) ;
    buf_clk cell_1978 ( .C (CLK), .D (signal_3389), .Q (signal_3390) ) ;
    buf_clk cell_1982 ( .C (CLK), .D (signal_3393), .Q (signal_3394) ) ;
    buf_clk cell_1986 ( .C (CLK), .D (signal_3397), .Q (signal_3398) ) ;
    buf_clk cell_1990 ( .C (CLK), .D (signal_3401), .Q (signal_3402) ) ;
    buf_clk cell_1994 ( .C (CLK), .D (signal_3405), .Q (signal_3406) ) ;
    buf_clk cell_1998 ( .C (CLK), .D (signal_3409), .Q (signal_3410) ) ;
    buf_clk cell_2002 ( .C (CLK), .D (signal_3413), .Q (signal_3414) ) ;
    buf_clk cell_2006 ( .C (CLK), .D (signal_3417), .Q (signal_3418) ) ;
    buf_clk cell_2010 ( .C (CLK), .D (signal_3421), .Q (signal_3422) ) ;
    buf_clk cell_2014 ( .C (CLK), .D (signal_3425), .Q (signal_3426) ) ;
    buf_clk cell_2018 ( .C (CLK), .D (signal_3429), .Q (signal_3430) ) ;
    buf_clk cell_2022 ( .C (CLK), .D (signal_3433), .Q (signal_3434) ) ;
    buf_clk cell_2026 ( .C (CLK), .D (signal_3437), .Q (signal_3438) ) ;
    buf_clk cell_2030 ( .C (CLK), .D (signal_3441), .Q (signal_3442) ) ;
    buf_clk cell_2034 ( .C (CLK), .D (signal_3445), .Q (signal_3446) ) ;
    buf_clk cell_2038 ( .C (CLK), .D (signal_3449), .Q (signal_3450) ) ;
    buf_clk cell_2042 ( .C (CLK), .D (signal_3453), .Q (signal_3454) ) ;
    buf_clk cell_2046 ( .C (CLK), .D (signal_3457), .Q (signal_3458) ) ;
    buf_clk cell_2050 ( .C (CLK), .D (signal_3461), .Q (signal_3462) ) ;
    buf_clk cell_2054 ( .C (CLK), .D (signal_3465), .Q (signal_3466) ) ;
    buf_clk cell_2058 ( .C (CLK), .D (signal_3469), .Q (signal_3470) ) ;
    buf_clk cell_2062 ( .C (CLK), .D (signal_3473), .Q (signal_3474) ) ;
    buf_clk cell_2066 ( .C (CLK), .D (signal_3477), .Q (signal_3478) ) ;
    buf_clk cell_2070 ( .C (CLK), .D (signal_3481), .Q (signal_3482) ) ;
    buf_clk cell_2074 ( .C (CLK), .D (signal_3485), .Q (signal_3486) ) ;
    buf_clk cell_2078 ( .C (CLK), .D (signal_3489), .Q (signal_3490) ) ;
    buf_clk cell_2082 ( .C (CLK), .D (signal_3493), .Q (signal_3494) ) ;
    buf_clk cell_2086 ( .C (CLK), .D (signal_3497), .Q (signal_3498) ) ;
    buf_clk cell_2090 ( .C (CLK), .D (signal_3501), .Q (signal_3502) ) ;
    buf_clk cell_2094 ( .C (CLK), .D (signal_3505), .Q (signal_3506) ) ;
    buf_clk cell_2098 ( .C (CLK), .D (signal_3509), .Q (signal_3510) ) ;
    buf_clk cell_2102 ( .C (CLK), .D (signal_3513), .Q (signal_3514) ) ;
    buf_clk cell_2106 ( .C (CLK), .D (signal_3517), .Q (signal_3518) ) ;
    buf_clk cell_2110 ( .C (CLK), .D (signal_3521), .Q (signal_3522) ) ;
    buf_clk cell_2114 ( .C (CLK), .D (signal_3525), .Q (signal_3526) ) ;
    buf_clk cell_2118 ( .C (CLK), .D (signal_3529), .Q (signal_3530) ) ;
    buf_clk cell_2122 ( .C (CLK), .D (signal_3533), .Q (signal_3534) ) ;
    buf_clk cell_2126 ( .C (CLK), .D (signal_3537), .Q (signal_3538) ) ;
    buf_clk cell_2130 ( .C (CLK), .D (signal_3541), .Q (signal_3542) ) ;
    buf_clk cell_2134 ( .C (CLK), .D (signal_3545), .Q (signal_3546) ) ;
    buf_clk cell_2138 ( .C (CLK), .D (signal_3549), .Q (signal_3550) ) ;
    buf_clk cell_2142 ( .C (CLK), .D (signal_3553), .Q (signal_3554) ) ;
    buf_clk cell_2146 ( .C (CLK), .D (signal_3557), .Q (signal_3558) ) ;
    buf_clk cell_2150 ( .C (CLK), .D (signal_3561), .Q (signal_3562) ) ;
    buf_clk cell_2154 ( .C (CLK), .D (signal_3565), .Q (signal_3566) ) ;
    buf_clk cell_2158 ( .C (CLK), .D (signal_3569), .Q (signal_3570) ) ;
    buf_clk cell_2162 ( .C (CLK), .D (signal_3573), .Q (signal_3574) ) ;
    buf_clk cell_2166 ( .C (CLK), .D (signal_3577), .Q (signal_3578) ) ;
    buf_clk cell_2170 ( .C (CLK), .D (signal_3581), .Q (signal_3582) ) ;
    buf_clk cell_2174 ( .C (CLK), .D (signal_3585), .Q (signal_3586) ) ;
    buf_clk cell_2178 ( .C (CLK), .D (signal_3589), .Q (signal_3590) ) ;
    buf_clk cell_2182 ( .C (CLK), .D (signal_3593), .Q (signal_3594) ) ;
    buf_clk cell_2186 ( .C (CLK), .D (signal_3597), .Q (signal_3598) ) ;
    buf_clk cell_2190 ( .C (CLK), .D (signal_3601), .Q (signal_3602) ) ;
    buf_clk cell_2194 ( .C (CLK), .D (signal_3605), .Q (signal_3606) ) ;
    buf_clk cell_2198 ( .C (CLK), .D (signal_3609), .Q (signal_3610) ) ;
    buf_clk cell_2202 ( .C (CLK), .D (signal_3613), .Q (signal_3614) ) ;
    buf_clk cell_2206 ( .C (CLK), .D (signal_3617), .Q (signal_3618) ) ;
    buf_clk cell_2210 ( .C (CLK), .D (signal_3621), .Q (signal_3622) ) ;
    buf_clk cell_2214 ( .C (CLK), .D (signal_3625), .Q (signal_3626) ) ;
    buf_clk cell_2218 ( .C (CLK), .D (signal_3629), .Q (signal_3630) ) ;
    buf_clk cell_2222 ( .C (CLK), .D (signal_3633), .Q (signal_3634) ) ;
    buf_clk cell_2226 ( .C (CLK), .D (signal_3637), .Q (signal_3638) ) ;
    buf_clk cell_2230 ( .C (CLK), .D (signal_3641), .Q (signal_3642) ) ;
    buf_clk cell_2234 ( .C (CLK), .D (signal_3645), .Q (signal_3646) ) ;
    buf_clk cell_2238 ( .C (CLK), .D (signal_3649), .Q (signal_3650) ) ;
    buf_clk cell_2242 ( .C (CLK), .D (signal_3653), .Q (signal_3654) ) ;
    buf_clk cell_2246 ( .C (CLK), .D (signal_3657), .Q (signal_3658) ) ;
    buf_clk cell_2250 ( .C (CLK), .D (signal_3661), .Q (signal_3662) ) ;
    buf_clk cell_2254 ( .C (CLK), .D (signal_3665), .Q (signal_3666) ) ;
    buf_clk cell_2258 ( .C (CLK), .D (signal_3669), .Q (signal_3670) ) ;
    buf_clk cell_2262 ( .C (CLK), .D (signal_3673), .Q (signal_3674) ) ;
    buf_clk cell_2266 ( .C (CLK), .D (signal_3677), .Q (signal_3678) ) ;
    buf_clk cell_2270 ( .C (CLK), .D (signal_3681), .Q (signal_3682) ) ;
    buf_clk cell_2274 ( .C (CLK), .D (signal_3685), .Q (signal_3686) ) ;
    buf_clk cell_2278 ( .C (CLK), .D (signal_3689), .Q (signal_3690) ) ;
    buf_clk cell_2282 ( .C (CLK), .D (signal_3693), .Q (signal_3694) ) ;
    buf_clk cell_2286 ( .C (CLK), .D (signal_3697), .Q (signal_3698) ) ;
    buf_clk cell_2290 ( .C (CLK), .D (signal_3701), .Q (signal_3702) ) ;
    buf_clk cell_2294 ( .C (CLK), .D (signal_3705), .Q (signal_3706) ) ;
    buf_clk cell_2298 ( .C (CLK), .D (signal_3709), .Q (signal_3710) ) ;
    buf_clk cell_2302 ( .C (CLK), .D (signal_3713), .Q (signal_3714) ) ;
    buf_clk cell_2306 ( .C (CLK), .D (signal_3717), .Q (signal_3718) ) ;
    buf_clk cell_2310 ( .C (CLK), .D (signal_3721), .Q (signal_3722) ) ;
    buf_clk cell_2314 ( .C (CLK), .D (signal_3725), .Q (signal_3726) ) ;
    buf_clk cell_2318 ( .C (CLK), .D (signal_3729), .Q (signal_3730) ) ;
    buf_clk cell_2322 ( .C (CLK), .D (signal_3733), .Q (signal_3734) ) ;
    buf_clk cell_2326 ( .C (CLK), .D (signal_3737), .Q (signal_3738) ) ;
    buf_clk cell_2330 ( .C (CLK), .D (signal_3741), .Q (signal_3742) ) ;
    buf_clk cell_2334 ( .C (CLK), .D (signal_3745), .Q (signal_3746) ) ;
    buf_clk cell_2338 ( .C (CLK), .D (signal_3749), .Q (signal_3750) ) ;
    buf_clk cell_2342 ( .C (CLK), .D (signal_3753), .Q (signal_3754) ) ;
    buf_clk cell_2346 ( .C (CLK), .D (signal_3757), .Q (signal_3758) ) ;
    buf_clk cell_2350 ( .C (CLK), .D (signal_3761), .Q (signal_3762) ) ;
    buf_clk cell_2354 ( .C (CLK), .D (signal_3765), .Q (signal_3766) ) ;
    buf_clk cell_2358 ( .C (CLK), .D (signal_3769), .Q (signal_3770) ) ;
    buf_clk cell_2362 ( .C (CLK), .D (signal_3773), .Q (signal_3774) ) ;
    buf_clk cell_2366 ( .C (CLK), .D (signal_3777), .Q (signal_3778) ) ;
    buf_clk cell_2370 ( .C (CLK), .D (signal_3781), .Q (signal_3782) ) ;
    buf_clk cell_2374 ( .C (CLK), .D (signal_3785), .Q (signal_3786) ) ;
    buf_clk cell_2378 ( .C (CLK), .D (signal_3789), .Q (signal_3790) ) ;
    buf_clk cell_2382 ( .C (CLK), .D (signal_3793), .Q (signal_3794) ) ;
    buf_clk cell_2386 ( .C (CLK), .D (signal_3797), .Q (signal_3798) ) ;
    buf_clk cell_2390 ( .C (CLK), .D (signal_3801), .Q (signal_3802) ) ;
    buf_clk cell_2394 ( .C (CLK), .D (signal_3805), .Q (signal_3806) ) ;
    buf_clk cell_2398 ( .C (CLK), .D (signal_3809), .Q (signal_3810) ) ;
    buf_clk cell_2402 ( .C (CLK), .D (signal_3813), .Q (signal_3814) ) ;
    buf_clk cell_2406 ( .C (CLK), .D (signal_3817), .Q (signal_3818) ) ;
    buf_clk cell_2410 ( .C (CLK), .D (signal_3821), .Q (signal_3822) ) ;
    buf_clk cell_2414 ( .C (CLK), .D (signal_3825), .Q (signal_3826) ) ;
    buf_clk cell_2418 ( .C (CLK), .D (signal_3829), .Q (signal_3830) ) ;
    buf_clk cell_2422 ( .C (CLK), .D (signal_3833), .Q (signal_3834) ) ;
    buf_clk cell_2426 ( .C (CLK), .D (signal_3837), .Q (signal_3838) ) ;
    buf_clk cell_2430 ( .C (CLK), .D (signal_3841), .Q (signal_3842) ) ;
    buf_clk cell_2434 ( .C (CLK), .D (signal_3845), .Q (signal_3846) ) ;
    buf_clk cell_2438 ( .C (CLK), .D (signal_3849), .Q (signal_3850) ) ;
    buf_clk cell_2442 ( .C (CLK), .D (signal_3853), .Q (signal_3854) ) ;
    buf_clk cell_2446 ( .C (CLK), .D (signal_3857), .Q (signal_3858) ) ;
    buf_clk cell_2450 ( .C (CLK), .D (signal_3861), .Q (signal_3862) ) ;
    buf_clk cell_2454 ( .C (CLK), .D (signal_3865), .Q (signal_3866) ) ;
    buf_clk cell_2458 ( .C (CLK), .D (signal_3869), .Q (signal_3870) ) ;
    buf_clk cell_2462 ( .C (CLK), .D (signal_3873), .Q (signal_3874) ) ;
    buf_clk cell_2466 ( .C (CLK), .D (signal_3877), .Q (signal_3878) ) ;
    buf_clk cell_2470 ( .C (CLK), .D (signal_3881), .Q (signal_3882) ) ;
    buf_clk cell_2474 ( .C (CLK), .D (signal_3885), .Q (signal_3886) ) ;
    buf_clk cell_2478 ( .C (CLK), .D (signal_3889), .Q (signal_3890) ) ;
    buf_clk cell_2482 ( .C (CLK), .D (signal_3893), .Q (signal_3894) ) ;
    buf_clk cell_2486 ( .C (CLK), .D (signal_3897), .Q (signal_3898) ) ;
    buf_clk cell_2490 ( .C (CLK), .D (signal_3901), .Q (signal_3902) ) ;
    buf_clk cell_2494 ( .C (CLK), .D (signal_3905), .Q (signal_3906) ) ;
    buf_clk cell_2498 ( .C (CLK), .D (signal_3909), .Q (signal_3910) ) ;
    buf_clk cell_2502 ( .C (CLK), .D (signal_3913), .Q (signal_3914) ) ;
    buf_clk cell_2506 ( .C (CLK), .D (signal_3917), .Q (signal_3918) ) ;
    buf_clk cell_2510 ( .C (CLK), .D (signal_3921), .Q (signal_3922) ) ;
    buf_clk cell_2514 ( .C (CLK), .D (signal_3925), .Q (signal_3926) ) ;
    buf_clk cell_2518 ( .C (CLK), .D (signal_3929), .Q (signal_3930) ) ;
    buf_clk cell_2522 ( .C (CLK), .D (signal_3933), .Q (signal_3934) ) ;
    buf_clk cell_2526 ( .C (CLK), .D (signal_3937), .Q (signal_3938) ) ;
    buf_clk cell_2530 ( .C (CLK), .D (signal_3941), .Q (signal_3942) ) ;
    buf_clk cell_2534 ( .C (CLK), .D (signal_3945), .Q (signal_3946) ) ;
    buf_clk cell_2538 ( .C (CLK), .D (signal_3949), .Q (signal_3950) ) ;
    buf_clk cell_2542 ( .C (CLK), .D (signal_3953), .Q (signal_3954) ) ;
    buf_clk cell_2546 ( .C (CLK), .D (signal_3957), .Q (signal_3958) ) ;
    buf_clk cell_2550 ( .C (CLK), .D (signal_3961), .Q (signal_3962) ) ;
    buf_clk cell_2554 ( .C (CLK), .D (signal_3965), .Q (signal_3966) ) ;
    buf_clk cell_2558 ( .C (CLK), .D (signal_3969), .Q (signal_3970) ) ;
    buf_clk cell_2562 ( .C (CLK), .D (signal_3973), .Q (signal_3974) ) ;
    buf_clk cell_2566 ( .C (CLK), .D (signal_3977), .Q (signal_3978) ) ;
    buf_clk cell_2570 ( .C (CLK), .D (signal_3981), .Q (signal_3982) ) ;
    buf_clk cell_2574 ( .C (CLK), .D (signal_3985), .Q (signal_3986) ) ;
    buf_clk cell_2578 ( .C (CLK), .D (signal_3989), .Q (signal_3990) ) ;
    buf_clk cell_2582 ( .C (CLK), .D (signal_3993), .Q (signal_3994) ) ;
    buf_clk cell_2586 ( .C (CLK), .D (signal_3997), .Q (signal_3998) ) ;
    buf_clk cell_2590 ( .C (CLK), .D (signal_4001), .Q (signal_4002) ) ;
    buf_clk cell_2594 ( .C (CLK), .D (signal_4005), .Q (signal_4006) ) ;
    buf_clk cell_2598 ( .C (CLK), .D (signal_4009), .Q (signal_4010) ) ;
    buf_clk cell_2602 ( .C (CLK), .D (signal_4013), .Q (signal_4014) ) ;
    buf_clk cell_2606 ( .C (CLK), .D (signal_4017), .Q (signal_4018) ) ;
    buf_clk cell_2610 ( .C (CLK), .D (signal_4021), .Q (signal_4022) ) ;
    buf_clk cell_2614 ( .C (CLK), .D (signal_4025), .Q (signal_4026) ) ;
    buf_clk cell_2618 ( .C (CLK), .D (signal_4029), .Q (signal_4030) ) ;
    buf_clk cell_2622 ( .C (CLK), .D (signal_4033), .Q (signal_4034) ) ;
    buf_clk cell_2626 ( .C (CLK), .D (signal_4037), .Q (signal_4038) ) ;
    buf_clk cell_2630 ( .C (CLK), .D (signal_4041), .Q (signal_4042) ) ;
    buf_clk cell_2634 ( .C (CLK), .D (signal_4045), .Q (signal_4046) ) ;
    buf_clk cell_2638 ( .C (CLK), .D (signal_4049), .Q (signal_4050) ) ;
    buf_clk cell_2642 ( .C (CLK), .D (signal_4053), .Q (signal_4054) ) ;
    buf_clk cell_2646 ( .C (CLK), .D (signal_4057), .Q (signal_4058) ) ;
    buf_clk cell_2650 ( .C (CLK), .D (signal_4061), .Q (signal_4062) ) ;
    buf_clk cell_2654 ( .C (CLK), .D (signal_4065), .Q (signal_4066) ) ;
    buf_clk cell_2658 ( .C (CLK), .D (signal_4069), .Q (signal_4070) ) ;
    buf_clk cell_2662 ( .C (CLK), .D (signal_4073), .Q (signal_4074) ) ;
    buf_clk cell_2666 ( .C (CLK), .D (signal_4077), .Q (signal_4078) ) ;
    buf_clk cell_2670 ( .C (CLK), .D (signal_4081), .Q (signal_4082) ) ;
    buf_clk cell_2674 ( .C (CLK), .D (signal_4085), .Q (signal_4086) ) ;
    buf_clk cell_2678 ( .C (CLK), .D (signal_4089), .Q (signal_4090) ) ;
    buf_clk cell_2682 ( .C (CLK), .D (signal_4093), .Q (signal_4094) ) ;
    buf_clk cell_2686 ( .C (CLK), .D (signal_4097), .Q (signal_4098) ) ;
    buf_clk cell_2690 ( .C (CLK), .D (signal_4101), .Q (signal_4102) ) ;
    buf_clk cell_2694 ( .C (CLK), .D (signal_4105), .Q (signal_4106) ) ;
    buf_clk cell_2698 ( .C (CLK), .D (signal_4109), .Q (signal_4110) ) ;
    buf_clk cell_2702 ( .C (CLK), .D (signal_4113), .Q (signal_4114) ) ;
    buf_clk cell_2706 ( .C (CLK), .D (signal_4117), .Q (signal_4118) ) ;
    buf_clk cell_2710 ( .C (CLK), .D (signal_4121), .Q (signal_4122) ) ;
    buf_clk cell_2714 ( .C (CLK), .D (signal_4125), .Q (signal_4126) ) ;
    buf_clk cell_2718 ( .C (CLK), .D (signal_4129), .Q (signal_4130) ) ;
    buf_clk cell_2722 ( .C (CLK), .D (signal_4133), .Q (signal_4134) ) ;
    buf_clk cell_2726 ( .C (CLK), .D (signal_4137), .Q (signal_4138) ) ;
    buf_clk cell_2730 ( .C (CLK), .D (signal_4141), .Q (signal_4142) ) ;
    buf_clk cell_2734 ( .C (CLK), .D (signal_4145), .Q (signal_4146) ) ;
    buf_clk cell_2738 ( .C (CLK), .D (signal_4149), .Q (signal_4150) ) ;
    buf_clk cell_2742 ( .C (CLK), .D (signal_4153), .Q (signal_4154) ) ;
    buf_clk cell_2746 ( .C (CLK), .D (signal_4157), .Q (signal_4158) ) ;
    buf_clk cell_2750 ( .C (CLK), .D (signal_4161), .Q (signal_4162) ) ;
    buf_clk cell_2754 ( .C (CLK), .D (signal_4165), .Q (signal_4166) ) ;
    buf_clk cell_2758 ( .C (CLK), .D (signal_4169), .Q (signal_4170) ) ;
    buf_clk cell_2762 ( .C (CLK), .D (signal_4173), .Q (signal_4174) ) ;
    buf_clk cell_2766 ( .C (CLK), .D (signal_4177), .Q (signal_4178) ) ;
    buf_clk cell_2770 ( .C (CLK), .D (signal_4181), .Q (signal_4182) ) ;
    buf_clk cell_2774 ( .C (CLK), .D (signal_4185), .Q (signal_4186) ) ;
    buf_clk cell_2778 ( .C (CLK), .D (signal_4189), .Q (signal_4190) ) ;
    buf_clk cell_2782 ( .C (CLK), .D (signal_4193), .Q (signal_4194) ) ;
    buf_clk cell_2786 ( .C (CLK), .D (signal_4197), .Q (signal_4198) ) ;
    buf_clk cell_2790 ( .C (CLK), .D (signal_4201), .Q (signal_4202) ) ;
    buf_clk cell_2794 ( .C (CLK), .D (signal_4205), .Q (signal_4206) ) ;
    buf_clk cell_2798 ( .C (CLK), .D (signal_4209), .Q (signal_4210) ) ;
    buf_clk cell_2802 ( .C (CLK), .D (signal_4213), .Q (signal_4214) ) ;
    buf_clk cell_2806 ( .C (CLK), .D (signal_4217), .Q (signal_4218) ) ;
    buf_clk cell_2810 ( .C (CLK), .D (signal_4221), .Q (signal_4222) ) ;
    buf_clk cell_2814 ( .C (CLK), .D (signal_4225), .Q (signal_4226) ) ;
    buf_clk cell_2818 ( .C (CLK), .D (signal_4229), .Q (signal_4230) ) ;
    buf_clk cell_2822 ( .C (CLK), .D (signal_4233), .Q (signal_4234) ) ;
    buf_clk cell_2826 ( .C (CLK), .D (signal_4237), .Q (signal_4238) ) ;
    buf_clk cell_2828 ( .C (CLK), .D (signal_883), .Q (signal_4240) ) ;
    buf_clk cell_2830 ( .C (CLK), .D (signal_2259), .Q (signal_4242) ) ;
    buf_clk cell_2832 ( .C (CLK), .D (signal_923), .Q (signal_4244) ) ;
    buf_clk cell_2834 ( .C (CLK), .D (signal_2271), .Q (signal_4246) ) ;
    buf_clk cell_2836 ( .C (CLK), .D (signal_903), .Q (signal_4248) ) ;
    buf_clk cell_2838 ( .C (CLK), .D (signal_2256), .Q (signal_4250) ) ;
    buf_clk cell_2840 ( .C (CLK), .D (signal_895), .Q (signal_4252) ) ;
    buf_clk cell_2842 ( .C (CLK), .D (signal_2274), .Q (signal_4254) ) ;
    buf_clk cell_2844 ( .C (CLK), .D (signal_919), .Q (signal_4256) ) ;
    buf_clk cell_2846 ( .C (CLK), .D (signal_2254), .Q (signal_4258) ) ;
    buf_clk cell_2848 ( .C (CLK), .D (signal_899), .Q (signal_4260) ) ;
    buf_clk cell_2850 ( .C (CLK), .D (signal_2257), .Q (signal_4262) ) ;
    buf_clk cell_2852 ( .C (CLK), .D (signal_891), .Q (signal_4264) ) ;
    buf_clk cell_2854 ( .C (CLK), .D (signal_2275), .Q (signal_4266) ) ;
    buf_clk cell_2856 ( .C (CLK), .D (signal_915), .Q (signal_4268) ) ;
    buf_clk cell_2858 ( .C (CLK), .D (signal_2255), .Q (signal_4270) ) ;
    buf_clk cell_2860 ( .C (CLK), .D (signal_911), .Q (signal_4272) ) ;
    buf_clk cell_2862 ( .C (CLK), .D (signal_2272), .Q (signal_4274) ) ;
    buf_clk cell_2864 ( .C (CLK), .D (signal_887), .Q (signal_4276) ) ;
    buf_clk cell_2866 ( .C (CLK), .D (signal_2258), .Q (signal_4278) ) ;
    buf_clk cell_2868 ( .C (CLK), .D (signal_927), .Q (signal_4280) ) ;
    buf_clk cell_2870 ( .C (CLK), .D (signal_2270), .Q (signal_4282) ) ;
    buf_clk cell_2872 ( .C (CLK), .D (signal_907), .Q (signal_4284) ) ;
    buf_clk cell_2874 ( .C (CLK), .D (signal_2273), .Q (signal_4286) ) ;
    buf_clk cell_3004 ( .C (CLK), .D (signal_1525), .Q (signal_4416) ) ;
    buf_clk cell_3006 ( .C (CLK), .D (signal_2293), .Q (signal_4418) ) ;
    buf_clk cell_3008 ( .C (CLK), .D (signal_1527), .Q (signal_4420) ) ;
    buf_clk cell_3010 ( .C (CLK), .D (signal_2295), .Q (signal_4422) ) ;
    buf_clk cell_3012 ( .C (CLK), .D (signal_1529), .Q (signal_4424) ) ;
    buf_clk cell_3014 ( .C (CLK), .D (signal_2277), .Q (signal_4426) ) ;
    buf_clk cell_3016 ( .C (CLK), .D (signal_1531), .Q (signal_4428) ) ;
    buf_clk cell_3018 ( .C (CLK), .D (signal_2279), .Q (signal_4430) ) ;
    buf_clk cell_3020 ( .C (CLK), .D (signal_1533), .Q (signal_4432) ) ;
    buf_clk cell_3022 ( .C (CLK), .D (signal_2297), .Q (signal_4434) ) ;
    buf_clk cell_3024 ( .C (CLK), .D (signal_1535), .Q (signal_4436) ) ;
    buf_clk cell_3026 ( .C (CLK), .D (signal_2299), .Q (signal_4438) ) ;
    buf_clk cell_3028 ( .C (CLK), .D (signal_1537), .Q (signal_4440) ) ;
    buf_clk cell_3030 ( .C (CLK), .D (signal_2281), .Q (signal_4442) ) ;
    buf_clk cell_3032 ( .C (CLK), .D (signal_1539), .Q (signal_4444) ) ;
    buf_clk cell_3034 ( .C (CLK), .D (signal_2283), .Q (signal_4446) ) ;
    buf_clk cell_3036 ( .C (CLK), .D (signal_1541), .Q (signal_4448) ) ;
    buf_clk cell_3038 ( .C (CLK), .D (signal_2301), .Q (signal_4450) ) ;
    buf_clk cell_3040 ( .C (CLK), .D (signal_1543), .Q (signal_4452) ) ;
    buf_clk cell_3042 ( .C (CLK), .D (signal_2303), .Q (signal_4454) ) ;
    buf_clk cell_3044 ( .C (CLK), .D (signal_1545), .Q (signal_4456) ) ;
    buf_clk cell_3046 ( .C (CLK), .D (signal_2285), .Q (signal_4458) ) ;
    buf_clk cell_3048 ( .C (CLK), .D (signal_1547), .Q (signal_4460) ) ;
    buf_clk cell_3050 ( .C (CLK), .D (signal_2287), .Q (signal_4462) ) ;
    buf_clk cell_3052 ( .C (CLK), .D (signal_1549), .Q (signal_4464) ) ;
    buf_clk cell_3054 ( .C (CLK), .D (signal_2305), .Q (signal_4466) ) ;
    buf_clk cell_3056 ( .C (CLK), .D (signal_1551), .Q (signal_4468) ) ;
    buf_clk cell_3058 ( .C (CLK), .D (signal_2307), .Q (signal_4470) ) ;
    buf_clk cell_3060 ( .C (CLK), .D (signal_1553), .Q (signal_4472) ) ;
    buf_clk cell_3062 ( .C (CLK), .D (signal_2289), .Q (signal_4474) ) ;
    buf_clk cell_3064 ( .C (CLK), .D (signal_1555), .Q (signal_4476) ) ;
    buf_clk cell_3066 ( .C (CLK), .D (signal_2291), .Q (signal_4478) ) ;
    buf_clk cell_3070 ( .C (CLK), .D (signal_4481), .Q (signal_4482) ) ;
    buf_clk cell_3074 ( .C (CLK), .D (signal_4485), .Q (signal_4486) ) ;
    buf_clk cell_3076 ( .C (CLK), .D (signal_3069), .Q (signal_4488) ) ;
    buf_clk cell_3078 ( .C (CLK), .D (signal_3071), .Q (signal_4490) ) ;
    buf_clk cell_3082 ( .C (CLK), .D (signal_4493), .Q (signal_4494) ) ;
    buf_clk cell_3086 ( .C (CLK), .D (signal_4497), .Q (signal_4498) ) ;
    buf_clk cell_3088 ( .C (CLK), .D (signal_3073), .Q (signal_4500) ) ;
    buf_clk cell_3090 ( .C (CLK), .D (signal_3075), .Q (signal_4502) ) ;
    buf_clk cell_3094 ( .C (CLK), .D (signal_4505), .Q (signal_4506) ) ;
    buf_clk cell_3098 ( .C (CLK), .D (signal_4509), .Q (signal_4510) ) ;
    buf_clk cell_3100 ( .C (CLK), .D (signal_3077), .Q (signal_4512) ) ;
    buf_clk cell_3102 ( .C (CLK), .D (signal_3079), .Q (signal_4514) ) ;
    buf_clk cell_3106 ( .C (CLK), .D (signal_4517), .Q (signal_4518) ) ;
    buf_clk cell_3110 ( .C (CLK), .D (signal_4521), .Q (signal_4522) ) ;
    buf_clk cell_3112 ( .C (CLK), .D (signal_3081), .Q (signal_4524) ) ;
    buf_clk cell_3114 ( .C (CLK), .D (signal_3083), .Q (signal_4526) ) ;
    buf_clk cell_3118 ( .C (CLK), .D (signal_4529), .Q (signal_4530) ) ;
    buf_clk cell_3122 ( .C (CLK), .D (signal_4533), .Q (signal_4534) ) ;
    buf_clk cell_3124 ( .C (CLK), .D (signal_3085), .Q (signal_4536) ) ;
    buf_clk cell_3126 ( .C (CLK), .D (signal_3087), .Q (signal_4538) ) ;
    buf_clk cell_3130 ( .C (CLK), .D (signal_4541), .Q (signal_4542) ) ;
    buf_clk cell_3134 ( .C (CLK), .D (signal_4545), .Q (signal_4546) ) ;
    buf_clk cell_3136 ( .C (CLK), .D (signal_3089), .Q (signal_4548) ) ;
    buf_clk cell_3138 ( .C (CLK), .D (signal_3091), .Q (signal_4550) ) ;
    buf_clk cell_3142 ( .C (CLK), .D (signal_4553), .Q (signal_4554) ) ;
    buf_clk cell_3146 ( .C (CLK), .D (signal_4557), .Q (signal_4558) ) ;
    buf_clk cell_3148 ( .C (CLK), .D (signal_3093), .Q (signal_4560) ) ;
    buf_clk cell_3150 ( .C (CLK), .D (signal_3095), .Q (signal_4562) ) ;
    buf_clk cell_3154 ( .C (CLK), .D (signal_4565), .Q (signal_4566) ) ;
    buf_clk cell_3158 ( .C (CLK), .D (signal_4569), .Q (signal_4570) ) ;
    buf_clk cell_3160 ( .C (CLK), .D (signal_3097), .Q (signal_4572) ) ;
    buf_clk cell_3162 ( .C (CLK), .D (signal_3099), .Q (signal_4574) ) ;
    buf_clk cell_3166 ( .C (CLK), .D (signal_4577), .Q (signal_4578) ) ;
    buf_clk cell_3170 ( .C (CLK), .D (signal_4581), .Q (signal_4582) ) ;
    buf_clk cell_3172 ( .C (CLK), .D (signal_3101), .Q (signal_4584) ) ;
    buf_clk cell_3174 ( .C (CLK), .D (signal_3103), .Q (signal_4586) ) ;
    buf_clk cell_3178 ( .C (CLK), .D (signal_4589), .Q (signal_4590) ) ;
    buf_clk cell_3182 ( .C (CLK), .D (signal_4593), .Q (signal_4594) ) ;
    buf_clk cell_3184 ( .C (CLK), .D (signal_3105), .Q (signal_4596) ) ;
    buf_clk cell_3186 ( .C (CLK), .D (signal_3107), .Q (signal_4598) ) ;
    buf_clk cell_3190 ( .C (CLK), .D (signal_4601), .Q (signal_4602) ) ;
    buf_clk cell_3194 ( .C (CLK), .D (signal_4605), .Q (signal_4606) ) ;
    buf_clk cell_3196 ( .C (CLK), .D (signal_3109), .Q (signal_4608) ) ;
    buf_clk cell_3198 ( .C (CLK), .D (signal_3111), .Q (signal_4610) ) ;
    buf_clk cell_3202 ( .C (CLK), .D (signal_4613), .Q (signal_4614) ) ;
    buf_clk cell_3206 ( .C (CLK), .D (signal_4617), .Q (signal_4618) ) ;
    buf_clk cell_3208 ( .C (CLK), .D (signal_3113), .Q (signal_4620) ) ;
    buf_clk cell_3210 ( .C (CLK), .D (signal_3115), .Q (signal_4622) ) ;
    buf_clk cell_3214 ( .C (CLK), .D (signal_4625), .Q (signal_4626) ) ;
    buf_clk cell_3218 ( .C (CLK), .D (signal_4629), .Q (signal_4630) ) ;
    buf_clk cell_3220 ( .C (CLK), .D (signal_3117), .Q (signal_4632) ) ;
    buf_clk cell_3222 ( .C (CLK), .D (signal_3119), .Q (signal_4634) ) ;
    buf_clk cell_3226 ( .C (CLK), .D (signal_4637), .Q (signal_4638) ) ;
    buf_clk cell_3230 ( .C (CLK), .D (signal_4641), .Q (signal_4642) ) ;
    buf_clk cell_3232 ( .C (CLK), .D (signal_3121), .Q (signal_4644) ) ;
    buf_clk cell_3234 ( .C (CLK), .D (signal_3123), .Q (signal_4646) ) ;
    buf_clk cell_3238 ( .C (CLK), .D (signal_4649), .Q (signal_4650) ) ;
    buf_clk cell_3242 ( .C (CLK), .D (signal_4653), .Q (signal_4654) ) ;
    buf_clk cell_3244 ( .C (CLK), .D (signal_3125), .Q (signal_4656) ) ;
    buf_clk cell_3246 ( .C (CLK), .D (signal_3127), .Q (signal_4658) ) ;
    buf_clk cell_3250 ( .C (CLK), .D (signal_4661), .Q (signal_4662) ) ;
    buf_clk cell_3254 ( .C (CLK), .D (signal_4665), .Q (signal_4666) ) ;
    buf_clk cell_3256 ( .C (CLK), .D (signal_3129), .Q (signal_4668) ) ;
    buf_clk cell_3258 ( .C (CLK), .D (signal_3131), .Q (signal_4670) ) ;
    buf_clk cell_3260 ( .C (CLK), .D (signal_1520), .Q (signal_4672) ) ;
    buf_clk cell_3262 ( .C (CLK), .D (signal_2268), .Q (signal_4674) ) ;
    buf_clk cell_3264 ( .C (CLK), .D (signal_1521), .Q (signal_4676) ) ;
    buf_clk cell_3266 ( .C (CLK), .D (signal_2269), .Q (signal_4678) ) ;
    buf_clk cell_3268 ( .C (CLK), .D (signal_1522), .Q (signal_4680) ) ;
    buf_clk cell_3270 ( .C (CLK), .D (signal_2252), .Q (signal_4682) ) ;
    buf_clk cell_3272 ( .C (CLK), .D (signal_1523), .Q (signal_4684) ) ;
    buf_clk cell_3274 ( .C (CLK), .D (signal_2253), .Q (signal_4686) ) ;
    buf_clk cell_3278 ( .C (CLK), .D (signal_4689), .Q (signal_4690) ) ;
    buf_clk cell_3282 ( .C (CLK), .D (signal_4693), .Q (signal_4694) ) ;
    buf_clk cell_3286 ( .C (CLK), .D (signal_4697), .Q (signal_4698) ) ;
    buf_clk cell_3290 ( .C (CLK), .D (signal_4701), .Q (signal_4702) ) ;
    buf_clk cell_3294 ( .C (CLK), .D (signal_4705), .Q (signal_4706) ) ;
    buf_clk cell_3298 ( .C (CLK), .D (signal_4709), .Q (signal_4710) ) ;
    buf_clk cell_3302 ( .C (CLK), .D (signal_4713), .Q (signal_4714) ) ;
    buf_clk cell_3306 ( .C (CLK), .D (signal_4717), .Q (signal_4718) ) ;
    buf_clk cell_3310 ( .C (CLK), .D (signal_4721), .Q (signal_4722) ) ;
    buf_clk cell_3314 ( .C (CLK), .D (signal_4725), .Q (signal_4726) ) ;
    buf_clk cell_3318 ( .C (CLK), .D (signal_4729), .Q (signal_4730) ) ;

    /* cells in depth 4 */
    mux2_masked #(.security_order(1), .pipeline(1)) cell_39 ( .s (signal_3135), .b ({signal_2503, signal_1327}), .a ({signal_3143, signal_3139}), .c ({signal_2531, signal_1263}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_40 ( .s (signal_3135), .b ({signal_2606, signal_1326}), .a ({signal_3151, signal_3147}), .c ({signal_2628, signal_1262}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_41 ( .s (signal_3155), .b ({signal_2534, signal_1325}), .a ({signal_3163, signal_3159}), .c ({signal_2551, signal_1261}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_42 ( .s (signal_3167), .b ({signal_2565, signal_1324}), .a ({signal_3175, signal_3171}), .c ({signal_2582, signal_1260}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_43 ( .s (signal_3167), .b ({signal_2538, signal_1323}), .a ({signal_3183, signal_3179}), .c ({signal_2552, signal_1259}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_44 ( .s (signal_3167), .b ({signal_2610, signal_1322}), .a ({signal_3191, signal_3187}), .c ({signal_2629, signal_1258}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_45 ( .s (signal_3167), .b ({signal_2537, signal_1321}), .a ({signal_3199, signal_3195}), .c ({signal_2553, signal_1257}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_46 ( .s (signal_3167), .b ({signal_2539, signal_1320}), .a ({signal_3207, signal_3203}), .c ({signal_2554, signal_1256}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_47 ( .s (signal_3167), .b ({signal_2543, signal_1319}), .a ({signal_3215, signal_3211}), .c ({signal_2555, signal_1255}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_48 ( .s (signal_3167), .b ({signal_2575, signal_1318}), .a ({signal_3223, signal_3219}), .c ({signal_2583, signal_1254}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_49 ( .s (signal_3167), .b ({signal_2542, signal_1317}), .a ({signal_3231, signal_3227}), .c ({signal_2556, signal_1253}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_50 ( .s (signal_3167), .b ({signal_2544, signal_1316}), .a ({signal_3239, signal_3235}), .c ({signal_2557, signal_1252}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_51 ( .s (signal_3167), .b ({signal_2549, signal_1315}), .a ({signal_3247, signal_3243}), .c ({signal_2558, signal_1251}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_52 ( .s (signal_3167), .b ({signal_2579, signal_1314}), .a ({signal_3255, signal_3251}), .c ({signal_2584, signal_1250}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_53 ( .s (signal_3167), .b ({signal_2548, signal_1313}), .a ({signal_3263, signal_3259}), .c ({signal_2559, signal_1249}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_54 ( .s (signal_3167), .b ({signal_2581, signal_1312}), .a ({signal_3271, signal_3267}), .c ({signal_2585, signal_1248}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_55 ( .s (signal_3135), .b ({signal_2648, signal_1311}), .a ({signal_3279, signal_3275}), .c ({signal_2670, signal_1247}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_56 ( .s (signal_3135), .b ({signal_2700, signal_1310}), .a ({signal_3287, signal_3283}), .c ({signal_2715, signal_1246}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_57 ( .s (signal_3135), .b ({signal_2697, signal_1309}), .a ({signal_3295, signal_3291}), .c ({signal_2716, signal_1245}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_58 ( .s (signal_3135), .b ({signal_2608, signal_1308}), .a ({signal_3303, signal_3299}), .c ({signal_2630, signal_1244}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_59 ( .s (signal_3135), .b ({signal_2612, signal_1307}), .a ({signal_3311, signal_3307}), .c ({signal_2631, signal_1243}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_60 ( .s (signal_3135), .b ({signal_2657, signal_1306}), .a ({signal_3319, signal_3315}), .c ({signal_2671, signal_1242}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_61 ( .s (signal_3135), .b ({signal_2702, signal_1305}), .a ({signal_3327, signal_3323}), .c ({signal_2717, signal_1241}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_62 ( .s (signal_3135), .b ({signal_2613, signal_1304}), .a ({signal_3335, signal_3331}), .c ({signal_2632, signal_1240}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_63 ( .s (signal_3135), .b ({signal_2618, signal_1303}), .a ({signal_3343, signal_3339}), .c ({signal_2633, signal_1239}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_64 ( .s (signal_3135), .b ({signal_2664, signal_1302}), .a ({signal_3351, signal_3347}), .c ({signal_2672, signal_1238}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_65 ( .s (signal_3135), .b ({signal_2661, signal_1301}), .a ({signal_3359, signal_3355}), .c ({signal_2673, signal_1237}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_66 ( .s (signal_3135), .b ({signal_2619, signal_1300}), .a ({signal_3367, signal_3363}), .c ({signal_2634, signal_1236}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_67 ( .s (signal_3155), .b ({signal_2668, signal_1299}), .a ({signal_3375, signal_3371}), .c ({signal_2674, signal_1235}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_68 ( .s (signal_3155), .b ({signal_2714, signal_1298}), .a ({signal_3383, signal_3379}), .c ({signal_2718, signal_1234}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_69 ( .s (signal_3155), .b ({signal_2666, signal_1297}), .a ({signal_3391, signal_3387}), .c ({signal_2675, signal_1233}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_70 ( .s (signal_3155), .b ({signal_2626, signal_1296}), .a ({signal_3399, signal_3395}), .c ({signal_2635, signal_1232}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_71 ( .s (signal_3155), .b ({signal_2696, signal_1295}), .a ({signal_3407, signal_3403}), .c ({signal_2719, signal_1231}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_72 ( .s (signal_3155), .b ({signal_2745, signal_1294}), .a ({signal_3415, signal_3411}), .c ({signal_2755, signal_1230}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_73 ( .s (signal_3155), .b ({signal_2694, signal_1293}), .a ({signal_3423, signal_3419}), .c ({signal_2720, signal_1229}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_74 ( .s (signal_3155), .b ({signal_2788, signal_1292}), .a ({signal_3431, signal_3427}), .c ({signal_2795, signal_1228}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_75 ( .s (signal_3155), .b ({signal_2701, signal_1291}), .a ({signal_3439, signal_3435}), .c ({signal_2721, signal_1227}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_76 ( .s (signal_3155), .b ({signal_2703, signal_1290}), .a ({signal_3447, signal_3443}), .c ({signal_2722, signal_1226}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_77 ( .s (signal_3155), .b ({signal_2650, signal_1289}), .a ({signal_3455, signal_3451}), .c ({signal_2676, signal_1225}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_78 ( .s (signal_3155), .b ({signal_2790, signal_1288}), .a ({signal_3463, signal_3459}), .c ({signal_2796, signal_1224}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_79 ( .s (signal_3155), .b ({signal_2705, signal_1287}), .a ({signal_3471, signal_3467}), .c ({signal_2723, signal_1223}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_80 ( .s (signal_3135), .b ({signal_2707, signal_1286}), .a ({signal_3479, signal_3475}), .c ({signal_2724, signal_1222}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_81 ( .s (signal_3167), .b ({signal_2658, signal_1285}), .a ({signal_3487, signal_3483}), .c ({signal_2677, signal_1221}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_82 ( .s (signal_3491), .b ({signal_2751, signal_1284}), .a ({signal_3499, signal_3495}), .c ({signal_2756, signal_1220}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_83 ( .s (signal_3135), .b ({signal_2710, signal_1283}), .a ({signal_3507, signal_3503}), .c ({signal_2725, signal_1219}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_84 ( .s (signal_3167), .b ({signal_2754, signal_1282}), .a ({signal_3515, signal_3511}), .c ({signal_2757, signal_1218}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_85 ( .s (signal_3155), .b ({signal_2708, signal_1281}), .a ({signal_3523, signal_3519}), .c ({signal_2726, signal_1217}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_86 ( .s (signal_3491), .b ({signal_2753, signal_1280}), .a ({signal_3531, signal_3527}), .c ({signal_2758, signal_1216}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_87 ( .s (signal_3491), .b ({signal_2847, signal_1279}), .a ({signal_3539, signal_3535}), .c ({signal_2852, signal_1215}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_88 ( .s (signal_3491), .b ({signal_2860, signal_1278}), .a ({signal_3547, signal_3543}), .c ({signal_2862, signal_1214}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_89 ( .s (signal_3491), .b ({signal_2787, signal_1277}), .a ({signal_3555, signal_3551}), .c ({signal_2797, signal_1213}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_90 ( .s (signal_3491), .b ({signal_2786, signal_1276}), .a ({signal_3563, signal_3559}), .c ({signal_2798, signal_1212}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_91 ( .s (signal_3491), .b ({signal_2849, signal_1275}), .a ({signal_3571, signal_3567}), .c ({signal_2853, signal_1211}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_92 ( .s (signal_3491), .b ({signal_2861, signal_1274}), .a ({signal_3579, signal_3575}), .c ({signal_2863, signal_1210}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_93 ( .s (signal_3155), .b ({signal_2747, signal_1273}), .a ({signal_3587, signal_3583}), .c ({signal_2759, signal_1209}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_94 ( .s (signal_3135), .b ({signal_2789, signal_1272}), .a ({signal_3595, signal_3591}), .c ({signal_2799, signal_1208}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_95 ( .s (signal_3167), .b ({signal_2841, signal_1271}), .a ({signal_3603, signal_3599}), .c ({signal_2844, signal_1207}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_96 ( .s (signal_3155), .b ({signal_2850, signal_1270}), .a ({signal_3611, signal_3607}), .c ({signal_2854, signal_1206}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_97 ( .s (signal_3135), .b ({signal_2750, signal_1269}), .a ({signal_3619, signal_3615}), .c ({signal_2760, signal_1205}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_98 ( .s (signal_3167), .b ({signal_2749, signal_1268}), .a ({signal_3627, signal_3623}), .c ({signal_2761, signal_1204}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_99 ( .s (signal_3135), .b ({signal_2843, signal_1267}), .a ({signal_3635, signal_3631}), .c ({signal_2845, signal_1203}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_100 ( .s (signal_3167), .b ({signal_2851, signal_1266}), .a ({signal_3643, signal_3639}), .c ({signal_2855, signal_1202}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_101 ( .s (signal_3155), .b ({signal_2793, signal_1265}), .a ({signal_3651, signal_3647}), .c ({signal_2800, signal_1201}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_102 ( .s (signal_3155), .b ({signal_2792, signal_1264}), .a ({signal_3659, signal_3655}), .c ({signal_2801, signal_1200}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_103 ( .s (signal_3663), .b ({signal_2531, signal_1263}), .a ({signal_3671, signal_3667}), .c ({signal_2561, signal_1199}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_104 ( .s (signal_3663), .b ({signal_2628, signal_1262}), .a ({signal_3679, signal_3675}), .c ({signal_2679, signal_1198}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_105 ( .s (signal_3663), .b ({signal_2551, signal_1261}), .a ({signal_3687, signal_3683}), .c ({signal_2587, signal_1197}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_106 ( .s (signal_3663), .b ({signal_2582, signal_1260}), .a ({signal_3695, signal_3691}), .c ({signal_2637, signal_1196}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_107 ( .s (signal_3663), .b ({signal_2552, signal_1259}), .a ({signal_3703, signal_3699}), .c ({signal_2589, signal_1195}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_108 ( .s (signal_3663), .b ({signal_2629, signal_1258}), .a ({signal_3711, signal_3707}), .c ({signal_2681, signal_1194}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_109 ( .s (signal_3663), .b ({signal_2553, signal_1257}), .a ({signal_3719, signal_3715}), .c ({signal_2591, signal_1193}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_110 ( .s (signal_3663), .b ({signal_2554, signal_1256}), .a ({signal_3727, signal_3723}), .c ({signal_2593, signal_1192}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_111 ( .s (signal_3663), .b ({signal_2555, signal_1255}), .a ({signal_3735, signal_3731}), .c ({signal_2595, signal_1191}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_112 ( .s (signal_3663), .b ({signal_2583, signal_1254}), .a ({signal_3743, signal_3739}), .c ({signal_2639, signal_1190}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_113 ( .s (signal_3663), .b ({signal_2556, signal_1253}), .a ({signal_3751, signal_3747}), .c ({signal_2597, signal_1189}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_114 ( .s (signal_3663), .b ({signal_2557, signal_1252}), .a ({signal_3759, signal_3755}), .c ({signal_2599, signal_1188}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_115 ( .s (signal_3663), .b ({signal_2558, signal_1251}), .a ({signal_3767, signal_3763}), .c ({signal_2601, signal_1187}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_116 ( .s (signal_3663), .b ({signal_2584, signal_1250}), .a ({signal_3775, signal_3771}), .c ({signal_2641, signal_1186}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_117 ( .s (signal_3663), .b ({signal_2559, signal_1249}), .a ({signal_3783, signal_3779}), .c ({signal_2603, signal_1185}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_118 ( .s (signal_3663), .b ({signal_2585, signal_1248}), .a ({signal_3791, signal_3787}), .c ({signal_2643, signal_1184}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_119 ( .s (signal_3663), .b ({signal_2670, signal_1247}), .a ({signal_3799, signal_3795}), .c ({signal_2728, signal_1183}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_120 ( .s (signal_3663), .b ({signal_2715, signal_1246}), .a ({signal_3807, signal_3803}), .c ({signal_2763, signal_1182}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_121 ( .s (signal_3663), .b ({signal_2716, signal_1245}), .a ({signal_3815, signal_3811}), .c ({signal_2765, signal_1181}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_122 ( .s (signal_3663), .b ({signal_2630, signal_1244}), .a ({signal_3823, signal_3819}), .c ({signal_2683, signal_1180}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_123 ( .s (signal_3663), .b ({signal_2631, signal_1243}), .a ({signal_3831, signal_3827}), .c ({signal_2685, signal_1179}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_124 ( .s (signal_3663), .b ({signal_2671, signal_1242}), .a ({signal_3839, signal_3835}), .c ({signal_2730, signal_1178}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_125 ( .s (signal_3663), .b ({signal_2717, signal_1241}), .a ({signal_3847, signal_3843}), .c ({signal_2767, signal_1177}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_126 ( .s (signal_3663), .b ({signal_2632, signal_1240}), .a ({signal_3855, signal_3851}), .c ({signal_2687, signal_1176}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_127 ( .s (signal_3663), .b ({signal_2633, signal_1239}), .a ({signal_3863, signal_3859}), .c ({signal_2689, signal_1175}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_128 ( .s (signal_3663), .b ({signal_2672, signal_1238}), .a ({signal_3871, signal_3867}), .c ({signal_2732, signal_1174}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_129 ( .s (signal_3663), .b ({signal_2673, signal_1237}), .a ({signal_3879, signal_3875}), .c ({signal_2734, signal_1173}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_130 ( .s (signal_3663), .b ({signal_2634, signal_1236}), .a ({signal_3887, signal_3883}), .c ({signal_2691, signal_1172}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_131 ( .s (signal_3663), .b ({signal_2674, signal_1235}), .a ({signal_3895, signal_3891}), .c ({signal_2736, signal_1171}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_132 ( .s (signal_3663), .b ({signal_2718, signal_1234}), .a ({signal_3903, signal_3899}), .c ({signal_2769, signal_1170}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_133 ( .s (signal_3663), .b ({signal_2675, signal_1233}), .a ({signal_3911, signal_3907}), .c ({signal_2738, signal_1169}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_134 ( .s (signal_3663), .b ({signal_2635, signal_1232}), .a ({signal_3919, signal_3915}), .c ({signal_2693, signal_1168}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_135 ( .s (signal_3663), .b ({signal_2719, signal_1231}), .a ({signal_3927, signal_3923}), .c ({signal_2771, signal_1167}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_136 ( .s (signal_3663), .b ({signal_2755, signal_1230}), .a ({signal_3935, signal_3931}), .c ({signal_2803, signal_1166}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_137 ( .s (signal_3663), .b ({signal_2720, signal_1229}), .a ({signal_3943, signal_3939}), .c ({signal_2773, signal_1165}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_138 ( .s (signal_3663), .b ({signal_2795, signal_1228}), .a ({signal_3951, signal_3947}), .c ({signal_2823, signal_1164}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_139 ( .s (signal_3663), .b ({signal_2721, signal_1227}), .a ({signal_3959, signal_3955}), .c ({signal_2775, signal_1163}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_140 ( .s (signal_3663), .b ({signal_2722, signal_1226}), .a ({signal_3967, signal_3963}), .c ({signal_2777, signal_1162}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_141 ( .s (signal_3663), .b ({signal_2676, signal_1225}), .a ({signal_3975, signal_3971}), .c ({signal_2740, signal_1161}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_142 ( .s (signal_3663), .b ({signal_2796, signal_1224}), .a ({signal_3983, signal_3979}), .c ({signal_2825, signal_1160}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_143 ( .s (signal_3663), .b ({signal_2723, signal_1223}), .a ({signal_3991, signal_3987}), .c ({signal_2779, signal_1159}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_144 ( .s (signal_3663), .b ({signal_2724, signal_1222}), .a ({signal_3999, signal_3995}), .c ({signal_2781, signal_1158}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_145 ( .s (signal_3663), .b ({signal_2677, signal_1221}), .a ({signal_4007, signal_4003}), .c ({signal_2742, signal_1157}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_146 ( .s (signal_3663), .b ({signal_2756, signal_1220}), .a ({signal_4015, signal_4011}), .c ({signal_2805, signal_1156}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_147 ( .s (signal_3663), .b ({signal_2725, signal_1219}), .a ({signal_4023, signal_4019}), .c ({signal_2783, signal_1155}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_148 ( .s (signal_3663), .b ({signal_2757, signal_1218}), .a ({signal_4031, signal_4027}), .c ({signal_2807, signal_1154}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_149 ( .s (signal_3663), .b ({signal_2726, signal_1217}), .a ({signal_4039, signal_4035}), .c ({signal_2785, signal_1153}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_150 ( .s (signal_3663), .b ({signal_2758, signal_1216}), .a ({signal_4047, signal_4043}), .c ({signal_2809, signal_1152}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_151 ( .s (signal_3663), .b ({signal_2852, signal_1215}), .a ({signal_4055, signal_4051}), .c ({signal_2865, signal_1151}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_152 ( .s (signal_3663), .b ({signal_2862, signal_1214}), .a ({signal_4063, signal_4059}), .c ({signal_2873, signal_1150}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_153 ( .s (signal_3663), .b ({signal_2797, signal_1213}), .a ({signal_4071, signal_4067}), .c ({signal_2827, signal_1149}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_154 ( .s (signal_3663), .b ({signal_2798, signal_1212}), .a ({signal_4079, signal_4075}), .c ({signal_2829, signal_1148}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_155 ( .s (signal_3663), .b ({signal_2853, signal_1211}), .a ({signal_4087, signal_4083}), .c ({signal_2867, signal_1147}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_156 ( .s (signal_3663), .b ({signal_2863, signal_1210}), .a ({signal_4095, signal_4091}), .c ({signal_2875, signal_1146}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_157 ( .s (signal_3663), .b ({signal_2759, signal_1209}), .a ({signal_4103, signal_4099}), .c ({signal_2811, signal_1145}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_158 ( .s (signal_3663), .b ({signal_2799, signal_1208}), .a ({signal_4111, signal_4107}), .c ({signal_2831, signal_1144}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_159 ( .s (signal_3663), .b ({signal_2844, signal_1207}), .a ({signal_4119, signal_4115}), .c ({signal_2857, signal_1143}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_160 ( .s (signal_3663), .b ({signal_2854, signal_1206}), .a ({signal_4127, signal_4123}), .c ({signal_2869, signal_1142}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_161 ( .s (signal_3663), .b ({signal_2760, signal_1205}), .a ({signal_4135, signal_4131}), .c ({signal_2813, signal_1141}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_162 ( .s (signal_3663), .b ({signal_2761, signal_1204}), .a ({signal_4143, signal_4139}), .c ({signal_2815, signal_1140}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_163 ( .s (signal_3663), .b ({signal_2845, signal_1203}), .a ({signal_4151, signal_4147}), .c ({signal_2859, signal_1139}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_164 ( .s (signal_3663), .b ({signal_2855, signal_1202}), .a ({signal_4159, signal_4155}), .c ({signal_2871, signal_1138}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_165 ( .s (signal_3663), .b ({signal_2800, signal_1201}), .a ({signal_4167, signal_4163}), .c ({signal_2833, signal_1137}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_166 ( .s (signal_3663), .b ({signal_2801, signal_1200}), .a ({signal_4175, signal_4171}), .c ({signal_2835, signal_1136}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_412 ( .a ({signal_4183, signal_4179}), .b ({signal_2436, signal_356}), .c ({signal_2467, signal_940}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_435 ( .a ({signal_4191, signal_4187}), .b ({signal_2439, signal_375}), .c ({signal_2468, signal_936}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_458 ( .a ({signal_3215, signal_3211}), .b ({signal_2404, signal_394}), .c ({signal_2428, signal_932}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_481 ( .a ({signal_3247, signal_3243}), .b ({signal_2407, signal_413}), .c ({signal_2429, signal_928}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_504 ( .a ({signal_4199, signal_4195}), .b ({signal_2442, signal_432}), .c ({signal_2469, signal_924}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_527 ( .a ({signal_4207, signal_4203}), .b ({signal_2445, signal_451}), .c ({signal_2470, signal_920}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_550 ( .a ({signal_3343, signal_3339}), .b ({signal_2410, signal_470}), .c ({signal_2430, signal_916}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_573 ( .a ({signal_3375, signal_3371}), .b ({signal_2413, signal_489}), .c ({signal_2431, signal_912}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_596 ( .a ({signal_4215, signal_4211}), .b ({signal_2448, signal_508}), .c ({signal_2471, signal_908}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_619 ( .a ({signal_4223, signal_4219}), .b ({signal_2451, signal_527}), .c ({signal_2472, signal_904}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_642 ( .a ({signal_3471, signal_3467}), .b ({signal_2416, signal_546}), .c ({signal_2432, signal_900}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_665 ( .a ({signal_3507, signal_3503}), .b ({signal_2419, signal_565}), .c ({signal_2433, signal_896}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_688 ( .a ({signal_4231, signal_4227}), .b ({signal_2454, signal_584}), .c ({signal_2473, signal_892}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_711 ( .a ({signal_4239, signal_4235}), .b ({signal_2457, signal_603}), .c ({signal_2474, signal_888}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_734 ( .a ({signal_3603, signal_3599}), .b ({signal_2422, signal_622}), .c ({signal_2434, signal_884}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_757 ( .a ({signal_3635, signal_3631}), .b ({signal_2425, signal_641}), .c ({signal_2435, signal_880}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_762 ( .a ({signal_2743, signal_656}), .b ({signal_2604, signal_657}), .c ({signal_2786, signal_1276}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_763 ( .a ({signal_2565, signal_1324}), .b ({signal_2427, signal_882}), .c ({signal_2604, signal_657}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_764 ( .a ({signal_2694, signal_1293}), .b ({signal_2697, signal_1309}), .c ({signal_2743, signal_656}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_765 ( .a ({signal_2562, signal_658}), .b ({signal_2649, signal_659}), .c ({signal_2694, signal_1293}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_766 ( .a ({signal_2426, signal_881}), .b ({signal_2533, signal_660}), .c ({signal_2562, signal_658}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_767 ( .a ({signal_2695, signal_661}), .b ({signal_2745, signal_1294}), .c ({signal_2787, signal_1277}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_768 ( .a ({signal_2534, signal_1325}), .b ({signal_2649, signal_659}), .c ({signal_2695, signal_661}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_769 ( .a ({signal_2846, signal_662}), .b ({signal_2698, signal_663}), .c ({signal_2860, signal_1278}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_770 ( .a ({signal_2836, signal_664}), .b ({signal_2644, signal_665}), .c ({signal_2846, signal_662}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_771 ( .a ({signal_2435, signal_880}), .b ({signal_2606, signal_1326}), .c ({signal_2644, signal_665}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_772 ( .a ({signal_2696, signal_1295}), .b ({signal_2816, signal_666}), .c ({signal_2836, signal_664}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_773 ( .a ({signal_2645, signal_667}), .b ({signal_2605, signal_668}), .c ({signal_2696, signal_1295}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_774 ( .a ({signal_2417, signal_901}), .b ({signal_2565, signal_1324}), .c ({signal_2605, signal_668}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_775 ( .a ({signal_4243, signal_4241}), .b ({signal_2608, signal_1308}), .c ({signal_2645, signal_667}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_776 ( .a ({signal_2837, signal_669}), .b ({signal_2503, signal_1327}), .c ({signal_2847, signal_1279}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_777 ( .a ({signal_2608, signal_1308}), .b ({signal_2816, signal_666}), .c ({signal_2837, signal_669}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_778 ( .a ({signal_2426, signal_881}), .b ({signal_2788, signal_1292}), .c ({signal_2816, signal_666}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_779 ( .a ({signal_2744, signal_670}), .b ({signal_2475, signal_671}), .c ({signal_2788, signal_1292}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_780 ( .a ({signal_2435, signal_880}), .b ({signal_2418, signal_902}), .c ({signal_2475, signal_671}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_781 ( .a ({signal_2697, signal_1309}), .b ({signal_2534, signal_1325}), .c ({signal_2744, signal_670}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_782 ( .a ({signal_2646, signal_672}), .b ({signal_2532, signal_673}), .c ({signal_2697, signal_1309}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_783 ( .a ({signal_2504, signal_674}), .b ({signal_2427, signal_882}), .c ({signal_2532, signal_673}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_784 ( .a ({signal_2606, signal_1326}), .b ({signal_4247, signal_4245}), .c ({signal_2646, signal_672}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_785 ( .a ({signal_2563, signal_675}), .b ({signal_2476, signal_676}), .c ({signal_2606, signal_1326}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_786 ( .a ({signal_4251, signal_4249}), .b ({signal_2432, signal_900}), .c ({signal_2476, signal_676}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_787 ( .a ({signal_2479, signal_677}), .b ({signal_2533, signal_660}), .c ({signal_2563, signal_675}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_788 ( .a ({signal_2500, signal_678}), .b ({signal_2437, signal_941}), .c ({signal_2533, signal_660}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_789 ( .a ({signal_2447, signal_922}), .b ({signal_2467, signal_940}), .c ({signal_2500, signal_678}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_790 ( .a ({signal_2699, signal_679}), .b ({signal_2698, signal_663}), .c ({signal_2745, signal_1294}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_791 ( .a ({signal_2648, signal_1311}), .b ({signal_2608, signal_1308}), .c ({signal_2698, signal_663}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_792 ( .a ({signal_2647, signal_680}), .b ({signal_2477, signal_681}), .c ({signal_2699, signal_679}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_793 ( .a ({signal_2417, signal_901}), .b ({signal_2432, signal_900}), .c ({signal_2477, signal_681}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_794 ( .a ({signal_2609, signal_682}), .b ({signal_2427, signal_882}), .c ({signal_2647, signal_680}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_795 ( .a ({signal_2491, signal_683}), .b ({signal_2607, signal_684}), .c ({signal_2648, signal_1311}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_796 ( .a ({signal_2565, signal_1324}), .b ({signal_2435, signal_880}), .c ({signal_2607, signal_684}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_798 ( .a ({signal_2564, signal_685}), .b ({signal_2478, signal_686}), .c ({signal_2608, signal_1308}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_799 ( .a ({signal_2426, signal_881}), .b ({signal_2432, signal_900}), .c ({signal_2478, signal_686}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_800 ( .a ({signal_2534, signal_1325}), .b ({signal_2447, signal_922}), .c ({signal_2564, signal_685}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_801 ( .a ({signal_2460, signal_687}), .b ({signal_2501, signal_688}), .c ({signal_2534, signal_1325}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_802 ( .a ({signal_2492, signal_689}), .b ({signal_2467, signal_940}), .c ({signal_2501, signal_688}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_804 ( .a ({signal_2479, signal_677}), .b ({signal_2649, signal_659}), .c ({signal_2700, signal_1310}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_805 ( .a ({signal_2502, signal_690}), .b ({signal_2609, signal_682}), .c ({signal_2649, signal_659}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_806 ( .a ({signal_2565, signal_1324}), .b ({signal_2503, signal_1327}), .c ({signal_2609, signal_682}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_807 ( .a ({signal_2470, signal_920}), .b ({signal_2492, signal_689}), .c ({signal_2502, signal_690}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_809 ( .a ({signal_2435, signal_880}), .b ({signal_4243, signal_4241}), .c ({signal_2479, signal_677}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_810 ( .a ({signal_2493, signal_691}), .b ({signal_2480, signal_692}), .c ({signal_2503, signal_1327}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_811 ( .a ({signal_2435, signal_880}), .b ({signal_2432, signal_900}), .c ({signal_2480, signal_692}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_813 ( .a ({signal_2535, signal_693}), .b ({signal_2426, signal_881}), .c ({signal_2565, signal_1324}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_814 ( .a ({signal_2504, signal_674}), .b ({signal_2438, signal_942}), .c ({signal_2535, signal_693}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_815 ( .a ({signal_2417, signal_901}), .b ({signal_2470, signal_920}), .c ({signal_2504, signal_674}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_816 ( .a ({signal_2746, signal_694}), .b ({signal_2566, signal_695}), .c ({signal_2789, signal_1272}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_817 ( .a ({signal_2539, signal_1320}), .b ({signal_2456, signal_894}), .c ({signal_2566, signal_695}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_818 ( .a ({signal_2650, signal_1289}), .b ({signal_2702, signal_1305}), .c ({signal_2746, signal_694}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_819 ( .a ({signal_2567, signal_696}), .b ({signal_2614, signal_697}), .c ({signal_2650, signal_1289}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_820 ( .a ({signal_2455, signal_893}), .b ({signal_2536, signal_698}), .c ({signal_2567, signal_696}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_821 ( .a ({signal_2651, signal_699}), .b ({signal_2703, signal_1290}), .c ({signal_2747, signal_1273}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_822 ( .a ({signal_2537, signal_1321}), .b ({signal_2614, signal_697}), .c ({signal_2651, signal_699}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_823 ( .a ({signal_2848, signal_700}), .b ({signal_2655, signal_701}), .c ({signal_2861, signal_1274}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_824 ( .a ({signal_2838, signal_702}), .b ({signal_2652, signal_703}), .c ({signal_2848, signal_700}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_825 ( .a ({signal_2473, signal_892}), .b ({signal_2610, signal_1322}), .c ({signal_2652, signal_703}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_826 ( .a ({signal_2701, signal_1291}), .b ({signal_2817, signal_704}), .c ({signal_2838, signal_702}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_827 ( .a ({signal_2653, signal_705}), .b ({signal_2568, signal_706}), .c ({signal_2701, signal_1291}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_828 ( .a ({signal_2420, signal_897}), .b ({signal_2539, signal_1320}), .c ({signal_2568, signal_706}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_829 ( .a ({signal_4255, signal_4253}), .b ({signal_2613, signal_1304}), .c ({signal_2653, signal_705}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_830 ( .a ({signal_2839, signal_707}), .b ({signal_2538, signal_1323}), .c ({signal_2849, signal_1275}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_831 ( .a ({signal_2613, signal_1304}), .b ({signal_2817, signal_704}), .c ({signal_2839, signal_707}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_832 ( .a ({signal_2455, signal_893}), .b ({signal_2790, signal_1288}), .c ({signal_2817, signal_704}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_833 ( .a ({signal_2748, signal_708}), .b ({signal_2505, signal_709}), .c ({signal_2790, signal_1288}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_834 ( .a ({signal_2473, signal_892}), .b ({signal_2421, signal_898}), .c ({signal_2505, signal_709}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_835 ( .a ({signal_2702, signal_1305}), .b ({signal_2537, signal_1321}), .c ({signal_2748, signal_708}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_836 ( .a ({signal_2654, signal_710}), .b ({signal_2506, signal_711}), .c ({signal_2702, signal_1305}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_837 ( .a ({signal_2485, signal_712}), .b ({signal_2456, signal_894}), .c ({signal_2506, signal_711}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_838 ( .a ({signal_2610, signal_1322}), .b ({signal_4259, signal_4257}), .c ({signal_2654, signal_710}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_839 ( .a ({signal_2569, signal_713}), .b ({signal_2481, signal_714}), .c ({signal_2610, signal_1322}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_840 ( .a ({signal_4263, signal_4261}), .b ({signal_2433, signal_896}), .c ({signal_2481, signal_714}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_841 ( .a ({signal_2509, signal_715}), .b ({signal_2536, signal_698}), .c ({signal_2569, signal_713}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_842 ( .a ({signal_2507, signal_716}), .b ({signal_2440, signal_937}), .c ({signal_2536, signal_698}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_843 ( .a ({signal_2412, signal_918}), .b ({signal_2468, signal_936}), .c ({signal_2507, signal_716}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_844 ( .a ({signal_2656, signal_717}), .b ({signal_2655, signal_701}), .c ({signal_2703, signal_1290}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_845 ( .a ({signal_2612, signal_1307}), .b ({signal_2613, signal_1304}), .c ({signal_2655, signal_701}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_846 ( .a ({signal_2611, signal_718}), .b ({signal_2482, signal_719}), .c ({signal_2656, signal_717}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_847 ( .a ({signal_2420, signal_897}), .b ({signal_2433, signal_896}), .c ({signal_2482, signal_719}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_848 ( .a ({signal_2572, signal_720}), .b ({signal_2456, signal_894}), .c ({signal_2611, signal_718}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_849 ( .a ({signal_2461, signal_721}), .b ({signal_2570, signal_722}), .c ({signal_2612, signal_1307}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_850 ( .a ({signal_2539, signal_1320}), .b ({signal_2473, signal_892}), .c ({signal_2570, signal_722}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_852 ( .a ({signal_2571, signal_723}), .b ({signal_2483, signal_724}), .c ({signal_2613, signal_1304}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_853 ( .a ({signal_2455, signal_893}), .b ({signal_2433, signal_896}), .c ({signal_2483, signal_724}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_854 ( .a ({signal_2537, signal_1321}), .b ({signal_2412, signal_918}), .c ({signal_2571, signal_723}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_855 ( .a ({signal_2494, signal_725}), .b ({signal_2508, signal_726}), .c ({signal_2537, signal_1321}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_856 ( .a ({signal_2462, signal_727}), .b ({signal_2468, signal_936}), .c ({signal_2508, signal_726}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_858 ( .a ({signal_2509, signal_715}), .b ({signal_2614, signal_697}), .c ({signal_2657, signal_1306}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_859 ( .a ({signal_2484, signal_728}), .b ({signal_2572, signal_720}), .c ({signal_2614, signal_697}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_860 ( .a ({signal_2539, signal_1320}), .b ({signal_2538, signal_1323}), .c ({signal_2572, signal_720}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_861 ( .a ({signal_2430, signal_916}), .b ({signal_2462, signal_727}), .c ({signal_2484, signal_728}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_863 ( .a ({signal_2473, signal_892}), .b ({signal_4255, signal_4253}), .c ({signal_2509, signal_715}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_864 ( .a ({signal_2495, signal_729}), .b ({signal_2510, signal_730}), .c ({signal_2538, signal_1323}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_865 ( .a ({signal_2473, signal_892}), .b ({signal_2433, signal_896}), .c ({signal_2510, signal_730}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_867 ( .a ({signal_2511, signal_731}), .b ({signal_2455, signal_893}), .c ({signal_2539, signal_1320}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_868 ( .a ({signal_2485, signal_712}), .b ({signal_2441, signal_938}), .c ({signal_2511, signal_731}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_869 ( .a ({signal_2420, signal_897}), .b ({signal_2430, signal_916}), .c ({signal_2485, signal_712}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_870 ( .a ({signal_2704, signal_732}), .b ({signal_2573, signal_733}), .c ({signal_2749, signal_1268}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_871 ( .a ({signal_2544, signal_1316}), .b ({signal_2459, signal_890}), .c ({signal_2573, signal_733}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_872 ( .a ({signal_2658, signal_1285}), .b ({signal_2661, signal_1301}), .c ({signal_2704, signal_732}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_873 ( .a ({signal_2540, signal_734}), .b ({signal_2620, signal_735}), .c ({signal_2658, signal_1285}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_874 ( .a ({signal_2458, signal_889}), .b ({signal_2515, signal_736}), .c ({signal_2540, signal_734}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_875 ( .a ({signal_2659, signal_737}), .b ({signal_2707, signal_1286}), .c ({signal_2750, signal_1269}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_876 ( .a ({signal_2542, signal_1317}), .b ({signal_2620, signal_735}), .c ({signal_2659, signal_737}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_877 ( .a ({signal_2840, signal_738}), .b ({signal_2662, signal_739}), .c ({signal_2850, signal_1270}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_878 ( .a ({signal_2818, signal_740}), .b ({signal_2615, signal_741}), .c ({signal_2840, signal_738}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_879 ( .a ({signal_2474, signal_888}), .b ({signal_2575, signal_1318}), .c ({signal_2615, signal_741}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_880 ( .a ({signal_2705, signal_1287}), .b ({signal_2791, signal_742}), .c ({signal_2818, signal_740}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_881 ( .a ({signal_2660, signal_743}), .b ({signal_2574, signal_744}), .c ({signal_2705, signal_1287}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_882 ( .a ({signal_2449, signal_909}), .b ({signal_2544, signal_1316}), .c ({signal_2574, signal_744}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_883 ( .a ({signal_4267, signal_4265}), .b ({signal_2619, signal_1300}), .c ({signal_2660, signal_743}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_884 ( .a ({signal_2819, signal_745}), .b ({signal_2543, signal_1319}), .c ({signal_2841, signal_1271}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_885 ( .a ({signal_2619, signal_1300}), .b ({signal_2791, signal_742}), .c ({signal_2819, signal_745}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_886 ( .a ({signal_2458, signal_889}), .b ({signal_2751, signal_1284}), .c ({signal_2791, signal_742}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_887 ( .a ({signal_2706, signal_746}), .b ({signal_2512, signal_747}), .c ({signal_2751, signal_1284}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_888 ( .a ({signal_2474, signal_888}), .b ({signal_2450, signal_910}), .c ({signal_2512, signal_747}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_889 ( .a ({signal_2661, signal_1301}), .b ({signal_2542, signal_1317}), .c ({signal_2706, signal_746}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_890 ( .a ({signal_2616, signal_748}), .b ({signal_2513, signal_749}), .c ({signal_2661, signal_1301}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_891 ( .a ({signal_2487, signal_750}), .b ({signal_2459, signal_890}), .c ({signal_2513, signal_749}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_892 ( .a ({signal_2575, signal_1318}), .b ({signal_4271, signal_4269}), .c ({signal_2616, signal_748}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_893 ( .a ({signal_2541, signal_751}), .b ({signal_2514, signal_752}), .c ({signal_2575, signal_1318}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_894 ( .a ({signal_4275, signal_4273}), .b ({signal_2471, signal_908}), .c ({signal_2514, signal_752}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_895 ( .a ({signal_2520, signal_753}), .b ({signal_2515, signal_736}), .c ({signal_2541, signal_751}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_896 ( .a ({signal_2486, signal_754}), .b ({signal_2405, signal_933}), .c ({signal_2515, signal_736}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_897 ( .a ({signal_2415, signal_914}), .b ({signal_2428, signal_932}), .c ({signal_2486, signal_754}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_898 ( .a ({signal_2663, signal_755}), .b ({signal_2662, signal_739}), .c ({signal_2707, signal_1286}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_899 ( .a ({signal_2618, signal_1303}), .b ({signal_2619, signal_1300}), .c ({signal_2662, signal_739}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_900 ( .a ({signal_2617, signal_756}), .b ({signal_2516, signal_757}), .c ({signal_2663, signal_755}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_901 ( .a ({signal_2449, signal_909}), .b ({signal_2471, signal_908}), .c ({signal_2516, signal_757}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_902 ( .a ({signal_2578, signal_758}), .b ({signal_2459, signal_890}), .c ({signal_2617, signal_756}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_903 ( .a ({signal_2463, signal_759}), .b ({signal_2576, signal_760}), .c ({signal_2618, signal_1303}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_904 ( .a ({signal_2544, signal_1316}), .b ({signal_2474, signal_888}), .c ({signal_2576, signal_760}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_906 ( .a ({signal_2577, signal_761}), .b ({signal_2517, signal_762}), .c ({signal_2619, signal_1300}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_907 ( .a ({signal_2458, signal_889}), .b ({signal_2471, signal_908}), .c ({signal_2517, signal_762}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_908 ( .a ({signal_2542, signal_1317}), .b ({signal_2415, signal_914}), .c ({signal_2577, signal_761}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_909 ( .a ({signal_2496, signal_763}), .b ({signal_2518, signal_764}), .c ({signal_2542, signal_1317}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_910 ( .a ({signal_2497, signal_765}), .b ({signal_2428, signal_932}), .c ({signal_2518, signal_764}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_912 ( .a ({signal_2520, signal_753}), .b ({signal_2620, signal_735}), .c ({signal_2664, signal_1302}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_913 ( .a ({signal_2519, signal_766}), .b ({signal_2578, signal_758}), .c ({signal_2620, signal_735}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_914 ( .a ({signal_2544, signal_1316}), .b ({signal_2543, signal_1319}), .c ({signal_2578, signal_758}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_915 ( .a ({signal_2431, signal_912}), .b ({signal_2497, signal_765}), .c ({signal_2519, signal_766}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_917 ( .a ({signal_2474, signal_888}), .b ({signal_4267, signal_4265}), .c ({signal_2520, signal_753}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_918 ( .a ({signal_2464, signal_767}), .b ({signal_2521, signal_768}), .c ({signal_2543, signal_1319}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_919 ( .a ({signal_2474, signal_888}), .b ({signal_2471, signal_908}), .c ({signal_2521, signal_768}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_921 ( .a ({signal_2522, signal_769}), .b ({signal_2458, signal_889}), .c ({signal_2544, signal_1316}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_922 ( .a ({signal_2487, signal_750}), .b ({signal_2406, signal_934}), .c ({signal_2522, signal_769}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_923 ( .a ({signal_2449, signal_909}), .b ({signal_2431, signal_912}), .c ({signal_2487, signal_750}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_924 ( .a ({signal_2752, signal_770}), .b ({signal_2621, signal_771}), .c ({signal_2792, signal_1264}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_925 ( .a ({signal_2581, signal_1312}), .b ({signal_2424, signal_886}), .c ({signal_2621, signal_771}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_926 ( .a ({signal_2708, signal_1281}), .b ({signal_2666, signal_1297}), .c ({signal_2752, signal_770}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_927 ( .a ({signal_2545, signal_772}), .b ({signal_2669, signal_773}), .c ({signal_2708, signal_1281}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_928 ( .a ({signal_2423, signal_885}), .b ({signal_2524, signal_774}), .c ({signal_2545, signal_772}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_929 ( .a ({signal_2709, signal_775}), .b ({signal_2754, signal_1282}), .c ({signal_2793, signal_1265}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_930 ( .a ({signal_2548, signal_1313}), .b ({signal_2669, signal_773}), .c ({signal_2709, signal_775}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_931 ( .a ({signal_2842, signal_776}), .b ({signal_2712, signal_777}), .c ({signal_2851, signal_1266}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_932 ( .a ({signal_2820, signal_778}), .b ({signal_2622, signal_779}), .c ({signal_2842, signal_776}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_933 ( .a ({signal_2434, signal_884}), .b ({signal_2579, signal_1314}), .c ({signal_2622, signal_779}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_934 ( .a ({signal_2710, signal_1283}), .b ({signal_2794, signal_780}), .c ({signal_2820, signal_778}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_935 ( .a ({signal_2665, signal_781}), .b ({signal_2623, signal_782}), .c ({signal_2710, signal_1283}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_936 ( .a ({signal_2452, signal_905}), .b ({signal_2581, signal_1312}), .c ({signal_2623, signal_782}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_937 ( .a ({signal_4279, signal_4277}), .b ({signal_2626, signal_1296}), .c ({signal_2665, signal_781}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_938 ( .a ({signal_2821, signal_783}), .b ({signal_2549, signal_1315}), .c ({signal_2843, signal_1267}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_939 ( .a ({signal_2626, signal_1296}), .b ({signal_2794, signal_780}), .c ({signal_2821, signal_783}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_940 ( .a ({signal_2423, signal_885}), .b ({signal_2753, signal_1280}), .c ({signal_2794, signal_780}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_941 ( .a ({signal_2711, signal_784}), .b ({signal_2488, signal_785}), .c ({signal_2753, signal_1280}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_942 ( .a ({signal_2434, signal_884}), .b ({signal_2453, signal_906}), .c ({signal_2488, signal_785}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_943 ( .a ({signal_2666, signal_1297}), .b ({signal_2548, signal_1313}), .c ({signal_2711, signal_784}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_944 ( .a ({signal_2624, signal_786}), .b ({signal_2546, signal_787}), .c ({signal_2666, signal_1297}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_945 ( .a ({signal_2530, signal_788}), .b ({signal_2424, signal_886}), .c ({signal_2546, signal_787}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_946 ( .a ({signal_2579, signal_1314}), .b ({signal_4283, signal_4281}), .c ({signal_2624, signal_786}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_947 ( .a ({signal_2547, signal_789}), .b ({signal_2523, signal_790}), .c ({signal_2579, signal_1314}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_948 ( .a ({signal_4287, signal_4285}), .b ({signal_2472, signal_904}), .c ({signal_2523, signal_790}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_949 ( .a ({signal_2490, signal_791}), .b ({signal_2524, signal_774}), .c ({signal_2547, signal_789}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_950 ( .a ({signal_2489, signal_792}), .b ({signal_2408, signal_929}), .c ({signal_2524, signal_774}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_951 ( .a ({signal_2444, signal_926}), .b ({signal_2429, signal_928}), .c ({signal_2489, signal_792}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_952 ( .a ({signal_2713, signal_793}), .b ({signal_2712, signal_777}), .c ({signal_2754, signal_1282}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_953 ( .a ({signal_2668, signal_1299}), .b ({signal_2626, signal_1296}), .c ({signal_2712, signal_777}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_954 ( .a ({signal_2667, signal_794}), .b ({signal_2525, signal_795}), .c ({signal_2713, signal_793}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_955 ( .a ({signal_2452, signal_905}), .b ({signal_2472, signal_904}), .c ({signal_2525, signal_795}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_956 ( .a ({signal_2627, signal_796}), .b ({signal_2424, signal_886}), .c ({signal_2667, signal_794}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_957 ( .a ({signal_2498, signal_797}), .b ({signal_2625, signal_798}), .c ({signal_2668, signal_1299}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_958 ( .a ({signal_2581, signal_1312}), .b ({signal_2434, signal_884}), .c ({signal_2625, signal_798}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_960 ( .a ({signal_2580, signal_799}), .b ({signal_2526, signal_800}), .c ({signal_2626, signal_1296}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_961 ( .a ({signal_2423, signal_885}), .b ({signal_2472, signal_904}), .c ({signal_2526, signal_800}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_962 ( .a ({signal_2548, signal_1313}), .b ({signal_2444, signal_926}), .c ({signal_2580, signal_799}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_963 ( .a ({signal_2465, signal_801}), .b ({signal_2527, signal_802}), .c ({signal_2548, signal_1313}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_964 ( .a ({signal_2499, signal_803}), .b ({signal_2429, signal_928}), .c ({signal_2527, signal_802}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_966 ( .a ({signal_2490, signal_791}), .b ({signal_2669, signal_773}), .c ({signal_2714, signal_1298}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_967 ( .a ({signal_2528, signal_804}), .b ({signal_2627, signal_796}), .c ({signal_2669, signal_773}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_968 ( .a ({signal_2581, signal_1312}), .b ({signal_2549, signal_1315}), .c ({signal_2627, signal_796}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_969 ( .a ({signal_2469, signal_924}), .b ({signal_2499, signal_803}), .c ({signal_2528, signal_804}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_971 ( .a ({signal_2434, signal_884}), .b ({signal_4279, signal_4277}), .c ({signal_2490, signal_791}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_972 ( .a ({signal_2466, signal_805}), .b ({signal_2529, signal_806}), .c ({signal_2549, signal_1315}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_973 ( .a ({signal_2434, signal_884}), .b ({signal_2472, signal_904}), .c ({signal_2529, signal_806}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_975 ( .a ({signal_2550, signal_807}), .b ({signal_2423, signal_885}), .c ({signal_2581, signal_1312}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_976 ( .a ({signal_2530, signal_788}), .b ({signal_2409, signal_930}), .c ({signal_2550, signal_807}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_977 ( .a ({signal_2452, signal_905}), .b ({signal_2469, signal_924}), .c ({signal_2530, signal_788}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1416 ( .a ({signal_4291, signal_4289}), .b ({signal_2324, signal_1556}), .clk (CLK), .r (Fresh[32]), .c ({signal_2364, signal_1604}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1417 ( .a ({signal_4295, signal_4293}), .b ({signal_2325, signal_1557}), .clk (CLK), .r (Fresh[33]), .c ({signal_2365, signal_1605}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1418 ( .a ({signal_4299, signal_4297}), .b ({signal_2308, signal_1558}), .clk (CLK), .r (Fresh[34]), .c ({signal_2348, signal_1606}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1419 ( .a ({signal_4303, signal_4301}), .b ({signal_2309, signal_1559}), .clk (CLK), .r (Fresh[35]), .c ({signal_2349, signal_1607}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1420 ( .a ({signal_4307, signal_4305}), .b ({signal_2326, signal_1560}), .clk (CLK), .r (Fresh[36]), .c ({signal_2366, signal_1608}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1421 ( .a ({signal_4311, signal_4309}), .b ({signal_2327, signal_1561}), .clk (CLK), .r (Fresh[37]), .c ({signal_2367, signal_1609}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1422 ( .a ({signal_4315, signal_4313}), .b ({signal_2310, signal_1562}), .clk (CLK), .r (Fresh[38]), .c ({signal_2350, signal_1610}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1423 ( .a ({signal_4319, signal_4317}), .b ({signal_2311, signal_1563}), .clk (CLK), .r (Fresh[39]), .c ({signal_2351, signal_1611}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1424 ( .a ({signal_4323, signal_4321}), .b ({signal_2328, signal_1564}), .clk (CLK), .r (Fresh[40]), .c ({signal_2368, signal_1612}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1425 ( .a ({signal_4327, signal_4325}), .b ({signal_2329, signal_1565}), .clk (CLK), .r (Fresh[41]), .c ({signal_2369, signal_1613}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1426 ( .a ({signal_4331, signal_4329}), .b ({signal_2312, signal_1566}), .clk (CLK), .r (Fresh[42]), .c ({signal_2352, signal_1614}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1427 ( .a ({signal_4335, signal_4333}), .b ({signal_2313, signal_1567}), .clk (CLK), .r (Fresh[43]), .c ({signal_2353, signal_1615}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1428 ( .a ({signal_4339, signal_4337}), .b ({signal_2330, signal_1568}), .clk (CLK), .r (Fresh[44]), .c ({signal_2370, signal_1616}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1429 ( .a ({signal_4343, signal_4341}), .b ({signal_2331, signal_1569}), .clk (CLK), .r (Fresh[45]), .c ({signal_2371, signal_1617}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1430 ( .a ({signal_4347, signal_4345}), .b ({signal_2314, signal_1570}), .clk (CLK), .r (Fresh[46]), .c ({signal_2354, signal_1618}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1431 ( .a ({signal_4351, signal_4349}), .b ({signal_2315, signal_1571}), .clk (CLK), .r (Fresh[47]), .c ({signal_2355, signal_1619}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1432 ( .a ({signal_4355, signal_4353}), .b ({signal_2356, signal_1588}), .clk (CLK), .r (Fresh[48]), .c ({signal_2388, signal_1620}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1433 ( .a ({signal_4359, signal_4357}), .b ({signal_2357, signal_1589}), .clk (CLK), .r (Fresh[49]), .c ({signal_2389, signal_1621}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1434 ( .a ({signal_4363, signal_4361}), .b ({signal_2340, signal_1590}), .clk (CLK), .r (Fresh[50]), .c ({signal_2372, signal_1622}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1435 ( .a ({signal_4367, signal_4365}), .b ({signal_2341, signal_1591}), .clk (CLK), .r (Fresh[51]), .c ({signal_2373, signal_1623}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1436 ( .a ({signal_4371, signal_4369}), .b ({signal_2358, signal_1592}), .clk (CLK), .r (Fresh[52]), .c ({signal_2390, signal_1624}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1437 ( .a ({signal_4375, signal_4373}), .b ({signal_2359, signal_1593}), .clk (CLK), .r (Fresh[53]), .c ({signal_2391, signal_1625}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1438 ( .a ({signal_4379, signal_4377}), .b ({signal_2342, signal_1594}), .clk (CLK), .r (Fresh[54]), .c ({signal_2374, signal_1626}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1439 ( .a ({signal_4383, signal_4381}), .b ({signal_2343, signal_1595}), .clk (CLK), .r (Fresh[55]), .c ({signal_2375, signal_1627}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1440 ( .a ({signal_4387, signal_4385}), .b ({signal_2360, signal_1596}), .clk (CLK), .r (Fresh[56]), .c ({signal_2392, signal_1628}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1441 ( .a ({signal_4391, signal_4389}), .b ({signal_2361, signal_1597}), .clk (CLK), .r (Fresh[57]), .c ({signal_2393, signal_1629}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1442 ( .a ({signal_4395, signal_4393}), .b ({signal_2344, signal_1598}), .clk (CLK), .r (Fresh[58]), .c ({signal_2376, signal_1630}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1443 ( .a ({signal_4399, signal_4397}), .b ({signal_2345, signal_1599}), .clk (CLK), .r (Fresh[59]), .c ({signal_2377, signal_1631}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1444 ( .a ({signal_4403, signal_4401}), .b ({signal_2362, signal_1600}), .clk (CLK), .r (Fresh[60]), .c ({signal_2394, signal_1632}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1445 ( .a ({signal_4407, signal_4405}), .b ({signal_2363, signal_1601}), .clk (CLK), .r (Fresh[61]), .c ({signal_2395, signal_1633}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1446 ( .a ({signal_4411, signal_4409}), .b ({signal_2346, signal_1602}), .clk (CLK), .r (Fresh[62]), .c ({signal_2378, signal_1634}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1447 ( .a ({signal_4415, signal_4413}), .b ({signal_2347, signal_1603}), .clk (CLK), .r (Fresh[63]), .c ({signal_2379, signal_1635}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1448 ( .a ({signal_4419, signal_4417}), .b ({signal_2364, signal_1604}), .c ({signal_2396, signal_1636}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1449 ( .a ({signal_4423, signal_4421}), .b ({signal_2365, signal_1605}), .c ({signal_2397, signal_1637}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1450 ( .a ({signal_4427, signal_4425}), .b ({signal_2348, signal_1606}), .c ({signal_2380, signal_1638}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1451 ( .a ({signal_4431, signal_4429}), .b ({signal_2349, signal_1607}), .c ({signal_2381, signal_1639}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1452 ( .a ({signal_4435, signal_4433}), .b ({signal_2366, signal_1608}), .c ({signal_2398, signal_1640}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1453 ( .a ({signal_4439, signal_4437}), .b ({signal_2367, signal_1609}), .c ({signal_2399, signal_1641}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1454 ( .a ({signal_4443, signal_4441}), .b ({signal_2350, signal_1610}), .c ({signal_2382, signal_1642}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1455 ( .a ({signal_4447, signal_4445}), .b ({signal_2351, signal_1611}), .c ({signal_2383, signal_1643}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1456 ( .a ({signal_4451, signal_4449}), .b ({signal_2368, signal_1612}), .c ({signal_2400, signal_1644}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1457 ( .a ({signal_4455, signal_4453}), .b ({signal_2369, signal_1613}), .c ({signal_2401, signal_1645}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1458 ( .a ({signal_4459, signal_4457}), .b ({signal_2352, signal_1614}), .c ({signal_2384, signal_1646}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1459 ( .a ({signal_4463, signal_4461}), .b ({signal_2353, signal_1615}), .c ({signal_2385, signal_1647}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1460 ( .a ({signal_4467, signal_4465}), .b ({signal_2370, signal_1616}), .c ({signal_2402, signal_1648}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1461 ( .a ({signal_4471, signal_4469}), .b ({signal_2371, signal_1617}), .c ({signal_2403, signal_1649}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1462 ( .a ({signal_4475, signal_4473}), .b ({signal_2354, signal_1618}), .c ({signal_2386, signal_1650}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1463 ( .a ({signal_4479, signal_4477}), .b ({signal_2355, signal_1619}), .c ({signal_2387, signal_1651}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1464 ( .a ({signal_4419, signal_4417}), .b ({signal_2388, signal_1620}), .c ({signal_2436, signal_356}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1465 ( .a ({signal_4487, signal_4483}), .b ({signal_2396, signal_1636}), .c ({signal_2437, signal_941}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1466 ( .a ({signal_4491, signal_4489}), .b ({signal_2388, signal_1620}), .c ({signal_2438, signal_942}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1467 ( .a ({signal_4423, signal_4421}), .b ({signal_2389, signal_1621}), .c ({signal_2439, signal_375}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1468 ( .a ({signal_4499, signal_4495}), .b ({signal_2397, signal_1637}), .c ({signal_2440, signal_937}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1469 ( .a ({signal_4503, signal_4501}), .b ({signal_2389, signal_1621}), .c ({signal_2441, signal_938}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1470 ( .a ({signal_4427, signal_4425}), .b ({signal_2372, signal_1622}), .c ({signal_2404, signal_394}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1471 ( .a ({signal_4511, signal_4507}), .b ({signal_2380, signal_1638}), .c ({signal_2405, signal_933}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1472 ( .a ({signal_4515, signal_4513}), .b ({signal_2372, signal_1622}), .c ({signal_2406, signal_934}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1473 ( .a ({signal_4431, signal_4429}), .b ({signal_2373, signal_1623}), .c ({signal_2407, signal_413}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1474 ( .a ({signal_4523, signal_4519}), .b ({signal_2381, signal_1639}), .c ({signal_2408, signal_929}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1475 ( .a ({signal_4527, signal_4525}), .b ({signal_2373, signal_1623}), .c ({signal_2409, signal_930}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1476 ( .a ({signal_4435, signal_4433}), .b ({signal_2390, signal_1624}), .c ({signal_2442, signal_432}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1477 ( .a ({signal_4535, signal_4531}), .b ({signal_2398, signal_1640}), .c ({signal_2443, signal_1652}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1478 ( .a ({signal_4539, signal_4537}), .b ({signal_2390, signal_1624}), .c ({signal_2444, signal_926}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1479 ( .a ({signal_4439, signal_4437}), .b ({signal_2391, signal_1625}), .c ({signal_2445, signal_451}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1480 ( .a ({signal_4547, signal_4543}), .b ({signal_2399, signal_1641}), .c ({signal_2446, signal_1653}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1481 ( .a ({signal_4551, signal_4549}), .b ({signal_2391, signal_1625}), .c ({signal_2447, signal_922}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1482 ( .a ({signal_4443, signal_4441}), .b ({signal_2374, signal_1626}), .c ({signal_2410, signal_470}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1483 ( .a ({signal_4559, signal_4555}), .b ({signal_2382, signal_1642}), .c ({signal_2411, signal_1654}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1484 ( .a ({signal_4563, signal_4561}), .b ({signal_2374, signal_1626}), .c ({signal_2412, signal_918}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1485 ( .a ({signal_4447, signal_4445}), .b ({signal_2375, signal_1627}), .c ({signal_2413, signal_489}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1486 ( .a ({signal_4571, signal_4567}), .b ({signal_2383, signal_1643}), .c ({signal_2414, signal_1655}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1487 ( .a ({signal_4575, signal_4573}), .b ({signal_2375, signal_1627}), .c ({signal_2415, signal_914}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1488 ( .a ({signal_4451, signal_4449}), .b ({signal_2392, signal_1628}), .c ({signal_2448, signal_508}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1489 ( .a ({signal_4583, signal_4579}), .b ({signal_2400, signal_1644}), .c ({signal_2449, signal_909}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1490 ( .a ({signal_4587, signal_4585}), .b ({signal_2392, signal_1628}), .c ({signal_2450, signal_910}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1491 ( .a ({signal_4455, signal_4453}), .b ({signal_2393, signal_1629}), .c ({signal_2451, signal_527}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1492 ( .a ({signal_4595, signal_4591}), .b ({signal_2401, signal_1645}), .c ({signal_2452, signal_905}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1493 ( .a ({signal_4599, signal_4597}), .b ({signal_2393, signal_1629}), .c ({signal_2453, signal_906}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1494 ( .a ({signal_4459, signal_4457}), .b ({signal_2376, signal_1630}), .c ({signal_2416, signal_546}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1495 ( .a ({signal_4607, signal_4603}), .b ({signal_2384, signal_1646}), .c ({signal_2417, signal_901}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1496 ( .a ({signal_4611, signal_4609}), .b ({signal_2376, signal_1630}), .c ({signal_2418, signal_902}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1497 ( .a ({signal_4463, signal_4461}), .b ({signal_2377, signal_1631}), .c ({signal_2419, signal_565}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1498 ( .a ({signal_4619, signal_4615}), .b ({signal_2385, signal_1647}), .c ({signal_2420, signal_897}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1499 ( .a ({signal_4623, signal_4621}), .b ({signal_2377, signal_1631}), .c ({signal_2421, signal_898}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1500 ( .a ({signal_4467, signal_4465}), .b ({signal_2394, signal_1632}), .c ({signal_2454, signal_584}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1501 ( .a ({signal_4631, signal_4627}), .b ({signal_2402, signal_1648}), .c ({signal_2455, signal_893}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1502 ( .a ({signal_4635, signal_4633}), .b ({signal_2394, signal_1632}), .c ({signal_2456, signal_894}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1503 ( .a ({signal_4471, signal_4469}), .b ({signal_2395, signal_1633}), .c ({signal_2457, signal_603}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1504 ( .a ({signal_4643, signal_4639}), .b ({signal_2403, signal_1649}), .c ({signal_2458, signal_889}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1505 ( .a ({signal_4647, signal_4645}), .b ({signal_2395, signal_1633}), .c ({signal_2459, signal_890}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1506 ( .a ({signal_4475, signal_4473}), .b ({signal_2378, signal_1634}), .c ({signal_2422, signal_622}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1507 ( .a ({signal_4655, signal_4651}), .b ({signal_2386, signal_1650}), .c ({signal_2423, signal_885}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1508 ( .a ({signal_4659, signal_4657}), .b ({signal_2378, signal_1634}), .c ({signal_2424, signal_886}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1509 ( .a ({signal_4479, signal_4477}), .b ({signal_2379, signal_1635}), .c ({signal_2425, signal_641}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1510 ( .a ({signal_4667, signal_4663}), .b ({signal_2387, signal_1651}), .c ({signal_2426, signal_881}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1511 ( .a ({signal_4671, signal_4669}), .b ({signal_2379, signal_1635}), .c ({signal_2427, signal_882}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1512 ( .a ({signal_4251, signal_4249}), .b ({signal_2446, signal_1653}), .c ({signal_2491, signal_683}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1513 ( .a ({signal_4675, signal_4673}), .b ({signal_2427, signal_882}), .c ({signal_2460, signal_687}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1514 ( .a ({signal_2446, signal_1653}), .b ({signal_2418, signal_902}), .c ({signal_2492, signal_689}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1515 ( .a ({signal_4247, signal_4245}), .b ({signal_2437, signal_941}), .c ({signal_2493, signal_691}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1516 ( .a ({signal_4263, signal_4261}), .b ({signal_2411, signal_1654}), .c ({signal_2461, signal_721}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1517 ( .a ({signal_4679, signal_4677}), .b ({signal_2456, signal_894}), .c ({signal_2494, signal_725}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1518 ( .a ({signal_2411, signal_1654}), .b ({signal_2421, signal_898}), .c ({signal_2462, signal_727}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1519 ( .a ({signal_4259, signal_4257}), .b ({signal_2440, signal_937}), .c ({signal_2495, signal_729}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1520 ( .a ({signal_4275, signal_4273}), .b ({signal_2414, signal_1655}), .c ({signal_2463, signal_759}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1521 ( .a ({signal_4683, signal_4681}), .b ({signal_2459, signal_890}), .c ({signal_2496, signal_763}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1522 ( .a ({signal_2414, signal_1655}), .b ({signal_2450, signal_910}), .c ({signal_2497, signal_765}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1523 ( .a ({signal_4271, signal_4269}), .b ({signal_2405, signal_933}), .c ({signal_2464, signal_767}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1524 ( .a ({signal_4287, signal_4285}), .b ({signal_2443, signal_1652}), .c ({signal_2498, signal_797}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1525 ( .a ({signal_4687, signal_4685}), .b ({signal_2424, signal_886}), .c ({signal_2465, signal_801}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1526 ( .a ({signal_2443, signal_1652}), .b ({signal_2453, signal_906}), .c ({signal_2499, signal_803}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1527 ( .a ({signal_4283, signal_4281}), .b ({signal_2408, signal_929}), .c ({signal_2466, signal_805}) ) ;
    buf_clk cell_1723 ( .C (CLK), .D (signal_3134), .Q (signal_3135) ) ;
    buf_clk cell_1727 ( .C (CLK), .D (signal_3138), .Q (signal_3139) ) ;
    buf_clk cell_1731 ( .C (CLK), .D (signal_3142), .Q (signal_3143) ) ;
    buf_clk cell_1735 ( .C (CLK), .D (signal_3146), .Q (signal_3147) ) ;
    buf_clk cell_1739 ( .C (CLK), .D (signal_3150), .Q (signal_3151) ) ;
    buf_clk cell_1743 ( .C (CLK), .D (signal_3154), .Q (signal_3155) ) ;
    buf_clk cell_1747 ( .C (CLK), .D (signal_3158), .Q (signal_3159) ) ;
    buf_clk cell_1751 ( .C (CLK), .D (signal_3162), .Q (signal_3163) ) ;
    buf_clk cell_1755 ( .C (CLK), .D (signal_3166), .Q (signal_3167) ) ;
    buf_clk cell_1759 ( .C (CLK), .D (signal_3170), .Q (signal_3171) ) ;
    buf_clk cell_1763 ( .C (CLK), .D (signal_3174), .Q (signal_3175) ) ;
    buf_clk cell_1767 ( .C (CLK), .D (signal_3178), .Q (signal_3179) ) ;
    buf_clk cell_1771 ( .C (CLK), .D (signal_3182), .Q (signal_3183) ) ;
    buf_clk cell_1775 ( .C (CLK), .D (signal_3186), .Q (signal_3187) ) ;
    buf_clk cell_1779 ( .C (CLK), .D (signal_3190), .Q (signal_3191) ) ;
    buf_clk cell_1783 ( .C (CLK), .D (signal_3194), .Q (signal_3195) ) ;
    buf_clk cell_1787 ( .C (CLK), .D (signal_3198), .Q (signal_3199) ) ;
    buf_clk cell_1791 ( .C (CLK), .D (signal_3202), .Q (signal_3203) ) ;
    buf_clk cell_1795 ( .C (CLK), .D (signal_3206), .Q (signal_3207) ) ;
    buf_clk cell_1799 ( .C (CLK), .D (signal_3210), .Q (signal_3211) ) ;
    buf_clk cell_1803 ( .C (CLK), .D (signal_3214), .Q (signal_3215) ) ;
    buf_clk cell_1807 ( .C (CLK), .D (signal_3218), .Q (signal_3219) ) ;
    buf_clk cell_1811 ( .C (CLK), .D (signal_3222), .Q (signal_3223) ) ;
    buf_clk cell_1815 ( .C (CLK), .D (signal_3226), .Q (signal_3227) ) ;
    buf_clk cell_1819 ( .C (CLK), .D (signal_3230), .Q (signal_3231) ) ;
    buf_clk cell_1823 ( .C (CLK), .D (signal_3234), .Q (signal_3235) ) ;
    buf_clk cell_1827 ( .C (CLK), .D (signal_3238), .Q (signal_3239) ) ;
    buf_clk cell_1831 ( .C (CLK), .D (signal_3242), .Q (signal_3243) ) ;
    buf_clk cell_1835 ( .C (CLK), .D (signal_3246), .Q (signal_3247) ) ;
    buf_clk cell_1839 ( .C (CLK), .D (signal_3250), .Q (signal_3251) ) ;
    buf_clk cell_1843 ( .C (CLK), .D (signal_3254), .Q (signal_3255) ) ;
    buf_clk cell_1847 ( .C (CLK), .D (signal_3258), .Q (signal_3259) ) ;
    buf_clk cell_1851 ( .C (CLK), .D (signal_3262), .Q (signal_3263) ) ;
    buf_clk cell_1855 ( .C (CLK), .D (signal_3266), .Q (signal_3267) ) ;
    buf_clk cell_1859 ( .C (CLK), .D (signal_3270), .Q (signal_3271) ) ;
    buf_clk cell_1863 ( .C (CLK), .D (signal_3274), .Q (signal_3275) ) ;
    buf_clk cell_1867 ( .C (CLK), .D (signal_3278), .Q (signal_3279) ) ;
    buf_clk cell_1871 ( .C (CLK), .D (signal_3282), .Q (signal_3283) ) ;
    buf_clk cell_1875 ( .C (CLK), .D (signal_3286), .Q (signal_3287) ) ;
    buf_clk cell_1879 ( .C (CLK), .D (signal_3290), .Q (signal_3291) ) ;
    buf_clk cell_1883 ( .C (CLK), .D (signal_3294), .Q (signal_3295) ) ;
    buf_clk cell_1887 ( .C (CLK), .D (signal_3298), .Q (signal_3299) ) ;
    buf_clk cell_1891 ( .C (CLK), .D (signal_3302), .Q (signal_3303) ) ;
    buf_clk cell_1895 ( .C (CLK), .D (signal_3306), .Q (signal_3307) ) ;
    buf_clk cell_1899 ( .C (CLK), .D (signal_3310), .Q (signal_3311) ) ;
    buf_clk cell_1903 ( .C (CLK), .D (signal_3314), .Q (signal_3315) ) ;
    buf_clk cell_1907 ( .C (CLK), .D (signal_3318), .Q (signal_3319) ) ;
    buf_clk cell_1911 ( .C (CLK), .D (signal_3322), .Q (signal_3323) ) ;
    buf_clk cell_1915 ( .C (CLK), .D (signal_3326), .Q (signal_3327) ) ;
    buf_clk cell_1919 ( .C (CLK), .D (signal_3330), .Q (signal_3331) ) ;
    buf_clk cell_1923 ( .C (CLK), .D (signal_3334), .Q (signal_3335) ) ;
    buf_clk cell_1927 ( .C (CLK), .D (signal_3338), .Q (signal_3339) ) ;
    buf_clk cell_1931 ( .C (CLK), .D (signal_3342), .Q (signal_3343) ) ;
    buf_clk cell_1935 ( .C (CLK), .D (signal_3346), .Q (signal_3347) ) ;
    buf_clk cell_1939 ( .C (CLK), .D (signal_3350), .Q (signal_3351) ) ;
    buf_clk cell_1943 ( .C (CLK), .D (signal_3354), .Q (signal_3355) ) ;
    buf_clk cell_1947 ( .C (CLK), .D (signal_3358), .Q (signal_3359) ) ;
    buf_clk cell_1951 ( .C (CLK), .D (signal_3362), .Q (signal_3363) ) ;
    buf_clk cell_1955 ( .C (CLK), .D (signal_3366), .Q (signal_3367) ) ;
    buf_clk cell_1959 ( .C (CLK), .D (signal_3370), .Q (signal_3371) ) ;
    buf_clk cell_1963 ( .C (CLK), .D (signal_3374), .Q (signal_3375) ) ;
    buf_clk cell_1967 ( .C (CLK), .D (signal_3378), .Q (signal_3379) ) ;
    buf_clk cell_1971 ( .C (CLK), .D (signal_3382), .Q (signal_3383) ) ;
    buf_clk cell_1975 ( .C (CLK), .D (signal_3386), .Q (signal_3387) ) ;
    buf_clk cell_1979 ( .C (CLK), .D (signal_3390), .Q (signal_3391) ) ;
    buf_clk cell_1983 ( .C (CLK), .D (signal_3394), .Q (signal_3395) ) ;
    buf_clk cell_1987 ( .C (CLK), .D (signal_3398), .Q (signal_3399) ) ;
    buf_clk cell_1991 ( .C (CLK), .D (signal_3402), .Q (signal_3403) ) ;
    buf_clk cell_1995 ( .C (CLK), .D (signal_3406), .Q (signal_3407) ) ;
    buf_clk cell_1999 ( .C (CLK), .D (signal_3410), .Q (signal_3411) ) ;
    buf_clk cell_2003 ( .C (CLK), .D (signal_3414), .Q (signal_3415) ) ;
    buf_clk cell_2007 ( .C (CLK), .D (signal_3418), .Q (signal_3419) ) ;
    buf_clk cell_2011 ( .C (CLK), .D (signal_3422), .Q (signal_3423) ) ;
    buf_clk cell_2015 ( .C (CLK), .D (signal_3426), .Q (signal_3427) ) ;
    buf_clk cell_2019 ( .C (CLK), .D (signal_3430), .Q (signal_3431) ) ;
    buf_clk cell_2023 ( .C (CLK), .D (signal_3434), .Q (signal_3435) ) ;
    buf_clk cell_2027 ( .C (CLK), .D (signal_3438), .Q (signal_3439) ) ;
    buf_clk cell_2031 ( .C (CLK), .D (signal_3442), .Q (signal_3443) ) ;
    buf_clk cell_2035 ( .C (CLK), .D (signal_3446), .Q (signal_3447) ) ;
    buf_clk cell_2039 ( .C (CLK), .D (signal_3450), .Q (signal_3451) ) ;
    buf_clk cell_2043 ( .C (CLK), .D (signal_3454), .Q (signal_3455) ) ;
    buf_clk cell_2047 ( .C (CLK), .D (signal_3458), .Q (signal_3459) ) ;
    buf_clk cell_2051 ( .C (CLK), .D (signal_3462), .Q (signal_3463) ) ;
    buf_clk cell_2055 ( .C (CLK), .D (signal_3466), .Q (signal_3467) ) ;
    buf_clk cell_2059 ( .C (CLK), .D (signal_3470), .Q (signal_3471) ) ;
    buf_clk cell_2063 ( .C (CLK), .D (signal_3474), .Q (signal_3475) ) ;
    buf_clk cell_2067 ( .C (CLK), .D (signal_3478), .Q (signal_3479) ) ;
    buf_clk cell_2071 ( .C (CLK), .D (signal_3482), .Q (signal_3483) ) ;
    buf_clk cell_2075 ( .C (CLK), .D (signal_3486), .Q (signal_3487) ) ;
    buf_clk cell_2079 ( .C (CLK), .D (signal_3490), .Q (signal_3491) ) ;
    buf_clk cell_2083 ( .C (CLK), .D (signal_3494), .Q (signal_3495) ) ;
    buf_clk cell_2087 ( .C (CLK), .D (signal_3498), .Q (signal_3499) ) ;
    buf_clk cell_2091 ( .C (CLK), .D (signal_3502), .Q (signal_3503) ) ;
    buf_clk cell_2095 ( .C (CLK), .D (signal_3506), .Q (signal_3507) ) ;
    buf_clk cell_2099 ( .C (CLK), .D (signal_3510), .Q (signal_3511) ) ;
    buf_clk cell_2103 ( .C (CLK), .D (signal_3514), .Q (signal_3515) ) ;
    buf_clk cell_2107 ( .C (CLK), .D (signal_3518), .Q (signal_3519) ) ;
    buf_clk cell_2111 ( .C (CLK), .D (signal_3522), .Q (signal_3523) ) ;
    buf_clk cell_2115 ( .C (CLK), .D (signal_3526), .Q (signal_3527) ) ;
    buf_clk cell_2119 ( .C (CLK), .D (signal_3530), .Q (signal_3531) ) ;
    buf_clk cell_2123 ( .C (CLK), .D (signal_3534), .Q (signal_3535) ) ;
    buf_clk cell_2127 ( .C (CLK), .D (signal_3538), .Q (signal_3539) ) ;
    buf_clk cell_2131 ( .C (CLK), .D (signal_3542), .Q (signal_3543) ) ;
    buf_clk cell_2135 ( .C (CLK), .D (signal_3546), .Q (signal_3547) ) ;
    buf_clk cell_2139 ( .C (CLK), .D (signal_3550), .Q (signal_3551) ) ;
    buf_clk cell_2143 ( .C (CLK), .D (signal_3554), .Q (signal_3555) ) ;
    buf_clk cell_2147 ( .C (CLK), .D (signal_3558), .Q (signal_3559) ) ;
    buf_clk cell_2151 ( .C (CLK), .D (signal_3562), .Q (signal_3563) ) ;
    buf_clk cell_2155 ( .C (CLK), .D (signal_3566), .Q (signal_3567) ) ;
    buf_clk cell_2159 ( .C (CLK), .D (signal_3570), .Q (signal_3571) ) ;
    buf_clk cell_2163 ( .C (CLK), .D (signal_3574), .Q (signal_3575) ) ;
    buf_clk cell_2167 ( .C (CLK), .D (signal_3578), .Q (signal_3579) ) ;
    buf_clk cell_2171 ( .C (CLK), .D (signal_3582), .Q (signal_3583) ) ;
    buf_clk cell_2175 ( .C (CLK), .D (signal_3586), .Q (signal_3587) ) ;
    buf_clk cell_2179 ( .C (CLK), .D (signal_3590), .Q (signal_3591) ) ;
    buf_clk cell_2183 ( .C (CLK), .D (signal_3594), .Q (signal_3595) ) ;
    buf_clk cell_2187 ( .C (CLK), .D (signal_3598), .Q (signal_3599) ) ;
    buf_clk cell_2191 ( .C (CLK), .D (signal_3602), .Q (signal_3603) ) ;
    buf_clk cell_2195 ( .C (CLK), .D (signal_3606), .Q (signal_3607) ) ;
    buf_clk cell_2199 ( .C (CLK), .D (signal_3610), .Q (signal_3611) ) ;
    buf_clk cell_2203 ( .C (CLK), .D (signal_3614), .Q (signal_3615) ) ;
    buf_clk cell_2207 ( .C (CLK), .D (signal_3618), .Q (signal_3619) ) ;
    buf_clk cell_2211 ( .C (CLK), .D (signal_3622), .Q (signal_3623) ) ;
    buf_clk cell_2215 ( .C (CLK), .D (signal_3626), .Q (signal_3627) ) ;
    buf_clk cell_2219 ( .C (CLK), .D (signal_3630), .Q (signal_3631) ) ;
    buf_clk cell_2223 ( .C (CLK), .D (signal_3634), .Q (signal_3635) ) ;
    buf_clk cell_2227 ( .C (CLK), .D (signal_3638), .Q (signal_3639) ) ;
    buf_clk cell_2231 ( .C (CLK), .D (signal_3642), .Q (signal_3643) ) ;
    buf_clk cell_2235 ( .C (CLK), .D (signal_3646), .Q (signal_3647) ) ;
    buf_clk cell_2239 ( .C (CLK), .D (signal_3650), .Q (signal_3651) ) ;
    buf_clk cell_2243 ( .C (CLK), .D (signal_3654), .Q (signal_3655) ) ;
    buf_clk cell_2247 ( .C (CLK), .D (signal_3658), .Q (signal_3659) ) ;
    buf_clk cell_2251 ( .C (CLK), .D (signal_3662), .Q (signal_3663) ) ;
    buf_clk cell_2255 ( .C (CLK), .D (signal_3666), .Q (signal_3667) ) ;
    buf_clk cell_2259 ( .C (CLK), .D (signal_3670), .Q (signal_3671) ) ;
    buf_clk cell_2263 ( .C (CLK), .D (signal_3674), .Q (signal_3675) ) ;
    buf_clk cell_2267 ( .C (CLK), .D (signal_3678), .Q (signal_3679) ) ;
    buf_clk cell_2271 ( .C (CLK), .D (signal_3682), .Q (signal_3683) ) ;
    buf_clk cell_2275 ( .C (CLK), .D (signal_3686), .Q (signal_3687) ) ;
    buf_clk cell_2279 ( .C (CLK), .D (signal_3690), .Q (signal_3691) ) ;
    buf_clk cell_2283 ( .C (CLK), .D (signal_3694), .Q (signal_3695) ) ;
    buf_clk cell_2287 ( .C (CLK), .D (signal_3698), .Q (signal_3699) ) ;
    buf_clk cell_2291 ( .C (CLK), .D (signal_3702), .Q (signal_3703) ) ;
    buf_clk cell_2295 ( .C (CLK), .D (signal_3706), .Q (signal_3707) ) ;
    buf_clk cell_2299 ( .C (CLK), .D (signal_3710), .Q (signal_3711) ) ;
    buf_clk cell_2303 ( .C (CLK), .D (signal_3714), .Q (signal_3715) ) ;
    buf_clk cell_2307 ( .C (CLK), .D (signal_3718), .Q (signal_3719) ) ;
    buf_clk cell_2311 ( .C (CLK), .D (signal_3722), .Q (signal_3723) ) ;
    buf_clk cell_2315 ( .C (CLK), .D (signal_3726), .Q (signal_3727) ) ;
    buf_clk cell_2319 ( .C (CLK), .D (signal_3730), .Q (signal_3731) ) ;
    buf_clk cell_2323 ( .C (CLK), .D (signal_3734), .Q (signal_3735) ) ;
    buf_clk cell_2327 ( .C (CLK), .D (signal_3738), .Q (signal_3739) ) ;
    buf_clk cell_2331 ( .C (CLK), .D (signal_3742), .Q (signal_3743) ) ;
    buf_clk cell_2335 ( .C (CLK), .D (signal_3746), .Q (signal_3747) ) ;
    buf_clk cell_2339 ( .C (CLK), .D (signal_3750), .Q (signal_3751) ) ;
    buf_clk cell_2343 ( .C (CLK), .D (signal_3754), .Q (signal_3755) ) ;
    buf_clk cell_2347 ( .C (CLK), .D (signal_3758), .Q (signal_3759) ) ;
    buf_clk cell_2351 ( .C (CLK), .D (signal_3762), .Q (signal_3763) ) ;
    buf_clk cell_2355 ( .C (CLK), .D (signal_3766), .Q (signal_3767) ) ;
    buf_clk cell_2359 ( .C (CLK), .D (signal_3770), .Q (signal_3771) ) ;
    buf_clk cell_2363 ( .C (CLK), .D (signal_3774), .Q (signal_3775) ) ;
    buf_clk cell_2367 ( .C (CLK), .D (signal_3778), .Q (signal_3779) ) ;
    buf_clk cell_2371 ( .C (CLK), .D (signal_3782), .Q (signal_3783) ) ;
    buf_clk cell_2375 ( .C (CLK), .D (signal_3786), .Q (signal_3787) ) ;
    buf_clk cell_2379 ( .C (CLK), .D (signal_3790), .Q (signal_3791) ) ;
    buf_clk cell_2383 ( .C (CLK), .D (signal_3794), .Q (signal_3795) ) ;
    buf_clk cell_2387 ( .C (CLK), .D (signal_3798), .Q (signal_3799) ) ;
    buf_clk cell_2391 ( .C (CLK), .D (signal_3802), .Q (signal_3803) ) ;
    buf_clk cell_2395 ( .C (CLK), .D (signal_3806), .Q (signal_3807) ) ;
    buf_clk cell_2399 ( .C (CLK), .D (signal_3810), .Q (signal_3811) ) ;
    buf_clk cell_2403 ( .C (CLK), .D (signal_3814), .Q (signal_3815) ) ;
    buf_clk cell_2407 ( .C (CLK), .D (signal_3818), .Q (signal_3819) ) ;
    buf_clk cell_2411 ( .C (CLK), .D (signal_3822), .Q (signal_3823) ) ;
    buf_clk cell_2415 ( .C (CLK), .D (signal_3826), .Q (signal_3827) ) ;
    buf_clk cell_2419 ( .C (CLK), .D (signal_3830), .Q (signal_3831) ) ;
    buf_clk cell_2423 ( .C (CLK), .D (signal_3834), .Q (signal_3835) ) ;
    buf_clk cell_2427 ( .C (CLK), .D (signal_3838), .Q (signal_3839) ) ;
    buf_clk cell_2431 ( .C (CLK), .D (signal_3842), .Q (signal_3843) ) ;
    buf_clk cell_2435 ( .C (CLK), .D (signal_3846), .Q (signal_3847) ) ;
    buf_clk cell_2439 ( .C (CLK), .D (signal_3850), .Q (signal_3851) ) ;
    buf_clk cell_2443 ( .C (CLK), .D (signal_3854), .Q (signal_3855) ) ;
    buf_clk cell_2447 ( .C (CLK), .D (signal_3858), .Q (signal_3859) ) ;
    buf_clk cell_2451 ( .C (CLK), .D (signal_3862), .Q (signal_3863) ) ;
    buf_clk cell_2455 ( .C (CLK), .D (signal_3866), .Q (signal_3867) ) ;
    buf_clk cell_2459 ( .C (CLK), .D (signal_3870), .Q (signal_3871) ) ;
    buf_clk cell_2463 ( .C (CLK), .D (signal_3874), .Q (signal_3875) ) ;
    buf_clk cell_2467 ( .C (CLK), .D (signal_3878), .Q (signal_3879) ) ;
    buf_clk cell_2471 ( .C (CLK), .D (signal_3882), .Q (signal_3883) ) ;
    buf_clk cell_2475 ( .C (CLK), .D (signal_3886), .Q (signal_3887) ) ;
    buf_clk cell_2479 ( .C (CLK), .D (signal_3890), .Q (signal_3891) ) ;
    buf_clk cell_2483 ( .C (CLK), .D (signal_3894), .Q (signal_3895) ) ;
    buf_clk cell_2487 ( .C (CLK), .D (signal_3898), .Q (signal_3899) ) ;
    buf_clk cell_2491 ( .C (CLK), .D (signal_3902), .Q (signal_3903) ) ;
    buf_clk cell_2495 ( .C (CLK), .D (signal_3906), .Q (signal_3907) ) ;
    buf_clk cell_2499 ( .C (CLK), .D (signal_3910), .Q (signal_3911) ) ;
    buf_clk cell_2503 ( .C (CLK), .D (signal_3914), .Q (signal_3915) ) ;
    buf_clk cell_2507 ( .C (CLK), .D (signal_3918), .Q (signal_3919) ) ;
    buf_clk cell_2511 ( .C (CLK), .D (signal_3922), .Q (signal_3923) ) ;
    buf_clk cell_2515 ( .C (CLK), .D (signal_3926), .Q (signal_3927) ) ;
    buf_clk cell_2519 ( .C (CLK), .D (signal_3930), .Q (signal_3931) ) ;
    buf_clk cell_2523 ( .C (CLK), .D (signal_3934), .Q (signal_3935) ) ;
    buf_clk cell_2527 ( .C (CLK), .D (signal_3938), .Q (signal_3939) ) ;
    buf_clk cell_2531 ( .C (CLK), .D (signal_3942), .Q (signal_3943) ) ;
    buf_clk cell_2535 ( .C (CLK), .D (signal_3946), .Q (signal_3947) ) ;
    buf_clk cell_2539 ( .C (CLK), .D (signal_3950), .Q (signal_3951) ) ;
    buf_clk cell_2543 ( .C (CLK), .D (signal_3954), .Q (signal_3955) ) ;
    buf_clk cell_2547 ( .C (CLK), .D (signal_3958), .Q (signal_3959) ) ;
    buf_clk cell_2551 ( .C (CLK), .D (signal_3962), .Q (signal_3963) ) ;
    buf_clk cell_2555 ( .C (CLK), .D (signal_3966), .Q (signal_3967) ) ;
    buf_clk cell_2559 ( .C (CLK), .D (signal_3970), .Q (signal_3971) ) ;
    buf_clk cell_2563 ( .C (CLK), .D (signal_3974), .Q (signal_3975) ) ;
    buf_clk cell_2567 ( .C (CLK), .D (signal_3978), .Q (signal_3979) ) ;
    buf_clk cell_2571 ( .C (CLK), .D (signal_3982), .Q (signal_3983) ) ;
    buf_clk cell_2575 ( .C (CLK), .D (signal_3986), .Q (signal_3987) ) ;
    buf_clk cell_2579 ( .C (CLK), .D (signal_3990), .Q (signal_3991) ) ;
    buf_clk cell_2583 ( .C (CLK), .D (signal_3994), .Q (signal_3995) ) ;
    buf_clk cell_2587 ( .C (CLK), .D (signal_3998), .Q (signal_3999) ) ;
    buf_clk cell_2591 ( .C (CLK), .D (signal_4002), .Q (signal_4003) ) ;
    buf_clk cell_2595 ( .C (CLK), .D (signal_4006), .Q (signal_4007) ) ;
    buf_clk cell_2599 ( .C (CLK), .D (signal_4010), .Q (signal_4011) ) ;
    buf_clk cell_2603 ( .C (CLK), .D (signal_4014), .Q (signal_4015) ) ;
    buf_clk cell_2607 ( .C (CLK), .D (signal_4018), .Q (signal_4019) ) ;
    buf_clk cell_2611 ( .C (CLK), .D (signal_4022), .Q (signal_4023) ) ;
    buf_clk cell_2615 ( .C (CLK), .D (signal_4026), .Q (signal_4027) ) ;
    buf_clk cell_2619 ( .C (CLK), .D (signal_4030), .Q (signal_4031) ) ;
    buf_clk cell_2623 ( .C (CLK), .D (signal_4034), .Q (signal_4035) ) ;
    buf_clk cell_2627 ( .C (CLK), .D (signal_4038), .Q (signal_4039) ) ;
    buf_clk cell_2631 ( .C (CLK), .D (signal_4042), .Q (signal_4043) ) ;
    buf_clk cell_2635 ( .C (CLK), .D (signal_4046), .Q (signal_4047) ) ;
    buf_clk cell_2639 ( .C (CLK), .D (signal_4050), .Q (signal_4051) ) ;
    buf_clk cell_2643 ( .C (CLK), .D (signal_4054), .Q (signal_4055) ) ;
    buf_clk cell_2647 ( .C (CLK), .D (signal_4058), .Q (signal_4059) ) ;
    buf_clk cell_2651 ( .C (CLK), .D (signal_4062), .Q (signal_4063) ) ;
    buf_clk cell_2655 ( .C (CLK), .D (signal_4066), .Q (signal_4067) ) ;
    buf_clk cell_2659 ( .C (CLK), .D (signal_4070), .Q (signal_4071) ) ;
    buf_clk cell_2663 ( .C (CLK), .D (signal_4074), .Q (signal_4075) ) ;
    buf_clk cell_2667 ( .C (CLK), .D (signal_4078), .Q (signal_4079) ) ;
    buf_clk cell_2671 ( .C (CLK), .D (signal_4082), .Q (signal_4083) ) ;
    buf_clk cell_2675 ( .C (CLK), .D (signal_4086), .Q (signal_4087) ) ;
    buf_clk cell_2679 ( .C (CLK), .D (signal_4090), .Q (signal_4091) ) ;
    buf_clk cell_2683 ( .C (CLK), .D (signal_4094), .Q (signal_4095) ) ;
    buf_clk cell_2687 ( .C (CLK), .D (signal_4098), .Q (signal_4099) ) ;
    buf_clk cell_2691 ( .C (CLK), .D (signal_4102), .Q (signal_4103) ) ;
    buf_clk cell_2695 ( .C (CLK), .D (signal_4106), .Q (signal_4107) ) ;
    buf_clk cell_2699 ( .C (CLK), .D (signal_4110), .Q (signal_4111) ) ;
    buf_clk cell_2703 ( .C (CLK), .D (signal_4114), .Q (signal_4115) ) ;
    buf_clk cell_2707 ( .C (CLK), .D (signal_4118), .Q (signal_4119) ) ;
    buf_clk cell_2711 ( .C (CLK), .D (signal_4122), .Q (signal_4123) ) ;
    buf_clk cell_2715 ( .C (CLK), .D (signal_4126), .Q (signal_4127) ) ;
    buf_clk cell_2719 ( .C (CLK), .D (signal_4130), .Q (signal_4131) ) ;
    buf_clk cell_2723 ( .C (CLK), .D (signal_4134), .Q (signal_4135) ) ;
    buf_clk cell_2727 ( .C (CLK), .D (signal_4138), .Q (signal_4139) ) ;
    buf_clk cell_2731 ( .C (CLK), .D (signal_4142), .Q (signal_4143) ) ;
    buf_clk cell_2735 ( .C (CLK), .D (signal_4146), .Q (signal_4147) ) ;
    buf_clk cell_2739 ( .C (CLK), .D (signal_4150), .Q (signal_4151) ) ;
    buf_clk cell_2743 ( .C (CLK), .D (signal_4154), .Q (signal_4155) ) ;
    buf_clk cell_2747 ( .C (CLK), .D (signal_4158), .Q (signal_4159) ) ;
    buf_clk cell_2751 ( .C (CLK), .D (signal_4162), .Q (signal_4163) ) ;
    buf_clk cell_2755 ( .C (CLK), .D (signal_4166), .Q (signal_4167) ) ;
    buf_clk cell_2759 ( .C (CLK), .D (signal_4170), .Q (signal_4171) ) ;
    buf_clk cell_2763 ( .C (CLK), .D (signal_4174), .Q (signal_4175) ) ;
    buf_clk cell_2767 ( .C (CLK), .D (signal_4178), .Q (signal_4179) ) ;
    buf_clk cell_2771 ( .C (CLK), .D (signal_4182), .Q (signal_4183) ) ;
    buf_clk cell_2775 ( .C (CLK), .D (signal_4186), .Q (signal_4187) ) ;
    buf_clk cell_2779 ( .C (CLK), .D (signal_4190), .Q (signal_4191) ) ;
    buf_clk cell_2783 ( .C (CLK), .D (signal_4194), .Q (signal_4195) ) ;
    buf_clk cell_2787 ( .C (CLK), .D (signal_4198), .Q (signal_4199) ) ;
    buf_clk cell_2791 ( .C (CLK), .D (signal_4202), .Q (signal_4203) ) ;
    buf_clk cell_2795 ( .C (CLK), .D (signal_4206), .Q (signal_4207) ) ;
    buf_clk cell_2799 ( .C (CLK), .D (signal_4210), .Q (signal_4211) ) ;
    buf_clk cell_2803 ( .C (CLK), .D (signal_4214), .Q (signal_4215) ) ;
    buf_clk cell_2807 ( .C (CLK), .D (signal_4218), .Q (signal_4219) ) ;
    buf_clk cell_2811 ( .C (CLK), .D (signal_4222), .Q (signal_4223) ) ;
    buf_clk cell_2815 ( .C (CLK), .D (signal_4226), .Q (signal_4227) ) ;
    buf_clk cell_2819 ( .C (CLK), .D (signal_4230), .Q (signal_4231) ) ;
    buf_clk cell_2823 ( .C (CLK), .D (signal_4234), .Q (signal_4235) ) ;
    buf_clk cell_2827 ( .C (CLK), .D (signal_4238), .Q (signal_4239) ) ;
    buf_clk cell_2829 ( .C (CLK), .D (signal_4240), .Q (signal_4241) ) ;
    buf_clk cell_2831 ( .C (CLK), .D (signal_4242), .Q (signal_4243) ) ;
    buf_clk cell_2833 ( .C (CLK), .D (signal_4244), .Q (signal_4245) ) ;
    buf_clk cell_2835 ( .C (CLK), .D (signal_4246), .Q (signal_4247) ) ;
    buf_clk cell_2837 ( .C (CLK), .D (signal_4248), .Q (signal_4249) ) ;
    buf_clk cell_2839 ( .C (CLK), .D (signal_4250), .Q (signal_4251) ) ;
    buf_clk cell_2841 ( .C (CLK), .D (signal_4252), .Q (signal_4253) ) ;
    buf_clk cell_2843 ( .C (CLK), .D (signal_4254), .Q (signal_4255) ) ;
    buf_clk cell_2845 ( .C (CLK), .D (signal_4256), .Q (signal_4257) ) ;
    buf_clk cell_2847 ( .C (CLK), .D (signal_4258), .Q (signal_4259) ) ;
    buf_clk cell_2849 ( .C (CLK), .D (signal_4260), .Q (signal_4261) ) ;
    buf_clk cell_2851 ( .C (CLK), .D (signal_4262), .Q (signal_4263) ) ;
    buf_clk cell_2853 ( .C (CLK), .D (signal_4264), .Q (signal_4265) ) ;
    buf_clk cell_2855 ( .C (CLK), .D (signal_4266), .Q (signal_4267) ) ;
    buf_clk cell_2857 ( .C (CLK), .D (signal_4268), .Q (signal_4269) ) ;
    buf_clk cell_2859 ( .C (CLK), .D (signal_4270), .Q (signal_4271) ) ;
    buf_clk cell_2861 ( .C (CLK), .D (signal_4272), .Q (signal_4273) ) ;
    buf_clk cell_2863 ( .C (CLK), .D (signal_4274), .Q (signal_4275) ) ;
    buf_clk cell_2865 ( .C (CLK), .D (signal_4276), .Q (signal_4277) ) ;
    buf_clk cell_2867 ( .C (CLK), .D (signal_4278), .Q (signal_4279) ) ;
    buf_clk cell_2869 ( .C (CLK), .D (signal_4280), .Q (signal_4281) ) ;
    buf_clk cell_2871 ( .C (CLK), .D (signal_4282), .Q (signal_4283) ) ;
    buf_clk cell_2873 ( .C (CLK), .D (signal_4284), .Q (signal_4285) ) ;
    buf_clk cell_2875 ( .C (CLK), .D (signal_4286), .Q (signal_4287) ) ;
    buf_clk cell_3005 ( .C (CLK), .D (signal_4416), .Q (signal_4417) ) ;
    buf_clk cell_3007 ( .C (CLK), .D (signal_4418), .Q (signal_4419) ) ;
    buf_clk cell_3009 ( .C (CLK), .D (signal_4420), .Q (signal_4421) ) ;
    buf_clk cell_3011 ( .C (CLK), .D (signal_4422), .Q (signal_4423) ) ;
    buf_clk cell_3013 ( .C (CLK), .D (signal_4424), .Q (signal_4425) ) ;
    buf_clk cell_3015 ( .C (CLK), .D (signal_4426), .Q (signal_4427) ) ;
    buf_clk cell_3017 ( .C (CLK), .D (signal_4428), .Q (signal_4429) ) ;
    buf_clk cell_3019 ( .C (CLK), .D (signal_4430), .Q (signal_4431) ) ;
    buf_clk cell_3021 ( .C (CLK), .D (signal_4432), .Q (signal_4433) ) ;
    buf_clk cell_3023 ( .C (CLK), .D (signal_4434), .Q (signal_4435) ) ;
    buf_clk cell_3025 ( .C (CLK), .D (signal_4436), .Q (signal_4437) ) ;
    buf_clk cell_3027 ( .C (CLK), .D (signal_4438), .Q (signal_4439) ) ;
    buf_clk cell_3029 ( .C (CLK), .D (signal_4440), .Q (signal_4441) ) ;
    buf_clk cell_3031 ( .C (CLK), .D (signal_4442), .Q (signal_4443) ) ;
    buf_clk cell_3033 ( .C (CLK), .D (signal_4444), .Q (signal_4445) ) ;
    buf_clk cell_3035 ( .C (CLK), .D (signal_4446), .Q (signal_4447) ) ;
    buf_clk cell_3037 ( .C (CLK), .D (signal_4448), .Q (signal_4449) ) ;
    buf_clk cell_3039 ( .C (CLK), .D (signal_4450), .Q (signal_4451) ) ;
    buf_clk cell_3041 ( .C (CLK), .D (signal_4452), .Q (signal_4453) ) ;
    buf_clk cell_3043 ( .C (CLK), .D (signal_4454), .Q (signal_4455) ) ;
    buf_clk cell_3045 ( .C (CLK), .D (signal_4456), .Q (signal_4457) ) ;
    buf_clk cell_3047 ( .C (CLK), .D (signal_4458), .Q (signal_4459) ) ;
    buf_clk cell_3049 ( .C (CLK), .D (signal_4460), .Q (signal_4461) ) ;
    buf_clk cell_3051 ( .C (CLK), .D (signal_4462), .Q (signal_4463) ) ;
    buf_clk cell_3053 ( .C (CLK), .D (signal_4464), .Q (signal_4465) ) ;
    buf_clk cell_3055 ( .C (CLK), .D (signal_4466), .Q (signal_4467) ) ;
    buf_clk cell_3057 ( .C (CLK), .D (signal_4468), .Q (signal_4469) ) ;
    buf_clk cell_3059 ( .C (CLK), .D (signal_4470), .Q (signal_4471) ) ;
    buf_clk cell_3061 ( .C (CLK), .D (signal_4472), .Q (signal_4473) ) ;
    buf_clk cell_3063 ( .C (CLK), .D (signal_4474), .Q (signal_4475) ) ;
    buf_clk cell_3065 ( .C (CLK), .D (signal_4476), .Q (signal_4477) ) ;
    buf_clk cell_3067 ( .C (CLK), .D (signal_4478), .Q (signal_4479) ) ;
    buf_clk cell_3071 ( .C (CLK), .D (signal_4482), .Q (signal_4483) ) ;
    buf_clk cell_3075 ( .C (CLK), .D (signal_4486), .Q (signal_4487) ) ;
    buf_clk cell_3077 ( .C (CLK), .D (signal_4488), .Q (signal_4489) ) ;
    buf_clk cell_3079 ( .C (CLK), .D (signal_4490), .Q (signal_4491) ) ;
    buf_clk cell_3083 ( .C (CLK), .D (signal_4494), .Q (signal_4495) ) ;
    buf_clk cell_3087 ( .C (CLK), .D (signal_4498), .Q (signal_4499) ) ;
    buf_clk cell_3089 ( .C (CLK), .D (signal_4500), .Q (signal_4501) ) ;
    buf_clk cell_3091 ( .C (CLK), .D (signal_4502), .Q (signal_4503) ) ;
    buf_clk cell_3095 ( .C (CLK), .D (signal_4506), .Q (signal_4507) ) ;
    buf_clk cell_3099 ( .C (CLK), .D (signal_4510), .Q (signal_4511) ) ;
    buf_clk cell_3101 ( .C (CLK), .D (signal_4512), .Q (signal_4513) ) ;
    buf_clk cell_3103 ( .C (CLK), .D (signal_4514), .Q (signal_4515) ) ;
    buf_clk cell_3107 ( .C (CLK), .D (signal_4518), .Q (signal_4519) ) ;
    buf_clk cell_3111 ( .C (CLK), .D (signal_4522), .Q (signal_4523) ) ;
    buf_clk cell_3113 ( .C (CLK), .D (signal_4524), .Q (signal_4525) ) ;
    buf_clk cell_3115 ( .C (CLK), .D (signal_4526), .Q (signal_4527) ) ;
    buf_clk cell_3119 ( .C (CLK), .D (signal_4530), .Q (signal_4531) ) ;
    buf_clk cell_3123 ( .C (CLK), .D (signal_4534), .Q (signal_4535) ) ;
    buf_clk cell_3125 ( .C (CLK), .D (signal_4536), .Q (signal_4537) ) ;
    buf_clk cell_3127 ( .C (CLK), .D (signal_4538), .Q (signal_4539) ) ;
    buf_clk cell_3131 ( .C (CLK), .D (signal_4542), .Q (signal_4543) ) ;
    buf_clk cell_3135 ( .C (CLK), .D (signal_4546), .Q (signal_4547) ) ;
    buf_clk cell_3137 ( .C (CLK), .D (signal_4548), .Q (signal_4549) ) ;
    buf_clk cell_3139 ( .C (CLK), .D (signal_4550), .Q (signal_4551) ) ;
    buf_clk cell_3143 ( .C (CLK), .D (signal_4554), .Q (signal_4555) ) ;
    buf_clk cell_3147 ( .C (CLK), .D (signal_4558), .Q (signal_4559) ) ;
    buf_clk cell_3149 ( .C (CLK), .D (signal_4560), .Q (signal_4561) ) ;
    buf_clk cell_3151 ( .C (CLK), .D (signal_4562), .Q (signal_4563) ) ;
    buf_clk cell_3155 ( .C (CLK), .D (signal_4566), .Q (signal_4567) ) ;
    buf_clk cell_3159 ( .C (CLK), .D (signal_4570), .Q (signal_4571) ) ;
    buf_clk cell_3161 ( .C (CLK), .D (signal_4572), .Q (signal_4573) ) ;
    buf_clk cell_3163 ( .C (CLK), .D (signal_4574), .Q (signal_4575) ) ;
    buf_clk cell_3167 ( .C (CLK), .D (signal_4578), .Q (signal_4579) ) ;
    buf_clk cell_3171 ( .C (CLK), .D (signal_4582), .Q (signal_4583) ) ;
    buf_clk cell_3173 ( .C (CLK), .D (signal_4584), .Q (signal_4585) ) ;
    buf_clk cell_3175 ( .C (CLK), .D (signal_4586), .Q (signal_4587) ) ;
    buf_clk cell_3179 ( .C (CLK), .D (signal_4590), .Q (signal_4591) ) ;
    buf_clk cell_3183 ( .C (CLK), .D (signal_4594), .Q (signal_4595) ) ;
    buf_clk cell_3185 ( .C (CLK), .D (signal_4596), .Q (signal_4597) ) ;
    buf_clk cell_3187 ( .C (CLK), .D (signal_4598), .Q (signal_4599) ) ;
    buf_clk cell_3191 ( .C (CLK), .D (signal_4602), .Q (signal_4603) ) ;
    buf_clk cell_3195 ( .C (CLK), .D (signal_4606), .Q (signal_4607) ) ;
    buf_clk cell_3197 ( .C (CLK), .D (signal_4608), .Q (signal_4609) ) ;
    buf_clk cell_3199 ( .C (CLK), .D (signal_4610), .Q (signal_4611) ) ;
    buf_clk cell_3203 ( .C (CLK), .D (signal_4614), .Q (signal_4615) ) ;
    buf_clk cell_3207 ( .C (CLK), .D (signal_4618), .Q (signal_4619) ) ;
    buf_clk cell_3209 ( .C (CLK), .D (signal_4620), .Q (signal_4621) ) ;
    buf_clk cell_3211 ( .C (CLK), .D (signal_4622), .Q (signal_4623) ) ;
    buf_clk cell_3215 ( .C (CLK), .D (signal_4626), .Q (signal_4627) ) ;
    buf_clk cell_3219 ( .C (CLK), .D (signal_4630), .Q (signal_4631) ) ;
    buf_clk cell_3221 ( .C (CLK), .D (signal_4632), .Q (signal_4633) ) ;
    buf_clk cell_3223 ( .C (CLK), .D (signal_4634), .Q (signal_4635) ) ;
    buf_clk cell_3227 ( .C (CLK), .D (signal_4638), .Q (signal_4639) ) ;
    buf_clk cell_3231 ( .C (CLK), .D (signal_4642), .Q (signal_4643) ) ;
    buf_clk cell_3233 ( .C (CLK), .D (signal_4644), .Q (signal_4645) ) ;
    buf_clk cell_3235 ( .C (CLK), .D (signal_4646), .Q (signal_4647) ) ;
    buf_clk cell_3239 ( .C (CLK), .D (signal_4650), .Q (signal_4651) ) ;
    buf_clk cell_3243 ( .C (CLK), .D (signal_4654), .Q (signal_4655) ) ;
    buf_clk cell_3245 ( .C (CLK), .D (signal_4656), .Q (signal_4657) ) ;
    buf_clk cell_3247 ( .C (CLK), .D (signal_4658), .Q (signal_4659) ) ;
    buf_clk cell_3251 ( .C (CLK), .D (signal_4662), .Q (signal_4663) ) ;
    buf_clk cell_3255 ( .C (CLK), .D (signal_4666), .Q (signal_4667) ) ;
    buf_clk cell_3257 ( .C (CLK), .D (signal_4668), .Q (signal_4669) ) ;
    buf_clk cell_3259 ( .C (CLK), .D (signal_4670), .Q (signal_4671) ) ;
    buf_clk cell_3261 ( .C (CLK), .D (signal_4672), .Q (signal_4673) ) ;
    buf_clk cell_3263 ( .C (CLK), .D (signal_4674), .Q (signal_4675) ) ;
    buf_clk cell_3265 ( .C (CLK), .D (signal_4676), .Q (signal_4677) ) ;
    buf_clk cell_3267 ( .C (CLK), .D (signal_4678), .Q (signal_4679) ) ;
    buf_clk cell_3269 ( .C (CLK), .D (signal_4680), .Q (signal_4681) ) ;
    buf_clk cell_3271 ( .C (CLK), .D (signal_4682), .Q (signal_4683) ) ;
    buf_clk cell_3273 ( .C (CLK), .D (signal_4684), .Q (signal_4685) ) ;
    buf_clk cell_3275 ( .C (CLK), .D (signal_4686), .Q (signal_4687) ) ;
    buf_clk cell_3279 ( .C (CLK), .D (signal_4690), .Q (signal_4691) ) ;
    buf_clk cell_3283 ( .C (CLK), .D (signal_4694), .Q (signal_4695) ) ;
    buf_clk cell_3287 ( .C (CLK), .D (signal_4698), .Q (signal_4699) ) ;
    buf_clk cell_3291 ( .C (CLK), .D (signal_4702), .Q (signal_4703) ) ;
    buf_clk cell_3295 ( .C (CLK), .D (signal_4706), .Q (signal_4707) ) ;
    buf_clk cell_3299 ( .C (CLK), .D (signal_4710), .Q (signal_4711) ) ;
    buf_clk cell_3303 ( .C (CLK), .D (signal_4714), .Q (signal_4715) ) ;
    buf_clk cell_3307 ( .C (CLK), .D (signal_4718), .Q (signal_4719) ) ;
    buf_clk cell_3311 ( .C (CLK), .D (signal_4722), .Q (signal_4723) ) ;
    buf_clk cell_3315 ( .C (CLK), .D (signal_4726), .Q (signal_4727) ) ;
    buf_clk cell_3319 ( .C (CLK), .D (signal_4730), .Q (signal_4731) ) ;

    /* register cells */
    DFF_X1 cell_979 ( .CK (CLK), .D (signal_4691), .Q (signal_808), .QN () ) ;
    DFF_X1 cell_981 ( .CK (CLK), .D (signal_4695), .Q (signal_307), .QN () ) ;
    DFF_X1 cell_983 ( .CK (CLK), .D (signal_4699), .Q (signal_304), .QN () ) ;
    DFF_X1 cell_985 ( .CK (CLK), .D (signal_4703), .Q (signal_288), .QN () ) ;
    DFF_X1 cell_987 ( .CK (CLK), .D (signal_4707), .Q (signal_879), .QN () ) ;
    DFF_X1 cell_989 ( .CK (CLK), .D (signal_4711), .Q (signal_878), .QN () ) ;
    DFF_X1 cell_991 ( .CK (CLK), .D (signal_4715), .Q (signal_877), .QN () ) ;
    DFF_X1 cell_993 ( .CK (CLK), .D (signal_4719), .Q (signal_876), .QN () ) ;
    DFF_X1 cell_995 ( .CK (CLK), .D (signal_4723), .Q (signal_875), .QN () ) ;
    DFF_X1 cell_997 ( .CK (CLK), .D (signal_4727), .Q (signal_874), .QN () ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_999 ( .clk (CLK), .D ({signal_2561, signal_1199}), .Q ({OUT_ciphertext_s1[0], OUT_ciphertext_s0[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1001 ( .clk (CLK), .D ({signal_2679, signal_1198}), .Q ({OUT_ciphertext_s1[1], OUT_ciphertext_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1003 ( .clk (CLK), .D ({signal_2587, signal_1197}), .Q ({OUT_ciphertext_s1[2], OUT_ciphertext_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1005 ( .clk (CLK), .D ({signal_2637, signal_1196}), .Q ({OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1007 ( .clk (CLK), .D ({signal_2589, signal_1195}), .Q ({OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1009 ( .clk (CLK), .D ({signal_2681, signal_1194}), .Q ({OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1011 ( .clk (CLK), .D ({signal_2591, signal_1193}), .Q ({OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1013 ( .clk (CLK), .D ({signal_2593, signal_1192}), .Q ({OUT_ciphertext_s1[7], OUT_ciphertext_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1015 ( .clk (CLK), .D ({signal_2595, signal_1191}), .Q ({OUT_ciphertext_s1[8], OUT_ciphertext_s0[8]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1017 ( .clk (CLK), .D ({signal_2639, signal_1190}), .Q ({OUT_ciphertext_s1[9], OUT_ciphertext_s0[9]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1019 ( .clk (CLK), .D ({signal_2597, signal_1189}), .Q ({OUT_ciphertext_s1[10], OUT_ciphertext_s0[10]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1021 ( .clk (CLK), .D ({signal_2599, signal_1188}), .Q ({OUT_ciphertext_s1[11], OUT_ciphertext_s0[11]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1023 ( .clk (CLK), .D ({signal_2601, signal_1187}), .Q ({OUT_ciphertext_s1[12], OUT_ciphertext_s0[12]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1025 ( .clk (CLK), .D ({signal_2641, signal_1186}), .Q ({OUT_ciphertext_s1[13], OUT_ciphertext_s0[13]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1027 ( .clk (CLK), .D ({signal_2603, signal_1185}), .Q ({OUT_ciphertext_s1[14], OUT_ciphertext_s0[14]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1029 ( .clk (CLK), .D ({signal_2643, signal_1184}), .Q ({OUT_ciphertext_s1[15], OUT_ciphertext_s0[15]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1031 ( .clk (CLK), .D ({signal_2728, signal_1183}), .Q ({OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1033 ( .clk (CLK), .D ({signal_2763, signal_1182}), .Q ({OUT_ciphertext_s1[17], OUT_ciphertext_s0[17]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1035 ( .clk (CLK), .D ({signal_2765, signal_1181}), .Q ({OUT_ciphertext_s1[18], OUT_ciphertext_s0[18]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1037 ( .clk (CLK), .D ({signal_2683, signal_1180}), .Q ({OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1039 ( .clk (CLK), .D ({signal_2685, signal_1179}), .Q ({OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1041 ( .clk (CLK), .D ({signal_2730, signal_1178}), .Q ({OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1043 ( .clk (CLK), .D ({signal_2767, signal_1177}), .Q ({OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1045 ( .clk (CLK), .D ({signal_2687, signal_1176}), .Q ({OUT_ciphertext_s1[23], OUT_ciphertext_s0[23]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1047 ( .clk (CLK), .D ({signal_2689, signal_1175}), .Q ({OUT_ciphertext_s1[24], OUT_ciphertext_s0[24]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1049 ( .clk (CLK), .D ({signal_2732, signal_1174}), .Q ({OUT_ciphertext_s1[25], OUT_ciphertext_s0[25]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1051 ( .clk (CLK), .D ({signal_2734, signal_1173}), .Q ({OUT_ciphertext_s1[26], OUT_ciphertext_s0[26]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1053 ( .clk (CLK), .D ({signal_2691, signal_1172}), .Q ({OUT_ciphertext_s1[27], OUT_ciphertext_s0[27]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1055 ( .clk (CLK), .D ({signal_2736, signal_1171}), .Q ({OUT_ciphertext_s1[28], OUT_ciphertext_s0[28]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1057 ( .clk (CLK), .D ({signal_2769, signal_1170}), .Q ({OUT_ciphertext_s1[29], OUT_ciphertext_s0[29]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1059 ( .clk (CLK), .D ({signal_2738, signal_1169}), .Q ({OUT_ciphertext_s1[30], OUT_ciphertext_s0[30]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1061 ( .clk (CLK), .D ({signal_2693, signal_1168}), .Q ({OUT_ciphertext_s1[31], OUT_ciphertext_s0[31]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1063 ( .clk (CLK), .D ({signal_2771, signal_1167}), .Q ({OUT_ciphertext_s1[32], OUT_ciphertext_s0[32]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1065 ( .clk (CLK), .D ({signal_2803, signal_1166}), .Q ({OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1067 ( .clk (CLK), .D ({signal_2773, signal_1165}), .Q ({OUT_ciphertext_s1[34], OUT_ciphertext_s0[34]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1069 ( .clk (CLK), .D ({signal_2823, signal_1164}), .Q ({OUT_ciphertext_s1[35], OUT_ciphertext_s0[35]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1071 ( .clk (CLK), .D ({signal_2775, signal_1163}), .Q ({OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1073 ( .clk (CLK), .D ({signal_2777, signal_1162}), .Q ({OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1075 ( .clk (CLK), .D ({signal_2740, signal_1161}), .Q ({OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1077 ( .clk (CLK), .D ({signal_2825, signal_1160}), .Q ({OUT_ciphertext_s1[39], OUT_ciphertext_s0[39]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1079 ( .clk (CLK), .D ({signal_2779, signal_1159}), .Q ({OUT_ciphertext_s1[40], OUT_ciphertext_s0[40]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1081 ( .clk (CLK), .D ({signal_2781, signal_1158}), .Q ({OUT_ciphertext_s1[41], OUT_ciphertext_s0[41]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1083 ( .clk (CLK), .D ({signal_2742, signal_1157}), .Q ({OUT_ciphertext_s1[42], OUT_ciphertext_s0[42]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1085 ( .clk (CLK), .D ({signal_2805, signal_1156}), .Q ({OUT_ciphertext_s1[43], OUT_ciphertext_s0[43]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1087 ( .clk (CLK), .D ({signal_2783, signal_1155}), .Q ({OUT_ciphertext_s1[44], OUT_ciphertext_s0[44]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1089 ( .clk (CLK), .D ({signal_2807, signal_1154}), .Q ({OUT_ciphertext_s1[45], OUT_ciphertext_s0[45]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1091 ( .clk (CLK), .D ({signal_2785, signal_1153}), .Q ({OUT_ciphertext_s1[46], OUT_ciphertext_s0[46]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1093 ( .clk (CLK), .D ({signal_2809, signal_1152}), .Q ({OUT_ciphertext_s1[47], OUT_ciphertext_s0[47]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1095 ( .clk (CLK), .D ({signal_2865, signal_1151}), .Q ({OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1097 ( .clk (CLK), .D ({signal_2873, signal_1150}), .Q ({OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1099 ( .clk (CLK), .D ({signal_2827, signal_1149}), .Q ({OUT_ciphertext_s1[50], OUT_ciphertext_s0[50]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1101 ( .clk (CLK), .D ({signal_2829, signal_1148}), .Q ({OUT_ciphertext_s1[51], OUT_ciphertext_s0[51]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1103 ( .clk (CLK), .D ({signal_2867, signal_1147}), .Q ({OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1105 ( .clk (CLK), .D ({signal_2875, signal_1146}), .Q ({OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1107 ( .clk (CLK), .D ({signal_2811, signal_1145}), .Q ({OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1109 ( .clk (CLK), .D ({signal_2831, signal_1144}), .Q ({OUT_ciphertext_s1[55], OUT_ciphertext_s0[55]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1111 ( .clk (CLK), .D ({signal_2857, signal_1143}), .Q ({OUT_ciphertext_s1[56], OUT_ciphertext_s0[56]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1113 ( .clk (CLK), .D ({signal_2869, signal_1142}), .Q ({OUT_ciphertext_s1[57], OUT_ciphertext_s0[57]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1115 ( .clk (CLK), .D ({signal_2813, signal_1141}), .Q ({OUT_ciphertext_s1[58], OUT_ciphertext_s0[58]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1117 ( .clk (CLK), .D ({signal_2815, signal_1140}), .Q ({OUT_ciphertext_s1[59], OUT_ciphertext_s0[59]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1119 ( .clk (CLK), .D ({signal_2859, signal_1139}), .Q ({OUT_ciphertext_s1[60], OUT_ciphertext_s0[60]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1121 ( .clk (CLK), .D ({signal_2871, signal_1138}), .Q ({OUT_ciphertext_s1[61], OUT_ciphertext_s0[61]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1123 ( .clk (CLK), .D ({signal_2833, signal_1137}), .Q ({OUT_ciphertext_s1[62], OUT_ciphertext_s0[62]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1125 ( .clk (CLK), .D ({signal_2835, signal_1136}), .Q ({OUT_ciphertext_s1[63], OUT_ciphertext_s0[63]}) ) ;
    DFF_X1 cell_1127 ( .CK (CLK), .D (signal_4731), .Q (OUT_done), .QN () ) ;
endmodule
