/* modified netlist. Source: module sbox in file Designs/AESSbox/optBP2/AGEMA/sbox.v */
/* 8 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 9 register stage(s) in total */

module sbox_HPC1_Pipeline_d2 (X_s0, clk, X_s1, X_s2, Fresh, Y_s0, Y_s1, Y_s2);
    input [7:0] X_s0 ;
    input clk ;
    input [7:0] X_s1 ;
    input [7:0] X_s2 ;
    input [169:0] Fresh ;
    output [7:0] Y_s0 ;
    output [7:0] Y_s1 ;
    output [7:0] Y_s2 ;
    wire T1 ;
    wire T2 ;
    wire T3 ;
    wire T4 ;
    wire T5 ;
    wire T6 ;
    wire T7 ;
    wire T8 ;
    wire T9 ;
    wire T10 ;
    wire T11 ;
    wire T12 ;
    wire T13 ;
    wire T14 ;
    wire T15 ;
    wire T16 ;
    wire T17 ;
    wire T18 ;
    wire T19 ;
    wire T20 ;
    wire T21 ;
    wire T22 ;
    wire T23 ;
    wire T24 ;
    wire T25 ;
    wire T26 ;
    wire T27 ;
    wire M1 ;
    wire M2 ;
    wire M3 ;
    wire M4 ;
    wire M5 ;
    wire M6 ;
    wire M7 ;
    wire M8 ;
    wire M9 ;
    wire M10 ;
    wire M11 ;
    wire M12 ;
    wire M13 ;
    wire M14 ;
    wire M15 ;
    wire M16 ;
    wire M17 ;
    wire M18 ;
    wire M19 ;
    wire M20 ;
    wire M21 ;
    wire M22 ;
    wire M23 ;
    wire M24 ;
    wire M25 ;
    wire M26 ;
    wire M27 ;
    wire M28 ;
    wire M29 ;
    wire M30 ;
    wire M31 ;
    wire M32 ;
    wire M33 ;
    wire M34 ;
    wire M35 ;
    wire M36 ;
    wire M37 ;
    wire M38 ;
    wire M39 ;
    wire M40 ;
    wire M41 ;
    wire M42 ;
    wire M43 ;
    wire M44 ;
    wire M45 ;
    wire M46 ;
    wire M47 ;
    wire M48 ;
    wire M49 ;
    wire M50 ;
    wire M51 ;
    wire M52 ;
    wire M53 ;
    wire M54 ;
    wire M55 ;
    wire M56 ;
    wire M57 ;
    wire M58 ;
    wire M59 ;
    wire M60 ;
    wire M61 ;
    wire M62 ;
    wire M63 ;
    wire L0 ;
    wire L1 ;
    wire L2 ;
    wire L3 ;
    wire L4 ;
    wire L5 ;
    wire L6 ;
    wire L7 ;
    wire L8 ;
    wire L9 ;
    wire L10 ;
    wire L11 ;
    wire L12 ;
    wire L13 ;
    wire L14 ;
    wire L15 ;
    wire L16 ;
    wire L17 ;
    wire L18 ;
    wire L19 ;
    wire L20 ;
    wire L21 ;
    wire L22 ;
    wire L23 ;
    wire L24 ;
    wire L25 ;
    wire L26 ;
    wire L27 ;
    wire L28 ;
    wire L29 ;
    wire [7:0] O ;
    wire new_AGEMA_signal_155 ;
    wire new_AGEMA_signal_156 ;
    wire new_AGEMA_signal_159 ;
    wire new_AGEMA_signal_160 ;
    wire new_AGEMA_signal_163 ;
    wire new_AGEMA_signal_164 ;
    wire new_AGEMA_signal_165 ;
    wire new_AGEMA_signal_166 ;
    wire new_AGEMA_signal_169 ;
    wire new_AGEMA_signal_170 ;
    wire new_AGEMA_signal_175 ;
    wire new_AGEMA_signal_176 ;
    wire new_AGEMA_signal_177 ;
    wire new_AGEMA_signal_178 ;
    wire new_AGEMA_signal_179 ;
    wire new_AGEMA_signal_180 ;
    wire new_AGEMA_signal_183 ;
    wire new_AGEMA_signal_184 ;
    wire new_AGEMA_signal_185 ;
    wire new_AGEMA_signal_186 ;
    wire new_AGEMA_signal_187 ;
    wire new_AGEMA_signal_188 ;
    wire new_AGEMA_signal_189 ;
    wire new_AGEMA_signal_190 ;
    wire new_AGEMA_signal_191 ;
    wire new_AGEMA_signal_192 ;
    wire new_AGEMA_signal_193 ;
    wire new_AGEMA_signal_194 ;
    wire new_AGEMA_signal_195 ;
    wire new_AGEMA_signal_196 ;
    wire new_AGEMA_signal_197 ;
    wire new_AGEMA_signal_198 ;
    wire new_AGEMA_signal_199 ;
    wire new_AGEMA_signal_200 ;
    wire new_AGEMA_signal_201 ;
    wire new_AGEMA_signal_202 ;
    wire new_AGEMA_signal_203 ;
    wire new_AGEMA_signal_204 ;
    wire new_AGEMA_signal_205 ;
    wire new_AGEMA_signal_206 ;
    wire new_AGEMA_signal_207 ;
    wire new_AGEMA_signal_208 ;
    wire new_AGEMA_signal_209 ;
    wire new_AGEMA_signal_210 ;
    wire new_AGEMA_signal_211 ;
    wire new_AGEMA_signal_212 ;
    wire new_AGEMA_signal_213 ;
    wire new_AGEMA_signal_214 ;
    wire new_AGEMA_signal_215 ;
    wire new_AGEMA_signal_216 ;
    wire new_AGEMA_signal_217 ;
    wire new_AGEMA_signal_218 ;
    wire new_AGEMA_signal_219 ;
    wire new_AGEMA_signal_220 ;
    wire new_AGEMA_signal_221 ;
    wire new_AGEMA_signal_222 ;
    wire new_AGEMA_signal_223 ;
    wire new_AGEMA_signal_224 ;
    wire new_AGEMA_signal_225 ;
    wire new_AGEMA_signal_226 ;
    wire new_AGEMA_signal_227 ;
    wire new_AGEMA_signal_228 ;
    wire new_AGEMA_signal_229 ;
    wire new_AGEMA_signal_230 ;
    wire new_AGEMA_signal_231 ;
    wire new_AGEMA_signal_232 ;
    wire new_AGEMA_signal_233 ;
    wire new_AGEMA_signal_234 ;
    wire new_AGEMA_signal_235 ;
    wire new_AGEMA_signal_236 ;
    wire new_AGEMA_signal_237 ;
    wire new_AGEMA_signal_238 ;
    wire new_AGEMA_signal_239 ;
    wire new_AGEMA_signal_240 ;
    wire new_AGEMA_signal_241 ;
    wire new_AGEMA_signal_242 ;
    wire new_AGEMA_signal_243 ;
    wire new_AGEMA_signal_244 ;
    wire new_AGEMA_signal_245 ;
    wire new_AGEMA_signal_246 ;
    wire new_AGEMA_signal_247 ;
    wire new_AGEMA_signal_248 ;
    wire new_AGEMA_signal_249 ;
    wire new_AGEMA_signal_250 ;
    wire new_AGEMA_signal_251 ;
    wire new_AGEMA_signal_252 ;
    wire new_AGEMA_signal_253 ;
    wire new_AGEMA_signal_254 ;
    wire new_AGEMA_signal_255 ;
    wire new_AGEMA_signal_256 ;
    wire new_AGEMA_signal_257 ;
    wire new_AGEMA_signal_258 ;
    wire new_AGEMA_signal_259 ;
    wire new_AGEMA_signal_260 ;
    wire new_AGEMA_signal_261 ;
    wire new_AGEMA_signal_262 ;
    wire new_AGEMA_signal_263 ;
    wire new_AGEMA_signal_264 ;
    wire new_AGEMA_signal_265 ;
    wire new_AGEMA_signal_266 ;
    wire new_AGEMA_signal_267 ;
    wire new_AGEMA_signal_268 ;
    wire new_AGEMA_signal_269 ;
    wire new_AGEMA_signal_270 ;
    wire new_AGEMA_signal_271 ;
    wire new_AGEMA_signal_272 ;
    wire new_AGEMA_signal_273 ;
    wire new_AGEMA_signal_274 ;
    wire new_AGEMA_signal_275 ;
    wire new_AGEMA_signal_276 ;
    wire new_AGEMA_signal_277 ;
    wire new_AGEMA_signal_278 ;
    wire new_AGEMA_signal_279 ;
    wire new_AGEMA_signal_280 ;
    wire new_AGEMA_signal_281 ;
    wire new_AGEMA_signal_282 ;
    wire new_AGEMA_signal_283 ;
    wire new_AGEMA_signal_284 ;
    wire new_AGEMA_signal_285 ;
    wire new_AGEMA_signal_286 ;
    wire new_AGEMA_signal_287 ;
    wire new_AGEMA_signal_288 ;
    wire new_AGEMA_signal_289 ;
    wire new_AGEMA_signal_290 ;
    wire new_AGEMA_signal_291 ;
    wire new_AGEMA_signal_292 ;
    wire new_AGEMA_signal_293 ;
    wire new_AGEMA_signal_294 ;
    wire new_AGEMA_signal_295 ;
    wire new_AGEMA_signal_296 ;
    wire new_AGEMA_signal_297 ;
    wire new_AGEMA_signal_298 ;
    wire new_AGEMA_signal_299 ;
    wire new_AGEMA_signal_300 ;
    wire new_AGEMA_signal_301 ;
    wire new_AGEMA_signal_302 ;
    wire new_AGEMA_signal_303 ;
    wire new_AGEMA_signal_304 ;
    wire new_AGEMA_signal_305 ;
    wire new_AGEMA_signal_306 ;
    wire new_AGEMA_signal_307 ;
    wire new_AGEMA_signal_308 ;
    wire new_AGEMA_signal_309 ;
    wire new_AGEMA_signal_310 ;
    wire new_AGEMA_signal_311 ;
    wire new_AGEMA_signal_312 ;
    wire new_AGEMA_signal_313 ;
    wire new_AGEMA_signal_314 ;
    wire new_AGEMA_signal_315 ;
    wire new_AGEMA_signal_316 ;
    wire new_AGEMA_signal_317 ;
    wire new_AGEMA_signal_318 ;
    wire new_AGEMA_signal_319 ;
    wire new_AGEMA_signal_320 ;
    wire new_AGEMA_signal_321 ;
    wire new_AGEMA_signal_322 ;
    wire new_AGEMA_signal_323 ;
    wire new_AGEMA_signal_324 ;
    wire new_AGEMA_signal_325 ;
    wire new_AGEMA_signal_326 ;
    wire new_AGEMA_signal_327 ;
    wire new_AGEMA_signal_328 ;
    wire new_AGEMA_signal_329 ;
    wire new_AGEMA_signal_330 ;
    wire new_AGEMA_signal_331 ;
    wire new_AGEMA_signal_332 ;
    wire new_AGEMA_signal_333 ;
    wire new_AGEMA_signal_334 ;
    wire new_AGEMA_signal_335 ;
    wire new_AGEMA_signal_336 ;
    wire new_AGEMA_signal_337 ;
    wire new_AGEMA_signal_338 ;
    wire new_AGEMA_signal_339 ;
    wire new_AGEMA_signal_340 ;
    wire new_AGEMA_signal_341 ;
    wire new_AGEMA_signal_342 ;
    wire new_AGEMA_signal_343 ;
    wire new_AGEMA_signal_344 ;
    wire new_AGEMA_signal_345 ;
    wire new_AGEMA_signal_346 ;
    wire new_AGEMA_signal_347 ;
    wire new_AGEMA_signal_348 ;
    wire new_AGEMA_signal_349 ;
    wire new_AGEMA_signal_350 ;
    wire new_AGEMA_signal_351 ;
    wire new_AGEMA_signal_352 ;
    wire new_AGEMA_signal_353 ;
    wire new_AGEMA_signal_354 ;
    wire new_AGEMA_signal_355 ;
    wire new_AGEMA_signal_356 ;
    wire new_AGEMA_signal_357 ;
    wire new_AGEMA_signal_358 ;
    wire new_AGEMA_signal_359 ;
    wire new_AGEMA_signal_360 ;
    wire new_AGEMA_signal_361 ;
    wire new_AGEMA_signal_362 ;
    wire new_AGEMA_signal_363 ;
    wire new_AGEMA_signal_364 ;
    wire new_AGEMA_signal_365 ;
    wire new_AGEMA_signal_366 ;
    wire new_AGEMA_signal_367 ;
    wire new_AGEMA_signal_368 ;
    wire new_AGEMA_signal_369 ;
    wire new_AGEMA_signal_370 ;
    wire new_AGEMA_signal_371 ;
    wire new_AGEMA_signal_372 ;
    wire new_AGEMA_signal_373 ;
    wire new_AGEMA_signal_374 ;
    wire new_AGEMA_signal_375 ;
    wire new_AGEMA_signal_376 ;
    wire new_AGEMA_signal_377 ;
    wire new_AGEMA_signal_378 ;
    wire new_AGEMA_signal_379 ;
    wire new_AGEMA_signal_380 ;
    wire new_AGEMA_signal_381 ;
    wire new_AGEMA_signal_382 ;
    wire new_AGEMA_signal_383 ;
    wire new_AGEMA_signal_384 ;
    wire new_AGEMA_signal_385 ;
    wire new_AGEMA_signal_386 ;
    wire new_AGEMA_signal_387 ;
    wire new_AGEMA_signal_388 ;
    wire new_AGEMA_signal_389 ;
    wire new_AGEMA_signal_390 ;
    wire new_AGEMA_signal_391 ;
    wire new_AGEMA_signal_392 ;
    wire new_AGEMA_signal_393 ;
    wire new_AGEMA_signal_394 ;
    wire new_AGEMA_signal_395 ;
    wire new_AGEMA_signal_396 ;
    wire new_AGEMA_signal_397 ;
    wire new_AGEMA_signal_398 ;
    wire new_AGEMA_signal_399 ;
    wire new_AGEMA_signal_400 ;
    wire new_AGEMA_signal_401 ;
    wire new_AGEMA_signal_402 ;
    wire new_AGEMA_signal_403 ;
    wire new_AGEMA_signal_404 ;
    wire new_AGEMA_signal_405 ;
    wire new_AGEMA_signal_406 ;
    wire new_AGEMA_signal_407 ;
    wire new_AGEMA_signal_408 ;
    wire new_AGEMA_signal_409 ;
    wire new_AGEMA_signal_410 ;
    wire new_AGEMA_signal_411 ;
    wire new_AGEMA_signal_412 ;
    wire new_AGEMA_signal_413 ;
    wire new_AGEMA_signal_414 ;
    wire new_AGEMA_signal_415 ;
    wire new_AGEMA_signal_416 ;
    wire new_AGEMA_signal_417 ;
    wire new_AGEMA_signal_418 ;
    wire new_AGEMA_signal_419 ;
    wire new_AGEMA_signal_420 ;
    wire new_AGEMA_signal_421 ;
    wire new_AGEMA_signal_422 ;
    wire new_AGEMA_signal_609 ;
    wire new_AGEMA_signal_610 ;
    wire new_AGEMA_signal_611 ;
    wire new_AGEMA_signal_612 ;
    wire new_AGEMA_signal_613 ;
    wire new_AGEMA_signal_614 ;
    wire new_AGEMA_signal_615 ;
    wire new_AGEMA_signal_616 ;
    wire new_AGEMA_signal_617 ;
    wire new_AGEMA_signal_618 ;
    wire new_AGEMA_signal_619 ;
    wire new_AGEMA_signal_620 ;
    wire new_AGEMA_signal_621 ;
    wire new_AGEMA_signal_622 ;
    wire new_AGEMA_signal_623 ;
    wire new_AGEMA_signal_624 ;
    wire new_AGEMA_signal_625 ;
    wire new_AGEMA_signal_626 ;
    wire new_AGEMA_signal_627 ;
    wire new_AGEMA_signal_628 ;
    wire new_AGEMA_signal_629 ;
    wire new_AGEMA_signal_630 ;
    wire new_AGEMA_signal_631 ;
    wire new_AGEMA_signal_632 ;
    wire new_AGEMA_signal_633 ;
    wire new_AGEMA_signal_634 ;
    wire new_AGEMA_signal_635 ;
    wire new_AGEMA_signal_636 ;
    wire new_AGEMA_signal_637 ;
    wire new_AGEMA_signal_638 ;
    wire new_AGEMA_signal_639 ;
    wire new_AGEMA_signal_640 ;
    wire new_AGEMA_signal_641 ;
    wire new_AGEMA_signal_642 ;
    wire new_AGEMA_signal_643 ;
    wire new_AGEMA_signal_644 ;
    wire new_AGEMA_signal_645 ;
    wire new_AGEMA_signal_646 ;
    wire new_AGEMA_signal_647 ;
    wire new_AGEMA_signal_648 ;
    wire new_AGEMA_signal_649 ;
    wire new_AGEMA_signal_650 ;
    wire new_AGEMA_signal_651 ;
    wire new_AGEMA_signal_652 ;
    wire new_AGEMA_signal_653 ;
    wire new_AGEMA_signal_654 ;
    wire new_AGEMA_signal_655 ;
    wire new_AGEMA_signal_656 ;
    wire new_AGEMA_signal_657 ;
    wire new_AGEMA_signal_658 ;
    wire new_AGEMA_signal_659 ;
    wire new_AGEMA_signal_660 ;
    wire new_AGEMA_signal_661 ;
    wire new_AGEMA_signal_662 ;
    wire new_AGEMA_signal_663 ;
    wire new_AGEMA_signal_664 ;
    wire new_AGEMA_signal_665 ;
    wire new_AGEMA_signal_666 ;
    wire new_AGEMA_signal_667 ;
    wire new_AGEMA_signal_668 ;
    wire new_AGEMA_signal_669 ;
    wire new_AGEMA_signal_670 ;
    wire new_AGEMA_signal_671 ;
    wire new_AGEMA_signal_672 ;
    wire new_AGEMA_signal_673 ;
    wire new_AGEMA_signal_674 ;
    wire new_AGEMA_signal_675 ;
    wire new_AGEMA_signal_676 ;
    wire new_AGEMA_signal_677 ;
    wire new_AGEMA_signal_678 ;
    wire new_AGEMA_signal_679 ;
    wire new_AGEMA_signal_680 ;
    wire new_AGEMA_signal_681 ;
    wire new_AGEMA_signal_682 ;
    wire new_AGEMA_signal_683 ;
    wire new_AGEMA_signal_684 ;
    wire new_AGEMA_signal_685 ;
    wire new_AGEMA_signal_686 ;
    wire new_AGEMA_signal_687 ;
    wire new_AGEMA_signal_688 ;
    wire new_AGEMA_signal_689 ;
    wire new_AGEMA_signal_690 ;
    wire new_AGEMA_signal_691 ;
    wire new_AGEMA_signal_692 ;
    wire new_AGEMA_signal_693 ;
    wire new_AGEMA_signal_694 ;
    wire new_AGEMA_signal_695 ;
    wire new_AGEMA_signal_696 ;
    wire new_AGEMA_signal_697 ;
    wire new_AGEMA_signal_698 ;
    wire new_AGEMA_signal_699 ;
    wire new_AGEMA_signal_700 ;
    wire new_AGEMA_signal_701 ;
    wire new_AGEMA_signal_702 ;
    wire new_AGEMA_signal_703 ;
    wire new_AGEMA_signal_704 ;
    wire new_AGEMA_signal_705 ;
    wire new_AGEMA_signal_706 ;
    wire new_AGEMA_signal_707 ;
    wire new_AGEMA_signal_708 ;
    wire new_AGEMA_signal_709 ;
    wire new_AGEMA_signal_710 ;
    wire new_AGEMA_signal_711 ;
    wire new_AGEMA_signal_712 ;
    wire new_AGEMA_signal_713 ;
    wire new_AGEMA_signal_714 ;
    wire new_AGEMA_signal_715 ;
    wire new_AGEMA_signal_716 ;
    wire new_AGEMA_signal_717 ;
    wire new_AGEMA_signal_718 ;
    wire new_AGEMA_signal_719 ;
    wire new_AGEMA_signal_720 ;
    wire new_AGEMA_signal_721 ;
    wire new_AGEMA_signal_722 ;
    wire new_AGEMA_signal_723 ;
    wire new_AGEMA_signal_724 ;
    wire new_AGEMA_signal_725 ;
    wire new_AGEMA_signal_726 ;
    wire new_AGEMA_signal_727 ;
    wire new_AGEMA_signal_728 ;
    wire new_AGEMA_signal_729 ;
    wire new_AGEMA_signal_730 ;
    wire new_AGEMA_signal_731 ;
    wire new_AGEMA_signal_732 ;
    wire new_AGEMA_signal_733 ;
    wire new_AGEMA_signal_734 ;
    wire new_AGEMA_signal_735 ;
    wire new_AGEMA_signal_736 ;
    wire new_AGEMA_signal_737 ;
    wire new_AGEMA_signal_738 ;
    wire new_AGEMA_signal_739 ;
    wire new_AGEMA_signal_740 ;
    wire new_AGEMA_signal_741 ;
    wire new_AGEMA_signal_742 ;
    wire new_AGEMA_signal_743 ;
    wire new_AGEMA_signal_744 ;
    wire new_AGEMA_signal_745 ;
    wire new_AGEMA_signal_746 ;
    wire new_AGEMA_signal_747 ;
    wire new_AGEMA_signal_748 ;
    wire new_AGEMA_signal_749 ;
    wire new_AGEMA_signal_750 ;
    wire new_AGEMA_signal_751 ;
    wire new_AGEMA_signal_752 ;
    wire new_AGEMA_signal_753 ;
    wire new_AGEMA_signal_754 ;
    wire new_AGEMA_signal_755 ;
    wire new_AGEMA_signal_756 ;
    wire new_AGEMA_signal_757 ;
    wire new_AGEMA_signal_758 ;
    wire new_AGEMA_signal_759 ;
    wire new_AGEMA_signal_760 ;
    wire new_AGEMA_signal_761 ;
    wire new_AGEMA_signal_762 ;
    wire new_AGEMA_signal_763 ;
    wire new_AGEMA_signal_764 ;
    wire new_AGEMA_signal_765 ;
    wire new_AGEMA_signal_766 ;
    wire new_AGEMA_signal_767 ;
    wire new_AGEMA_signal_768 ;
    wire new_AGEMA_signal_769 ;
    wire new_AGEMA_signal_770 ;
    wire new_AGEMA_signal_771 ;
    wire new_AGEMA_signal_772 ;
    wire new_AGEMA_signal_773 ;
    wire new_AGEMA_signal_774 ;
    wire new_AGEMA_signal_775 ;
    wire new_AGEMA_signal_776 ;
    wire new_AGEMA_signal_777 ;
    wire new_AGEMA_signal_778 ;
    wire new_AGEMA_signal_779 ;
    wire new_AGEMA_signal_780 ;
    wire new_AGEMA_signal_781 ;
    wire new_AGEMA_signal_782 ;
    wire new_AGEMA_signal_783 ;
    wire new_AGEMA_signal_784 ;
    wire new_AGEMA_signal_785 ;
    wire new_AGEMA_signal_786 ;
    wire new_AGEMA_signal_787 ;
    wire new_AGEMA_signal_788 ;
    wire new_AGEMA_signal_789 ;
    wire new_AGEMA_signal_790 ;
    wire new_AGEMA_signal_791 ;
    wire new_AGEMA_signal_792 ;
    wire new_AGEMA_signal_793 ;
    wire new_AGEMA_signal_794 ;
    wire new_AGEMA_signal_795 ;
    wire new_AGEMA_signal_796 ;
    wire new_AGEMA_signal_797 ;
    wire new_AGEMA_signal_798 ;
    wire new_AGEMA_signal_799 ;
    wire new_AGEMA_signal_800 ;
    wire new_AGEMA_signal_801 ;
    wire new_AGEMA_signal_802 ;
    wire new_AGEMA_signal_803 ;
    wire new_AGEMA_signal_804 ;
    wire new_AGEMA_signal_805 ;
    wire new_AGEMA_signal_806 ;
    wire new_AGEMA_signal_807 ;
    wire new_AGEMA_signal_808 ;
    wire new_AGEMA_signal_809 ;
    wire new_AGEMA_signal_810 ;
    wire new_AGEMA_signal_811 ;
    wire new_AGEMA_signal_812 ;
    wire new_AGEMA_signal_813 ;
    wire new_AGEMA_signal_814 ;
    wire new_AGEMA_signal_815 ;
    wire new_AGEMA_signal_816 ;
    wire new_AGEMA_signal_817 ;
    wire new_AGEMA_signal_818 ;
    wire new_AGEMA_signal_819 ;
    wire new_AGEMA_signal_820 ;
    wire new_AGEMA_signal_821 ;
    wire new_AGEMA_signal_822 ;
    wire new_AGEMA_signal_823 ;
    wire new_AGEMA_signal_824 ;
    wire new_AGEMA_signal_825 ;
    wire new_AGEMA_signal_826 ;
    wire new_AGEMA_signal_827 ;
    wire new_AGEMA_signal_828 ;
    wire new_AGEMA_signal_829 ;
    wire new_AGEMA_signal_830 ;
    wire new_AGEMA_signal_831 ;
    wire new_AGEMA_signal_832 ;
    wire new_AGEMA_signal_833 ;
    wire new_AGEMA_signal_834 ;
    wire new_AGEMA_signal_835 ;
    wire new_AGEMA_signal_836 ;
    wire new_AGEMA_signal_837 ;
    wire new_AGEMA_signal_838 ;
    wire new_AGEMA_signal_839 ;
    wire new_AGEMA_signal_840 ;
    wire new_AGEMA_signal_841 ;
    wire new_AGEMA_signal_842 ;
    wire new_AGEMA_signal_843 ;
    wire new_AGEMA_signal_844 ;
    wire new_AGEMA_signal_845 ;
    wire new_AGEMA_signal_846 ;
    wire new_AGEMA_signal_847 ;
    wire new_AGEMA_signal_848 ;
    wire new_AGEMA_signal_849 ;
    wire new_AGEMA_signal_850 ;
    wire new_AGEMA_signal_851 ;
    wire new_AGEMA_signal_852 ;
    wire new_AGEMA_signal_853 ;
    wire new_AGEMA_signal_854 ;
    wire new_AGEMA_signal_855 ;
    wire new_AGEMA_signal_856 ;
    wire new_AGEMA_signal_857 ;
    wire new_AGEMA_signal_858 ;
    wire new_AGEMA_signal_859 ;
    wire new_AGEMA_signal_860 ;
    wire new_AGEMA_signal_861 ;
    wire new_AGEMA_signal_862 ;
    wire new_AGEMA_signal_863 ;
    wire new_AGEMA_signal_864 ;
    wire new_AGEMA_signal_865 ;
    wire new_AGEMA_signal_866 ;
    wire new_AGEMA_signal_867 ;
    wire new_AGEMA_signal_868 ;
    wire new_AGEMA_signal_869 ;
    wire new_AGEMA_signal_870 ;
    wire new_AGEMA_signal_871 ;
    wire new_AGEMA_signal_872 ;
    wire new_AGEMA_signal_873 ;
    wire new_AGEMA_signal_874 ;
    wire new_AGEMA_signal_875 ;
    wire new_AGEMA_signal_876 ;
    wire new_AGEMA_signal_877 ;
    wire new_AGEMA_signal_878 ;
    wire new_AGEMA_signal_879 ;
    wire new_AGEMA_signal_880 ;
    wire new_AGEMA_signal_881 ;
    wire new_AGEMA_signal_882 ;
    wire new_AGEMA_signal_883 ;
    wire new_AGEMA_signal_884 ;
    wire new_AGEMA_signal_885 ;
    wire new_AGEMA_signal_886 ;
    wire new_AGEMA_signal_887 ;
    wire new_AGEMA_signal_888 ;
    wire new_AGEMA_signal_889 ;
    wire new_AGEMA_signal_890 ;
    wire new_AGEMA_signal_891 ;
    wire new_AGEMA_signal_892 ;
    wire new_AGEMA_signal_893 ;
    wire new_AGEMA_signal_894 ;
    wire new_AGEMA_signal_895 ;
    wire new_AGEMA_signal_896 ;
    wire new_AGEMA_signal_897 ;
    wire new_AGEMA_signal_898 ;
    wire new_AGEMA_signal_899 ;
    wire new_AGEMA_signal_900 ;
    wire new_AGEMA_signal_901 ;
    wire new_AGEMA_signal_902 ;
    wire new_AGEMA_signal_903 ;
    wire new_AGEMA_signal_904 ;
    wire new_AGEMA_signal_905 ;
    wire new_AGEMA_signal_906 ;
    wire new_AGEMA_signal_907 ;
    wire new_AGEMA_signal_908 ;
    wire new_AGEMA_signal_909 ;
    wire new_AGEMA_signal_910 ;
    wire new_AGEMA_signal_911 ;
    wire new_AGEMA_signal_912 ;
    wire new_AGEMA_signal_913 ;
    wire new_AGEMA_signal_914 ;
    wire new_AGEMA_signal_915 ;
    wire new_AGEMA_signal_916 ;
    wire new_AGEMA_signal_917 ;
    wire new_AGEMA_signal_918 ;
    wire new_AGEMA_signal_919 ;
    wire new_AGEMA_signal_920 ;
    wire new_AGEMA_signal_921 ;
    wire new_AGEMA_signal_922 ;
    wire new_AGEMA_signal_923 ;
    wire new_AGEMA_signal_924 ;
    wire new_AGEMA_signal_925 ;
    wire new_AGEMA_signal_926 ;
    wire new_AGEMA_signal_927 ;
    wire new_AGEMA_signal_928 ;
    wire new_AGEMA_signal_929 ;
    wire new_AGEMA_signal_930 ;
    wire new_AGEMA_signal_931 ;
    wire new_AGEMA_signal_932 ;
    wire new_AGEMA_signal_933 ;
    wire new_AGEMA_signal_934 ;
    wire new_AGEMA_signal_935 ;
    wire new_AGEMA_signal_936 ;
    wire new_AGEMA_signal_937 ;
    wire new_AGEMA_signal_938 ;
    wire new_AGEMA_signal_939 ;
    wire new_AGEMA_signal_940 ;
    wire new_AGEMA_signal_941 ;
    wire new_AGEMA_signal_942 ;
    wire new_AGEMA_signal_943 ;
    wire new_AGEMA_signal_944 ;
    wire new_AGEMA_signal_945 ;
    wire new_AGEMA_signal_946 ;
    wire new_AGEMA_signal_947 ;
    wire new_AGEMA_signal_948 ;
    wire new_AGEMA_signal_949 ;
    wire new_AGEMA_signal_950 ;
    wire new_AGEMA_signal_951 ;
    wire new_AGEMA_signal_952 ;
    wire new_AGEMA_signal_953 ;
    wire new_AGEMA_signal_954 ;
    wire new_AGEMA_signal_955 ;
    wire new_AGEMA_signal_956 ;
    wire new_AGEMA_signal_957 ;
    wire new_AGEMA_signal_958 ;
    wire new_AGEMA_signal_959 ;
    wire new_AGEMA_signal_960 ;
    wire new_AGEMA_signal_961 ;
    wire new_AGEMA_signal_962 ;
    wire new_AGEMA_signal_963 ;
    wire new_AGEMA_signal_964 ;
    wire new_AGEMA_signal_965 ;
    wire new_AGEMA_signal_966 ;
    wire new_AGEMA_signal_967 ;
    wire new_AGEMA_signal_968 ;
    wire new_AGEMA_signal_969 ;
    wire new_AGEMA_signal_970 ;
    wire new_AGEMA_signal_971 ;
    wire new_AGEMA_signal_972 ;
    wire new_AGEMA_signal_973 ;
    wire new_AGEMA_signal_974 ;
    wire new_AGEMA_signal_975 ;
    wire new_AGEMA_signal_976 ;
    wire new_AGEMA_signal_977 ;
    wire new_AGEMA_signal_978 ;
    wire new_AGEMA_signal_979 ;
    wire new_AGEMA_signal_980 ;
    wire new_AGEMA_signal_981 ;
    wire new_AGEMA_signal_982 ;
    wire new_AGEMA_signal_983 ;
    wire new_AGEMA_signal_984 ;
    wire new_AGEMA_signal_985 ;
    wire new_AGEMA_signal_986 ;
    wire new_AGEMA_signal_987 ;
    wire new_AGEMA_signal_988 ;
    wire new_AGEMA_signal_989 ;
    wire new_AGEMA_signal_990 ;
    wire new_AGEMA_signal_991 ;
    wire new_AGEMA_signal_992 ;
    wire new_AGEMA_signal_993 ;
    wire new_AGEMA_signal_994 ;
    wire new_AGEMA_signal_995 ;
    wire new_AGEMA_signal_996 ;
    wire new_AGEMA_signal_997 ;
    wire new_AGEMA_signal_998 ;
    wire new_AGEMA_signal_999 ;
    wire new_AGEMA_signal_1000 ;
    wire new_AGEMA_signal_1001 ;
    wire new_AGEMA_signal_1002 ;
    wire new_AGEMA_signal_1003 ;
    wire new_AGEMA_signal_1004 ;

    /* cells in depth 0 */
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_T1_U1 ( .a ({X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s2[4], X_s1[4], X_s0[4]}), .c ({new_AGEMA_signal_156, new_AGEMA_signal_155, T1}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_T2_U1 ( .a ({X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s2[2], X_s1[2], X_s0[2]}), .c ({new_AGEMA_signal_160, new_AGEMA_signal_159, T2}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_T3_U1 ( .a ({X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s2[1], X_s1[1], X_s0[1]}), .c ({new_AGEMA_signal_164, new_AGEMA_signal_163, T3}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_T4_U1 ( .a ({X_s2[4], X_s1[4], X_s0[4]}), .b ({X_s2[2], X_s1[2], X_s0[2]}), .c ({new_AGEMA_signal_166, new_AGEMA_signal_165, T4}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_T5_U1 ( .a ({X_s2[3], X_s1[3], X_s0[3]}), .b ({X_s2[1], X_s1[1], X_s0[1]}), .c ({new_AGEMA_signal_170, new_AGEMA_signal_169, T5}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_T6_U1 ( .a ({new_AGEMA_signal_156, new_AGEMA_signal_155, T1}), .b ({new_AGEMA_signal_170, new_AGEMA_signal_169, T5}), .c ({new_AGEMA_signal_188, new_AGEMA_signal_187, T6}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_T7_U1 ( .a ({X_s2[6], X_s1[6], X_s0[6]}), .b ({X_s2[5], X_s1[5], X_s0[5]}), .c ({new_AGEMA_signal_176, new_AGEMA_signal_175, T7}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_T8_U1 ( .a ({X_s2[0], X_s1[0], X_s0[0]}), .b ({new_AGEMA_signal_188, new_AGEMA_signal_187, T6}), .c ({new_AGEMA_signal_204, new_AGEMA_signal_203, T8}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_T9_U1 ( .a ({X_s2[0], X_s1[0], X_s0[0]}), .b ({new_AGEMA_signal_176, new_AGEMA_signal_175, T7}), .c ({new_AGEMA_signal_190, new_AGEMA_signal_189, T9}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_T10_U1 ( .a ({new_AGEMA_signal_188, new_AGEMA_signal_187, T6}), .b ({new_AGEMA_signal_176, new_AGEMA_signal_175, T7}), .c ({new_AGEMA_signal_206, new_AGEMA_signal_205, T10}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_T11_U1 ( .a ({X_s2[6], X_s1[6], X_s0[6]}), .b ({X_s2[2], X_s1[2], X_s0[2]}), .c ({new_AGEMA_signal_178, new_AGEMA_signal_177, T11}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_T12_U1 ( .a ({X_s2[5], X_s1[5], X_s0[5]}), .b ({X_s2[2], X_s1[2], X_s0[2]}), .c ({new_AGEMA_signal_180, new_AGEMA_signal_179, T12}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_T13_U1 ( .a ({new_AGEMA_signal_164, new_AGEMA_signal_163, T3}), .b ({new_AGEMA_signal_166, new_AGEMA_signal_165, T4}), .c ({new_AGEMA_signal_192, new_AGEMA_signal_191, T13}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_T14_U1 ( .a ({new_AGEMA_signal_188, new_AGEMA_signal_187, T6}), .b ({new_AGEMA_signal_178, new_AGEMA_signal_177, T11}), .c ({new_AGEMA_signal_208, new_AGEMA_signal_207, T14}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_T15_U1 ( .a ({new_AGEMA_signal_170, new_AGEMA_signal_169, T5}), .b ({new_AGEMA_signal_178, new_AGEMA_signal_177, T11}), .c ({new_AGEMA_signal_194, new_AGEMA_signal_193, T15}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_T16_U1 ( .a ({new_AGEMA_signal_170, new_AGEMA_signal_169, T5}), .b ({new_AGEMA_signal_180, new_AGEMA_signal_179, T12}), .c ({new_AGEMA_signal_196, new_AGEMA_signal_195, T16}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_T17_U1 ( .a ({new_AGEMA_signal_190, new_AGEMA_signal_189, T9}), .b ({new_AGEMA_signal_196, new_AGEMA_signal_195, T16}), .c ({new_AGEMA_signal_210, new_AGEMA_signal_209, T17}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_T18_U1 ( .a ({X_s2[4], X_s1[4], X_s0[4]}), .b ({X_s2[0], X_s1[0], X_s0[0]}), .c ({new_AGEMA_signal_184, new_AGEMA_signal_183, T18}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_T19_U1 ( .a ({new_AGEMA_signal_176, new_AGEMA_signal_175, T7}), .b ({new_AGEMA_signal_184, new_AGEMA_signal_183, T18}), .c ({new_AGEMA_signal_198, new_AGEMA_signal_197, T19}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_T20_U1 ( .a ({new_AGEMA_signal_156, new_AGEMA_signal_155, T1}), .b ({new_AGEMA_signal_198, new_AGEMA_signal_197, T19}), .c ({new_AGEMA_signal_212, new_AGEMA_signal_211, T20}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_T21_U1 ( .a ({X_s2[1], X_s1[1], X_s0[1]}), .b ({X_s2[0], X_s1[0], X_s0[0]}), .c ({new_AGEMA_signal_186, new_AGEMA_signal_185, T21}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_T22_U1 ( .a ({new_AGEMA_signal_176, new_AGEMA_signal_175, T7}), .b ({new_AGEMA_signal_186, new_AGEMA_signal_185, T21}), .c ({new_AGEMA_signal_200, new_AGEMA_signal_199, T22}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_T23_U1 ( .a ({new_AGEMA_signal_160, new_AGEMA_signal_159, T2}), .b ({new_AGEMA_signal_200, new_AGEMA_signal_199, T22}), .c ({new_AGEMA_signal_214, new_AGEMA_signal_213, T23}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_T24_U1 ( .a ({new_AGEMA_signal_160, new_AGEMA_signal_159, T2}), .b ({new_AGEMA_signal_206, new_AGEMA_signal_205, T10}), .c ({new_AGEMA_signal_230, new_AGEMA_signal_229, T24}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_T25_U1 ( .a ({new_AGEMA_signal_212, new_AGEMA_signal_211, T20}), .b ({new_AGEMA_signal_210, new_AGEMA_signal_209, T17}), .c ({new_AGEMA_signal_232, new_AGEMA_signal_231, T25}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_T26_U1 ( .a ({new_AGEMA_signal_164, new_AGEMA_signal_163, T3}), .b ({new_AGEMA_signal_196, new_AGEMA_signal_195, T16}), .c ({new_AGEMA_signal_216, new_AGEMA_signal_215, T26}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_T27_U1 ( .a ({new_AGEMA_signal_156, new_AGEMA_signal_155, T1}), .b ({new_AGEMA_signal_180, new_AGEMA_signal_179, T12}), .c ({new_AGEMA_signal_202, new_AGEMA_signal_201, T27}) ) ;

    /* cells in depth 1 */
    buf_clk new_AGEMA_reg_buffer_136 ( .C (clk), .D (T14), .Q (new_AGEMA_signal_609) ) ;
    buf_clk new_AGEMA_reg_buffer_138 ( .C (clk), .D (new_AGEMA_signal_207), .Q (new_AGEMA_signal_611) ) ;
    buf_clk new_AGEMA_reg_buffer_140 ( .C (clk), .D (new_AGEMA_signal_208), .Q (new_AGEMA_signal_613) ) ;
    buf_clk new_AGEMA_reg_buffer_142 ( .C (clk), .D (T26), .Q (new_AGEMA_signal_615) ) ;
    buf_clk new_AGEMA_reg_buffer_144 ( .C (clk), .D (new_AGEMA_signal_215), .Q (new_AGEMA_signal_617) ) ;
    buf_clk new_AGEMA_reg_buffer_146 ( .C (clk), .D (new_AGEMA_signal_216), .Q (new_AGEMA_signal_619) ) ;
    buf_clk new_AGEMA_reg_buffer_148 ( .C (clk), .D (T24), .Q (new_AGEMA_signal_621) ) ;
    buf_clk new_AGEMA_reg_buffer_150 ( .C (clk), .D (new_AGEMA_signal_229), .Q (new_AGEMA_signal_623) ) ;
    buf_clk new_AGEMA_reg_buffer_152 ( .C (clk), .D (new_AGEMA_signal_230), .Q (new_AGEMA_signal_625) ) ;
    buf_clk new_AGEMA_reg_buffer_154 ( .C (clk), .D (T25), .Q (new_AGEMA_signal_627) ) ;
    buf_clk new_AGEMA_reg_buffer_156 ( .C (clk), .D (new_AGEMA_signal_231), .Q (new_AGEMA_signal_629) ) ;
    buf_clk new_AGEMA_reg_buffer_158 ( .C (clk), .D (new_AGEMA_signal_232), .Q (new_AGEMA_signal_631) ) ;
    buf_clk new_AGEMA_reg_buffer_208 ( .C (clk), .D (T6), .Q (new_AGEMA_signal_681) ) ;
    buf_clk new_AGEMA_reg_buffer_214 ( .C (clk), .D (new_AGEMA_signal_187), .Q (new_AGEMA_signal_687) ) ;
    buf_clk new_AGEMA_reg_buffer_220 ( .C (clk), .D (new_AGEMA_signal_188), .Q (new_AGEMA_signal_693) ) ;
    buf_clk new_AGEMA_reg_buffer_226 ( .C (clk), .D (T8), .Q (new_AGEMA_signal_699) ) ;
    buf_clk new_AGEMA_reg_buffer_232 ( .C (clk), .D (new_AGEMA_signal_203), .Q (new_AGEMA_signal_705) ) ;
    buf_clk new_AGEMA_reg_buffer_238 ( .C (clk), .D (new_AGEMA_signal_204), .Q (new_AGEMA_signal_711) ) ;
    buf_clk new_AGEMA_reg_buffer_244 ( .C (clk), .D (X_s0[0]), .Q (new_AGEMA_signal_717) ) ;
    buf_clk new_AGEMA_reg_buffer_250 ( .C (clk), .D (X_s1[0]), .Q (new_AGEMA_signal_723) ) ;
    buf_clk new_AGEMA_reg_buffer_256 ( .C (clk), .D (X_s2[0]), .Q (new_AGEMA_signal_729) ) ;
    buf_clk new_AGEMA_reg_buffer_262 ( .C (clk), .D (T16), .Q (new_AGEMA_signal_735) ) ;
    buf_clk new_AGEMA_reg_buffer_268 ( .C (clk), .D (new_AGEMA_signal_195), .Q (new_AGEMA_signal_741) ) ;
    buf_clk new_AGEMA_reg_buffer_274 ( .C (clk), .D (new_AGEMA_signal_196), .Q (new_AGEMA_signal_747) ) ;
    buf_clk new_AGEMA_reg_buffer_280 ( .C (clk), .D (T9), .Q (new_AGEMA_signal_753) ) ;
    buf_clk new_AGEMA_reg_buffer_286 ( .C (clk), .D (new_AGEMA_signal_189), .Q (new_AGEMA_signal_759) ) ;
    buf_clk new_AGEMA_reg_buffer_292 ( .C (clk), .D (new_AGEMA_signal_190), .Q (new_AGEMA_signal_765) ) ;
    buf_clk new_AGEMA_reg_buffer_298 ( .C (clk), .D (T17), .Q (new_AGEMA_signal_771) ) ;
    buf_clk new_AGEMA_reg_buffer_304 ( .C (clk), .D (new_AGEMA_signal_209), .Q (new_AGEMA_signal_777) ) ;
    buf_clk new_AGEMA_reg_buffer_310 ( .C (clk), .D (new_AGEMA_signal_210), .Q (new_AGEMA_signal_783) ) ;
    buf_clk new_AGEMA_reg_buffer_316 ( .C (clk), .D (T15), .Q (new_AGEMA_signal_789) ) ;
    buf_clk new_AGEMA_reg_buffer_322 ( .C (clk), .D (new_AGEMA_signal_193), .Q (new_AGEMA_signal_795) ) ;
    buf_clk new_AGEMA_reg_buffer_328 ( .C (clk), .D (new_AGEMA_signal_194), .Q (new_AGEMA_signal_801) ) ;
    buf_clk new_AGEMA_reg_buffer_334 ( .C (clk), .D (T27), .Q (new_AGEMA_signal_807) ) ;
    buf_clk new_AGEMA_reg_buffer_340 ( .C (clk), .D (new_AGEMA_signal_201), .Q (new_AGEMA_signal_813) ) ;
    buf_clk new_AGEMA_reg_buffer_346 ( .C (clk), .D (new_AGEMA_signal_202), .Q (new_AGEMA_signal_819) ) ;
    buf_clk new_AGEMA_reg_buffer_352 ( .C (clk), .D (T10), .Q (new_AGEMA_signal_825) ) ;
    buf_clk new_AGEMA_reg_buffer_358 ( .C (clk), .D (new_AGEMA_signal_205), .Q (new_AGEMA_signal_831) ) ;
    buf_clk new_AGEMA_reg_buffer_364 ( .C (clk), .D (new_AGEMA_signal_206), .Q (new_AGEMA_signal_837) ) ;
    buf_clk new_AGEMA_reg_buffer_370 ( .C (clk), .D (T13), .Q (new_AGEMA_signal_843) ) ;
    buf_clk new_AGEMA_reg_buffer_376 ( .C (clk), .D (new_AGEMA_signal_191), .Q (new_AGEMA_signal_849) ) ;
    buf_clk new_AGEMA_reg_buffer_382 ( .C (clk), .D (new_AGEMA_signal_192), .Q (new_AGEMA_signal_855) ) ;
    buf_clk new_AGEMA_reg_buffer_388 ( .C (clk), .D (T23), .Q (new_AGEMA_signal_861) ) ;
    buf_clk new_AGEMA_reg_buffer_394 ( .C (clk), .D (new_AGEMA_signal_213), .Q (new_AGEMA_signal_867) ) ;
    buf_clk new_AGEMA_reg_buffer_400 ( .C (clk), .D (new_AGEMA_signal_214), .Q (new_AGEMA_signal_873) ) ;
    buf_clk new_AGEMA_reg_buffer_406 ( .C (clk), .D (T19), .Q (new_AGEMA_signal_879) ) ;
    buf_clk new_AGEMA_reg_buffer_412 ( .C (clk), .D (new_AGEMA_signal_197), .Q (new_AGEMA_signal_885) ) ;
    buf_clk new_AGEMA_reg_buffer_418 ( .C (clk), .D (new_AGEMA_signal_198), .Q (new_AGEMA_signal_891) ) ;
    buf_clk new_AGEMA_reg_buffer_424 ( .C (clk), .D (T3), .Q (new_AGEMA_signal_897) ) ;
    buf_clk new_AGEMA_reg_buffer_430 ( .C (clk), .D (new_AGEMA_signal_163), .Q (new_AGEMA_signal_903) ) ;
    buf_clk new_AGEMA_reg_buffer_436 ( .C (clk), .D (new_AGEMA_signal_164), .Q (new_AGEMA_signal_909) ) ;
    buf_clk new_AGEMA_reg_buffer_442 ( .C (clk), .D (T22), .Q (new_AGEMA_signal_915) ) ;
    buf_clk new_AGEMA_reg_buffer_448 ( .C (clk), .D (new_AGEMA_signal_199), .Q (new_AGEMA_signal_921) ) ;
    buf_clk new_AGEMA_reg_buffer_454 ( .C (clk), .D (new_AGEMA_signal_200), .Q (new_AGEMA_signal_927) ) ;
    buf_clk new_AGEMA_reg_buffer_460 ( .C (clk), .D (T20), .Q (new_AGEMA_signal_933) ) ;
    buf_clk new_AGEMA_reg_buffer_466 ( .C (clk), .D (new_AGEMA_signal_211), .Q (new_AGEMA_signal_939) ) ;
    buf_clk new_AGEMA_reg_buffer_472 ( .C (clk), .D (new_AGEMA_signal_212), .Q (new_AGEMA_signal_945) ) ;
    buf_clk new_AGEMA_reg_buffer_478 ( .C (clk), .D (T1), .Q (new_AGEMA_signal_951) ) ;
    buf_clk new_AGEMA_reg_buffer_484 ( .C (clk), .D (new_AGEMA_signal_155), .Q (new_AGEMA_signal_957) ) ;
    buf_clk new_AGEMA_reg_buffer_490 ( .C (clk), .D (new_AGEMA_signal_156), .Q (new_AGEMA_signal_963) ) ;
    buf_clk new_AGEMA_reg_buffer_496 ( .C (clk), .D (T4), .Q (new_AGEMA_signal_969) ) ;
    buf_clk new_AGEMA_reg_buffer_502 ( .C (clk), .D (new_AGEMA_signal_165), .Q (new_AGEMA_signal_975) ) ;
    buf_clk new_AGEMA_reg_buffer_508 ( .C (clk), .D (new_AGEMA_signal_166), .Q (new_AGEMA_signal_981) ) ;
    buf_clk new_AGEMA_reg_buffer_514 ( .C (clk), .D (T2), .Q (new_AGEMA_signal_987) ) ;
    buf_clk new_AGEMA_reg_buffer_520 ( .C (clk), .D (new_AGEMA_signal_159), .Q (new_AGEMA_signal_993) ) ;
    buf_clk new_AGEMA_reg_buffer_526 ( .C (clk), .D (new_AGEMA_signal_160), .Q (new_AGEMA_signal_999) ) ;

    /* cells in depth 2 */
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M1_U1 ( .ina ({new_AGEMA_signal_192, new_AGEMA_signal_191, T13}), .inb ({new_AGEMA_signal_188, new_AGEMA_signal_187, T6}), .clk (clk), .rnd ({Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .outt ({new_AGEMA_signal_218, new_AGEMA_signal_217, M1}) ) ;
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M2_U1 ( .ina ({new_AGEMA_signal_214, new_AGEMA_signal_213, T23}), .inb ({new_AGEMA_signal_204, new_AGEMA_signal_203, T8}), .clk (clk), .rnd ({Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5]}), .outt ({new_AGEMA_signal_234, new_AGEMA_signal_233, M2}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_M3_U1 ( .a ({new_AGEMA_signal_614, new_AGEMA_signal_612, new_AGEMA_signal_610}), .b ({new_AGEMA_signal_218, new_AGEMA_signal_217, M1}), .c ({new_AGEMA_signal_236, new_AGEMA_signal_235, M3}) ) ;
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M4_U1 ( .ina ({new_AGEMA_signal_198, new_AGEMA_signal_197, T19}), .inb ({X_s2[0], X_s1[0], X_s0[0]}), .clk (clk), .rnd ({Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10]}), .outt ({new_AGEMA_signal_220, new_AGEMA_signal_219, M4}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_M5_U1 ( .a ({new_AGEMA_signal_220, new_AGEMA_signal_219, M4}), .b ({new_AGEMA_signal_218, new_AGEMA_signal_217, M1}), .c ({new_AGEMA_signal_238, new_AGEMA_signal_237, M5}) ) ;
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M6_U1 ( .ina ({new_AGEMA_signal_164, new_AGEMA_signal_163, T3}), .inb ({new_AGEMA_signal_196, new_AGEMA_signal_195, T16}), .clk (clk), .rnd ({Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15]}), .outt ({new_AGEMA_signal_222, new_AGEMA_signal_221, M6}) ) ;
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M7_U1 ( .ina ({new_AGEMA_signal_200, new_AGEMA_signal_199, T22}), .inb ({new_AGEMA_signal_190, new_AGEMA_signal_189, T9}), .clk (clk), .rnd ({Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20]}), .outt ({new_AGEMA_signal_224, new_AGEMA_signal_223, M7}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_M8_U1 ( .a ({new_AGEMA_signal_620, new_AGEMA_signal_618, new_AGEMA_signal_616}), .b ({new_AGEMA_signal_222, new_AGEMA_signal_221, M6}), .c ({new_AGEMA_signal_240, new_AGEMA_signal_239, M8}) ) ;
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M9_U1 ( .ina ({new_AGEMA_signal_212, new_AGEMA_signal_211, T20}), .inb ({new_AGEMA_signal_210, new_AGEMA_signal_209, T17}), .clk (clk), .rnd ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25]}), .outt ({new_AGEMA_signal_242, new_AGEMA_signal_241, M9}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_M10_U1 ( .a ({new_AGEMA_signal_242, new_AGEMA_signal_241, M9}), .b ({new_AGEMA_signal_222, new_AGEMA_signal_221, M6}), .c ({new_AGEMA_signal_248, new_AGEMA_signal_247, M10}) ) ;
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M11_U1 ( .ina ({new_AGEMA_signal_156, new_AGEMA_signal_155, T1}), .inb ({new_AGEMA_signal_194, new_AGEMA_signal_193, T15}), .clk (clk), .rnd ({Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .outt ({new_AGEMA_signal_226, new_AGEMA_signal_225, M11}) ) ;
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M12_U1 ( .ina ({new_AGEMA_signal_166, new_AGEMA_signal_165, T4}), .inb ({new_AGEMA_signal_202, new_AGEMA_signal_201, T27}), .clk (clk), .rnd ({Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35]}), .outt ({new_AGEMA_signal_228, new_AGEMA_signal_227, M12}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_M13_U1 ( .a ({new_AGEMA_signal_228, new_AGEMA_signal_227, M12}), .b ({new_AGEMA_signal_226, new_AGEMA_signal_225, M11}), .c ({new_AGEMA_signal_244, new_AGEMA_signal_243, M13}) ) ;
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M14_U1 ( .ina ({new_AGEMA_signal_160, new_AGEMA_signal_159, T2}), .inb ({new_AGEMA_signal_206, new_AGEMA_signal_205, T10}), .clk (clk), .rnd ({Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40]}), .outt ({new_AGEMA_signal_246, new_AGEMA_signal_245, M14}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_M15_U1 ( .a ({new_AGEMA_signal_246, new_AGEMA_signal_245, M14}), .b ({new_AGEMA_signal_226, new_AGEMA_signal_225, M11}), .c ({new_AGEMA_signal_250, new_AGEMA_signal_249, M15}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_M16_U1 ( .a ({new_AGEMA_signal_236, new_AGEMA_signal_235, M3}), .b ({new_AGEMA_signal_234, new_AGEMA_signal_233, M2}), .c ({new_AGEMA_signal_252, new_AGEMA_signal_251, M16}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_M17_U1 ( .a ({new_AGEMA_signal_238, new_AGEMA_signal_237, M5}), .b ({new_AGEMA_signal_626, new_AGEMA_signal_624, new_AGEMA_signal_622}), .c ({new_AGEMA_signal_254, new_AGEMA_signal_253, M17}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_M18_U1 ( .a ({new_AGEMA_signal_240, new_AGEMA_signal_239, M8}), .b ({new_AGEMA_signal_224, new_AGEMA_signal_223, M7}), .c ({new_AGEMA_signal_256, new_AGEMA_signal_255, M18}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_M19_U1 ( .a ({new_AGEMA_signal_248, new_AGEMA_signal_247, M10}), .b ({new_AGEMA_signal_250, new_AGEMA_signal_249, M15}), .c ({new_AGEMA_signal_258, new_AGEMA_signal_257, M19}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_M20_U1 ( .a ({new_AGEMA_signal_252, new_AGEMA_signal_251, M16}), .b ({new_AGEMA_signal_244, new_AGEMA_signal_243, M13}), .c ({new_AGEMA_signal_260, new_AGEMA_signal_259, M20}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_M21_U1 ( .a ({new_AGEMA_signal_254, new_AGEMA_signal_253, M17}), .b ({new_AGEMA_signal_250, new_AGEMA_signal_249, M15}), .c ({new_AGEMA_signal_262, new_AGEMA_signal_261, M21}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_M22_U1 ( .a ({new_AGEMA_signal_256, new_AGEMA_signal_255, M18}), .b ({new_AGEMA_signal_244, new_AGEMA_signal_243, M13}), .c ({new_AGEMA_signal_264, new_AGEMA_signal_263, M22}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_M23_U1 ( .a ({new_AGEMA_signal_258, new_AGEMA_signal_257, M19}), .b ({new_AGEMA_signal_632, new_AGEMA_signal_630, new_AGEMA_signal_628}), .c ({new_AGEMA_signal_266, new_AGEMA_signal_265, M23}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_M24_U1 ( .a ({new_AGEMA_signal_264, new_AGEMA_signal_263, M22}), .b ({new_AGEMA_signal_266, new_AGEMA_signal_265, M23}), .c ({new_AGEMA_signal_274, new_AGEMA_signal_273, M24}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_M27_U1 ( .a ({new_AGEMA_signal_260, new_AGEMA_signal_259, M20}), .b ({new_AGEMA_signal_262, new_AGEMA_signal_261, M21}), .c ({new_AGEMA_signal_270, new_AGEMA_signal_269, M27}) ) ;
    buf_clk new_AGEMA_reg_buffer_137 ( .C (clk), .D (new_AGEMA_signal_609), .Q (new_AGEMA_signal_610) ) ;
    buf_clk new_AGEMA_reg_buffer_139 ( .C (clk), .D (new_AGEMA_signal_611), .Q (new_AGEMA_signal_612) ) ;
    buf_clk new_AGEMA_reg_buffer_141 ( .C (clk), .D (new_AGEMA_signal_613), .Q (new_AGEMA_signal_614) ) ;
    buf_clk new_AGEMA_reg_buffer_143 ( .C (clk), .D (new_AGEMA_signal_615), .Q (new_AGEMA_signal_616) ) ;
    buf_clk new_AGEMA_reg_buffer_145 ( .C (clk), .D (new_AGEMA_signal_617), .Q (new_AGEMA_signal_618) ) ;
    buf_clk new_AGEMA_reg_buffer_147 ( .C (clk), .D (new_AGEMA_signal_619), .Q (new_AGEMA_signal_620) ) ;
    buf_clk new_AGEMA_reg_buffer_149 ( .C (clk), .D (new_AGEMA_signal_621), .Q (new_AGEMA_signal_622) ) ;
    buf_clk new_AGEMA_reg_buffer_151 ( .C (clk), .D (new_AGEMA_signal_623), .Q (new_AGEMA_signal_624) ) ;
    buf_clk new_AGEMA_reg_buffer_153 ( .C (clk), .D (new_AGEMA_signal_625), .Q (new_AGEMA_signal_626) ) ;
    buf_clk new_AGEMA_reg_buffer_155 ( .C (clk), .D (new_AGEMA_signal_627), .Q (new_AGEMA_signal_628) ) ;
    buf_clk new_AGEMA_reg_buffer_157 ( .C (clk), .D (new_AGEMA_signal_629), .Q (new_AGEMA_signal_630) ) ;
    buf_clk new_AGEMA_reg_buffer_159 ( .C (clk), .D (new_AGEMA_signal_631), .Q (new_AGEMA_signal_632) ) ;
    buf_clk new_AGEMA_reg_buffer_209 ( .C (clk), .D (new_AGEMA_signal_681), .Q (new_AGEMA_signal_682) ) ;
    buf_clk new_AGEMA_reg_buffer_215 ( .C (clk), .D (new_AGEMA_signal_687), .Q (new_AGEMA_signal_688) ) ;
    buf_clk new_AGEMA_reg_buffer_221 ( .C (clk), .D (new_AGEMA_signal_693), .Q (new_AGEMA_signal_694) ) ;
    buf_clk new_AGEMA_reg_buffer_227 ( .C (clk), .D (new_AGEMA_signal_699), .Q (new_AGEMA_signal_700) ) ;
    buf_clk new_AGEMA_reg_buffer_233 ( .C (clk), .D (new_AGEMA_signal_705), .Q (new_AGEMA_signal_706) ) ;
    buf_clk new_AGEMA_reg_buffer_239 ( .C (clk), .D (new_AGEMA_signal_711), .Q (new_AGEMA_signal_712) ) ;
    buf_clk new_AGEMA_reg_buffer_245 ( .C (clk), .D (new_AGEMA_signal_717), .Q (new_AGEMA_signal_718) ) ;
    buf_clk new_AGEMA_reg_buffer_251 ( .C (clk), .D (new_AGEMA_signal_723), .Q (new_AGEMA_signal_724) ) ;
    buf_clk new_AGEMA_reg_buffer_257 ( .C (clk), .D (new_AGEMA_signal_729), .Q (new_AGEMA_signal_730) ) ;
    buf_clk new_AGEMA_reg_buffer_263 ( .C (clk), .D (new_AGEMA_signal_735), .Q (new_AGEMA_signal_736) ) ;
    buf_clk new_AGEMA_reg_buffer_269 ( .C (clk), .D (new_AGEMA_signal_741), .Q (new_AGEMA_signal_742) ) ;
    buf_clk new_AGEMA_reg_buffer_275 ( .C (clk), .D (new_AGEMA_signal_747), .Q (new_AGEMA_signal_748) ) ;
    buf_clk new_AGEMA_reg_buffer_281 ( .C (clk), .D (new_AGEMA_signal_753), .Q (new_AGEMA_signal_754) ) ;
    buf_clk new_AGEMA_reg_buffer_287 ( .C (clk), .D (new_AGEMA_signal_759), .Q (new_AGEMA_signal_760) ) ;
    buf_clk new_AGEMA_reg_buffer_293 ( .C (clk), .D (new_AGEMA_signal_765), .Q (new_AGEMA_signal_766) ) ;
    buf_clk new_AGEMA_reg_buffer_299 ( .C (clk), .D (new_AGEMA_signal_771), .Q (new_AGEMA_signal_772) ) ;
    buf_clk new_AGEMA_reg_buffer_305 ( .C (clk), .D (new_AGEMA_signal_777), .Q (new_AGEMA_signal_778) ) ;
    buf_clk new_AGEMA_reg_buffer_311 ( .C (clk), .D (new_AGEMA_signal_783), .Q (new_AGEMA_signal_784) ) ;
    buf_clk new_AGEMA_reg_buffer_317 ( .C (clk), .D (new_AGEMA_signal_789), .Q (new_AGEMA_signal_790) ) ;
    buf_clk new_AGEMA_reg_buffer_323 ( .C (clk), .D (new_AGEMA_signal_795), .Q (new_AGEMA_signal_796) ) ;
    buf_clk new_AGEMA_reg_buffer_329 ( .C (clk), .D (new_AGEMA_signal_801), .Q (new_AGEMA_signal_802) ) ;
    buf_clk new_AGEMA_reg_buffer_335 ( .C (clk), .D (new_AGEMA_signal_807), .Q (new_AGEMA_signal_808) ) ;
    buf_clk new_AGEMA_reg_buffer_341 ( .C (clk), .D (new_AGEMA_signal_813), .Q (new_AGEMA_signal_814) ) ;
    buf_clk new_AGEMA_reg_buffer_347 ( .C (clk), .D (new_AGEMA_signal_819), .Q (new_AGEMA_signal_820) ) ;
    buf_clk new_AGEMA_reg_buffer_353 ( .C (clk), .D (new_AGEMA_signal_825), .Q (new_AGEMA_signal_826) ) ;
    buf_clk new_AGEMA_reg_buffer_359 ( .C (clk), .D (new_AGEMA_signal_831), .Q (new_AGEMA_signal_832) ) ;
    buf_clk new_AGEMA_reg_buffer_365 ( .C (clk), .D (new_AGEMA_signal_837), .Q (new_AGEMA_signal_838) ) ;
    buf_clk new_AGEMA_reg_buffer_371 ( .C (clk), .D (new_AGEMA_signal_843), .Q (new_AGEMA_signal_844) ) ;
    buf_clk new_AGEMA_reg_buffer_377 ( .C (clk), .D (new_AGEMA_signal_849), .Q (new_AGEMA_signal_850) ) ;
    buf_clk new_AGEMA_reg_buffer_383 ( .C (clk), .D (new_AGEMA_signal_855), .Q (new_AGEMA_signal_856) ) ;
    buf_clk new_AGEMA_reg_buffer_389 ( .C (clk), .D (new_AGEMA_signal_861), .Q (new_AGEMA_signal_862) ) ;
    buf_clk new_AGEMA_reg_buffer_395 ( .C (clk), .D (new_AGEMA_signal_867), .Q (new_AGEMA_signal_868) ) ;
    buf_clk new_AGEMA_reg_buffer_401 ( .C (clk), .D (new_AGEMA_signal_873), .Q (new_AGEMA_signal_874) ) ;
    buf_clk new_AGEMA_reg_buffer_407 ( .C (clk), .D (new_AGEMA_signal_879), .Q (new_AGEMA_signal_880) ) ;
    buf_clk new_AGEMA_reg_buffer_413 ( .C (clk), .D (new_AGEMA_signal_885), .Q (new_AGEMA_signal_886) ) ;
    buf_clk new_AGEMA_reg_buffer_419 ( .C (clk), .D (new_AGEMA_signal_891), .Q (new_AGEMA_signal_892) ) ;
    buf_clk new_AGEMA_reg_buffer_425 ( .C (clk), .D (new_AGEMA_signal_897), .Q (new_AGEMA_signal_898) ) ;
    buf_clk new_AGEMA_reg_buffer_431 ( .C (clk), .D (new_AGEMA_signal_903), .Q (new_AGEMA_signal_904) ) ;
    buf_clk new_AGEMA_reg_buffer_437 ( .C (clk), .D (new_AGEMA_signal_909), .Q (new_AGEMA_signal_910) ) ;
    buf_clk new_AGEMA_reg_buffer_443 ( .C (clk), .D (new_AGEMA_signal_915), .Q (new_AGEMA_signal_916) ) ;
    buf_clk new_AGEMA_reg_buffer_449 ( .C (clk), .D (new_AGEMA_signal_921), .Q (new_AGEMA_signal_922) ) ;
    buf_clk new_AGEMA_reg_buffer_455 ( .C (clk), .D (new_AGEMA_signal_927), .Q (new_AGEMA_signal_928) ) ;
    buf_clk new_AGEMA_reg_buffer_461 ( .C (clk), .D (new_AGEMA_signal_933), .Q (new_AGEMA_signal_934) ) ;
    buf_clk new_AGEMA_reg_buffer_467 ( .C (clk), .D (new_AGEMA_signal_939), .Q (new_AGEMA_signal_940) ) ;
    buf_clk new_AGEMA_reg_buffer_473 ( .C (clk), .D (new_AGEMA_signal_945), .Q (new_AGEMA_signal_946) ) ;
    buf_clk new_AGEMA_reg_buffer_479 ( .C (clk), .D (new_AGEMA_signal_951), .Q (new_AGEMA_signal_952) ) ;
    buf_clk new_AGEMA_reg_buffer_485 ( .C (clk), .D (new_AGEMA_signal_957), .Q (new_AGEMA_signal_958) ) ;
    buf_clk new_AGEMA_reg_buffer_491 ( .C (clk), .D (new_AGEMA_signal_963), .Q (new_AGEMA_signal_964) ) ;
    buf_clk new_AGEMA_reg_buffer_497 ( .C (clk), .D (new_AGEMA_signal_969), .Q (new_AGEMA_signal_970) ) ;
    buf_clk new_AGEMA_reg_buffer_503 ( .C (clk), .D (new_AGEMA_signal_975), .Q (new_AGEMA_signal_976) ) ;
    buf_clk new_AGEMA_reg_buffer_509 ( .C (clk), .D (new_AGEMA_signal_981), .Q (new_AGEMA_signal_982) ) ;
    buf_clk new_AGEMA_reg_buffer_515 ( .C (clk), .D (new_AGEMA_signal_987), .Q (new_AGEMA_signal_988) ) ;
    buf_clk new_AGEMA_reg_buffer_521 ( .C (clk), .D (new_AGEMA_signal_993), .Q (new_AGEMA_signal_994) ) ;
    buf_clk new_AGEMA_reg_buffer_527 ( .C (clk), .D (new_AGEMA_signal_999), .Q (new_AGEMA_signal_1000) ) ;

    /* cells in depth 3 */
    buf_clk new_AGEMA_reg_buffer_160 ( .C (clk), .D (M21), .Q (new_AGEMA_signal_633) ) ;
    buf_clk new_AGEMA_reg_buffer_162 ( .C (clk), .D (new_AGEMA_signal_261), .Q (new_AGEMA_signal_635) ) ;
    buf_clk new_AGEMA_reg_buffer_164 ( .C (clk), .D (new_AGEMA_signal_262), .Q (new_AGEMA_signal_637) ) ;
    buf_clk new_AGEMA_reg_buffer_166 ( .C (clk), .D (M23), .Q (new_AGEMA_signal_639) ) ;
    buf_clk new_AGEMA_reg_buffer_168 ( .C (clk), .D (new_AGEMA_signal_265), .Q (new_AGEMA_signal_641) ) ;
    buf_clk new_AGEMA_reg_buffer_170 ( .C (clk), .D (new_AGEMA_signal_266), .Q (new_AGEMA_signal_643) ) ;
    buf_clk new_AGEMA_reg_buffer_172 ( .C (clk), .D (M27), .Q (new_AGEMA_signal_645) ) ;
    buf_clk new_AGEMA_reg_buffer_174 ( .C (clk), .D (new_AGEMA_signal_269), .Q (new_AGEMA_signal_647) ) ;
    buf_clk new_AGEMA_reg_buffer_176 ( .C (clk), .D (new_AGEMA_signal_270), .Q (new_AGEMA_signal_649) ) ;
    buf_clk new_AGEMA_reg_buffer_178 ( .C (clk), .D (M24), .Q (new_AGEMA_signal_651) ) ;
    buf_clk new_AGEMA_reg_buffer_180 ( .C (clk), .D (new_AGEMA_signal_273), .Q (new_AGEMA_signal_653) ) ;
    buf_clk new_AGEMA_reg_buffer_182 ( .C (clk), .D (new_AGEMA_signal_274), .Q (new_AGEMA_signal_655) ) ;
    buf_clk new_AGEMA_reg_buffer_210 ( .C (clk), .D (new_AGEMA_signal_682), .Q (new_AGEMA_signal_683) ) ;
    buf_clk new_AGEMA_reg_buffer_216 ( .C (clk), .D (new_AGEMA_signal_688), .Q (new_AGEMA_signal_689) ) ;
    buf_clk new_AGEMA_reg_buffer_222 ( .C (clk), .D (new_AGEMA_signal_694), .Q (new_AGEMA_signal_695) ) ;
    buf_clk new_AGEMA_reg_buffer_228 ( .C (clk), .D (new_AGEMA_signal_700), .Q (new_AGEMA_signal_701) ) ;
    buf_clk new_AGEMA_reg_buffer_234 ( .C (clk), .D (new_AGEMA_signal_706), .Q (new_AGEMA_signal_707) ) ;
    buf_clk new_AGEMA_reg_buffer_240 ( .C (clk), .D (new_AGEMA_signal_712), .Q (new_AGEMA_signal_713) ) ;
    buf_clk new_AGEMA_reg_buffer_246 ( .C (clk), .D (new_AGEMA_signal_718), .Q (new_AGEMA_signal_719) ) ;
    buf_clk new_AGEMA_reg_buffer_252 ( .C (clk), .D (new_AGEMA_signal_724), .Q (new_AGEMA_signal_725) ) ;
    buf_clk new_AGEMA_reg_buffer_258 ( .C (clk), .D (new_AGEMA_signal_730), .Q (new_AGEMA_signal_731) ) ;
    buf_clk new_AGEMA_reg_buffer_264 ( .C (clk), .D (new_AGEMA_signal_736), .Q (new_AGEMA_signal_737) ) ;
    buf_clk new_AGEMA_reg_buffer_270 ( .C (clk), .D (new_AGEMA_signal_742), .Q (new_AGEMA_signal_743) ) ;
    buf_clk new_AGEMA_reg_buffer_276 ( .C (clk), .D (new_AGEMA_signal_748), .Q (new_AGEMA_signal_749) ) ;
    buf_clk new_AGEMA_reg_buffer_282 ( .C (clk), .D (new_AGEMA_signal_754), .Q (new_AGEMA_signal_755) ) ;
    buf_clk new_AGEMA_reg_buffer_288 ( .C (clk), .D (new_AGEMA_signal_760), .Q (new_AGEMA_signal_761) ) ;
    buf_clk new_AGEMA_reg_buffer_294 ( .C (clk), .D (new_AGEMA_signal_766), .Q (new_AGEMA_signal_767) ) ;
    buf_clk new_AGEMA_reg_buffer_300 ( .C (clk), .D (new_AGEMA_signal_772), .Q (new_AGEMA_signal_773) ) ;
    buf_clk new_AGEMA_reg_buffer_306 ( .C (clk), .D (new_AGEMA_signal_778), .Q (new_AGEMA_signal_779) ) ;
    buf_clk new_AGEMA_reg_buffer_312 ( .C (clk), .D (new_AGEMA_signal_784), .Q (new_AGEMA_signal_785) ) ;
    buf_clk new_AGEMA_reg_buffer_318 ( .C (clk), .D (new_AGEMA_signal_790), .Q (new_AGEMA_signal_791) ) ;
    buf_clk new_AGEMA_reg_buffer_324 ( .C (clk), .D (new_AGEMA_signal_796), .Q (new_AGEMA_signal_797) ) ;
    buf_clk new_AGEMA_reg_buffer_330 ( .C (clk), .D (new_AGEMA_signal_802), .Q (new_AGEMA_signal_803) ) ;
    buf_clk new_AGEMA_reg_buffer_336 ( .C (clk), .D (new_AGEMA_signal_808), .Q (new_AGEMA_signal_809) ) ;
    buf_clk new_AGEMA_reg_buffer_342 ( .C (clk), .D (new_AGEMA_signal_814), .Q (new_AGEMA_signal_815) ) ;
    buf_clk new_AGEMA_reg_buffer_348 ( .C (clk), .D (new_AGEMA_signal_820), .Q (new_AGEMA_signal_821) ) ;
    buf_clk new_AGEMA_reg_buffer_354 ( .C (clk), .D (new_AGEMA_signal_826), .Q (new_AGEMA_signal_827) ) ;
    buf_clk new_AGEMA_reg_buffer_360 ( .C (clk), .D (new_AGEMA_signal_832), .Q (new_AGEMA_signal_833) ) ;
    buf_clk new_AGEMA_reg_buffer_366 ( .C (clk), .D (new_AGEMA_signal_838), .Q (new_AGEMA_signal_839) ) ;
    buf_clk new_AGEMA_reg_buffer_372 ( .C (clk), .D (new_AGEMA_signal_844), .Q (new_AGEMA_signal_845) ) ;
    buf_clk new_AGEMA_reg_buffer_378 ( .C (clk), .D (new_AGEMA_signal_850), .Q (new_AGEMA_signal_851) ) ;
    buf_clk new_AGEMA_reg_buffer_384 ( .C (clk), .D (new_AGEMA_signal_856), .Q (new_AGEMA_signal_857) ) ;
    buf_clk new_AGEMA_reg_buffer_390 ( .C (clk), .D (new_AGEMA_signal_862), .Q (new_AGEMA_signal_863) ) ;
    buf_clk new_AGEMA_reg_buffer_396 ( .C (clk), .D (new_AGEMA_signal_868), .Q (new_AGEMA_signal_869) ) ;
    buf_clk new_AGEMA_reg_buffer_402 ( .C (clk), .D (new_AGEMA_signal_874), .Q (new_AGEMA_signal_875) ) ;
    buf_clk new_AGEMA_reg_buffer_408 ( .C (clk), .D (new_AGEMA_signal_880), .Q (new_AGEMA_signal_881) ) ;
    buf_clk new_AGEMA_reg_buffer_414 ( .C (clk), .D (new_AGEMA_signal_886), .Q (new_AGEMA_signal_887) ) ;
    buf_clk new_AGEMA_reg_buffer_420 ( .C (clk), .D (new_AGEMA_signal_892), .Q (new_AGEMA_signal_893) ) ;
    buf_clk new_AGEMA_reg_buffer_426 ( .C (clk), .D (new_AGEMA_signal_898), .Q (new_AGEMA_signal_899) ) ;
    buf_clk new_AGEMA_reg_buffer_432 ( .C (clk), .D (new_AGEMA_signal_904), .Q (new_AGEMA_signal_905) ) ;
    buf_clk new_AGEMA_reg_buffer_438 ( .C (clk), .D (new_AGEMA_signal_910), .Q (new_AGEMA_signal_911) ) ;
    buf_clk new_AGEMA_reg_buffer_444 ( .C (clk), .D (new_AGEMA_signal_916), .Q (new_AGEMA_signal_917) ) ;
    buf_clk new_AGEMA_reg_buffer_450 ( .C (clk), .D (new_AGEMA_signal_922), .Q (new_AGEMA_signal_923) ) ;
    buf_clk new_AGEMA_reg_buffer_456 ( .C (clk), .D (new_AGEMA_signal_928), .Q (new_AGEMA_signal_929) ) ;
    buf_clk new_AGEMA_reg_buffer_462 ( .C (clk), .D (new_AGEMA_signal_934), .Q (new_AGEMA_signal_935) ) ;
    buf_clk new_AGEMA_reg_buffer_468 ( .C (clk), .D (new_AGEMA_signal_940), .Q (new_AGEMA_signal_941) ) ;
    buf_clk new_AGEMA_reg_buffer_474 ( .C (clk), .D (new_AGEMA_signal_946), .Q (new_AGEMA_signal_947) ) ;
    buf_clk new_AGEMA_reg_buffer_480 ( .C (clk), .D (new_AGEMA_signal_952), .Q (new_AGEMA_signal_953) ) ;
    buf_clk new_AGEMA_reg_buffer_486 ( .C (clk), .D (new_AGEMA_signal_958), .Q (new_AGEMA_signal_959) ) ;
    buf_clk new_AGEMA_reg_buffer_492 ( .C (clk), .D (new_AGEMA_signal_964), .Q (new_AGEMA_signal_965) ) ;
    buf_clk new_AGEMA_reg_buffer_498 ( .C (clk), .D (new_AGEMA_signal_970), .Q (new_AGEMA_signal_971) ) ;
    buf_clk new_AGEMA_reg_buffer_504 ( .C (clk), .D (new_AGEMA_signal_976), .Q (new_AGEMA_signal_977) ) ;
    buf_clk new_AGEMA_reg_buffer_510 ( .C (clk), .D (new_AGEMA_signal_982), .Q (new_AGEMA_signal_983) ) ;
    buf_clk new_AGEMA_reg_buffer_516 ( .C (clk), .D (new_AGEMA_signal_988), .Q (new_AGEMA_signal_989) ) ;
    buf_clk new_AGEMA_reg_buffer_522 ( .C (clk), .D (new_AGEMA_signal_994), .Q (new_AGEMA_signal_995) ) ;
    buf_clk new_AGEMA_reg_buffer_528 ( .C (clk), .D (new_AGEMA_signal_1000), .Q (new_AGEMA_signal_1001) ) ;

    /* cells in depth 4 */
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M25_U1 ( .ina ({new_AGEMA_signal_264, new_AGEMA_signal_263, M22}), .inb ({new_AGEMA_signal_260, new_AGEMA_signal_259, M20}), .clk (clk), .rnd ({Fresh[49], Fresh[48], Fresh[47], Fresh[46], Fresh[45]}), .outt ({new_AGEMA_signal_268, new_AGEMA_signal_267, M25}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_M26_U1 ( .a ({new_AGEMA_signal_638, new_AGEMA_signal_636, new_AGEMA_signal_634}), .b ({new_AGEMA_signal_268, new_AGEMA_signal_267, M25}), .c ({new_AGEMA_signal_276, new_AGEMA_signal_275, M26}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_M28_U1 ( .a ({new_AGEMA_signal_644, new_AGEMA_signal_642, new_AGEMA_signal_640}), .b ({new_AGEMA_signal_268, new_AGEMA_signal_267, M25}), .c ({new_AGEMA_signal_278, new_AGEMA_signal_277, M28}) ) ;
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M31_U1 ( .ina ({new_AGEMA_signal_260, new_AGEMA_signal_259, M20}), .inb ({new_AGEMA_signal_266, new_AGEMA_signal_265, M23}), .clk (clk), .rnd ({Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50]}), .outt ({new_AGEMA_signal_280, new_AGEMA_signal_279, M31}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_M33_U1 ( .a ({new_AGEMA_signal_650, new_AGEMA_signal_648, new_AGEMA_signal_646}), .b ({new_AGEMA_signal_268, new_AGEMA_signal_267, M25}), .c ({new_AGEMA_signal_282, new_AGEMA_signal_281, M33}) ) ;
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M34_U1 ( .ina ({new_AGEMA_signal_262, new_AGEMA_signal_261, M21}), .inb ({new_AGEMA_signal_264, new_AGEMA_signal_263, M22}), .clk (clk), .rnd ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55]}), .outt ({new_AGEMA_signal_272, new_AGEMA_signal_271, M34}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_M36_U1 ( .a ({new_AGEMA_signal_656, new_AGEMA_signal_654, new_AGEMA_signal_652}), .b ({new_AGEMA_signal_268, new_AGEMA_signal_267, M25}), .c ({new_AGEMA_signal_292, new_AGEMA_signal_291, M36}) ) ;
    buf_clk new_AGEMA_reg_buffer_161 ( .C (clk), .D (new_AGEMA_signal_633), .Q (new_AGEMA_signal_634) ) ;
    buf_clk new_AGEMA_reg_buffer_163 ( .C (clk), .D (new_AGEMA_signal_635), .Q (new_AGEMA_signal_636) ) ;
    buf_clk new_AGEMA_reg_buffer_165 ( .C (clk), .D (new_AGEMA_signal_637), .Q (new_AGEMA_signal_638) ) ;
    buf_clk new_AGEMA_reg_buffer_167 ( .C (clk), .D (new_AGEMA_signal_639), .Q (new_AGEMA_signal_640) ) ;
    buf_clk new_AGEMA_reg_buffer_169 ( .C (clk), .D (new_AGEMA_signal_641), .Q (new_AGEMA_signal_642) ) ;
    buf_clk new_AGEMA_reg_buffer_171 ( .C (clk), .D (new_AGEMA_signal_643), .Q (new_AGEMA_signal_644) ) ;
    buf_clk new_AGEMA_reg_buffer_173 ( .C (clk), .D (new_AGEMA_signal_645), .Q (new_AGEMA_signal_646) ) ;
    buf_clk new_AGEMA_reg_buffer_175 ( .C (clk), .D (new_AGEMA_signal_647), .Q (new_AGEMA_signal_648) ) ;
    buf_clk new_AGEMA_reg_buffer_177 ( .C (clk), .D (new_AGEMA_signal_649), .Q (new_AGEMA_signal_650) ) ;
    buf_clk new_AGEMA_reg_buffer_179 ( .C (clk), .D (new_AGEMA_signal_651), .Q (new_AGEMA_signal_652) ) ;
    buf_clk new_AGEMA_reg_buffer_181 ( .C (clk), .D (new_AGEMA_signal_653), .Q (new_AGEMA_signal_654) ) ;
    buf_clk new_AGEMA_reg_buffer_183 ( .C (clk), .D (new_AGEMA_signal_655), .Q (new_AGEMA_signal_656) ) ;
    buf_clk new_AGEMA_reg_buffer_211 ( .C (clk), .D (new_AGEMA_signal_683), .Q (new_AGEMA_signal_684) ) ;
    buf_clk new_AGEMA_reg_buffer_217 ( .C (clk), .D (new_AGEMA_signal_689), .Q (new_AGEMA_signal_690) ) ;
    buf_clk new_AGEMA_reg_buffer_223 ( .C (clk), .D (new_AGEMA_signal_695), .Q (new_AGEMA_signal_696) ) ;
    buf_clk new_AGEMA_reg_buffer_229 ( .C (clk), .D (new_AGEMA_signal_701), .Q (new_AGEMA_signal_702) ) ;
    buf_clk new_AGEMA_reg_buffer_235 ( .C (clk), .D (new_AGEMA_signal_707), .Q (new_AGEMA_signal_708) ) ;
    buf_clk new_AGEMA_reg_buffer_241 ( .C (clk), .D (new_AGEMA_signal_713), .Q (new_AGEMA_signal_714) ) ;
    buf_clk new_AGEMA_reg_buffer_247 ( .C (clk), .D (new_AGEMA_signal_719), .Q (new_AGEMA_signal_720) ) ;
    buf_clk new_AGEMA_reg_buffer_253 ( .C (clk), .D (new_AGEMA_signal_725), .Q (new_AGEMA_signal_726) ) ;
    buf_clk new_AGEMA_reg_buffer_259 ( .C (clk), .D (new_AGEMA_signal_731), .Q (new_AGEMA_signal_732) ) ;
    buf_clk new_AGEMA_reg_buffer_265 ( .C (clk), .D (new_AGEMA_signal_737), .Q (new_AGEMA_signal_738) ) ;
    buf_clk new_AGEMA_reg_buffer_271 ( .C (clk), .D (new_AGEMA_signal_743), .Q (new_AGEMA_signal_744) ) ;
    buf_clk new_AGEMA_reg_buffer_277 ( .C (clk), .D (new_AGEMA_signal_749), .Q (new_AGEMA_signal_750) ) ;
    buf_clk new_AGEMA_reg_buffer_283 ( .C (clk), .D (new_AGEMA_signal_755), .Q (new_AGEMA_signal_756) ) ;
    buf_clk new_AGEMA_reg_buffer_289 ( .C (clk), .D (new_AGEMA_signal_761), .Q (new_AGEMA_signal_762) ) ;
    buf_clk new_AGEMA_reg_buffer_295 ( .C (clk), .D (new_AGEMA_signal_767), .Q (new_AGEMA_signal_768) ) ;
    buf_clk new_AGEMA_reg_buffer_301 ( .C (clk), .D (new_AGEMA_signal_773), .Q (new_AGEMA_signal_774) ) ;
    buf_clk new_AGEMA_reg_buffer_307 ( .C (clk), .D (new_AGEMA_signal_779), .Q (new_AGEMA_signal_780) ) ;
    buf_clk new_AGEMA_reg_buffer_313 ( .C (clk), .D (new_AGEMA_signal_785), .Q (new_AGEMA_signal_786) ) ;
    buf_clk new_AGEMA_reg_buffer_319 ( .C (clk), .D (new_AGEMA_signal_791), .Q (new_AGEMA_signal_792) ) ;
    buf_clk new_AGEMA_reg_buffer_325 ( .C (clk), .D (new_AGEMA_signal_797), .Q (new_AGEMA_signal_798) ) ;
    buf_clk new_AGEMA_reg_buffer_331 ( .C (clk), .D (new_AGEMA_signal_803), .Q (new_AGEMA_signal_804) ) ;
    buf_clk new_AGEMA_reg_buffer_337 ( .C (clk), .D (new_AGEMA_signal_809), .Q (new_AGEMA_signal_810) ) ;
    buf_clk new_AGEMA_reg_buffer_343 ( .C (clk), .D (new_AGEMA_signal_815), .Q (new_AGEMA_signal_816) ) ;
    buf_clk new_AGEMA_reg_buffer_349 ( .C (clk), .D (new_AGEMA_signal_821), .Q (new_AGEMA_signal_822) ) ;
    buf_clk new_AGEMA_reg_buffer_355 ( .C (clk), .D (new_AGEMA_signal_827), .Q (new_AGEMA_signal_828) ) ;
    buf_clk new_AGEMA_reg_buffer_361 ( .C (clk), .D (new_AGEMA_signal_833), .Q (new_AGEMA_signal_834) ) ;
    buf_clk new_AGEMA_reg_buffer_367 ( .C (clk), .D (new_AGEMA_signal_839), .Q (new_AGEMA_signal_840) ) ;
    buf_clk new_AGEMA_reg_buffer_373 ( .C (clk), .D (new_AGEMA_signal_845), .Q (new_AGEMA_signal_846) ) ;
    buf_clk new_AGEMA_reg_buffer_379 ( .C (clk), .D (new_AGEMA_signal_851), .Q (new_AGEMA_signal_852) ) ;
    buf_clk new_AGEMA_reg_buffer_385 ( .C (clk), .D (new_AGEMA_signal_857), .Q (new_AGEMA_signal_858) ) ;
    buf_clk new_AGEMA_reg_buffer_391 ( .C (clk), .D (new_AGEMA_signal_863), .Q (new_AGEMA_signal_864) ) ;
    buf_clk new_AGEMA_reg_buffer_397 ( .C (clk), .D (new_AGEMA_signal_869), .Q (new_AGEMA_signal_870) ) ;
    buf_clk new_AGEMA_reg_buffer_403 ( .C (clk), .D (new_AGEMA_signal_875), .Q (new_AGEMA_signal_876) ) ;
    buf_clk new_AGEMA_reg_buffer_409 ( .C (clk), .D (new_AGEMA_signal_881), .Q (new_AGEMA_signal_882) ) ;
    buf_clk new_AGEMA_reg_buffer_415 ( .C (clk), .D (new_AGEMA_signal_887), .Q (new_AGEMA_signal_888) ) ;
    buf_clk new_AGEMA_reg_buffer_421 ( .C (clk), .D (new_AGEMA_signal_893), .Q (new_AGEMA_signal_894) ) ;
    buf_clk new_AGEMA_reg_buffer_427 ( .C (clk), .D (new_AGEMA_signal_899), .Q (new_AGEMA_signal_900) ) ;
    buf_clk new_AGEMA_reg_buffer_433 ( .C (clk), .D (new_AGEMA_signal_905), .Q (new_AGEMA_signal_906) ) ;
    buf_clk new_AGEMA_reg_buffer_439 ( .C (clk), .D (new_AGEMA_signal_911), .Q (new_AGEMA_signal_912) ) ;
    buf_clk new_AGEMA_reg_buffer_445 ( .C (clk), .D (new_AGEMA_signal_917), .Q (new_AGEMA_signal_918) ) ;
    buf_clk new_AGEMA_reg_buffer_451 ( .C (clk), .D (new_AGEMA_signal_923), .Q (new_AGEMA_signal_924) ) ;
    buf_clk new_AGEMA_reg_buffer_457 ( .C (clk), .D (new_AGEMA_signal_929), .Q (new_AGEMA_signal_930) ) ;
    buf_clk new_AGEMA_reg_buffer_463 ( .C (clk), .D (new_AGEMA_signal_935), .Q (new_AGEMA_signal_936) ) ;
    buf_clk new_AGEMA_reg_buffer_469 ( .C (clk), .D (new_AGEMA_signal_941), .Q (new_AGEMA_signal_942) ) ;
    buf_clk new_AGEMA_reg_buffer_475 ( .C (clk), .D (new_AGEMA_signal_947), .Q (new_AGEMA_signal_948) ) ;
    buf_clk new_AGEMA_reg_buffer_481 ( .C (clk), .D (new_AGEMA_signal_953), .Q (new_AGEMA_signal_954) ) ;
    buf_clk new_AGEMA_reg_buffer_487 ( .C (clk), .D (new_AGEMA_signal_959), .Q (new_AGEMA_signal_960) ) ;
    buf_clk new_AGEMA_reg_buffer_493 ( .C (clk), .D (new_AGEMA_signal_965), .Q (new_AGEMA_signal_966) ) ;
    buf_clk new_AGEMA_reg_buffer_499 ( .C (clk), .D (new_AGEMA_signal_971), .Q (new_AGEMA_signal_972) ) ;
    buf_clk new_AGEMA_reg_buffer_505 ( .C (clk), .D (new_AGEMA_signal_977), .Q (new_AGEMA_signal_978) ) ;
    buf_clk new_AGEMA_reg_buffer_511 ( .C (clk), .D (new_AGEMA_signal_983), .Q (new_AGEMA_signal_984) ) ;
    buf_clk new_AGEMA_reg_buffer_517 ( .C (clk), .D (new_AGEMA_signal_989), .Q (new_AGEMA_signal_990) ) ;
    buf_clk new_AGEMA_reg_buffer_523 ( .C (clk), .D (new_AGEMA_signal_995), .Q (new_AGEMA_signal_996) ) ;
    buf_clk new_AGEMA_reg_buffer_529 ( .C (clk), .D (new_AGEMA_signal_1001), .Q (new_AGEMA_signal_1002) ) ;

    /* cells in depth 5 */
    buf_clk new_AGEMA_reg_buffer_184 ( .C (clk), .D (new_AGEMA_signal_634), .Q (new_AGEMA_signal_657) ) ;
    buf_clk new_AGEMA_reg_buffer_186 ( .C (clk), .D (new_AGEMA_signal_636), .Q (new_AGEMA_signal_659) ) ;
    buf_clk new_AGEMA_reg_buffer_188 ( .C (clk), .D (new_AGEMA_signal_638), .Q (new_AGEMA_signal_661) ) ;
    buf_clk new_AGEMA_reg_buffer_190 ( .C (clk), .D (M33), .Q (new_AGEMA_signal_663) ) ;
    buf_clk new_AGEMA_reg_buffer_192 ( .C (clk), .D (new_AGEMA_signal_281), .Q (new_AGEMA_signal_665) ) ;
    buf_clk new_AGEMA_reg_buffer_194 ( .C (clk), .D (new_AGEMA_signal_282), .Q (new_AGEMA_signal_667) ) ;
    buf_clk new_AGEMA_reg_buffer_196 ( .C (clk), .D (new_AGEMA_signal_640), .Q (new_AGEMA_signal_669) ) ;
    buf_clk new_AGEMA_reg_buffer_198 ( .C (clk), .D (new_AGEMA_signal_642), .Q (new_AGEMA_signal_671) ) ;
    buf_clk new_AGEMA_reg_buffer_200 ( .C (clk), .D (new_AGEMA_signal_644), .Q (new_AGEMA_signal_673) ) ;
    buf_clk new_AGEMA_reg_buffer_202 ( .C (clk), .D (M36), .Q (new_AGEMA_signal_675) ) ;
    buf_clk new_AGEMA_reg_buffer_204 ( .C (clk), .D (new_AGEMA_signal_291), .Q (new_AGEMA_signal_677) ) ;
    buf_clk new_AGEMA_reg_buffer_206 ( .C (clk), .D (new_AGEMA_signal_292), .Q (new_AGEMA_signal_679) ) ;
    buf_clk new_AGEMA_reg_buffer_212 ( .C (clk), .D (new_AGEMA_signal_684), .Q (new_AGEMA_signal_685) ) ;
    buf_clk new_AGEMA_reg_buffer_218 ( .C (clk), .D (new_AGEMA_signal_690), .Q (new_AGEMA_signal_691) ) ;
    buf_clk new_AGEMA_reg_buffer_224 ( .C (clk), .D (new_AGEMA_signal_696), .Q (new_AGEMA_signal_697) ) ;
    buf_clk new_AGEMA_reg_buffer_230 ( .C (clk), .D (new_AGEMA_signal_702), .Q (new_AGEMA_signal_703) ) ;
    buf_clk new_AGEMA_reg_buffer_236 ( .C (clk), .D (new_AGEMA_signal_708), .Q (new_AGEMA_signal_709) ) ;
    buf_clk new_AGEMA_reg_buffer_242 ( .C (clk), .D (new_AGEMA_signal_714), .Q (new_AGEMA_signal_715) ) ;
    buf_clk new_AGEMA_reg_buffer_248 ( .C (clk), .D (new_AGEMA_signal_720), .Q (new_AGEMA_signal_721) ) ;
    buf_clk new_AGEMA_reg_buffer_254 ( .C (clk), .D (new_AGEMA_signal_726), .Q (new_AGEMA_signal_727) ) ;
    buf_clk new_AGEMA_reg_buffer_260 ( .C (clk), .D (new_AGEMA_signal_732), .Q (new_AGEMA_signal_733) ) ;
    buf_clk new_AGEMA_reg_buffer_266 ( .C (clk), .D (new_AGEMA_signal_738), .Q (new_AGEMA_signal_739) ) ;
    buf_clk new_AGEMA_reg_buffer_272 ( .C (clk), .D (new_AGEMA_signal_744), .Q (new_AGEMA_signal_745) ) ;
    buf_clk new_AGEMA_reg_buffer_278 ( .C (clk), .D (new_AGEMA_signal_750), .Q (new_AGEMA_signal_751) ) ;
    buf_clk new_AGEMA_reg_buffer_284 ( .C (clk), .D (new_AGEMA_signal_756), .Q (new_AGEMA_signal_757) ) ;
    buf_clk new_AGEMA_reg_buffer_290 ( .C (clk), .D (new_AGEMA_signal_762), .Q (new_AGEMA_signal_763) ) ;
    buf_clk new_AGEMA_reg_buffer_296 ( .C (clk), .D (new_AGEMA_signal_768), .Q (new_AGEMA_signal_769) ) ;
    buf_clk new_AGEMA_reg_buffer_302 ( .C (clk), .D (new_AGEMA_signal_774), .Q (new_AGEMA_signal_775) ) ;
    buf_clk new_AGEMA_reg_buffer_308 ( .C (clk), .D (new_AGEMA_signal_780), .Q (new_AGEMA_signal_781) ) ;
    buf_clk new_AGEMA_reg_buffer_314 ( .C (clk), .D (new_AGEMA_signal_786), .Q (new_AGEMA_signal_787) ) ;
    buf_clk new_AGEMA_reg_buffer_320 ( .C (clk), .D (new_AGEMA_signal_792), .Q (new_AGEMA_signal_793) ) ;
    buf_clk new_AGEMA_reg_buffer_326 ( .C (clk), .D (new_AGEMA_signal_798), .Q (new_AGEMA_signal_799) ) ;
    buf_clk new_AGEMA_reg_buffer_332 ( .C (clk), .D (new_AGEMA_signal_804), .Q (new_AGEMA_signal_805) ) ;
    buf_clk new_AGEMA_reg_buffer_338 ( .C (clk), .D (new_AGEMA_signal_810), .Q (new_AGEMA_signal_811) ) ;
    buf_clk new_AGEMA_reg_buffer_344 ( .C (clk), .D (new_AGEMA_signal_816), .Q (new_AGEMA_signal_817) ) ;
    buf_clk new_AGEMA_reg_buffer_350 ( .C (clk), .D (new_AGEMA_signal_822), .Q (new_AGEMA_signal_823) ) ;
    buf_clk new_AGEMA_reg_buffer_356 ( .C (clk), .D (new_AGEMA_signal_828), .Q (new_AGEMA_signal_829) ) ;
    buf_clk new_AGEMA_reg_buffer_362 ( .C (clk), .D (new_AGEMA_signal_834), .Q (new_AGEMA_signal_835) ) ;
    buf_clk new_AGEMA_reg_buffer_368 ( .C (clk), .D (new_AGEMA_signal_840), .Q (new_AGEMA_signal_841) ) ;
    buf_clk new_AGEMA_reg_buffer_374 ( .C (clk), .D (new_AGEMA_signal_846), .Q (new_AGEMA_signal_847) ) ;
    buf_clk new_AGEMA_reg_buffer_380 ( .C (clk), .D (new_AGEMA_signal_852), .Q (new_AGEMA_signal_853) ) ;
    buf_clk new_AGEMA_reg_buffer_386 ( .C (clk), .D (new_AGEMA_signal_858), .Q (new_AGEMA_signal_859) ) ;
    buf_clk new_AGEMA_reg_buffer_392 ( .C (clk), .D (new_AGEMA_signal_864), .Q (new_AGEMA_signal_865) ) ;
    buf_clk new_AGEMA_reg_buffer_398 ( .C (clk), .D (new_AGEMA_signal_870), .Q (new_AGEMA_signal_871) ) ;
    buf_clk new_AGEMA_reg_buffer_404 ( .C (clk), .D (new_AGEMA_signal_876), .Q (new_AGEMA_signal_877) ) ;
    buf_clk new_AGEMA_reg_buffer_410 ( .C (clk), .D (new_AGEMA_signal_882), .Q (new_AGEMA_signal_883) ) ;
    buf_clk new_AGEMA_reg_buffer_416 ( .C (clk), .D (new_AGEMA_signal_888), .Q (new_AGEMA_signal_889) ) ;
    buf_clk new_AGEMA_reg_buffer_422 ( .C (clk), .D (new_AGEMA_signal_894), .Q (new_AGEMA_signal_895) ) ;
    buf_clk new_AGEMA_reg_buffer_428 ( .C (clk), .D (new_AGEMA_signal_900), .Q (new_AGEMA_signal_901) ) ;
    buf_clk new_AGEMA_reg_buffer_434 ( .C (clk), .D (new_AGEMA_signal_906), .Q (new_AGEMA_signal_907) ) ;
    buf_clk new_AGEMA_reg_buffer_440 ( .C (clk), .D (new_AGEMA_signal_912), .Q (new_AGEMA_signal_913) ) ;
    buf_clk new_AGEMA_reg_buffer_446 ( .C (clk), .D (new_AGEMA_signal_918), .Q (new_AGEMA_signal_919) ) ;
    buf_clk new_AGEMA_reg_buffer_452 ( .C (clk), .D (new_AGEMA_signal_924), .Q (new_AGEMA_signal_925) ) ;
    buf_clk new_AGEMA_reg_buffer_458 ( .C (clk), .D (new_AGEMA_signal_930), .Q (new_AGEMA_signal_931) ) ;
    buf_clk new_AGEMA_reg_buffer_464 ( .C (clk), .D (new_AGEMA_signal_936), .Q (new_AGEMA_signal_937) ) ;
    buf_clk new_AGEMA_reg_buffer_470 ( .C (clk), .D (new_AGEMA_signal_942), .Q (new_AGEMA_signal_943) ) ;
    buf_clk new_AGEMA_reg_buffer_476 ( .C (clk), .D (new_AGEMA_signal_948), .Q (new_AGEMA_signal_949) ) ;
    buf_clk new_AGEMA_reg_buffer_482 ( .C (clk), .D (new_AGEMA_signal_954), .Q (new_AGEMA_signal_955) ) ;
    buf_clk new_AGEMA_reg_buffer_488 ( .C (clk), .D (new_AGEMA_signal_960), .Q (new_AGEMA_signal_961) ) ;
    buf_clk new_AGEMA_reg_buffer_494 ( .C (clk), .D (new_AGEMA_signal_966), .Q (new_AGEMA_signal_967) ) ;
    buf_clk new_AGEMA_reg_buffer_500 ( .C (clk), .D (new_AGEMA_signal_972), .Q (new_AGEMA_signal_973) ) ;
    buf_clk new_AGEMA_reg_buffer_506 ( .C (clk), .D (new_AGEMA_signal_978), .Q (new_AGEMA_signal_979) ) ;
    buf_clk new_AGEMA_reg_buffer_512 ( .C (clk), .D (new_AGEMA_signal_984), .Q (new_AGEMA_signal_985) ) ;
    buf_clk new_AGEMA_reg_buffer_518 ( .C (clk), .D (new_AGEMA_signal_990), .Q (new_AGEMA_signal_991) ) ;
    buf_clk new_AGEMA_reg_buffer_524 ( .C (clk), .D (new_AGEMA_signal_996), .Q (new_AGEMA_signal_997) ) ;
    buf_clk new_AGEMA_reg_buffer_530 ( .C (clk), .D (new_AGEMA_signal_1002), .Q (new_AGEMA_signal_1003) ) ;

    /* cells in depth 6 */
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M29_U1 ( .ina ({new_AGEMA_signal_278, new_AGEMA_signal_277, M28}), .inb ({new_AGEMA_signal_650, new_AGEMA_signal_648, new_AGEMA_signal_646}), .clk (clk), .rnd ({Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .outt ({new_AGEMA_signal_284, new_AGEMA_signal_283, M29}) ) ;
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M30_U1 ( .ina ({new_AGEMA_signal_276, new_AGEMA_signal_275, M26}), .inb ({new_AGEMA_signal_656, new_AGEMA_signal_654, new_AGEMA_signal_652}), .clk (clk), .rnd ({Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65]}), .outt ({new_AGEMA_signal_286, new_AGEMA_signal_285, M30}) ) ;
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M32_U1 ( .ina ({new_AGEMA_signal_650, new_AGEMA_signal_648, new_AGEMA_signal_646}), .inb ({new_AGEMA_signal_280, new_AGEMA_signal_279, M31}), .clk (clk), .rnd ({Fresh[74], Fresh[73], Fresh[72], Fresh[71], Fresh[70]}), .outt ({new_AGEMA_signal_288, new_AGEMA_signal_287, M32}) ) ;
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M35_U1 ( .ina ({new_AGEMA_signal_656, new_AGEMA_signal_654, new_AGEMA_signal_652}), .inb ({new_AGEMA_signal_272, new_AGEMA_signal_271, M34}), .clk (clk), .rnd ({Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75]}), .outt ({new_AGEMA_signal_290, new_AGEMA_signal_289, M35}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_M37_U1 ( .a ({new_AGEMA_signal_662, new_AGEMA_signal_660, new_AGEMA_signal_658}), .b ({new_AGEMA_signal_284, new_AGEMA_signal_283, M29}), .c ({new_AGEMA_signal_294, new_AGEMA_signal_293, M37}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_M38_U1 ( .a ({new_AGEMA_signal_288, new_AGEMA_signal_287, M32}), .b ({new_AGEMA_signal_668, new_AGEMA_signal_666, new_AGEMA_signal_664}), .c ({new_AGEMA_signal_296, new_AGEMA_signal_295, M38}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_M39_U1 ( .a ({new_AGEMA_signal_674, new_AGEMA_signal_672, new_AGEMA_signal_670}), .b ({new_AGEMA_signal_286, new_AGEMA_signal_285, M30}), .c ({new_AGEMA_signal_298, new_AGEMA_signal_297, M39}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_M40_U1 ( .a ({new_AGEMA_signal_290, new_AGEMA_signal_289, M35}), .b ({new_AGEMA_signal_680, new_AGEMA_signal_678, new_AGEMA_signal_676}), .c ({new_AGEMA_signal_300, new_AGEMA_signal_299, M40}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_M41_U1 ( .a ({new_AGEMA_signal_296, new_AGEMA_signal_295, M38}), .b ({new_AGEMA_signal_300, new_AGEMA_signal_299, M40}), .c ({new_AGEMA_signal_302, new_AGEMA_signal_301, M41}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_M42_U1 ( .a ({new_AGEMA_signal_294, new_AGEMA_signal_293, M37}), .b ({new_AGEMA_signal_298, new_AGEMA_signal_297, M39}), .c ({new_AGEMA_signal_304, new_AGEMA_signal_303, M42}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_M43_U1 ( .a ({new_AGEMA_signal_294, new_AGEMA_signal_293, M37}), .b ({new_AGEMA_signal_296, new_AGEMA_signal_295, M38}), .c ({new_AGEMA_signal_306, new_AGEMA_signal_305, M43}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_M44_U1 ( .a ({new_AGEMA_signal_298, new_AGEMA_signal_297, M39}), .b ({new_AGEMA_signal_300, new_AGEMA_signal_299, M40}), .c ({new_AGEMA_signal_308, new_AGEMA_signal_307, M44}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_M45_U1 ( .a ({new_AGEMA_signal_304, new_AGEMA_signal_303, M42}), .b ({new_AGEMA_signal_302, new_AGEMA_signal_301, M41}), .c ({new_AGEMA_signal_326, new_AGEMA_signal_325, M45}) ) ;
    buf_clk new_AGEMA_reg_buffer_185 ( .C (clk), .D (new_AGEMA_signal_657), .Q (new_AGEMA_signal_658) ) ;
    buf_clk new_AGEMA_reg_buffer_187 ( .C (clk), .D (new_AGEMA_signal_659), .Q (new_AGEMA_signal_660) ) ;
    buf_clk new_AGEMA_reg_buffer_189 ( .C (clk), .D (new_AGEMA_signal_661), .Q (new_AGEMA_signal_662) ) ;
    buf_clk new_AGEMA_reg_buffer_191 ( .C (clk), .D (new_AGEMA_signal_663), .Q (new_AGEMA_signal_664) ) ;
    buf_clk new_AGEMA_reg_buffer_193 ( .C (clk), .D (new_AGEMA_signal_665), .Q (new_AGEMA_signal_666) ) ;
    buf_clk new_AGEMA_reg_buffer_195 ( .C (clk), .D (new_AGEMA_signal_667), .Q (new_AGEMA_signal_668) ) ;
    buf_clk new_AGEMA_reg_buffer_197 ( .C (clk), .D (new_AGEMA_signal_669), .Q (new_AGEMA_signal_670) ) ;
    buf_clk new_AGEMA_reg_buffer_199 ( .C (clk), .D (new_AGEMA_signal_671), .Q (new_AGEMA_signal_672) ) ;
    buf_clk new_AGEMA_reg_buffer_201 ( .C (clk), .D (new_AGEMA_signal_673), .Q (new_AGEMA_signal_674) ) ;
    buf_clk new_AGEMA_reg_buffer_203 ( .C (clk), .D (new_AGEMA_signal_675), .Q (new_AGEMA_signal_676) ) ;
    buf_clk new_AGEMA_reg_buffer_205 ( .C (clk), .D (new_AGEMA_signal_677), .Q (new_AGEMA_signal_678) ) ;
    buf_clk new_AGEMA_reg_buffer_207 ( .C (clk), .D (new_AGEMA_signal_679), .Q (new_AGEMA_signal_680) ) ;
    buf_clk new_AGEMA_reg_buffer_213 ( .C (clk), .D (new_AGEMA_signal_685), .Q (new_AGEMA_signal_686) ) ;
    buf_clk new_AGEMA_reg_buffer_219 ( .C (clk), .D (new_AGEMA_signal_691), .Q (new_AGEMA_signal_692) ) ;
    buf_clk new_AGEMA_reg_buffer_225 ( .C (clk), .D (new_AGEMA_signal_697), .Q (new_AGEMA_signal_698) ) ;
    buf_clk new_AGEMA_reg_buffer_231 ( .C (clk), .D (new_AGEMA_signal_703), .Q (new_AGEMA_signal_704) ) ;
    buf_clk new_AGEMA_reg_buffer_237 ( .C (clk), .D (new_AGEMA_signal_709), .Q (new_AGEMA_signal_710) ) ;
    buf_clk new_AGEMA_reg_buffer_243 ( .C (clk), .D (new_AGEMA_signal_715), .Q (new_AGEMA_signal_716) ) ;
    buf_clk new_AGEMA_reg_buffer_249 ( .C (clk), .D (new_AGEMA_signal_721), .Q (new_AGEMA_signal_722) ) ;
    buf_clk new_AGEMA_reg_buffer_255 ( .C (clk), .D (new_AGEMA_signal_727), .Q (new_AGEMA_signal_728) ) ;
    buf_clk new_AGEMA_reg_buffer_261 ( .C (clk), .D (new_AGEMA_signal_733), .Q (new_AGEMA_signal_734) ) ;
    buf_clk new_AGEMA_reg_buffer_267 ( .C (clk), .D (new_AGEMA_signal_739), .Q (new_AGEMA_signal_740) ) ;
    buf_clk new_AGEMA_reg_buffer_273 ( .C (clk), .D (new_AGEMA_signal_745), .Q (new_AGEMA_signal_746) ) ;
    buf_clk new_AGEMA_reg_buffer_279 ( .C (clk), .D (new_AGEMA_signal_751), .Q (new_AGEMA_signal_752) ) ;
    buf_clk new_AGEMA_reg_buffer_285 ( .C (clk), .D (new_AGEMA_signal_757), .Q (new_AGEMA_signal_758) ) ;
    buf_clk new_AGEMA_reg_buffer_291 ( .C (clk), .D (new_AGEMA_signal_763), .Q (new_AGEMA_signal_764) ) ;
    buf_clk new_AGEMA_reg_buffer_297 ( .C (clk), .D (new_AGEMA_signal_769), .Q (new_AGEMA_signal_770) ) ;
    buf_clk new_AGEMA_reg_buffer_303 ( .C (clk), .D (new_AGEMA_signal_775), .Q (new_AGEMA_signal_776) ) ;
    buf_clk new_AGEMA_reg_buffer_309 ( .C (clk), .D (new_AGEMA_signal_781), .Q (new_AGEMA_signal_782) ) ;
    buf_clk new_AGEMA_reg_buffer_315 ( .C (clk), .D (new_AGEMA_signal_787), .Q (new_AGEMA_signal_788) ) ;
    buf_clk new_AGEMA_reg_buffer_321 ( .C (clk), .D (new_AGEMA_signal_793), .Q (new_AGEMA_signal_794) ) ;
    buf_clk new_AGEMA_reg_buffer_327 ( .C (clk), .D (new_AGEMA_signal_799), .Q (new_AGEMA_signal_800) ) ;
    buf_clk new_AGEMA_reg_buffer_333 ( .C (clk), .D (new_AGEMA_signal_805), .Q (new_AGEMA_signal_806) ) ;
    buf_clk new_AGEMA_reg_buffer_339 ( .C (clk), .D (new_AGEMA_signal_811), .Q (new_AGEMA_signal_812) ) ;
    buf_clk new_AGEMA_reg_buffer_345 ( .C (clk), .D (new_AGEMA_signal_817), .Q (new_AGEMA_signal_818) ) ;
    buf_clk new_AGEMA_reg_buffer_351 ( .C (clk), .D (new_AGEMA_signal_823), .Q (new_AGEMA_signal_824) ) ;
    buf_clk new_AGEMA_reg_buffer_357 ( .C (clk), .D (new_AGEMA_signal_829), .Q (new_AGEMA_signal_830) ) ;
    buf_clk new_AGEMA_reg_buffer_363 ( .C (clk), .D (new_AGEMA_signal_835), .Q (new_AGEMA_signal_836) ) ;
    buf_clk new_AGEMA_reg_buffer_369 ( .C (clk), .D (new_AGEMA_signal_841), .Q (new_AGEMA_signal_842) ) ;
    buf_clk new_AGEMA_reg_buffer_375 ( .C (clk), .D (new_AGEMA_signal_847), .Q (new_AGEMA_signal_848) ) ;
    buf_clk new_AGEMA_reg_buffer_381 ( .C (clk), .D (new_AGEMA_signal_853), .Q (new_AGEMA_signal_854) ) ;
    buf_clk new_AGEMA_reg_buffer_387 ( .C (clk), .D (new_AGEMA_signal_859), .Q (new_AGEMA_signal_860) ) ;
    buf_clk new_AGEMA_reg_buffer_393 ( .C (clk), .D (new_AGEMA_signal_865), .Q (new_AGEMA_signal_866) ) ;
    buf_clk new_AGEMA_reg_buffer_399 ( .C (clk), .D (new_AGEMA_signal_871), .Q (new_AGEMA_signal_872) ) ;
    buf_clk new_AGEMA_reg_buffer_405 ( .C (clk), .D (new_AGEMA_signal_877), .Q (new_AGEMA_signal_878) ) ;
    buf_clk new_AGEMA_reg_buffer_411 ( .C (clk), .D (new_AGEMA_signal_883), .Q (new_AGEMA_signal_884) ) ;
    buf_clk new_AGEMA_reg_buffer_417 ( .C (clk), .D (new_AGEMA_signal_889), .Q (new_AGEMA_signal_890) ) ;
    buf_clk new_AGEMA_reg_buffer_423 ( .C (clk), .D (new_AGEMA_signal_895), .Q (new_AGEMA_signal_896) ) ;
    buf_clk new_AGEMA_reg_buffer_429 ( .C (clk), .D (new_AGEMA_signal_901), .Q (new_AGEMA_signal_902) ) ;
    buf_clk new_AGEMA_reg_buffer_435 ( .C (clk), .D (new_AGEMA_signal_907), .Q (new_AGEMA_signal_908) ) ;
    buf_clk new_AGEMA_reg_buffer_441 ( .C (clk), .D (new_AGEMA_signal_913), .Q (new_AGEMA_signal_914) ) ;
    buf_clk new_AGEMA_reg_buffer_447 ( .C (clk), .D (new_AGEMA_signal_919), .Q (new_AGEMA_signal_920) ) ;
    buf_clk new_AGEMA_reg_buffer_453 ( .C (clk), .D (new_AGEMA_signal_925), .Q (new_AGEMA_signal_926) ) ;
    buf_clk new_AGEMA_reg_buffer_459 ( .C (clk), .D (new_AGEMA_signal_931), .Q (new_AGEMA_signal_932) ) ;
    buf_clk new_AGEMA_reg_buffer_465 ( .C (clk), .D (new_AGEMA_signal_937), .Q (new_AGEMA_signal_938) ) ;
    buf_clk new_AGEMA_reg_buffer_471 ( .C (clk), .D (new_AGEMA_signal_943), .Q (new_AGEMA_signal_944) ) ;
    buf_clk new_AGEMA_reg_buffer_477 ( .C (clk), .D (new_AGEMA_signal_949), .Q (new_AGEMA_signal_950) ) ;
    buf_clk new_AGEMA_reg_buffer_483 ( .C (clk), .D (new_AGEMA_signal_955), .Q (new_AGEMA_signal_956) ) ;
    buf_clk new_AGEMA_reg_buffer_489 ( .C (clk), .D (new_AGEMA_signal_961), .Q (new_AGEMA_signal_962) ) ;
    buf_clk new_AGEMA_reg_buffer_495 ( .C (clk), .D (new_AGEMA_signal_967), .Q (new_AGEMA_signal_968) ) ;
    buf_clk new_AGEMA_reg_buffer_501 ( .C (clk), .D (new_AGEMA_signal_973), .Q (new_AGEMA_signal_974) ) ;
    buf_clk new_AGEMA_reg_buffer_507 ( .C (clk), .D (new_AGEMA_signal_979), .Q (new_AGEMA_signal_980) ) ;
    buf_clk new_AGEMA_reg_buffer_513 ( .C (clk), .D (new_AGEMA_signal_985), .Q (new_AGEMA_signal_986) ) ;
    buf_clk new_AGEMA_reg_buffer_519 ( .C (clk), .D (new_AGEMA_signal_991), .Q (new_AGEMA_signal_992) ) ;
    buf_clk new_AGEMA_reg_buffer_525 ( .C (clk), .D (new_AGEMA_signal_997), .Q (new_AGEMA_signal_998) ) ;
    buf_clk new_AGEMA_reg_buffer_531 ( .C (clk), .D (new_AGEMA_signal_1003), .Q (new_AGEMA_signal_1004) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M46_U1 ( .ina ({new_AGEMA_signal_308, new_AGEMA_signal_307, M44}), .inb ({new_AGEMA_signal_698, new_AGEMA_signal_692, new_AGEMA_signal_686}), .clk (clk), .rnd ({Fresh[84], Fresh[83], Fresh[82], Fresh[81], Fresh[80]}), .outt ({new_AGEMA_signal_328, new_AGEMA_signal_327, M46}) ) ;
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M47_U1 ( .ina ({new_AGEMA_signal_300, new_AGEMA_signal_299, M40}), .inb ({new_AGEMA_signal_716, new_AGEMA_signal_710, new_AGEMA_signal_704}), .clk (clk), .rnd ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85]}), .outt ({new_AGEMA_signal_310, new_AGEMA_signal_309, M47}) ) ;
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M48_U1 ( .ina ({new_AGEMA_signal_298, new_AGEMA_signal_297, M39}), .inb ({new_AGEMA_signal_734, new_AGEMA_signal_728, new_AGEMA_signal_722}), .clk (clk), .rnd ({Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .outt ({new_AGEMA_signal_312, new_AGEMA_signal_311, M48}) ) ;
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M49_U1 ( .ina ({new_AGEMA_signal_306, new_AGEMA_signal_305, M43}), .inb ({new_AGEMA_signal_752, new_AGEMA_signal_746, new_AGEMA_signal_740}), .clk (clk), .rnd ({Fresh[99], Fresh[98], Fresh[97], Fresh[96], Fresh[95]}), .outt ({new_AGEMA_signal_330, new_AGEMA_signal_329, M49}) ) ;
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M50_U1 ( .ina ({new_AGEMA_signal_296, new_AGEMA_signal_295, M38}), .inb ({new_AGEMA_signal_770, new_AGEMA_signal_764, new_AGEMA_signal_758}), .clk (clk), .rnd ({Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100]}), .outt ({new_AGEMA_signal_314, new_AGEMA_signal_313, M50}) ) ;
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M51_U1 ( .ina ({new_AGEMA_signal_294, new_AGEMA_signal_293, M37}), .inb ({new_AGEMA_signal_788, new_AGEMA_signal_782, new_AGEMA_signal_776}), .clk (clk), .rnd ({Fresh[109], Fresh[108], Fresh[107], Fresh[106], Fresh[105]}), .outt ({new_AGEMA_signal_316, new_AGEMA_signal_315, M51}) ) ;
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M52_U1 ( .ina ({new_AGEMA_signal_304, new_AGEMA_signal_303, M42}), .inb ({new_AGEMA_signal_806, new_AGEMA_signal_800, new_AGEMA_signal_794}), .clk (clk), .rnd ({Fresh[114], Fresh[113], Fresh[112], Fresh[111], Fresh[110]}), .outt ({new_AGEMA_signal_332, new_AGEMA_signal_331, M52}) ) ;
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M53_U1 ( .ina ({new_AGEMA_signal_326, new_AGEMA_signal_325, M45}), .inb ({new_AGEMA_signal_824, new_AGEMA_signal_818, new_AGEMA_signal_812}), .clk (clk), .rnd ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115]}), .outt ({new_AGEMA_signal_350, new_AGEMA_signal_349, M53}) ) ;
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M54_U1 ( .ina ({new_AGEMA_signal_302, new_AGEMA_signal_301, M41}), .inb ({new_AGEMA_signal_842, new_AGEMA_signal_836, new_AGEMA_signal_830}), .clk (clk), .rnd ({Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .outt ({new_AGEMA_signal_334, new_AGEMA_signal_333, M54}) ) ;
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M55_U1 ( .ina ({new_AGEMA_signal_308, new_AGEMA_signal_307, M44}), .inb ({new_AGEMA_signal_860, new_AGEMA_signal_854, new_AGEMA_signal_848}), .clk (clk), .rnd ({Fresh[129], Fresh[128], Fresh[127], Fresh[126], Fresh[125]}), .outt ({new_AGEMA_signal_336, new_AGEMA_signal_335, M55}) ) ;
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M56_U1 ( .ina ({new_AGEMA_signal_300, new_AGEMA_signal_299, M40}), .inb ({new_AGEMA_signal_878, new_AGEMA_signal_872, new_AGEMA_signal_866}), .clk (clk), .rnd ({Fresh[134], Fresh[133], Fresh[132], Fresh[131], Fresh[130]}), .outt ({new_AGEMA_signal_318, new_AGEMA_signal_317, M56}) ) ;
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M57_U1 ( .ina ({new_AGEMA_signal_298, new_AGEMA_signal_297, M39}), .inb ({new_AGEMA_signal_896, new_AGEMA_signal_890, new_AGEMA_signal_884}), .clk (clk), .rnd ({Fresh[139], Fresh[138], Fresh[137], Fresh[136], Fresh[135]}), .outt ({new_AGEMA_signal_320, new_AGEMA_signal_319, M57}) ) ;
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M58_U1 ( .ina ({new_AGEMA_signal_306, new_AGEMA_signal_305, M43}), .inb ({new_AGEMA_signal_914, new_AGEMA_signal_908, new_AGEMA_signal_902}), .clk (clk), .rnd ({Fresh[144], Fresh[143], Fresh[142], Fresh[141], Fresh[140]}), .outt ({new_AGEMA_signal_338, new_AGEMA_signal_337, M58}) ) ;
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M59_U1 ( .ina ({new_AGEMA_signal_296, new_AGEMA_signal_295, M38}), .inb ({new_AGEMA_signal_932, new_AGEMA_signal_926, new_AGEMA_signal_920}), .clk (clk), .rnd ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145]}), .outt ({new_AGEMA_signal_322, new_AGEMA_signal_321, M59}) ) ;
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M60_U1 ( .ina ({new_AGEMA_signal_294, new_AGEMA_signal_293, M37}), .inb ({new_AGEMA_signal_950, new_AGEMA_signal_944, new_AGEMA_signal_938}), .clk (clk), .rnd ({Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .outt ({new_AGEMA_signal_324, new_AGEMA_signal_323, M60}) ) ;
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M61_U1 ( .ina ({new_AGEMA_signal_304, new_AGEMA_signal_303, M42}), .inb ({new_AGEMA_signal_968, new_AGEMA_signal_962, new_AGEMA_signal_956}), .clk (clk), .rnd ({Fresh[159], Fresh[158], Fresh[157], Fresh[156], Fresh[155]}), .outt ({new_AGEMA_signal_340, new_AGEMA_signal_339, M61}) ) ;
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M62_U1 ( .ina ({new_AGEMA_signal_326, new_AGEMA_signal_325, M45}), .inb ({new_AGEMA_signal_986, new_AGEMA_signal_980, new_AGEMA_signal_974}), .clk (clk), .rnd ({Fresh[164], Fresh[163], Fresh[162], Fresh[161], Fresh[160]}), .outt ({new_AGEMA_signal_352, new_AGEMA_signal_351, M62}) ) ;
    and_HPC1 #(.security_order(2), .pipeline(1)) AND_M63_U1 ( .ina ({new_AGEMA_signal_302, new_AGEMA_signal_301, M41}), .inb ({new_AGEMA_signal_1004, new_AGEMA_signal_998, new_AGEMA_signal_992}), .clk (clk), .rnd ({Fresh[169], Fresh[168], Fresh[167], Fresh[166], Fresh[165]}), .outt ({new_AGEMA_signal_342, new_AGEMA_signal_341, M63}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_L0_U1 ( .a ({new_AGEMA_signal_340, new_AGEMA_signal_339, M61}), .b ({new_AGEMA_signal_352, new_AGEMA_signal_351, M62}), .c ({new_AGEMA_signal_370, new_AGEMA_signal_369, L0}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_L1_U1 ( .a ({new_AGEMA_signal_314, new_AGEMA_signal_313, M50}), .b ({new_AGEMA_signal_318, new_AGEMA_signal_317, M56}), .c ({new_AGEMA_signal_344, new_AGEMA_signal_343, L1}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_L2_U1 ( .a ({new_AGEMA_signal_328, new_AGEMA_signal_327, M46}), .b ({new_AGEMA_signal_312, new_AGEMA_signal_311, M48}), .c ({new_AGEMA_signal_354, new_AGEMA_signal_353, L2}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_L3_U1 ( .a ({new_AGEMA_signal_310, new_AGEMA_signal_309, M47}), .b ({new_AGEMA_signal_336, new_AGEMA_signal_335, M55}), .c ({new_AGEMA_signal_356, new_AGEMA_signal_355, L3}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_L4_U1 ( .a ({new_AGEMA_signal_334, new_AGEMA_signal_333, M54}), .b ({new_AGEMA_signal_338, new_AGEMA_signal_337, M58}), .c ({new_AGEMA_signal_358, new_AGEMA_signal_357, L4}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_L5_U1 ( .a ({new_AGEMA_signal_330, new_AGEMA_signal_329, M49}), .b ({new_AGEMA_signal_340, new_AGEMA_signal_339, M61}), .c ({new_AGEMA_signal_360, new_AGEMA_signal_359, L5}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_L6_U1 ( .a ({new_AGEMA_signal_352, new_AGEMA_signal_351, M62}), .b ({new_AGEMA_signal_360, new_AGEMA_signal_359, L5}), .c ({new_AGEMA_signal_372, new_AGEMA_signal_371, L6}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_L7_U1 ( .a ({new_AGEMA_signal_328, new_AGEMA_signal_327, M46}), .b ({new_AGEMA_signal_356, new_AGEMA_signal_355, L3}), .c ({new_AGEMA_signal_374, new_AGEMA_signal_373, L7}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_L8_U1 ( .a ({new_AGEMA_signal_316, new_AGEMA_signal_315, M51}), .b ({new_AGEMA_signal_322, new_AGEMA_signal_321, M59}), .c ({new_AGEMA_signal_346, new_AGEMA_signal_345, L8}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_L9_U1 ( .a ({new_AGEMA_signal_332, new_AGEMA_signal_331, M52}), .b ({new_AGEMA_signal_350, new_AGEMA_signal_349, M53}), .c ({new_AGEMA_signal_376, new_AGEMA_signal_375, L9}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_L10_U1 ( .a ({new_AGEMA_signal_350, new_AGEMA_signal_349, M53}), .b ({new_AGEMA_signal_358, new_AGEMA_signal_357, L4}), .c ({new_AGEMA_signal_378, new_AGEMA_signal_377, L10}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_L11_U1 ( .a ({new_AGEMA_signal_324, new_AGEMA_signal_323, M60}), .b ({new_AGEMA_signal_354, new_AGEMA_signal_353, L2}), .c ({new_AGEMA_signal_380, new_AGEMA_signal_379, L11}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_L12_U1 ( .a ({new_AGEMA_signal_312, new_AGEMA_signal_311, M48}), .b ({new_AGEMA_signal_316, new_AGEMA_signal_315, M51}), .c ({new_AGEMA_signal_348, new_AGEMA_signal_347, L12}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_L13_U1 ( .a ({new_AGEMA_signal_314, new_AGEMA_signal_313, M50}), .b ({new_AGEMA_signal_370, new_AGEMA_signal_369, L0}), .c ({new_AGEMA_signal_388, new_AGEMA_signal_387, L13}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_L14_U1 ( .a ({new_AGEMA_signal_332, new_AGEMA_signal_331, M52}), .b ({new_AGEMA_signal_340, new_AGEMA_signal_339, M61}), .c ({new_AGEMA_signal_362, new_AGEMA_signal_361, L14}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_L15_U1 ( .a ({new_AGEMA_signal_336, new_AGEMA_signal_335, M55}), .b ({new_AGEMA_signal_344, new_AGEMA_signal_343, L1}), .c ({new_AGEMA_signal_364, new_AGEMA_signal_363, L15}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_L16_U1 ( .a ({new_AGEMA_signal_318, new_AGEMA_signal_317, M56}), .b ({new_AGEMA_signal_370, new_AGEMA_signal_369, L0}), .c ({new_AGEMA_signal_390, new_AGEMA_signal_389, L16}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_L17_U1 ( .a ({new_AGEMA_signal_320, new_AGEMA_signal_319, M57}), .b ({new_AGEMA_signal_344, new_AGEMA_signal_343, L1}), .c ({new_AGEMA_signal_366, new_AGEMA_signal_365, L17}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_L18_U1 ( .a ({new_AGEMA_signal_338, new_AGEMA_signal_337, M58}), .b ({new_AGEMA_signal_346, new_AGEMA_signal_345, L8}), .c ({new_AGEMA_signal_368, new_AGEMA_signal_367, L18}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_L19_U1 ( .a ({new_AGEMA_signal_342, new_AGEMA_signal_341, M63}), .b ({new_AGEMA_signal_358, new_AGEMA_signal_357, L4}), .c ({new_AGEMA_signal_382, new_AGEMA_signal_381, L19}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_L20_U1 ( .a ({new_AGEMA_signal_370, new_AGEMA_signal_369, L0}), .b ({new_AGEMA_signal_344, new_AGEMA_signal_343, L1}), .c ({new_AGEMA_signal_392, new_AGEMA_signal_391, L20}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_L21_U1 ( .a ({new_AGEMA_signal_344, new_AGEMA_signal_343, L1}), .b ({new_AGEMA_signal_374, new_AGEMA_signal_373, L7}), .c ({new_AGEMA_signal_394, new_AGEMA_signal_393, L21}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_L22_U1 ( .a ({new_AGEMA_signal_356, new_AGEMA_signal_355, L3}), .b ({new_AGEMA_signal_348, new_AGEMA_signal_347, L12}), .c ({new_AGEMA_signal_384, new_AGEMA_signal_383, L22}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_L23_U1 ( .a ({new_AGEMA_signal_368, new_AGEMA_signal_367, L18}), .b ({new_AGEMA_signal_354, new_AGEMA_signal_353, L2}), .c ({new_AGEMA_signal_386, new_AGEMA_signal_385, L23}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_L24_U1 ( .a ({new_AGEMA_signal_364, new_AGEMA_signal_363, L15}), .b ({new_AGEMA_signal_376, new_AGEMA_signal_375, L9}), .c ({new_AGEMA_signal_396, new_AGEMA_signal_395, L24}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_L25_U1 ( .a ({new_AGEMA_signal_372, new_AGEMA_signal_371, L6}), .b ({new_AGEMA_signal_378, new_AGEMA_signal_377, L10}), .c ({new_AGEMA_signal_398, new_AGEMA_signal_397, L25}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_L26_U1 ( .a ({new_AGEMA_signal_374, new_AGEMA_signal_373, L7}), .b ({new_AGEMA_signal_376, new_AGEMA_signal_375, L9}), .c ({new_AGEMA_signal_400, new_AGEMA_signal_399, L26}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_L27_U1 ( .a ({new_AGEMA_signal_346, new_AGEMA_signal_345, L8}), .b ({new_AGEMA_signal_378, new_AGEMA_signal_377, L10}), .c ({new_AGEMA_signal_402, new_AGEMA_signal_401, L27}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_L28_U1 ( .a ({new_AGEMA_signal_380, new_AGEMA_signal_379, L11}), .b ({new_AGEMA_signal_362, new_AGEMA_signal_361, L14}), .c ({new_AGEMA_signal_404, new_AGEMA_signal_403, L28}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_L29_U1 ( .a ({new_AGEMA_signal_380, new_AGEMA_signal_379, L11}), .b ({new_AGEMA_signal_366, new_AGEMA_signal_365, L17}), .c ({new_AGEMA_signal_406, new_AGEMA_signal_405, L29}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_S0_U1 ( .a ({new_AGEMA_signal_372, new_AGEMA_signal_371, L6}), .b ({new_AGEMA_signal_396, new_AGEMA_signal_395, L24}), .c ({new_AGEMA_signal_410, new_AGEMA_signal_409, O[7]}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) XOR_S1_U1 ( .a ({new_AGEMA_signal_390, new_AGEMA_signal_389, L16}), .b ({new_AGEMA_signal_400, new_AGEMA_signal_399, L26}), .c ({new_AGEMA_signal_412, new_AGEMA_signal_411, O[6]}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) XOR_S2_U1 ( .a ({new_AGEMA_signal_382, new_AGEMA_signal_381, L19}), .b ({new_AGEMA_signal_404, new_AGEMA_signal_403, L28}), .c ({new_AGEMA_signal_414, new_AGEMA_signal_413, O[5]}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_S3_U1 ( .a ({new_AGEMA_signal_372, new_AGEMA_signal_371, L6}), .b ({new_AGEMA_signal_394, new_AGEMA_signal_393, L21}), .c ({new_AGEMA_signal_416, new_AGEMA_signal_415, O[4]}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_S4_U1 ( .a ({new_AGEMA_signal_392, new_AGEMA_signal_391, L20}), .b ({new_AGEMA_signal_384, new_AGEMA_signal_383, L22}), .c ({new_AGEMA_signal_418, new_AGEMA_signal_417, O[3]}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) XOR_S5_U1 ( .a ({new_AGEMA_signal_398, new_AGEMA_signal_397, L25}), .b ({new_AGEMA_signal_406, new_AGEMA_signal_405, L29}), .c ({new_AGEMA_signal_420, new_AGEMA_signal_419, O[2]}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) XOR_S6_U1 ( .a ({new_AGEMA_signal_388, new_AGEMA_signal_387, L13}), .b ({new_AGEMA_signal_402, new_AGEMA_signal_401, L27}), .c ({new_AGEMA_signal_422, new_AGEMA_signal_421, O[1]}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) XOR_S7_U1 ( .a ({new_AGEMA_signal_372, new_AGEMA_signal_371, L6}), .b ({new_AGEMA_signal_386, new_AGEMA_signal_385, L23}), .c ({new_AGEMA_signal_408, new_AGEMA_signal_407, O[0]}) ) ;

    /* register cells */
    reg_masked #(.security_order(2), .pipeline(1)) Y_reg_7_ ( .clk (clk), .D ({new_AGEMA_signal_410, new_AGEMA_signal_409, O[7]}), .Q ({Y_s2[7], Y_s1[7], Y_s0[7]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Y_reg_6_ ( .clk (clk), .D ({new_AGEMA_signal_412, new_AGEMA_signal_411, O[6]}), .Q ({Y_s2[6], Y_s1[6], Y_s0[6]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Y_reg_5_ ( .clk (clk), .D ({new_AGEMA_signal_414, new_AGEMA_signal_413, O[5]}), .Q ({Y_s2[5], Y_s1[5], Y_s0[5]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Y_reg_4_ ( .clk (clk), .D ({new_AGEMA_signal_416, new_AGEMA_signal_415, O[4]}), .Q ({Y_s2[4], Y_s1[4], Y_s0[4]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Y_reg_3_ ( .clk (clk), .D ({new_AGEMA_signal_418, new_AGEMA_signal_417, O[3]}), .Q ({Y_s2[3], Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Y_reg_2_ ( .clk (clk), .D ({new_AGEMA_signal_420, new_AGEMA_signal_419, O[2]}), .Q ({Y_s2[2], Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Y_reg_1_ ( .clk (clk), .D ({new_AGEMA_signal_422, new_AGEMA_signal_421, O[1]}), .Q ({Y_s2[1], Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Y_reg_0_ ( .clk (clk), .D ({new_AGEMA_signal_408, new_AGEMA_signal_407, O[0]}), .Q ({Y_s2[0], Y_s1[0], Y_s0[0]}) ) ;
endmodule
