/* modified netlist. Source: module SkinnyTop in file Designs/Skinny64_64_round-based/AGEMA/SkinnyTop.v */
/* 2 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 3 register stage(s) in total */

module SkinnyTop_GHPC_ANF_Pipeline_d1 (Plaintext_s0, Key_s0, clk, rst, Key_s1, Plaintext_s1, Fresh, Ciphertext_s0, done, Ciphertext_s1);
    input [63:0] Plaintext_s0 ;
    input [63:0] Key_s0 ;
    input clk ;
    input rst ;
    input [63:0] Key_s1 ;
    input [63:0] Plaintext_s1 ;
    input [63:0] Fresh ;
    output [63:0] Ciphertext_s0 ;
    output done ;
    output [63:0] Ciphertext_s1 ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_768 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_771 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_774 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_777 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_780 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_783 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_786 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_789 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_792 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_809 ;
    wire signal_810 ;
    wire signal_811 ;
    wire signal_812 ;
    wire signal_813 ;
    wire signal_814 ;
    wire signal_815 ;
    wire signal_816 ;
    wire signal_817 ;
    wire signal_818 ;
    wire signal_819 ;
    wire signal_820 ;
    wire signal_821 ;
    wire signal_822 ;
    wire signal_823 ;
    wire signal_824 ;
    wire signal_825 ;
    wire signal_826 ;
    wire signal_827 ;
    wire signal_828 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_831 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_834 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_837 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_840 ;
    wire signal_841 ;
    wire signal_842 ;
    wire signal_843 ;
    wire signal_844 ;
    wire signal_845 ;
    wire signal_846 ;
    wire signal_847 ;
    wire signal_848 ;
    wire signal_849 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_852 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_855 ;
    wire signal_856 ;
    wire signal_857 ;
    wire signal_858 ;
    wire signal_859 ;
    wire signal_860 ;
    wire signal_861 ;
    wire signal_862 ;
    wire signal_863 ;
    wire signal_864 ;
    wire signal_865 ;
    wire signal_866 ;
    wire signal_867 ;
    wire signal_868 ;
    wire signal_869 ;
    wire signal_870 ;
    wire signal_871 ;
    wire signal_872 ;
    wire signal_873 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_879 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_885 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_888 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_891 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_894 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_897 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_900 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_903 ;
    wire signal_939 ;
    wire signal_940 ;
    wire signal_943 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1355 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1485 ;
    wire signal_1487 ;
    wire signal_1489 ;
    wire signal_1491 ;
    wire signal_1493 ;
    wire signal_1495 ;
    wire signal_1497 ;
    wire signal_1499 ;
    wire signal_1501 ;
    wire signal_1503 ;
    wire signal_1505 ;
    wire signal_1507 ;
    wire signal_1509 ;
    wire signal_1511 ;
    wire signal_1513 ;
    wire signal_1515 ;
    wire signal_1517 ;
    wire signal_1519 ;
    wire signal_1521 ;
    wire signal_1523 ;
    wire signal_1525 ;
    wire signal_1527 ;
    wire signal_1529 ;
    wire signal_1531 ;
    wire signal_1533 ;
    wire signal_1535 ;
    wire signal_1537 ;
    wire signal_1539 ;
    wire signal_1541 ;
    wire signal_1543 ;
    wire signal_1545 ;
    wire signal_1547 ;
    wire signal_1549 ;
    wire signal_1551 ;
    wire signal_1553 ;
    wire signal_1555 ;
    wire signal_1557 ;
    wire signal_1559 ;
    wire signal_1561 ;
    wire signal_1563 ;
    wire signal_1565 ;
    wire signal_1567 ;
    wire signal_1569 ;
    wire signal_1571 ;
    wire signal_1573 ;
    wire signal_1575 ;
    wire signal_1577 ;
    wire signal_1579 ;
    wire signal_1581 ;
    wire signal_1583 ;
    wire signal_1585 ;
    wire signal_1587 ;
    wire signal_1589 ;
    wire signal_1591 ;
    wire signal_1593 ;
    wire signal_1595 ;
    wire signal_1597 ;
    wire signal_1599 ;
    wire signal_1601 ;
    wire signal_1603 ;
    wire signal_1605 ;
    wire signal_1607 ;
    wire signal_1609 ;
    wire signal_1611 ;
    wire signal_1676 ;
    wire signal_1677 ;
    wire signal_1678 ;
    wire signal_1679 ;
    wire signal_1680 ;
    wire signal_1681 ;
    wire signal_1682 ;
    wire signal_1683 ;
    wire signal_1684 ;
    wire signal_1685 ;
    wire signal_1686 ;
    wire signal_1687 ;
    wire signal_1688 ;
    wire signal_1689 ;
    wire signal_1690 ;
    wire signal_1691 ;
    wire signal_1692 ;
    wire signal_1693 ;
    wire signal_1694 ;
    wire signal_1695 ;
    wire signal_1696 ;
    wire signal_1697 ;
    wire signal_1698 ;
    wire signal_1699 ;
    wire signal_1700 ;
    wire signal_1701 ;
    wire signal_1702 ;
    wire signal_1703 ;
    wire signal_1704 ;
    wire signal_1705 ;
    wire signal_1706 ;
    wire signal_1707 ;
    wire signal_1708 ;
    wire signal_1709 ;
    wire signal_1710 ;
    wire signal_1711 ;
    wire signal_1712 ;
    wire signal_1713 ;
    wire signal_1714 ;
    wire signal_1715 ;
    wire signal_1716 ;
    wire signal_1717 ;
    wire signal_1718 ;
    wire signal_1719 ;
    wire signal_1720 ;
    wire signal_1721 ;
    wire signal_1722 ;
    wire signal_1723 ;
    wire signal_1724 ;
    wire signal_1725 ;
    wire signal_1726 ;
    wire signal_1727 ;
    wire signal_1728 ;
    wire signal_1729 ;
    wire signal_1730 ;
    wire signal_1731 ;
    wire signal_1732 ;
    wire signal_1733 ;
    wire signal_1734 ;
    wire signal_1735 ;
    wire signal_1736 ;
    wire signal_1737 ;
    wire signal_1738 ;
    wire signal_1739 ;
    wire signal_1740 ;
    wire signal_1741 ;
    wire signal_1742 ;
    wire signal_1743 ;
    wire signal_1744 ;
    wire signal_1745 ;
    wire signal_1746 ;
    wire signal_1747 ;
    wire signal_1748 ;
    wire signal_1749 ;
    wire signal_1750 ;
    wire signal_1751 ;
    wire signal_1752 ;
    wire signal_1753 ;
    wire signal_1754 ;
    wire signal_1755 ;
    wire signal_1756 ;
    wire signal_1757 ;
    wire signal_1758 ;
    wire signal_1759 ;
    wire signal_1760 ;
    wire signal_1761 ;
    wire signal_1762 ;
    wire signal_1763 ;
    wire signal_1764 ;
    wire signal_1765 ;
    wire signal_1766 ;
    wire signal_1767 ;
    wire signal_1768 ;
    wire signal_1769 ;
    wire signal_1770 ;
    wire signal_1771 ;
    wire signal_1772 ;
    wire signal_1773 ;
    wire signal_1774 ;
    wire signal_1775 ;
    wire signal_1776 ;
    wire signal_1777 ;
    wire signal_1778 ;
    wire signal_1779 ;
    wire signal_1780 ;
    wire signal_1781 ;
    wire signal_1782 ;
    wire signal_1783 ;
    wire signal_1784 ;
    wire signal_1785 ;
    wire signal_1786 ;
    wire signal_1787 ;
    wire signal_1788 ;
    wire signal_1789 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1792 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1795 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1813 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1844 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1854 ;
    wire signal_1855 ;
    wire signal_1856 ;
    wire signal_1857 ;
    wire signal_1858 ;
    wire signal_1859 ;
    wire signal_1860 ;
    wire signal_1861 ;
    wire signal_1862 ;
    wire signal_1863 ;
    wire signal_1864 ;
    wire signal_1865 ;
    wire signal_1866 ;
    wire signal_1867 ;
    wire signal_1868 ;
    wire signal_1869 ;
    wire signal_1870 ;
    wire signal_1871 ;
    wire signal_1872 ;
    wire signal_1873 ;
    wire signal_1874 ;
    wire signal_1875 ;
    wire signal_1876 ;
    wire signal_1877 ;
    wire signal_1878 ;
    wire signal_1879 ;
    wire signal_1880 ;
    wire signal_1881 ;
    wire signal_1882 ;
    wire signal_1883 ;
    wire signal_1884 ;
    wire signal_1885 ;
    wire signal_1886 ;
    wire signal_1887 ;
    wire signal_1888 ;
    wire signal_1889 ;
    wire signal_1890 ;
    wire signal_1891 ;
    wire signal_1892 ;
    wire signal_1893 ;
    wire signal_1894 ;
    wire signal_1895 ;
    wire signal_1896 ;
    wire signal_1897 ;
    wire signal_1898 ;
    wire signal_1899 ;
    wire signal_1900 ;
    wire signal_1901 ;
    wire signal_1902 ;
    wire signal_1903 ;
    wire signal_1904 ;
    wire signal_1905 ;
    wire signal_1906 ;
    wire signal_1907 ;
    wire signal_1908 ;
    wire signal_1909 ;
    wire signal_1910 ;
    wire signal_1911 ;
    wire signal_1912 ;
    wire signal_1913 ;
    wire signal_1914 ;
    wire signal_1915 ;
    wire signal_1916 ;
    wire signal_1917 ;
    wire signal_1918 ;
    wire signal_1919 ;
    wire signal_1920 ;
    wire signal_1921 ;
    wire signal_1922 ;
    wire signal_1923 ;
    wire signal_1924 ;
    wire signal_1925 ;
    wire signal_1926 ;
    wire signal_1927 ;
    wire signal_1928 ;
    wire signal_1929 ;
    wire signal_1930 ;
    wire signal_1931 ;
    wire signal_1932 ;
    wire signal_1933 ;
    wire signal_1934 ;
    wire signal_1935 ;
    wire signal_1936 ;
    wire signal_1937 ;
    wire signal_1938 ;
    wire signal_1939 ;
    wire signal_1940 ;
    wire signal_1941 ;
    wire signal_1942 ;
    wire signal_1943 ;
    wire signal_1944 ;
    wire signal_1945 ;
    wire signal_1946 ;
    wire signal_1947 ;
    wire signal_1948 ;
    wire signal_1949 ;
    wire signal_1950 ;
    wire signal_1951 ;
    wire signal_1952 ;
    wire signal_1953 ;
    wire signal_1954 ;
    wire signal_1955 ;
    wire signal_1956 ;
    wire signal_1957 ;
    wire signal_1958 ;
    wire signal_1959 ;
    wire signal_1960 ;
    wire signal_1961 ;
    wire signal_1962 ;
    wire signal_1963 ;
    wire signal_1964 ;
    wire signal_1965 ;
    wire signal_1966 ;
    wire signal_1967 ;
    wire signal_1968 ;
    wire signal_1969 ;
    wire signal_1970 ;
    wire signal_1971 ;
    wire signal_1972 ;
    wire signal_1973 ;
    wire signal_1974 ;
    wire signal_1975 ;
    wire signal_1976 ;
    wire signal_1977 ;
    wire signal_1978 ;
    wire signal_1979 ;
    wire signal_1980 ;
    wire signal_1981 ;
    wire signal_1982 ;
    wire signal_1983 ;
    wire signal_1984 ;
    wire signal_1985 ;
    wire signal_1986 ;
    wire signal_1987 ;
    wire signal_1988 ;
    wire signal_1989 ;
    wire signal_1990 ;
    wire signal_1991 ;
    wire signal_1992 ;
    wire signal_1993 ;
    wire signal_1994 ;
    wire signal_1995 ;
    wire signal_1996 ;
    wire signal_1997 ;
    wire signal_1998 ;
    wire signal_1999 ;
    wire signal_2000 ;
    wire signal_2001 ;
    wire signal_2002 ;
    wire signal_2003 ;
    wire signal_2004 ;
    wire signal_2005 ;
    wire signal_2006 ;
    wire signal_2007 ;
    wire signal_2008 ;
    wire signal_2009 ;
    wire signal_2010 ;
    wire signal_2011 ;
    wire signal_2012 ;
    wire signal_2013 ;
    wire signal_2014 ;
    wire signal_2015 ;
    wire signal_2016 ;
    wire signal_2017 ;
    wire signal_2018 ;
    wire signal_2019 ;
    wire signal_2020 ;
    wire signal_2021 ;
    wire signal_2022 ;
    wire signal_2023 ;
    wire signal_2024 ;
    wire signal_2025 ;
    wire signal_2026 ;
    wire signal_2027 ;
    wire signal_2028 ;
    wire signal_2029 ;
    wire signal_2030 ;
    wire signal_2031 ;
    wire signal_2032 ;
    wire signal_2033 ;
    wire signal_2034 ;
    wire signal_2035 ;
    wire signal_2036 ;
    wire signal_2037 ;
    wire signal_2038 ;
    wire signal_2039 ;
    wire signal_2040 ;
    wire signal_2041 ;
    wire signal_2042 ;
    wire signal_2043 ;
    wire signal_2044 ;
    wire signal_2045 ;
    wire signal_2046 ;
    wire signal_2047 ;
    wire signal_2048 ;
    wire signal_2049 ;
    wire signal_2050 ;
    wire signal_2051 ;
    wire signal_2052 ;
    wire signal_2053 ;
    wire signal_2054 ;
    wire signal_2055 ;
    wire signal_2056 ;
    wire signal_2057 ;
    wire signal_2058 ;
    wire signal_2059 ;
    wire signal_2060 ;
    wire signal_2061 ;
    wire signal_2062 ;
    wire signal_2063 ;
    wire signal_2064 ;
    wire signal_2065 ;
    wire signal_2066 ;
    wire signal_2067 ;
    wire signal_2068 ;
    wire signal_2069 ;
    wire signal_2070 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2079 ;
    wire signal_2080 ;
    wire signal_2081 ;
    wire signal_2082 ;
    wire signal_2083 ;
    wire signal_2084 ;
    wire signal_2085 ;
    wire signal_2086 ;
    wire signal_2087 ;
    wire signal_2088 ;
    wire signal_2089 ;
    wire signal_2090 ;
    wire signal_2091 ;
    wire signal_2092 ;
    wire signal_2093 ;
    wire signal_2094 ;
    wire signal_2095 ;
    wire signal_2096 ;
    wire signal_2097 ;
    wire signal_2098 ;
    wire signal_2099 ;
    wire signal_2100 ;
    wire signal_2101 ;
    wire signal_2102 ;
    wire signal_2103 ;
    wire signal_2104 ;
    wire signal_2105 ;
    wire signal_2106 ;
    wire signal_2107 ;
    wire signal_2108 ;
    wire signal_2109 ;
    wire signal_2110 ;
    wire signal_2111 ;
    wire signal_2112 ;
    wire signal_2113 ;
    wire signal_2114 ;
    wire signal_2115 ;
    wire signal_2116 ;
    wire signal_2117 ;
    wire signal_2118 ;
    wire signal_2119 ;
    wire signal_2120 ;
    wire signal_2121 ;
    wire signal_2122 ;
    wire signal_2123 ;
    wire signal_2124 ;
    wire signal_2125 ;
    wire signal_2126 ;
    wire signal_2127 ;
    wire signal_2128 ;
    wire signal_2129 ;
    wire signal_2130 ;
    wire signal_2131 ;
    wire signal_2132 ;
    wire signal_2133 ;
    wire signal_2134 ;
    wire signal_2135 ;
    wire signal_2136 ;
    wire signal_2137 ;
    wire signal_2138 ;
    wire signal_2139 ;
    wire signal_2140 ;
    wire signal_2141 ;
    wire signal_2142 ;
    wire signal_2143 ;
    wire signal_2144 ;
    wire signal_2145 ;
    wire signal_2146 ;
    wire signal_2147 ;
    wire signal_2148 ;
    wire signal_2149 ;
    wire signal_2150 ;
    wire signal_2151 ;
    wire signal_2152 ;
    wire signal_2153 ;
    wire signal_2154 ;
    wire signal_2155 ;
    wire signal_2156 ;
    wire signal_2157 ;
    wire signal_2158 ;
    wire signal_2159 ;
    wire signal_2160 ;
    wire signal_2161 ;
    wire signal_2162 ;
    wire signal_2163 ;
    wire signal_2164 ;
    wire signal_2165 ;
    wire signal_2166 ;
    wire signal_2167 ;
    wire signal_2168 ;
    wire signal_2169 ;
    wire signal_2170 ;
    wire signal_2171 ;
    wire signal_2172 ;
    wire signal_2173 ;
    wire signal_2174 ;
    wire signal_2175 ;
    wire signal_2176 ;
    wire signal_2177 ;
    wire signal_2178 ;
    wire signal_2179 ;
    wire signal_2180 ;
    wire signal_2181 ;
    wire signal_2182 ;
    wire signal_2183 ;
    wire signal_2184 ;
    wire signal_2185 ;
    wire signal_2186 ;
    wire signal_2187 ;
    wire signal_2188 ;
    wire signal_2189 ;
    wire signal_2190 ;
    wire signal_2191 ;
    wire signal_2192 ;
    wire signal_2193 ;
    wire signal_2194 ;
    wire signal_2195 ;
    wire signal_2196 ;
    wire signal_2197 ;
    wire signal_2198 ;
    wire signal_2199 ;
    wire signal_2200 ;
    wire signal_2201 ;

    /* cells in depth 0 */
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_769 ( .s (rst), .b ({signal_1164, signal_1163}), .a ({Key_s1[0], Key_s0[0]}), .c ({signal_1166, signal_1099}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_770 ( .s (rst), .b ({signal_1167, signal_1162}), .a ({Key_s1[1], Key_s0[1]}), .c ({signal_1169, signal_1098}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_771 ( .s (rst), .b ({signal_1170, signal_1161}), .a ({Key_s1[2], Key_s0[2]}), .c ({signal_1172, signal_1097}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_772 ( .s (rst), .b ({signal_1173, signal_1160}), .a ({Key_s1[3], Key_s0[3]}), .c ({signal_1175, signal_1096}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_773 ( .s (rst), .b ({signal_1176, signal_1159}), .a ({Key_s1[4], Key_s0[4]}), .c ({signal_1178, signal_1095}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_774 ( .s (rst), .b ({signal_1179, signal_1158}), .a ({Key_s1[5], Key_s0[5]}), .c ({signal_1181, signal_1094}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_775 ( .s (rst), .b ({signal_1182, signal_1157}), .a ({Key_s1[6], Key_s0[6]}), .c ({signal_1184, signal_1093}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_776 ( .s (rst), .b ({signal_1185, signal_1156}), .a ({Key_s1[7], Key_s0[7]}), .c ({signal_1187, signal_1092}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_777 ( .s (rst), .b ({signal_1188, signal_1155}), .a ({Key_s1[8], Key_s0[8]}), .c ({signal_1190, signal_1091}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_778 ( .s (rst), .b ({signal_1191, signal_1154}), .a ({Key_s1[9], Key_s0[9]}), .c ({signal_1193, signal_1090}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_779 ( .s (rst), .b ({signal_1194, signal_1153}), .a ({Key_s1[10], Key_s0[10]}), .c ({signal_1196, signal_1089}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_780 ( .s (rst), .b ({signal_1197, signal_1152}), .a ({Key_s1[11], Key_s0[11]}), .c ({signal_1199, signal_1088}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_781 ( .s (rst), .b ({signal_1200, signal_1151}), .a ({Key_s1[12], Key_s0[12]}), .c ({signal_1202, signal_1087}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_782 ( .s (rst), .b ({signal_1203, signal_1150}), .a ({Key_s1[13], Key_s0[13]}), .c ({signal_1205, signal_1086}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_783 ( .s (rst), .b ({signal_1206, signal_1149}), .a ({Key_s1[14], Key_s0[14]}), .c ({signal_1208, signal_1085}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_784 ( .s (rst), .b ({signal_1209, signal_1148}), .a ({Key_s1[15], Key_s0[15]}), .c ({signal_1211, signal_1084}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_785 ( .s (rst), .b ({signal_1212, signal_1147}), .a ({Key_s1[16], Key_s0[16]}), .c ({signal_1214, signal_1083}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_786 ( .s (rst), .b ({signal_1215, signal_1146}), .a ({Key_s1[17], Key_s0[17]}), .c ({signal_1217, signal_1082}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_787 ( .s (rst), .b ({signal_1218, signal_1145}), .a ({Key_s1[18], Key_s0[18]}), .c ({signal_1220, signal_1081}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_788 ( .s (rst), .b ({signal_1221, signal_1144}), .a ({Key_s1[19], Key_s0[19]}), .c ({signal_1223, signal_1080}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_789 ( .s (rst), .b ({signal_1224, signal_1143}), .a ({Key_s1[20], Key_s0[20]}), .c ({signal_1226, signal_1079}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_790 ( .s (rst), .b ({signal_1227, signal_1142}), .a ({Key_s1[21], Key_s0[21]}), .c ({signal_1229, signal_1078}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_791 ( .s (rst), .b ({signal_1230, signal_1141}), .a ({Key_s1[22], Key_s0[22]}), .c ({signal_1232, signal_1077}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_792 ( .s (rst), .b ({signal_1233, signal_1140}), .a ({Key_s1[23], Key_s0[23]}), .c ({signal_1235, signal_1076}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_793 ( .s (rst), .b ({signal_1236, signal_1139}), .a ({Key_s1[24], Key_s0[24]}), .c ({signal_1238, signal_1075}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_794 ( .s (rst), .b ({signal_1239, signal_1138}), .a ({Key_s1[25], Key_s0[25]}), .c ({signal_1241, signal_1074}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_795 ( .s (rst), .b ({signal_1242, signal_1137}), .a ({Key_s1[26], Key_s0[26]}), .c ({signal_1244, signal_1073}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_796 ( .s (rst), .b ({signal_1245, signal_1136}), .a ({Key_s1[27], Key_s0[27]}), .c ({signal_1247, signal_1072}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_797 ( .s (rst), .b ({signal_1248, signal_1135}), .a ({Key_s1[28], Key_s0[28]}), .c ({signal_1250, signal_1071}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_798 ( .s (rst), .b ({signal_1251, signal_1134}), .a ({Key_s1[29], Key_s0[29]}), .c ({signal_1253, signal_1070}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_799 ( .s (rst), .b ({signal_1254, signal_1133}), .a ({Key_s1[30], Key_s0[30]}), .c ({signal_1256, signal_1069}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_800 ( .s (rst), .b ({signal_1257, signal_1132}), .a ({Key_s1[31], Key_s0[31]}), .c ({signal_1259, signal_1068}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_801 ( .s (rst), .b ({signal_1260, signal_1131}), .a ({Key_s1[32], Key_s0[32]}), .c ({signal_1262, signal_1067}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_802 ( .s (rst), .b ({signal_1263, signal_1130}), .a ({Key_s1[33], Key_s0[33]}), .c ({signal_1265, signal_1066}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_803 ( .s (rst), .b ({signal_1266, signal_1129}), .a ({Key_s1[34], Key_s0[34]}), .c ({signal_1268, signal_1065}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_804 ( .s (rst), .b ({signal_1269, signal_1128}), .a ({Key_s1[35], Key_s0[35]}), .c ({signal_1271, signal_1064}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_805 ( .s (rst), .b ({signal_1272, signal_1127}), .a ({Key_s1[36], Key_s0[36]}), .c ({signal_1274, signal_1063}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_806 ( .s (rst), .b ({signal_1275, signal_1126}), .a ({Key_s1[37], Key_s0[37]}), .c ({signal_1277, signal_1062}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_807 ( .s (rst), .b ({signal_1278, signal_1125}), .a ({Key_s1[38], Key_s0[38]}), .c ({signal_1280, signal_1061}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_808 ( .s (rst), .b ({signal_1281, signal_1124}), .a ({Key_s1[39], Key_s0[39]}), .c ({signal_1283, signal_1060}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_809 ( .s (rst), .b ({signal_1284, signal_1123}), .a ({Key_s1[40], Key_s0[40]}), .c ({signal_1286, signal_1059}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_810 ( .s (rst), .b ({signal_1287, signal_1122}), .a ({Key_s1[41], Key_s0[41]}), .c ({signal_1289, signal_1058}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_811 ( .s (rst), .b ({signal_1290, signal_1121}), .a ({Key_s1[42], Key_s0[42]}), .c ({signal_1292, signal_1057}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_812 ( .s (rst), .b ({signal_1293, signal_1120}), .a ({Key_s1[43], Key_s0[43]}), .c ({signal_1295, signal_1056}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_813 ( .s (rst), .b ({signal_1296, signal_1119}), .a ({Key_s1[44], Key_s0[44]}), .c ({signal_1298, signal_1055}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_814 ( .s (rst), .b ({signal_1299, signal_1118}), .a ({Key_s1[45], Key_s0[45]}), .c ({signal_1301, signal_1054}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_815 ( .s (rst), .b ({signal_1302, signal_1117}), .a ({Key_s1[46], Key_s0[46]}), .c ({signal_1304, signal_1053}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_816 ( .s (rst), .b ({signal_1305, signal_1116}), .a ({Key_s1[47], Key_s0[47]}), .c ({signal_1307, signal_1052}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_817 ( .s (rst), .b ({signal_1308, signal_1115}), .a ({Key_s1[48], Key_s0[48]}), .c ({signal_1310, signal_1051}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_818 ( .s (rst), .b ({signal_1311, signal_1114}), .a ({Key_s1[49], Key_s0[49]}), .c ({signal_1313, signal_1050}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_819 ( .s (rst), .b ({signal_1314, signal_1113}), .a ({Key_s1[50], Key_s0[50]}), .c ({signal_1316, signal_1049}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_820 ( .s (rst), .b ({signal_1317, signal_1112}), .a ({Key_s1[51], Key_s0[51]}), .c ({signal_1319, signal_1048}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_821 ( .s (rst), .b ({signal_1320, signal_1111}), .a ({Key_s1[52], Key_s0[52]}), .c ({signal_1322, signal_1047}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_822 ( .s (rst), .b ({signal_1323, signal_1110}), .a ({Key_s1[53], Key_s0[53]}), .c ({signal_1325, signal_1046}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_823 ( .s (rst), .b ({signal_1326, signal_1109}), .a ({Key_s1[54], Key_s0[54]}), .c ({signal_1328, signal_1045}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_824 ( .s (rst), .b ({signal_1329, signal_1108}), .a ({Key_s1[55], Key_s0[55]}), .c ({signal_1331, signal_1044}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_825 ( .s (rst), .b ({signal_1332, signal_1107}), .a ({Key_s1[56], Key_s0[56]}), .c ({signal_1334, signal_1043}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_826 ( .s (rst), .b ({signal_1335, signal_1106}), .a ({Key_s1[57], Key_s0[57]}), .c ({signal_1337, signal_1042}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_827 ( .s (rst), .b ({signal_1338, signal_1105}), .a ({Key_s1[58], Key_s0[58]}), .c ({signal_1340, signal_1041}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_828 ( .s (rst), .b ({signal_1341, signal_1104}), .a ({Key_s1[59], Key_s0[59]}), .c ({signal_1343, signal_1040}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_829 ( .s (rst), .b ({signal_1344, signal_1103}), .a ({Key_s1[60], Key_s0[60]}), .c ({signal_1346, signal_1039}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_830 ( .s (rst), .b ({signal_1347, signal_1102}), .a ({Key_s1[61], Key_s0[61]}), .c ({signal_1349, signal_1038}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_831 ( .s (rst), .b ({signal_1350, signal_1101}), .a ({Key_s1[62], Key_s0[62]}), .c ({signal_1352, signal_1037}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_832 ( .s (rst), .b ({signal_1353, signal_1100}), .a ({Key_s1[63], Key_s0[63]}), .c ({signal_1355, signal_1036}) ) ;
    MUX2_X1 cell_961 ( .S (rst), .A (signal_1029), .B (1'b1), .Z (signal_1035) ) ;
    MUX2_X1 cell_962 ( .S (rst), .A (signal_1028), .B (1'b0), .Z (signal_1034) ) ;
    MUX2_X1 cell_963 ( .S (rst), .A (signal_1027), .B (1'b0), .Z (signal_1033) ) ;
    MUX2_X1 cell_964 ( .S (rst), .A (signal_1026), .B (1'b0), .Z (signal_1032) ) ;
    MUX2_X1 cell_965 ( .S (rst), .A (signal_1025), .B (1'b0), .Z (signal_1031) ) ;
    MUX2_X1 cell_966 ( .S (rst), .A (signal_1024), .B (1'b0), .Z (signal_1030) ) ;
    MUX2_X1 cell_979 ( .S (signal_940), .A (signal_759), .B (signal_939), .Z (signal_1029) ) ;
    NAND2_X1 cell_980 ( .A1 (signal_939), .A2 (signal_760), .ZN (signal_759) ) ;
    NAND2_X1 cell_981 ( .A1 (signal_761), .A2 (signal_762), .ZN (signal_760) ) ;
    NOR2_X1 cell_982 ( .A1 (signal_1026), .A2 (signal_1025), .ZN (signal_762) ) ;
    AND2_X1 cell_983 ( .A1 (signal_1028), .A2 (signal_943), .ZN (signal_761) ) ;
    AND2_X1 cell_984 ( .A1 (signal_763), .A2 (signal_943), .ZN (signal_1027) ) ;
    NAND2_X1 cell_985 ( .A1 (signal_764), .A2 (signal_939), .ZN (signal_763) ) ;
    NOR2_X1 cell_986 ( .A1 (signal_940), .A2 (signal_765), .ZN (signal_764) ) ;
    NAND2_X1 cell_987 ( .A1 (signal_1028), .A2 (signal_766), .ZN (signal_765) ) ;
    NOR2_X1 cell_988 ( .A1 (signal_1026), .A2 (signal_1025), .ZN (signal_766) ) ;
    OR2_X1 cell_989 ( .A1 (signal_940), .A2 (signal_767), .ZN (signal_1024) ) ;
    NOR2_X1 cell_990 ( .A1 (signal_1025), .A2 (signal_768), .ZN (signal_767) ) ;
    NAND2_X1 cell_991 ( .A1 (signal_939), .A2 (signal_769), .ZN (signal_768) ) ;
    NOR2_X1 cell_992 ( .A1 (signal_1026), .A2 (signal_770), .ZN (signal_769) ) ;
    NAND2_X1 cell_993 ( .A1 (signal_1028), .A2 (signal_943), .ZN (signal_770) ) ;
    NOR2_X1 cell_994 ( .A1 (signal_771), .A2 (signal_772), .ZN (done) ) ;
    NAND2_X1 cell_995 ( .A1 (signal_940), .A2 (signal_939), .ZN (signal_772) ) ;
    NAND2_X1 cell_996 ( .A1 (signal_773), .A2 (signal_774), .ZN (signal_771) ) ;
    NOR2_X1 cell_997 ( .A1 (signal_1025), .A2 (signal_775), .ZN (signal_774) ) ;
    INV_X1 cell_998 ( .A (signal_1028), .ZN (signal_775) ) ;
    NOR2_X1 cell_999 ( .A1 (signal_943), .A2 (signal_1026), .ZN (signal_773) ) ;

    /* cells in depth 1 */
    buf_clk cell_1001 ( .C (clk), .D (rst), .Q (signal_1676) ) ;
    buf_clk cell_1003 ( .C (clk), .D (Plaintext_s0[0]), .Q (signal_1678) ) ;
    buf_clk cell_1005 ( .C (clk), .D (Plaintext_s1[0]), .Q (signal_1680) ) ;
    buf_clk cell_1007 ( .C (clk), .D (Plaintext_s0[1]), .Q (signal_1682) ) ;
    buf_clk cell_1009 ( .C (clk), .D (Plaintext_s1[1]), .Q (signal_1684) ) ;
    buf_clk cell_1011 ( .C (clk), .D (Plaintext_s0[2]), .Q (signal_1686) ) ;
    buf_clk cell_1013 ( .C (clk), .D (Plaintext_s1[2]), .Q (signal_1688) ) ;
    buf_clk cell_1015 ( .C (clk), .D (Plaintext_s0[3]), .Q (signal_1690) ) ;
    buf_clk cell_1017 ( .C (clk), .D (Plaintext_s1[3]), .Q (signal_1692) ) ;
    buf_clk cell_1019 ( .C (clk), .D (Plaintext_s0[4]), .Q (signal_1694) ) ;
    buf_clk cell_1021 ( .C (clk), .D (Plaintext_s1[4]), .Q (signal_1696) ) ;
    buf_clk cell_1023 ( .C (clk), .D (Plaintext_s0[5]), .Q (signal_1698) ) ;
    buf_clk cell_1025 ( .C (clk), .D (Plaintext_s1[5]), .Q (signal_1700) ) ;
    buf_clk cell_1027 ( .C (clk), .D (Plaintext_s0[6]), .Q (signal_1702) ) ;
    buf_clk cell_1029 ( .C (clk), .D (Plaintext_s1[6]), .Q (signal_1704) ) ;
    buf_clk cell_1031 ( .C (clk), .D (Plaintext_s0[7]), .Q (signal_1706) ) ;
    buf_clk cell_1033 ( .C (clk), .D (Plaintext_s1[7]), .Q (signal_1708) ) ;
    buf_clk cell_1035 ( .C (clk), .D (Plaintext_s0[8]), .Q (signal_1710) ) ;
    buf_clk cell_1037 ( .C (clk), .D (Plaintext_s1[8]), .Q (signal_1712) ) ;
    buf_clk cell_1039 ( .C (clk), .D (Plaintext_s0[9]), .Q (signal_1714) ) ;
    buf_clk cell_1041 ( .C (clk), .D (Plaintext_s1[9]), .Q (signal_1716) ) ;
    buf_clk cell_1043 ( .C (clk), .D (Plaintext_s0[10]), .Q (signal_1718) ) ;
    buf_clk cell_1045 ( .C (clk), .D (Plaintext_s1[10]), .Q (signal_1720) ) ;
    buf_clk cell_1047 ( .C (clk), .D (Plaintext_s0[11]), .Q (signal_1722) ) ;
    buf_clk cell_1049 ( .C (clk), .D (Plaintext_s1[11]), .Q (signal_1724) ) ;
    buf_clk cell_1051 ( .C (clk), .D (Plaintext_s0[12]), .Q (signal_1726) ) ;
    buf_clk cell_1053 ( .C (clk), .D (Plaintext_s1[12]), .Q (signal_1728) ) ;
    buf_clk cell_1055 ( .C (clk), .D (Plaintext_s0[13]), .Q (signal_1730) ) ;
    buf_clk cell_1057 ( .C (clk), .D (Plaintext_s1[13]), .Q (signal_1732) ) ;
    buf_clk cell_1059 ( .C (clk), .D (Plaintext_s0[14]), .Q (signal_1734) ) ;
    buf_clk cell_1061 ( .C (clk), .D (Plaintext_s1[14]), .Q (signal_1736) ) ;
    buf_clk cell_1063 ( .C (clk), .D (Plaintext_s0[15]), .Q (signal_1738) ) ;
    buf_clk cell_1065 ( .C (clk), .D (Plaintext_s1[15]), .Q (signal_1740) ) ;
    buf_clk cell_1067 ( .C (clk), .D (Plaintext_s0[16]), .Q (signal_1742) ) ;
    buf_clk cell_1069 ( .C (clk), .D (Plaintext_s1[16]), .Q (signal_1744) ) ;
    buf_clk cell_1071 ( .C (clk), .D (Plaintext_s0[17]), .Q (signal_1746) ) ;
    buf_clk cell_1073 ( .C (clk), .D (Plaintext_s1[17]), .Q (signal_1748) ) ;
    buf_clk cell_1075 ( .C (clk), .D (Plaintext_s0[18]), .Q (signal_1750) ) ;
    buf_clk cell_1077 ( .C (clk), .D (Plaintext_s1[18]), .Q (signal_1752) ) ;
    buf_clk cell_1079 ( .C (clk), .D (Plaintext_s0[19]), .Q (signal_1754) ) ;
    buf_clk cell_1081 ( .C (clk), .D (Plaintext_s1[19]), .Q (signal_1756) ) ;
    buf_clk cell_1083 ( .C (clk), .D (Plaintext_s0[20]), .Q (signal_1758) ) ;
    buf_clk cell_1085 ( .C (clk), .D (Plaintext_s1[20]), .Q (signal_1760) ) ;
    buf_clk cell_1087 ( .C (clk), .D (Plaintext_s0[21]), .Q (signal_1762) ) ;
    buf_clk cell_1089 ( .C (clk), .D (Plaintext_s1[21]), .Q (signal_1764) ) ;
    buf_clk cell_1091 ( .C (clk), .D (Plaintext_s0[22]), .Q (signal_1766) ) ;
    buf_clk cell_1093 ( .C (clk), .D (Plaintext_s1[22]), .Q (signal_1768) ) ;
    buf_clk cell_1095 ( .C (clk), .D (Plaintext_s0[23]), .Q (signal_1770) ) ;
    buf_clk cell_1097 ( .C (clk), .D (Plaintext_s1[23]), .Q (signal_1772) ) ;
    buf_clk cell_1099 ( .C (clk), .D (Plaintext_s0[24]), .Q (signal_1774) ) ;
    buf_clk cell_1101 ( .C (clk), .D (Plaintext_s1[24]), .Q (signal_1776) ) ;
    buf_clk cell_1103 ( .C (clk), .D (Plaintext_s0[25]), .Q (signal_1778) ) ;
    buf_clk cell_1105 ( .C (clk), .D (Plaintext_s1[25]), .Q (signal_1780) ) ;
    buf_clk cell_1107 ( .C (clk), .D (Plaintext_s0[26]), .Q (signal_1782) ) ;
    buf_clk cell_1109 ( .C (clk), .D (Plaintext_s1[26]), .Q (signal_1784) ) ;
    buf_clk cell_1111 ( .C (clk), .D (Plaintext_s0[27]), .Q (signal_1786) ) ;
    buf_clk cell_1113 ( .C (clk), .D (Plaintext_s1[27]), .Q (signal_1788) ) ;
    buf_clk cell_1115 ( .C (clk), .D (Plaintext_s0[28]), .Q (signal_1790) ) ;
    buf_clk cell_1117 ( .C (clk), .D (Plaintext_s1[28]), .Q (signal_1792) ) ;
    buf_clk cell_1119 ( .C (clk), .D (Plaintext_s0[29]), .Q (signal_1794) ) ;
    buf_clk cell_1121 ( .C (clk), .D (Plaintext_s1[29]), .Q (signal_1796) ) ;
    buf_clk cell_1123 ( .C (clk), .D (Plaintext_s0[30]), .Q (signal_1798) ) ;
    buf_clk cell_1125 ( .C (clk), .D (Plaintext_s1[30]), .Q (signal_1800) ) ;
    buf_clk cell_1127 ( .C (clk), .D (Plaintext_s0[31]), .Q (signal_1802) ) ;
    buf_clk cell_1129 ( .C (clk), .D (Plaintext_s1[31]), .Q (signal_1804) ) ;
    buf_clk cell_1131 ( .C (clk), .D (Plaintext_s0[32]), .Q (signal_1806) ) ;
    buf_clk cell_1133 ( .C (clk), .D (Plaintext_s1[32]), .Q (signal_1808) ) ;
    buf_clk cell_1135 ( .C (clk), .D (Plaintext_s0[33]), .Q (signal_1810) ) ;
    buf_clk cell_1137 ( .C (clk), .D (Plaintext_s1[33]), .Q (signal_1812) ) ;
    buf_clk cell_1139 ( .C (clk), .D (Plaintext_s0[34]), .Q (signal_1814) ) ;
    buf_clk cell_1141 ( .C (clk), .D (Plaintext_s1[34]), .Q (signal_1816) ) ;
    buf_clk cell_1143 ( .C (clk), .D (Plaintext_s0[35]), .Q (signal_1818) ) ;
    buf_clk cell_1145 ( .C (clk), .D (Plaintext_s1[35]), .Q (signal_1820) ) ;
    buf_clk cell_1147 ( .C (clk), .D (Plaintext_s0[36]), .Q (signal_1822) ) ;
    buf_clk cell_1149 ( .C (clk), .D (Plaintext_s1[36]), .Q (signal_1824) ) ;
    buf_clk cell_1151 ( .C (clk), .D (Plaintext_s0[37]), .Q (signal_1826) ) ;
    buf_clk cell_1153 ( .C (clk), .D (Plaintext_s1[37]), .Q (signal_1828) ) ;
    buf_clk cell_1155 ( .C (clk), .D (Plaintext_s0[38]), .Q (signal_1830) ) ;
    buf_clk cell_1157 ( .C (clk), .D (Plaintext_s1[38]), .Q (signal_1832) ) ;
    buf_clk cell_1159 ( .C (clk), .D (Plaintext_s0[39]), .Q (signal_1834) ) ;
    buf_clk cell_1161 ( .C (clk), .D (Plaintext_s1[39]), .Q (signal_1836) ) ;
    buf_clk cell_1163 ( .C (clk), .D (Plaintext_s0[40]), .Q (signal_1838) ) ;
    buf_clk cell_1165 ( .C (clk), .D (Plaintext_s1[40]), .Q (signal_1840) ) ;
    buf_clk cell_1167 ( .C (clk), .D (Plaintext_s0[41]), .Q (signal_1842) ) ;
    buf_clk cell_1169 ( .C (clk), .D (Plaintext_s1[41]), .Q (signal_1844) ) ;
    buf_clk cell_1171 ( .C (clk), .D (Plaintext_s0[42]), .Q (signal_1846) ) ;
    buf_clk cell_1173 ( .C (clk), .D (Plaintext_s1[42]), .Q (signal_1848) ) ;
    buf_clk cell_1175 ( .C (clk), .D (Plaintext_s0[43]), .Q (signal_1850) ) ;
    buf_clk cell_1177 ( .C (clk), .D (Plaintext_s1[43]), .Q (signal_1852) ) ;
    buf_clk cell_1179 ( .C (clk), .D (Plaintext_s0[44]), .Q (signal_1854) ) ;
    buf_clk cell_1181 ( .C (clk), .D (Plaintext_s1[44]), .Q (signal_1856) ) ;
    buf_clk cell_1183 ( .C (clk), .D (Plaintext_s0[45]), .Q (signal_1858) ) ;
    buf_clk cell_1185 ( .C (clk), .D (Plaintext_s1[45]), .Q (signal_1860) ) ;
    buf_clk cell_1187 ( .C (clk), .D (Plaintext_s0[46]), .Q (signal_1862) ) ;
    buf_clk cell_1189 ( .C (clk), .D (Plaintext_s1[46]), .Q (signal_1864) ) ;
    buf_clk cell_1191 ( .C (clk), .D (Plaintext_s0[47]), .Q (signal_1866) ) ;
    buf_clk cell_1193 ( .C (clk), .D (Plaintext_s1[47]), .Q (signal_1868) ) ;
    buf_clk cell_1195 ( .C (clk), .D (Plaintext_s0[48]), .Q (signal_1870) ) ;
    buf_clk cell_1197 ( .C (clk), .D (Plaintext_s1[48]), .Q (signal_1872) ) ;
    buf_clk cell_1199 ( .C (clk), .D (Plaintext_s0[49]), .Q (signal_1874) ) ;
    buf_clk cell_1201 ( .C (clk), .D (Plaintext_s1[49]), .Q (signal_1876) ) ;
    buf_clk cell_1203 ( .C (clk), .D (Plaintext_s0[50]), .Q (signal_1878) ) ;
    buf_clk cell_1205 ( .C (clk), .D (Plaintext_s1[50]), .Q (signal_1880) ) ;
    buf_clk cell_1207 ( .C (clk), .D (Plaintext_s0[51]), .Q (signal_1882) ) ;
    buf_clk cell_1209 ( .C (clk), .D (Plaintext_s1[51]), .Q (signal_1884) ) ;
    buf_clk cell_1211 ( .C (clk), .D (Plaintext_s0[52]), .Q (signal_1886) ) ;
    buf_clk cell_1213 ( .C (clk), .D (Plaintext_s1[52]), .Q (signal_1888) ) ;
    buf_clk cell_1215 ( .C (clk), .D (Plaintext_s0[53]), .Q (signal_1890) ) ;
    buf_clk cell_1217 ( .C (clk), .D (Plaintext_s1[53]), .Q (signal_1892) ) ;
    buf_clk cell_1219 ( .C (clk), .D (Plaintext_s0[54]), .Q (signal_1894) ) ;
    buf_clk cell_1221 ( .C (clk), .D (Plaintext_s1[54]), .Q (signal_1896) ) ;
    buf_clk cell_1223 ( .C (clk), .D (Plaintext_s0[55]), .Q (signal_1898) ) ;
    buf_clk cell_1225 ( .C (clk), .D (Plaintext_s1[55]), .Q (signal_1900) ) ;
    buf_clk cell_1227 ( .C (clk), .D (Plaintext_s0[56]), .Q (signal_1902) ) ;
    buf_clk cell_1229 ( .C (clk), .D (Plaintext_s1[56]), .Q (signal_1904) ) ;
    buf_clk cell_1231 ( .C (clk), .D (Plaintext_s0[57]), .Q (signal_1906) ) ;
    buf_clk cell_1233 ( .C (clk), .D (Plaintext_s1[57]), .Q (signal_1908) ) ;
    buf_clk cell_1235 ( .C (clk), .D (Plaintext_s0[58]), .Q (signal_1910) ) ;
    buf_clk cell_1237 ( .C (clk), .D (Plaintext_s1[58]), .Q (signal_1912) ) ;
    buf_clk cell_1239 ( .C (clk), .D (Plaintext_s0[59]), .Q (signal_1914) ) ;
    buf_clk cell_1241 ( .C (clk), .D (Plaintext_s1[59]), .Q (signal_1916) ) ;
    buf_clk cell_1243 ( .C (clk), .D (Plaintext_s0[60]), .Q (signal_1918) ) ;
    buf_clk cell_1245 ( .C (clk), .D (Plaintext_s1[60]), .Q (signal_1920) ) ;
    buf_clk cell_1247 ( .C (clk), .D (Plaintext_s0[61]), .Q (signal_1922) ) ;
    buf_clk cell_1249 ( .C (clk), .D (Plaintext_s1[61]), .Q (signal_1924) ) ;
    buf_clk cell_1251 ( .C (clk), .D (Plaintext_s0[62]), .Q (signal_1926) ) ;
    buf_clk cell_1253 ( .C (clk), .D (Plaintext_s1[62]), .Q (signal_1928) ) ;
    buf_clk cell_1255 ( .C (clk), .D (Plaintext_s0[63]), .Q (signal_1930) ) ;
    buf_clk cell_1257 ( .C (clk), .D (Plaintext_s1[63]), .Q (signal_1932) ) ;
    buf_clk cell_1259 ( .C (clk), .D (signal_1036), .Q (signal_1934) ) ;
    buf_clk cell_1261 ( .C (clk), .D (signal_1355), .Q (signal_1936) ) ;
    buf_clk cell_1263 ( .C (clk), .D (signal_1037), .Q (signal_1938) ) ;
    buf_clk cell_1265 ( .C (clk), .D (signal_1352), .Q (signal_1940) ) ;
    buf_clk cell_1267 ( .C (clk), .D (signal_1038), .Q (signal_1942) ) ;
    buf_clk cell_1269 ( .C (clk), .D (signal_1349), .Q (signal_1944) ) ;
    buf_clk cell_1271 ( .C (clk), .D (signal_1039), .Q (signal_1946) ) ;
    buf_clk cell_1273 ( .C (clk), .D (signal_1346), .Q (signal_1948) ) ;
    buf_clk cell_1275 ( .C (clk), .D (signal_1040), .Q (signal_1950) ) ;
    buf_clk cell_1277 ( .C (clk), .D (signal_1343), .Q (signal_1952) ) ;
    buf_clk cell_1279 ( .C (clk), .D (signal_1041), .Q (signal_1954) ) ;
    buf_clk cell_1281 ( .C (clk), .D (signal_1340), .Q (signal_1956) ) ;
    buf_clk cell_1283 ( .C (clk), .D (signal_1042), .Q (signal_1958) ) ;
    buf_clk cell_1285 ( .C (clk), .D (signal_1337), .Q (signal_1960) ) ;
    buf_clk cell_1287 ( .C (clk), .D (signal_1043), .Q (signal_1962) ) ;
    buf_clk cell_1289 ( .C (clk), .D (signal_1334), .Q (signal_1964) ) ;
    buf_clk cell_1291 ( .C (clk), .D (signal_1044), .Q (signal_1966) ) ;
    buf_clk cell_1293 ( .C (clk), .D (signal_1331), .Q (signal_1968) ) ;
    buf_clk cell_1295 ( .C (clk), .D (signal_1045), .Q (signal_1970) ) ;
    buf_clk cell_1297 ( .C (clk), .D (signal_1328), .Q (signal_1972) ) ;
    buf_clk cell_1299 ( .C (clk), .D (signal_1046), .Q (signal_1974) ) ;
    buf_clk cell_1301 ( .C (clk), .D (signal_1325), .Q (signal_1976) ) ;
    buf_clk cell_1303 ( .C (clk), .D (signal_1047), .Q (signal_1978) ) ;
    buf_clk cell_1305 ( .C (clk), .D (signal_1322), .Q (signal_1980) ) ;
    buf_clk cell_1307 ( .C (clk), .D (signal_1048), .Q (signal_1982) ) ;
    buf_clk cell_1309 ( .C (clk), .D (signal_1319), .Q (signal_1984) ) ;
    buf_clk cell_1311 ( .C (clk), .D (signal_1049), .Q (signal_1986) ) ;
    buf_clk cell_1313 ( .C (clk), .D (signal_1316), .Q (signal_1988) ) ;
    buf_clk cell_1315 ( .C (clk), .D (signal_1050), .Q (signal_1990) ) ;
    buf_clk cell_1317 ( .C (clk), .D (signal_1313), .Q (signal_1992) ) ;
    buf_clk cell_1319 ( .C (clk), .D (signal_1051), .Q (signal_1994) ) ;
    buf_clk cell_1321 ( .C (clk), .D (signal_1310), .Q (signal_1996) ) ;
    buf_clk cell_1323 ( .C (clk), .D (signal_1052), .Q (signal_1998) ) ;
    buf_clk cell_1325 ( .C (clk), .D (signal_1307), .Q (signal_2000) ) ;
    buf_clk cell_1327 ( .C (clk), .D (signal_1053), .Q (signal_2002) ) ;
    buf_clk cell_1329 ( .C (clk), .D (signal_1304), .Q (signal_2004) ) ;
    buf_clk cell_1331 ( .C (clk), .D (signal_1054), .Q (signal_2006) ) ;
    buf_clk cell_1333 ( .C (clk), .D (signal_1301), .Q (signal_2008) ) ;
    buf_clk cell_1335 ( .C (clk), .D (signal_1055), .Q (signal_2010) ) ;
    buf_clk cell_1337 ( .C (clk), .D (signal_1298), .Q (signal_2012) ) ;
    buf_clk cell_1339 ( .C (clk), .D (signal_1056), .Q (signal_2014) ) ;
    buf_clk cell_1341 ( .C (clk), .D (signal_1295), .Q (signal_2016) ) ;
    buf_clk cell_1343 ( .C (clk), .D (signal_1057), .Q (signal_2018) ) ;
    buf_clk cell_1345 ( .C (clk), .D (signal_1292), .Q (signal_2020) ) ;
    buf_clk cell_1347 ( .C (clk), .D (signal_1058), .Q (signal_2022) ) ;
    buf_clk cell_1349 ( .C (clk), .D (signal_1289), .Q (signal_2024) ) ;
    buf_clk cell_1351 ( .C (clk), .D (signal_1059), .Q (signal_2026) ) ;
    buf_clk cell_1353 ( .C (clk), .D (signal_1286), .Q (signal_2028) ) ;
    buf_clk cell_1355 ( .C (clk), .D (signal_1060), .Q (signal_2030) ) ;
    buf_clk cell_1357 ( .C (clk), .D (signal_1283), .Q (signal_2032) ) ;
    buf_clk cell_1359 ( .C (clk), .D (signal_1061), .Q (signal_2034) ) ;
    buf_clk cell_1361 ( .C (clk), .D (signal_1280), .Q (signal_2036) ) ;
    buf_clk cell_1363 ( .C (clk), .D (signal_1062), .Q (signal_2038) ) ;
    buf_clk cell_1365 ( .C (clk), .D (signal_1277), .Q (signal_2040) ) ;
    buf_clk cell_1367 ( .C (clk), .D (signal_1063), .Q (signal_2042) ) ;
    buf_clk cell_1369 ( .C (clk), .D (signal_1274), .Q (signal_2044) ) ;
    buf_clk cell_1371 ( .C (clk), .D (signal_1064), .Q (signal_2046) ) ;
    buf_clk cell_1373 ( .C (clk), .D (signal_1271), .Q (signal_2048) ) ;
    buf_clk cell_1375 ( .C (clk), .D (signal_1065), .Q (signal_2050) ) ;
    buf_clk cell_1377 ( .C (clk), .D (signal_1268), .Q (signal_2052) ) ;
    buf_clk cell_1379 ( .C (clk), .D (signal_1066), .Q (signal_2054) ) ;
    buf_clk cell_1381 ( .C (clk), .D (signal_1265), .Q (signal_2056) ) ;
    buf_clk cell_1383 ( .C (clk), .D (signal_1067), .Q (signal_2058) ) ;
    buf_clk cell_1385 ( .C (clk), .D (signal_1262), .Q (signal_2060) ) ;
    buf_clk cell_1387 ( .C (clk), .D (signal_1068), .Q (signal_2062) ) ;
    buf_clk cell_1389 ( .C (clk), .D (signal_1259), .Q (signal_2064) ) ;
    buf_clk cell_1391 ( .C (clk), .D (signal_1069), .Q (signal_2066) ) ;
    buf_clk cell_1393 ( .C (clk), .D (signal_1256), .Q (signal_2068) ) ;
    buf_clk cell_1395 ( .C (clk), .D (signal_1070), .Q (signal_2070) ) ;
    buf_clk cell_1397 ( .C (clk), .D (signal_1253), .Q (signal_2072) ) ;
    buf_clk cell_1399 ( .C (clk), .D (signal_1071), .Q (signal_2074) ) ;
    buf_clk cell_1401 ( .C (clk), .D (signal_1250), .Q (signal_2076) ) ;
    buf_clk cell_1403 ( .C (clk), .D (signal_1072), .Q (signal_2078) ) ;
    buf_clk cell_1405 ( .C (clk), .D (signal_1247), .Q (signal_2080) ) ;
    buf_clk cell_1407 ( .C (clk), .D (signal_1073), .Q (signal_2082) ) ;
    buf_clk cell_1409 ( .C (clk), .D (signal_1244), .Q (signal_2084) ) ;
    buf_clk cell_1411 ( .C (clk), .D (signal_1074), .Q (signal_2086) ) ;
    buf_clk cell_1413 ( .C (clk), .D (signal_1241), .Q (signal_2088) ) ;
    buf_clk cell_1415 ( .C (clk), .D (signal_1075), .Q (signal_2090) ) ;
    buf_clk cell_1417 ( .C (clk), .D (signal_1238), .Q (signal_2092) ) ;
    buf_clk cell_1419 ( .C (clk), .D (signal_1076), .Q (signal_2094) ) ;
    buf_clk cell_1421 ( .C (clk), .D (signal_1235), .Q (signal_2096) ) ;
    buf_clk cell_1423 ( .C (clk), .D (signal_1077), .Q (signal_2098) ) ;
    buf_clk cell_1425 ( .C (clk), .D (signal_1232), .Q (signal_2100) ) ;
    buf_clk cell_1427 ( .C (clk), .D (signal_1078), .Q (signal_2102) ) ;
    buf_clk cell_1429 ( .C (clk), .D (signal_1229), .Q (signal_2104) ) ;
    buf_clk cell_1431 ( .C (clk), .D (signal_1079), .Q (signal_2106) ) ;
    buf_clk cell_1433 ( .C (clk), .D (signal_1226), .Q (signal_2108) ) ;
    buf_clk cell_1435 ( .C (clk), .D (signal_1080), .Q (signal_2110) ) ;
    buf_clk cell_1437 ( .C (clk), .D (signal_1223), .Q (signal_2112) ) ;
    buf_clk cell_1439 ( .C (clk), .D (signal_1081), .Q (signal_2114) ) ;
    buf_clk cell_1441 ( .C (clk), .D (signal_1220), .Q (signal_2116) ) ;
    buf_clk cell_1443 ( .C (clk), .D (signal_1082), .Q (signal_2118) ) ;
    buf_clk cell_1445 ( .C (clk), .D (signal_1217), .Q (signal_2120) ) ;
    buf_clk cell_1447 ( .C (clk), .D (signal_1083), .Q (signal_2122) ) ;
    buf_clk cell_1449 ( .C (clk), .D (signal_1214), .Q (signal_2124) ) ;
    buf_clk cell_1451 ( .C (clk), .D (signal_1084), .Q (signal_2126) ) ;
    buf_clk cell_1453 ( .C (clk), .D (signal_1211), .Q (signal_2128) ) ;
    buf_clk cell_1455 ( .C (clk), .D (signal_1085), .Q (signal_2130) ) ;
    buf_clk cell_1457 ( .C (clk), .D (signal_1208), .Q (signal_2132) ) ;
    buf_clk cell_1459 ( .C (clk), .D (signal_1086), .Q (signal_2134) ) ;
    buf_clk cell_1461 ( .C (clk), .D (signal_1205), .Q (signal_2136) ) ;
    buf_clk cell_1463 ( .C (clk), .D (signal_1087), .Q (signal_2138) ) ;
    buf_clk cell_1465 ( .C (clk), .D (signal_1202), .Q (signal_2140) ) ;
    buf_clk cell_1467 ( .C (clk), .D (signal_1088), .Q (signal_2142) ) ;
    buf_clk cell_1469 ( .C (clk), .D (signal_1199), .Q (signal_2144) ) ;
    buf_clk cell_1471 ( .C (clk), .D (signal_1089), .Q (signal_2146) ) ;
    buf_clk cell_1473 ( .C (clk), .D (signal_1196), .Q (signal_2148) ) ;
    buf_clk cell_1475 ( .C (clk), .D (signal_1090), .Q (signal_2150) ) ;
    buf_clk cell_1477 ( .C (clk), .D (signal_1193), .Q (signal_2152) ) ;
    buf_clk cell_1479 ( .C (clk), .D (signal_1091), .Q (signal_2154) ) ;
    buf_clk cell_1481 ( .C (clk), .D (signal_1190), .Q (signal_2156) ) ;
    buf_clk cell_1483 ( .C (clk), .D (signal_1092), .Q (signal_2158) ) ;
    buf_clk cell_1485 ( .C (clk), .D (signal_1187), .Q (signal_2160) ) ;
    buf_clk cell_1487 ( .C (clk), .D (signal_1093), .Q (signal_2162) ) ;
    buf_clk cell_1489 ( .C (clk), .D (signal_1184), .Q (signal_2164) ) ;
    buf_clk cell_1491 ( .C (clk), .D (signal_1094), .Q (signal_2166) ) ;
    buf_clk cell_1493 ( .C (clk), .D (signal_1181), .Q (signal_2168) ) ;
    buf_clk cell_1495 ( .C (clk), .D (signal_1095), .Q (signal_2170) ) ;
    buf_clk cell_1497 ( .C (clk), .D (signal_1178), .Q (signal_2172) ) ;
    buf_clk cell_1499 ( .C (clk), .D (signal_1096), .Q (signal_2174) ) ;
    buf_clk cell_1501 ( .C (clk), .D (signal_1175), .Q (signal_2176) ) ;
    buf_clk cell_1503 ( .C (clk), .D (signal_1097), .Q (signal_2178) ) ;
    buf_clk cell_1505 ( .C (clk), .D (signal_1172), .Q (signal_2180) ) ;
    buf_clk cell_1507 ( .C (clk), .D (signal_1098), .Q (signal_2182) ) ;
    buf_clk cell_1509 ( .C (clk), .D (signal_1169), .Q (signal_2184) ) ;
    buf_clk cell_1511 ( .C (clk), .D (signal_1099), .Q (signal_2186) ) ;
    buf_clk cell_1513 ( .C (clk), .D (signal_1166), .Q (signal_2188) ) ;
    buf_clk cell_1515 ( .C (clk), .D (signal_1030), .Q (signal_2190) ) ;
    buf_clk cell_1517 ( .C (clk), .D (signal_1031), .Q (signal_2192) ) ;
    buf_clk cell_1519 ( .C (clk), .D (signal_1032), .Q (signal_2194) ) ;
    buf_clk cell_1521 ( .C (clk), .D (signal_1033), .Q (signal_2196) ) ;
    buf_clk cell_1523 ( .C (clk), .D (signal_1034), .Q (signal_2198) ) ;
    buf_clk cell_1525 ( .C (clk), .D (signal_1035), .Q (signal_2200) ) ;

    /* cells in depth 2 */
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_0 ( .s (signal_1677), .b ({signal_1483, signal_839}), .a ({signal_1681, signal_1679}), .c ({signal_1485, signal_903}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1 ( .s (signal_1677), .b ({signal_1482, signal_838}), .a ({signal_1685, signal_1683}), .c ({signal_1487, signal_902}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_2 ( .s (signal_1677), .b ({signal_1481, signal_837}), .a ({signal_1689, signal_1687}), .c ({signal_1489, signal_901}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3 ( .s (signal_1677), .b ({signal_1480, signal_836}), .a ({signal_1693, signal_1691}), .c ({signal_1491, signal_900}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_4 ( .s (signal_1677), .b ({signal_1479, signal_835}), .a ({signal_1697, signal_1695}), .c ({signal_1493, signal_899}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_5 ( .s (signal_1677), .b ({signal_1478, signal_834}), .a ({signal_1701, signal_1699}), .c ({signal_1495, signal_898}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_6 ( .s (signal_1677), .b ({signal_1477, signal_833}), .a ({signal_1705, signal_1703}), .c ({signal_1497, signal_897}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_7 ( .s (signal_1677), .b ({signal_1476, signal_832}), .a ({signal_1709, signal_1707}), .c ({signal_1499, signal_896}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_8 ( .s (signal_1677), .b ({signal_1475, signal_831}), .a ({signal_1713, signal_1711}), .c ({signal_1501, signal_895}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_9 ( .s (signal_1677), .b ({signal_1474, signal_830}), .a ({signal_1717, signal_1715}), .c ({signal_1503, signal_894}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_10 ( .s (signal_1677), .b ({signal_1473, signal_829}), .a ({signal_1721, signal_1719}), .c ({signal_1505, signal_893}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_11 ( .s (signal_1677), .b ({signal_1472, signal_828}), .a ({signal_1725, signal_1723}), .c ({signal_1507, signal_892}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_12 ( .s (signal_1677), .b ({signal_1471, signal_827}), .a ({signal_1729, signal_1727}), .c ({signal_1509, signal_891}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_13 ( .s (signal_1677), .b ({signal_1470, signal_826}), .a ({signal_1733, signal_1731}), .c ({signal_1511, signal_890}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_14 ( .s (signal_1677), .b ({signal_1469, signal_825}), .a ({signal_1737, signal_1735}), .c ({signal_1513, signal_889}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_15 ( .s (signal_1677), .b ({signal_1468, signal_824}), .a ({signal_1741, signal_1739}), .c ({signal_1515, signal_888}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_16 ( .s (signal_1677), .b ({signal_1467, signal_823}), .a ({signal_1745, signal_1743}), .c ({signal_1517, signal_887}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_17 ( .s (signal_1677), .b ({signal_1466, signal_822}), .a ({signal_1749, signal_1747}), .c ({signal_1519, signal_886}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_18 ( .s (signal_1677), .b ({signal_1465, signal_821}), .a ({signal_1753, signal_1751}), .c ({signal_1521, signal_885}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_19 ( .s (signal_1677), .b ({signal_1464, signal_820}), .a ({signal_1757, signal_1755}), .c ({signal_1523, signal_884}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_20 ( .s (signal_1677), .b ({signal_1463, signal_819}), .a ({signal_1761, signal_1759}), .c ({signal_1525, signal_883}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_21 ( .s (signal_1677), .b ({signal_1462, signal_818}), .a ({signal_1765, signal_1763}), .c ({signal_1527, signal_882}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_22 ( .s (signal_1677), .b ({signal_1461, signal_817}), .a ({signal_1769, signal_1767}), .c ({signal_1529, signal_881}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_23 ( .s (signal_1677), .b ({signal_1460, signal_816}), .a ({signal_1773, signal_1771}), .c ({signal_1531, signal_880}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_24 ( .s (signal_1677), .b ({signal_1459, signal_815}), .a ({signal_1777, signal_1775}), .c ({signal_1533, signal_879}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_25 ( .s (signal_1677), .b ({signal_1458, signal_814}), .a ({signal_1781, signal_1779}), .c ({signal_1535, signal_878}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_26 ( .s (signal_1677), .b ({signal_1457, signal_813}), .a ({signal_1785, signal_1783}), .c ({signal_1537, signal_877}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_27 ( .s (signal_1677), .b ({signal_1456, signal_812}), .a ({signal_1789, signal_1787}), .c ({signal_1539, signal_876}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_28 ( .s (signal_1677), .b ({signal_1455, signal_811}), .a ({signal_1793, signal_1791}), .c ({signal_1541, signal_875}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_29 ( .s (signal_1677), .b ({signal_1454, signal_810}), .a ({signal_1797, signal_1795}), .c ({signal_1543, signal_874}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_30 ( .s (signal_1677), .b ({signal_1453, signal_809}), .a ({signal_1801, signal_1799}), .c ({signal_1545, signal_873}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_31 ( .s (signal_1677), .b ({signal_1452, signal_808}), .a ({signal_1805, signal_1803}), .c ({signal_1547, signal_872}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_32 ( .s (signal_1677), .b ({signal_1451, signal_807}), .a ({signal_1809, signal_1807}), .c ({signal_1549, signal_871}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_33 ( .s (signal_1677), .b ({signal_1450, signal_806}), .a ({signal_1813, signal_1811}), .c ({signal_1551, signal_870}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_34 ( .s (signal_1677), .b ({signal_1449, signal_805}), .a ({signal_1817, signal_1815}), .c ({signal_1553, signal_869}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_35 ( .s (signal_1677), .b ({signal_1448, signal_804}), .a ({signal_1821, signal_1819}), .c ({signal_1555, signal_868}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_36 ( .s (signal_1677), .b ({signal_1447, signal_803}), .a ({signal_1825, signal_1823}), .c ({signal_1557, signal_867}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_37 ( .s (signal_1677), .b ({signal_1446, signal_802}), .a ({signal_1829, signal_1827}), .c ({signal_1559, signal_866}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_38 ( .s (signal_1677), .b ({signal_1445, signal_801}), .a ({signal_1833, signal_1831}), .c ({signal_1561, signal_865}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_39 ( .s (signal_1677), .b ({signal_1444, signal_800}), .a ({signal_1837, signal_1835}), .c ({signal_1563, signal_864}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_40 ( .s (signal_1677), .b ({signal_1443, signal_799}), .a ({signal_1841, signal_1839}), .c ({signal_1565, signal_863}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_41 ( .s (signal_1677), .b ({signal_1442, signal_798}), .a ({signal_1845, signal_1843}), .c ({signal_1567, signal_862}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_42 ( .s (signal_1677), .b ({signal_1441, signal_797}), .a ({signal_1849, signal_1847}), .c ({signal_1569, signal_861}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_43 ( .s (signal_1677), .b ({signal_1440, signal_796}), .a ({signal_1853, signal_1851}), .c ({signal_1571, signal_860}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_44 ( .s (signal_1677), .b ({signal_1439, signal_795}), .a ({signal_1857, signal_1855}), .c ({signal_1573, signal_859}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_45 ( .s (signal_1677), .b ({signal_1438, signal_794}), .a ({signal_1861, signal_1859}), .c ({signal_1575, signal_858}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_46 ( .s (signal_1677), .b ({signal_1437, signal_793}), .a ({signal_1865, signal_1863}), .c ({signal_1577, signal_857}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_47 ( .s (signal_1677), .b ({signal_1436, signal_792}), .a ({signal_1869, signal_1867}), .c ({signal_1579, signal_856}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_48 ( .s (signal_1677), .b ({signal_1435, signal_791}), .a ({signal_1873, signal_1871}), .c ({signal_1581, signal_855}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_49 ( .s (signal_1677), .b ({signal_1434, signal_790}), .a ({signal_1877, signal_1875}), .c ({signal_1583, signal_854}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_50 ( .s (signal_1677), .b ({signal_1433, signal_789}), .a ({signal_1881, signal_1879}), .c ({signal_1585, signal_853}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_51 ( .s (signal_1677), .b ({signal_1432, signal_788}), .a ({signal_1885, signal_1883}), .c ({signal_1587, signal_852}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_52 ( .s (signal_1677), .b ({signal_1431, signal_787}), .a ({signal_1889, signal_1887}), .c ({signal_1589, signal_851}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_53 ( .s (signal_1677), .b ({signal_1430, signal_786}), .a ({signal_1893, signal_1891}), .c ({signal_1591, signal_850}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_54 ( .s (signal_1677), .b ({signal_1429, signal_785}), .a ({signal_1897, signal_1895}), .c ({signal_1593, signal_849}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_55 ( .s (signal_1677), .b ({signal_1428, signal_784}), .a ({signal_1901, signal_1899}), .c ({signal_1595, signal_848}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_56 ( .s (signal_1677), .b ({signal_1427, signal_783}), .a ({signal_1905, signal_1903}), .c ({signal_1597, signal_847}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_57 ( .s (signal_1677), .b ({signal_1426, signal_782}), .a ({signal_1909, signal_1907}), .c ({signal_1599, signal_846}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_58 ( .s (signal_1677), .b ({signal_1425, signal_781}), .a ({signal_1913, signal_1911}), .c ({signal_1601, signal_845}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_59 ( .s (signal_1677), .b ({signal_1424, signal_780}), .a ({signal_1917, signal_1915}), .c ({signal_1603, signal_844}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_60 ( .s (signal_1677), .b ({signal_1423, signal_779}), .a ({signal_1921, signal_1919}), .c ({signal_1605, signal_843}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_61 ( .s (signal_1677), .b ({signal_1422, signal_778}), .a ({signal_1925, signal_1923}), .c ({signal_1607, signal_842}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_62 ( .s (signal_1677), .b ({signal_1421, signal_777}), .a ({signal_1929, signal_1927}), .c ({signal_1609, signal_841}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_63 ( .s (signal_1677), .b ({signal_1420, signal_776}), .a ({signal_1933, signal_1931}), .c ({signal_1611, signal_840}) ) ;
    SkinnyTop_step2_ANF #(.low_latency(0), .pipeline(1)) cell_1000 ( .in0 ({signal_943, signal_940, signal_939, Ciphertext_s0[0], Ciphertext_s0[1], Ciphertext_s0[2], Ciphertext_s0[3], Ciphertext_s0[4], Ciphertext_s0[5], Ciphertext_s0[6], Ciphertext_s0[7], Ciphertext_s0[8], Ciphertext_s0[9], Ciphertext_s0[10], Ciphertext_s0[11], Ciphertext_s0[12], Ciphertext_s0[13], Ciphertext_s0[14], Ciphertext_s0[15], Ciphertext_s0[16], Ciphertext_s0[17], Ciphertext_s0[18], Ciphertext_s0[19], Ciphertext_s0[20], Ciphertext_s0[21], Ciphertext_s0[22], Ciphertext_s0[23], Ciphertext_s0[24], Ciphertext_s0[25], Ciphertext_s0[26], Ciphertext_s0[27], Ciphertext_s0[28], Ciphertext_s0[29], Ciphertext_s0[30], Ciphertext_s0[31], Ciphertext_s0[32], Ciphertext_s0[33], Ciphertext_s0[34], Ciphertext_s0[35], Ciphertext_s0[36], Ciphertext_s0[37], Ciphertext_s0[38], Ciphertext_s0[39], Ciphertext_s0[40], Ciphertext_s0[41], Ciphertext_s0[42], Ciphertext_s0[43], Ciphertext_s0[44], Ciphertext_s0[45], Ciphertext_s0[46], Ciphertext_s0[47], Ciphertext_s0[48], Ciphertext_s0[49], Ciphertext_s0[50], Ciphertext_s0[51], Ciphertext_s0[52], Ciphertext_s0[53], Ciphertext_s0[54], Ciphertext_s0[55], Ciphertext_s0[56], Ciphertext_s0[57], Ciphertext_s0[58], Ciphertext_s0[59], Ciphertext_s0[60], Ciphertext_s0[61], Ciphertext_s0[62], Ciphertext_s0[63], signal_1163, signal_1162, signal_1161, signal_1160, signal_1159, signal_1158, signal_1157, signal_1156, signal_1155, signal_1154, signal_1153, signal_1152, signal_1151, signal_1150, signal_1149, signal_1148, signal_1147, signal_1146, signal_1145, signal_1144, signal_1143, signal_1142, signal_1141, signal_1140, signal_1139, signal_1138, signal_1137, signal_1136, signal_1135, signal_1134, signal_1133, signal_1132, signal_1028, signal_1026, signal_1025, 1'b0}), .in1 ({1'b0, 1'b0, 1'b0, Ciphertext_s1[0], Ciphertext_s1[1], Ciphertext_s1[2], Ciphertext_s1[3], Ciphertext_s1[4], Ciphertext_s1[5], Ciphertext_s1[6], Ciphertext_s1[7], Ciphertext_s1[8], Ciphertext_s1[9], Ciphertext_s1[10], Ciphertext_s1[11], Ciphertext_s1[12], Ciphertext_s1[13], Ciphertext_s1[14], Ciphertext_s1[15], Ciphertext_s1[16], Ciphertext_s1[17], Ciphertext_s1[18], Ciphertext_s1[19], Ciphertext_s1[20], Ciphertext_s1[21], Ciphertext_s1[22], Ciphertext_s1[23], Ciphertext_s1[24], Ciphertext_s1[25], Ciphertext_s1[26], Ciphertext_s1[27], Ciphertext_s1[28], Ciphertext_s1[29], Ciphertext_s1[30], Ciphertext_s1[31], Ciphertext_s1[32], Ciphertext_s1[33], Ciphertext_s1[34], Ciphertext_s1[35], Ciphertext_s1[36], Ciphertext_s1[37], Ciphertext_s1[38], Ciphertext_s1[39], Ciphertext_s1[40], Ciphertext_s1[41], Ciphertext_s1[42], Ciphertext_s1[43], Ciphertext_s1[44], Ciphertext_s1[45], Ciphertext_s1[46], Ciphertext_s1[47], Ciphertext_s1[48], Ciphertext_s1[49], Ciphertext_s1[50], Ciphertext_s1[51], Ciphertext_s1[52], Ciphertext_s1[53], Ciphertext_s1[54], Ciphertext_s1[55], Ciphertext_s1[56], Ciphertext_s1[57], Ciphertext_s1[58], Ciphertext_s1[59], Ciphertext_s1[60], Ciphertext_s1[61], Ciphertext_s1[62], Ciphertext_s1[63], signal_1164, signal_1167, signal_1170, signal_1173, signal_1176, signal_1179, signal_1182, signal_1185, signal_1188, signal_1191, signal_1194, signal_1197, signal_1200, signal_1203, signal_1206, signal_1209, signal_1212, signal_1215, signal_1218, signal_1221, signal_1224, signal_1227, signal_1230, signal_1233, signal_1236, signal_1239, signal_1242, signal_1245, signal_1248, signal_1251, signal_1254, signal_1257, 1'b0, 1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[63], Fresh[62], Fresh[61], Fresh[60], Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48], Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30], Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .out0 ({signal_839, signal_838, signal_837, signal_836, signal_835, signal_834, signal_833, signal_832, signal_831, signal_830, signal_829, signal_828, signal_827, signal_826, signal_825, signal_824, signal_823, signal_822, signal_821, signal_820, signal_819, signal_818, signal_817, signal_816, signal_815, signal_814, signal_813, signal_812, signal_811, signal_810, signal_809, signal_808, signal_807, signal_806, signal_805, signal_804, signal_803, signal_802, signal_801, signal_800, signal_799, signal_798, signal_797, signal_796, signal_795, signal_794, signal_793, signal_792, signal_791, signal_790, signal_789, signal_788, signal_787, signal_786, signal_785, signal_784, signal_783, signal_782, signal_781, signal_780, signal_779, signal_778, signal_777, signal_776}), .out1 ({signal_1483, signal_1482, signal_1481, signal_1480, signal_1479, signal_1478, signal_1477, signal_1476, signal_1475, signal_1474, signal_1473, signal_1472, signal_1471, signal_1470, signal_1469, signal_1468, signal_1467, signal_1466, signal_1465, signal_1464, signal_1463, signal_1462, signal_1461, signal_1460, signal_1459, signal_1458, signal_1457, signal_1456, signal_1455, signal_1454, signal_1453, signal_1452, signal_1451, signal_1450, signal_1449, signal_1448, signal_1447, signal_1446, signal_1445, signal_1444, signal_1443, signal_1442, signal_1441, signal_1440, signal_1439, signal_1438, signal_1437, signal_1436, signal_1435, signal_1434, signal_1433, signal_1432, signal_1431, signal_1430, signal_1429, signal_1428, signal_1427, signal_1426, signal_1425, signal_1424, signal_1423, signal_1422, signal_1421, signal_1420}) ) ;
    buf_clk cell_1002 ( .C (clk), .D (signal_1676), .Q (signal_1677) ) ;
    buf_clk cell_1004 ( .C (clk), .D (signal_1678), .Q (signal_1679) ) ;
    buf_clk cell_1006 ( .C (clk), .D (signal_1680), .Q (signal_1681) ) ;
    buf_clk cell_1008 ( .C (clk), .D (signal_1682), .Q (signal_1683) ) ;
    buf_clk cell_1010 ( .C (clk), .D (signal_1684), .Q (signal_1685) ) ;
    buf_clk cell_1012 ( .C (clk), .D (signal_1686), .Q (signal_1687) ) ;
    buf_clk cell_1014 ( .C (clk), .D (signal_1688), .Q (signal_1689) ) ;
    buf_clk cell_1016 ( .C (clk), .D (signal_1690), .Q (signal_1691) ) ;
    buf_clk cell_1018 ( .C (clk), .D (signal_1692), .Q (signal_1693) ) ;
    buf_clk cell_1020 ( .C (clk), .D (signal_1694), .Q (signal_1695) ) ;
    buf_clk cell_1022 ( .C (clk), .D (signal_1696), .Q (signal_1697) ) ;
    buf_clk cell_1024 ( .C (clk), .D (signal_1698), .Q (signal_1699) ) ;
    buf_clk cell_1026 ( .C (clk), .D (signal_1700), .Q (signal_1701) ) ;
    buf_clk cell_1028 ( .C (clk), .D (signal_1702), .Q (signal_1703) ) ;
    buf_clk cell_1030 ( .C (clk), .D (signal_1704), .Q (signal_1705) ) ;
    buf_clk cell_1032 ( .C (clk), .D (signal_1706), .Q (signal_1707) ) ;
    buf_clk cell_1034 ( .C (clk), .D (signal_1708), .Q (signal_1709) ) ;
    buf_clk cell_1036 ( .C (clk), .D (signal_1710), .Q (signal_1711) ) ;
    buf_clk cell_1038 ( .C (clk), .D (signal_1712), .Q (signal_1713) ) ;
    buf_clk cell_1040 ( .C (clk), .D (signal_1714), .Q (signal_1715) ) ;
    buf_clk cell_1042 ( .C (clk), .D (signal_1716), .Q (signal_1717) ) ;
    buf_clk cell_1044 ( .C (clk), .D (signal_1718), .Q (signal_1719) ) ;
    buf_clk cell_1046 ( .C (clk), .D (signal_1720), .Q (signal_1721) ) ;
    buf_clk cell_1048 ( .C (clk), .D (signal_1722), .Q (signal_1723) ) ;
    buf_clk cell_1050 ( .C (clk), .D (signal_1724), .Q (signal_1725) ) ;
    buf_clk cell_1052 ( .C (clk), .D (signal_1726), .Q (signal_1727) ) ;
    buf_clk cell_1054 ( .C (clk), .D (signal_1728), .Q (signal_1729) ) ;
    buf_clk cell_1056 ( .C (clk), .D (signal_1730), .Q (signal_1731) ) ;
    buf_clk cell_1058 ( .C (clk), .D (signal_1732), .Q (signal_1733) ) ;
    buf_clk cell_1060 ( .C (clk), .D (signal_1734), .Q (signal_1735) ) ;
    buf_clk cell_1062 ( .C (clk), .D (signal_1736), .Q (signal_1737) ) ;
    buf_clk cell_1064 ( .C (clk), .D (signal_1738), .Q (signal_1739) ) ;
    buf_clk cell_1066 ( .C (clk), .D (signal_1740), .Q (signal_1741) ) ;
    buf_clk cell_1068 ( .C (clk), .D (signal_1742), .Q (signal_1743) ) ;
    buf_clk cell_1070 ( .C (clk), .D (signal_1744), .Q (signal_1745) ) ;
    buf_clk cell_1072 ( .C (clk), .D (signal_1746), .Q (signal_1747) ) ;
    buf_clk cell_1074 ( .C (clk), .D (signal_1748), .Q (signal_1749) ) ;
    buf_clk cell_1076 ( .C (clk), .D (signal_1750), .Q (signal_1751) ) ;
    buf_clk cell_1078 ( .C (clk), .D (signal_1752), .Q (signal_1753) ) ;
    buf_clk cell_1080 ( .C (clk), .D (signal_1754), .Q (signal_1755) ) ;
    buf_clk cell_1082 ( .C (clk), .D (signal_1756), .Q (signal_1757) ) ;
    buf_clk cell_1084 ( .C (clk), .D (signal_1758), .Q (signal_1759) ) ;
    buf_clk cell_1086 ( .C (clk), .D (signal_1760), .Q (signal_1761) ) ;
    buf_clk cell_1088 ( .C (clk), .D (signal_1762), .Q (signal_1763) ) ;
    buf_clk cell_1090 ( .C (clk), .D (signal_1764), .Q (signal_1765) ) ;
    buf_clk cell_1092 ( .C (clk), .D (signal_1766), .Q (signal_1767) ) ;
    buf_clk cell_1094 ( .C (clk), .D (signal_1768), .Q (signal_1769) ) ;
    buf_clk cell_1096 ( .C (clk), .D (signal_1770), .Q (signal_1771) ) ;
    buf_clk cell_1098 ( .C (clk), .D (signal_1772), .Q (signal_1773) ) ;
    buf_clk cell_1100 ( .C (clk), .D (signal_1774), .Q (signal_1775) ) ;
    buf_clk cell_1102 ( .C (clk), .D (signal_1776), .Q (signal_1777) ) ;
    buf_clk cell_1104 ( .C (clk), .D (signal_1778), .Q (signal_1779) ) ;
    buf_clk cell_1106 ( .C (clk), .D (signal_1780), .Q (signal_1781) ) ;
    buf_clk cell_1108 ( .C (clk), .D (signal_1782), .Q (signal_1783) ) ;
    buf_clk cell_1110 ( .C (clk), .D (signal_1784), .Q (signal_1785) ) ;
    buf_clk cell_1112 ( .C (clk), .D (signal_1786), .Q (signal_1787) ) ;
    buf_clk cell_1114 ( .C (clk), .D (signal_1788), .Q (signal_1789) ) ;
    buf_clk cell_1116 ( .C (clk), .D (signal_1790), .Q (signal_1791) ) ;
    buf_clk cell_1118 ( .C (clk), .D (signal_1792), .Q (signal_1793) ) ;
    buf_clk cell_1120 ( .C (clk), .D (signal_1794), .Q (signal_1795) ) ;
    buf_clk cell_1122 ( .C (clk), .D (signal_1796), .Q (signal_1797) ) ;
    buf_clk cell_1124 ( .C (clk), .D (signal_1798), .Q (signal_1799) ) ;
    buf_clk cell_1126 ( .C (clk), .D (signal_1800), .Q (signal_1801) ) ;
    buf_clk cell_1128 ( .C (clk), .D (signal_1802), .Q (signal_1803) ) ;
    buf_clk cell_1130 ( .C (clk), .D (signal_1804), .Q (signal_1805) ) ;
    buf_clk cell_1132 ( .C (clk), .D (signal_1806), .Q (signal_1807) ) ;
    buf_clk cell_1134 ( .C (clk), .D (signal_1808), .Q (signal_1809) ) ;
    buf_clk cell_1136 ( .C (clk), .D (signal_1810), .Q (signal_1811) ) ;
    buf_clk cell_1138 ( .C (clk), .D (signal_1812), .Q (signal_1813) ) ;
    buf_clk cell_1140 ( .C (clk), .D (signal_1814), .Q (signal_1815) ) ;
    buf_clk cell_1142 ( .C (clk), .D (signal_1816), .Q (signal_1817) ) ;
    buf_clk cell_1144 ( .C (clk), .D (signal_1818), .Q (signal_1819) ) ;
    buf_clk cell_1146 ( .C (clk), .D (signal_1820), .Q (signal_1821) ) ;
    buf_clk cell_1148 ( .C (clk), .D (signal_1822), .Q (signal_1823) ) ;
    buf_clk cell_1150 ( .C (clk), .D (signal_1824), .Q (signal_1825) ) ;
    buf_clk cell_1152 ( .C (clk), .D (signal_1826), .Q (signal_1827) ) ;
    buf_clk cell_1154 ( .C (clk), .D (signal_1828), .Q (signal_1829) ) ;
    buf_clk cell_1156 ( .C (clk), .D (signal_1830), .Q (signal_1831) ) ;
    buf_clk cell_1158 ( .C (clk), .D (signal_1832), .Q (signal_1833) ) ;
    buf_clk cell_1160 ( .C (clk), .D (signal_1834), .Q (signal_1835) ) ;
    buf_clk cell_1162 ( .C (clk), .D (signal_1836), .Q (signal_1837) ) ;
    buf_clk cell_1164 ( .C (clk), .D (signal_1838), .Q (signal_1839) ) ;
    buf_clk cell_1166 ( .C (clk), .D (signal_1840), .Q (signal_1841) ) ;
    buf_clk cell_1168 ( .C (clk), .D (signal_1842), .Q (signal_1843) ) ;
    buf_clk cell_1170 ( .C (clk), .D (signal_1844), .Q (signal_1845) ) ;
    buf_clk cell_1172 ( .C (clk), .D (signal_1846), .Q (signal_1847) ) ;
    buf_clk cell_1174 ( .C (clk), .D (signal_1848), .Q (signal_1849) ) ;
    buf_clk cell_1176 ( .C (clk), .D (signal_1850), .Q (signal_1851) ) ;
    buf_clk cell_1178 ( .C (clk), .D (signal_1852), .Q (signal_1853) ) ;
    buf_clk cell_1180 ( .C (clk), .D (signal_1854), .Q (signal_1855) ) ;
    buf_clk cell_1182 ( .C (clk), .D (signal_1856), .Q (signal_1857) ) ;
    buf_clk cell_1184 ( .C (clk), .D (signal_1858), .Q (signal_1859) ) ;
    buf_clk cell_1186 ( .C (clk), .D (signal_1860), .Q (signal_1861) ) ;
    buf_clk cell_1188 ( .C (clk), .D (signal_1862), .Q (signal_1863) ) ;
    buf_clk cell_1190 ( .C (clk), .D (signal_1864), .Q (signal_1865) ) ;
    buf_clk cell_1192 ( .C (clk), .D (signal_1866), .Q (signal_1867) ) ;
    buf_clk cell_1194 ( .C (clk), .D (signal_1868), .Q (signal_1869) ) ;
    buf_clk cell_1196 ( .C (clk), .D (signal_1870), .Q (signal_1871) ) ;
    buf_clk cell_1198 ( .C (clk), .D (signal_1872), .Q (signal_1873) ) ;
    buf_clk cell_1200 ( .C (clk), .D (signal_1874), .Q (signal_1875) ) ;
    buf_clk cell_1202 ( .C (clk), .D (signal_1876), .Q (signal_1877) ) ;
    buf_clk cell_1204 ( .C (clk), .D (signal_1878), .Q (signal_1879) ) ;
    buf_clk cell_1206 ( .C (clk), .D (signal_1880), .Q (signal_1881) ) ;
    buf_clk cell_1208 ( .C (clk), .D (signal_1882), .Q (signal_1883) ) ;
    buf_clk cell_1210 ( .C (clk), .D (signal_1884), .Q (signal_1885) ) ;
    buf_clk cell_1212 ( .C (clk), .D (signal_1886), .Q (signal_1887) ) ;
    buf_clk cell_1214 ( .C (clk), .D (signal_1888), .Q (signal_1889) ) ;
    buf_clk cell_1216 ( .C (clk), .D (signal_1890), .Q (signal_1891) ) ;
    buf_clk cell_1218 ( .C (clk), .D (signal_1892), .Q (signal_1893) ) ;
    buf_clk cell_1220 ( .C (clk), .D (signal_1894), .Q (signal_1895) ) ;
    buf_clk cell_1222 ( .C (clk), .D (signal_1896), .Q (signal_1897) ) ;
    buf_clk cell_1224 ( .C (clk), .D (signal_1898), .Q (signal_1899) ) ;
    buf_clk cell_1226 ( .C (clk), .D (signal_1900), .Q (signal_1901) ) ;
    buf_clk cell_1228 ( .C (clk), .D (signal_1902), .Q (signal_1903) ) ;
    buf_clk cell_1230 ( .C (clk), .D (signal_1904), .Q (signal_1905) ) ;
    buf_clk cell_1232 ( .C (clk), .D (signal_1906), .Q (signal_1907) ) ;
    buf_clk cell_1234 ( .C (clk), .D (signal_1908), .Q (signal_1909) ) ;
    buf_clk cell_1236 ( .C (clk), .D (signal_1910), .Q (signal_1911) ) ;
    buf_clk cell_1238 ( .C (clk), .D (signal_1912), .Q (signal_1913) ) ;
    buf_clk cell_1240 ( .C (clk), .D (signal_1914), .Q (signal_1915) ) ;
    buf_clk cell_1242 ( .C (clk), .D (signal_1916), .Q (signal_1917) ) ;
    buf_clk cell_1244 ( .C (clk), .D (signal_1918), .Q (signal_1919) ) ;
    buf_clk cell_1246 ( .C (clk), .D (signal_1920), .Q (signal_1921) ) ;
    buf_clk cell_1248 ( .C (clk), .D (signal_1922), .Q (signal_1923) ) ;
    buf_clk cell_1250 ( .C (clk), .D (signal_1924), .Q (signal_1925) ) ;
    buf_clk cell_1252 ( .C (clk), .D (signal_1926), .Q (signal_1927) ) ;
    buf_clk cell_1254 ( .C (clk), .D (signal_1928), .Q (signal_1929) ) ;
    buf_clk cell_1256 ( .C (clk), .D (signal_1930), .Q (signal_1931) ) ;
    buf_clk cell_1258 ( .C (clk), .D (signal_1932), .Q (signal_1933) ) ;
    buf_clk cell_1260 ( .C (clk), .D (signal_1934), .Q (signal_1935) ) ;
    buf_clk cell_1262 ( .C (clk), .D (signal_1936), .Q (signal_1937) ) ;
    buf_clk cell_1264 ( .C (clk), .D (signal_1938), .Q (signal_1939) ) ;
    buf_clk cell_1266 ( .C (clk), .D (signal_1940), .Q (signal_1941) ) ;
    buf_clk cell_1268 ( .C (clk), .D (signal_1942), .Q (signal_1943) ) ;
    buf_clk cell_1270 ( .C (clk), .D (signal_1944), .Q (signal_1945) ) ;
    buf_clk cell_1272 ( .C (clk), .D (signal_1946), .Q (signal_1947) ) ;
    buf_clk cell_1274 ( .C (clk), .D (signal_1948), .Q (signal_1949) ) ;
    buf_clk cell_1276 ( .C (clk), .D (signal_1950), .Q (signal_1951) ) ;
    buf_clk cell_1278 ( .C (clk), .D (signal_1952), .Q (signal_1953) ) ;
    buf_clk cell_1280 ( .C (clk), .D (signal_1954), .Q (signal_1955) ) ;
    buf_clk cell_1282 ( .C (clk), .D (signal_1956), .Q (signal_1957) ) ;
    buf_clk cell_1284 ( .C (clk), .D (signal_1958), .Q (signal_1959) ) ;
    buf_clk cell_1286 ( .C (clk), .D (signal_1960), .Q (signal_1961) ) ;
    buf_clk cell_1288 ( .C (clk), .D (signal_1962), .Q (signal_1963) ) ;
    buf_clk cell_1290 ( .C (clk), .D (signal_1964), .Q (signal_1965) ) ;
    buf_clk cell_1292 ( .C (clk), .D (signal_1966), .Q (signal_1967) ) ;
    buf_clk cell_1294 ( .C (clk), .D (signal_1968), .Q (signal_1969) ) ;
    buf_clk cell_1296 ( .C (clk), .D (signal_1970), .Q (signal_1971) ) ;
    buf_clk cell_1298 ( .C (clk), .D (signal_1972), .Q (signal_1973) ) ;
    buf_clk cell_1300 ( .C (clk), .D (signal_1974), .Q (signal_1975) ) ;
    buf_clk cell_1302 ( .C (clk), .D (signal_1976), .Q (signal_1977) ) ;
    buf_clk cell_1304 ( .C (clk), .D (signal_1978), .Q (signal_1979) ) ;
    buf_clk cell_1306 ( .C (clk), .D (signal_1980), .Q (signal_1981) ) ;
    buf_clk cell_1308 ( .C (clk), .D (signal_1982), .Q (signal_1983) ) ;
    buf_clk cell_1310 ( .C (clk), .D (signal_1984), .Q (signal_1985) ) ;
    buf_clk cell_1312 ( .C (clk), .D (signal_1986), .Q (signal_1987) ) ;
    buf_clk cell_1314 ( .C (clk), .D (signal_1988), .Q (signal_1989) ) ;
    buf_clk cell_1316 ( .C (clk), .D (signal_1990), .Q (signal_1991) ) ;
    buf_clk cell_1318 ( .C (clk), .D (signal_1992), .Q (signal_1993) ) ;
    buf_clk cell_1320 ( .C (clk), .D (signal_1994), .Q (signal_1995) ) ;
    buf_clk cell_1322 ( .C (clk), .D (signal_1996), .Q (signal_1997) ) ;
    buf_clk cell_1324 ( .C (clk), .D (signal_1998), .Q (signal_1999) ) ;
    buf_clk cell_1326 ( .C (clk), .D (signal_2000), .Q (signal_2001) ) ;
    buf_clk cell_1328 ( .C (clk), .D (signal_2002), .Q (signal_2003) ) ;
    buf_clk cell_1330 ( .C (clk), .D (signal_2004), .Q (signal_2005) ) ;
    buf_clk cell_1332 ( .C (clk), .D (signal_2006), .Q (signal_2007) ) ;
    buf_clk cell_1334 ( .C (clk), .D (signal_2008), .Q (signal_2009) ) ;
    buf_clk cell_1336 ( .C (clk), .D (signal_2010), .Q (signal_2011) ) ;
    buf_clk cell_1338 ( .C (clk), .D (signal_2012), .Q (signal_2013) ) ;
    buf_clk cell_1340 ( .C (clk), .D (signal_2014), .Q (signal_2015) ) ;
    buf_clk cell_1342 ( .C (clk), .D (signal_2016), .Q (signal_2017) ) ;
    buf_clk cell_1344 ( .C (clk), .D (signal_2018), .Q (signal_2019) ) ;
    buf_clk cell_1346 ( .C (clk), .D (signal_2020), .Q (signal_2021) ) ;
    buf_clk cell_1348 ( .C (clk), .D (signal_2022), .Q (signal_2023) ) ;
    buf_clk cell_1350 ( .C (clk), .D (signal_2024), .Q (signal_2025) ) ;
    buf_clk cell_1352 ( .C (clk), .D (signal_2026), .Q (signal_2027) ) ;
    buf_clk cell_1354 ( .C (clk), .D (signal_2028), .Q (signal_2029) ) ;
    buf_clk cell_1356 ( .C (clk), .D (signal_2030), .Q (signal_2031) ) ;
    buf_clk cell_1358 ( .C (clk), .D (signal_2032), .Q (signal_2033) ) ;
    buf_clk cell_1360 ( .C (clk), .D (signal_2034), .Q (signal_2035) ) ;
    buf_clk cell_1362 ( .C (clk), .D (signal_2036), .Q (signal_2037) ) ;
    buf_clk cell_1364 ( .C (clk), .D (signal_2038), .Q (signal_2039) ) ;
    buf_clk cell_1366 ( .C (clk), .D (signal_2040), .Q (signal_2041) ) ;
    buf_clk cell_1368 ( .C (clk), .D (signal_2042), .Q (signal_2043) ) ;
    buf_clk cell_1370 ( .C (clk), .D (signal_2044), .Q (signal_2045) ) ;
    buf_clk cell_1372 ( .C (clk), .D (signal_2046), .Q (signal_2047) ) ;
    buf_clk cell_1374 ( .C (clk), .D (signal_2048), .Q (signal_2049) ) ;
    buf_clk cell_1376 ( .C (clk), .D (signal_2050), .Q (signal_2051) ) ;
    buf_clk cell_1378 ( .C (clk), .D (signal_2052), .Q (signal_2053) ) ;
    buf_clk cell_1380 ( .C (clk), .D (signal_2054), .Q (signal_2055) ) ;
    buf_clk cell_1382 ( .C (clk), .D (signal_2056), .Q (signal_2057) ) ;
    buf_clk cell_1384 ( .C (clk), .D (signal_2058), .Q (signal_2059) ) ;
    buf_clk cell_1386 ( .C (clk), .D (signal_2060), .Q (signal_2061) ) ;
    buf_clk cell_1388 ( .C (clk), .D (signal_2062), .Q (signal_2063) ) ;
    buf_clk cell_1390 ( .C (clk), .D (signal_2064), .Q (signal_2065) ) ;
    buf_clk cell_1392 ( .C (clk), .D (signal_2066), .Q (signal_2067) ) ;
    buf_clk cell_1394 ( .C (clk), .D (signal_2068), .Q (signal_2069) ) ;
    buf_clk cell_1396 ( .C (clk), .D (signal_2070), .Q (signal_2071) ) ;
    buf_clk cell_1398 ( .C (clk), .D (signal_2072), .Q (signal_2073) ) ;
    buf_clk cell_1400 ( .C (clk), .D (signal_2074), .Q (signal_2075) ) ;
    buf_clk cell_1402 ( .C (clk), .D (signal_2076), .Q (signal_2077) ) ;
    buf_clk cell_1404 ( .C (clk), .D (signal_2078), .Q (signal_2079) ) ;
    buf_clk cell_1406 ( .C (clk), .D (signal_2080), .Q (signal_2081) ) ;
    buf_clk cell_1408 ( .C (clk), .D (signal_2082), .Q (signal_2083) ) ;
    buf_clk cell_1410 ( .C (clk), .D (signal_2084), .Q (signal_2085) ) ;
    buf_clk cell_1412 ( .C (clk), .D (signal_2086), .Q (signal_2087) ) ;
    buf_clk cell_1414 ( .C (clk), .D (signal_2088), .Q (signal_2089) ) ;
    buf_clk cell_1416 ( .C (clk), .D (signal_2090), .Q (signal_2091) ) ;
    buf_clk cell_1418 ( .C (clk), .D (signal_2092), .Q (signal_2093) ) ;
    buf_clk cell_1420 ( .C (clk), .D (signal_2094), .Q (signal_2095) ) ;
    buf_clk cell_1422 ( .C (clk), .D (signal_2096), .Q (signal_2097) ) ;
    buf_clk cell_1424 ( .C (clk), .D (signal_2098), .Q (signal_2099) ) ;
    buf_clk cell_1426 ( .C (clk), .D (signal_2100), .Q (signal_2101) ) ;
    buf_clk cell_1428 ( .C (clk), .D (signal_2102), .Q (signal_2103) ) ;
    buf_clk cell_1430 ( .C (clk), .D (signal_2104), .Q (signal_2105) ) ;
    buf_clk cell_1432 ( .C (clk), .D (signal_2106), .Q (signal_2107) ) ;
    buf_clk cell_1434 ( .C (clk), .D (signal_2108), .Q (signal_2109) ) ;
    buf_clk cell_1436 ( .C (clk), .D (signal_2110), .Q (signal_2111) ) ;
    buf_clk cell_1438 ( .C (clk), .D (signal_2112), .Q (signal_2113) ) ;
    buf_clk cell_1440 ( .C (clk), .D (signal_2114), .Q (signal_2115) ) ;
    buf_clk cell_1442 ( .C (clk), .D (signal_2116), .Q (signal_2117) ) ;
    buf_clk cell_1444 ( .C (clk), .D (signal_2118), .Q (signal_2119) ) ;
    buf_clk cell_1446 ( .C (clk), .D (signal_2120), .Q (signal_2121) ) ;
    buf_clk cell_1448 ( .C (clk), .D (signal_2122), .Q (signal_2123) ) ;
    buf_clk cell_1450 ( .C (clk), .D (signal_2124), .Q (signal_2125) ) ;
    buf_clk cell_1452 ( .C (clk), .D (signal_2126), .Q (signal_2127) ) ;
    buf_clk cell_1454 ( .C (clk), .D (signal_2128), .Q (signal_2129) ) ;
    buf_clk cell_1456 ( .C (clk), .D (signal_2130), .Q (signal_2131) ) ;
    buf_clk cell_1458 ( .C (clk), .D (signal_2132), .Q (signal_2133) ) ;
    buf_clk cell_1460 ( .C (clk), .D (signal_2134), .Q (signal_2135) ) ;
    buf_clk cell_1462 ( .C (clk), .D (signal_2136), .Q (signal_2137) ) ;
    buf_clk cell_1464 ( .C (clk), .D (signal_2138), .Q (signal_2139) ) ;
    buf_clk cell_1466 ( .C (clk), .D (signal_2140), .Q (signal_2141) ) ;
    buf_clk cell_1468 ( .C (clk), .D (signal_2142), .Q (signal_2143) ) ;
    buf_clk cell_1470 ( .C (clk), .D (signal_2144), .Q (signal_2145) ) ;
    buf_clk cell_1472 ( .C (clk), .D (signal_2146), .Q (signal_2147) ) ;
    buf_clk cell_1474 ( .C (clk), .D (signal_2148), .Q (signal_2149) ) ;
    buf_clk cell_1476 ( .C (clk), .D (signal_2150), .Q (signal_2151) ) ;
    buf_clk cell_1478 ( .C (clk), .D (signal_2152), .Q (signal_2153) ) ;
    buf_clk cell_1480 ( .C (clk), .D (signal_2154), .Q (signal_2155) ) ;
    buf_clk cell_1482 ( .C (clk), .D (signal_2156), .Q (signal_2157) ) ;
    buf_clk cell_1484 ( .C (clk), .D (signal_2158), .Q (signal_2159) ) ;
    buf_clk cell_1486 ( .C (clk), .D (signal_2160), .Q (signal_2161) ) ;
    buf_clk cell_1488 ( .C (clk), .D (signal_2162), .Q (signal_2163) ) ;
    buf_clk cell_1490 ( .C (clk), .D (signal_2164), .Q (signal_2165) ) ;
    buf_clk cell_1492 ( .C (clk), .D (signal_2166), .Q (signal_2167) ) ;
    buf_clk cell_1494 ( .C (clk), .D (signal_2168), .Q (signal_2169) ) ;
    buf_clk cell_1496 ( .C (clk), .D (signal_2170), .Q (signal_2171) ) ;
    buf_clk cell_1498 ( .C (clk), .D (signal_2172), .Q (signal_2173) ) ;
    buf_clk cell_1500 ( .C (clk), .D (signal_2174), .Q (signal_2175) ) ;
    buf_clk cell_1502 ( .C (clk), .D (signal_2176), .Q (signal_2177) ) ;
    buf_clk cell_1504 ( .C (clk), .D (signal_2178), .Q (signal_2179) ) ;
    buf_clk cell_1506 ( .C (clk), .D (signal_2180), .Q (signal_2181) ) ;
    buf_clk cell_1508 ( .C (clk), .D (signal_2182), .Q (signal_2183) ) ;
    buf_clk cell_1510 ( .C (clk), .D (signal_2184), .Q (signal_2185) ) ;
    buf_clk cell_1512 ( .C (clk), .D (signal_2186), .Q (signal_2187) ) ;
    buf_clk cell_1514 ( .C (clk), .D (signal_2188), .Q (signal_2189) ) ;
    buf_clk cell_1516 ( .C (clk), .D (signal_2190), .Q (signal_2191) ) ;
    buf_clk cell_1518 ( .C (clk), .D (signal_2192), .Q (signal_2193) ) ;
    buf_clk cell_1520 ( .C (clk), .D (signal_2194), .Q (signal_2195) ) ;
    buf_clk cell_1522 ( .C (clk), .D (signal_2196), .Q (signal_2197) ) ;
    buf_clk cell_1524 ( .C (clk), .D (signal_2198), .Q (signal_2199) ) ;
    buf_clk cell_1526 ( .C (clk), .D (signal_2200), .Q (signal_2201) ) ;

    /* register cells */
    reg_masked #(.low_latency(0), .pipeline(1)) cell_65 ( .clk (clk), .D ({signal_1611, signal_840}), .Q ({Ciphertext_s1[63], Ciphertext_s0[63]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_67 ( .clk (clk), .D ({signal_1609, signal_841}), .Q ({Ciphertext_s1[62], Ciphertext_s0[62]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_69 ( .clk (clk), .D ({signal_1607, signal_842}), .Q ({Ciphertext_s1[61], Ciphertext_s0[61]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_71 ( .clk (clk), .D ({signal_1605, signal_843}), .Q ({Ciphertext_s1[60], Ciphertext_s0[60]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_73 ( .clk (clk), .D ({signal_1603, signal_844}), .Q ({Ciphertext_s1[59], Ciphertext_s0[59]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_75 ( .clk (clk), .D ({signal_1601, signal_845}), .Q ({Ciphertext_s1[58], Ciphertext_s0[58]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_77 ( .clk (clk), .D ({signal_1599, signal_846}), .Q ({Ciphertext_s1[57], Ciphertext_s0[57]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_79 ( .clk (clk), .D ({signal_1597, signal_847}), .Q ({Ciphertext_s1[56], Ciphertext_s0[56]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_81 ( .clk (clk), .D ({signal_1595, signal_848}), .Q ({Ciphertext_s1[55], Ciphertext_s0[55]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_83 ( .clk (clk), .D ({signal_1593, signal_849}), .Q ({Ciphertext_s1[54], Ciphertext_s0[54]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_85 ( .clk (clk), .D ({signal_1591, signal_850}), .Q ({Ciphertext_s1[53], Ciphertext_s0[53]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_87 ( .clk (clk), .D ({signal_1589, signal_851}), .Q ({Ciphertext_s1[52], Ciphertext_s0[52]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_89 ( .clk (clk), .D ({signal_1587, signal_852}), .Q ({Ciphertext_s1[51], Ciphertext_s0[51]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_91 ( .clk (clk), .D ({signal_1585, signal_853}), .Q ({Ciphertext_s1[50], Ciphertext_s0[50]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_93 ( .clk (clk), .D ({signal_1583, signal_854}), .Q ({Ciphertext_s1[49], Ciphertext_s0[49]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_95 ( .clk (clk), .D ({signal_1581, signal_855}), .Q ({Ciphertext_s1[48], Ciphertext_s0[48]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_97 ( .clk (clk), .D ({signal_1579, signal_856}), .Q ({Ciphertext_s1[47], Ciphertext_s0[47]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_99 ( .clk (clk), .D ({signal_1577, signal_857}), .Q ({Ciphertext_s1[46], Ciphertext_s0[46]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_101 ( .clk (clk), .D ({signal_1575, signal_858}), .Q ({Ciphertext_s1[45], Ciphertext_s0[45]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_103 ( .clk (clk), .D ({signal_1573, signal_859}), .Q ({Ciphertext_s1[44], Ciphertext_s0[44]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_105 ( .clk (clk), .D ({signal_1571, signal_860}), .Q ({Ciphertext_s1[43], Ciphertext_s0[43]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_107 ( .clk (clk), .D ({signal_1569, signal_861}), .Q ({Ciphertext_s1[42], Ciphertext_s0[42]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_109 ( .clk (clk), .D ({signal_1567, signal_862}), .Q ({Ciphertext_s1[41], Ciphertext_s0[41]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_111 ( .clk (clk), .D ({signal_1565, signal_863}), .Q ({Ciphertext_s1[40], Ciphertext_s0[40]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_113 ( .clk (clk), .D ({signal_1563, signal_864}), .Q ({Ciphertext_s1[39], Ciphertext_s0[39]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_115 ( .clk (clk), .D ({signal_1561, signal_865}), .Q ({Ciphertext_s1[38], Ciphertext_s0[38]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_117 ( .clk (clk), .D ({signal_1559, signal_866}), .Q ({Ciphertext_s1[37], Ciphertext_s0[37]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_119 ( .clk (clk), .D ({signal_1557, signal_867}), .Q ({Ciphertext_s1[36], Ciphertext_s0[36]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_121 ( .clk (clk), .D ({signal_1555, signal_868}), .Q ({Ciphertext_s1[35], Ciphertext_s0[35]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_123 ( .clk (clk), .D ({signal_1553, signal_869}), .Q ({Ciphertext_s1[34], Ciphertext_s0[34]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_125 ( .clk (clk), .D ({signal_1551, signal_870}), .Q ({Ciphertext_s1[33], Ciphertext_s0[33]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_127 ( .clk (clk), .D ({signal_1549, signal_871}), .Q ({Ciphertext_s1[32], Ciphertext_s0[32]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_129 ( .clk (clk), .D ({signal_1547, signal_872}), .Q ({Ciphertext_s1[31], Ciphertext_s0[31]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_131 ( .clk (clk), .D ({signal_1545, signal_873}), .Q ({Ciphertext_s1[30], Ciphertext_s0[30]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_133 ( .clk (clk), .D ({signal_1543, signal_874}), .Q ({Ciphertext_s1[29], Ciphertext_s0[29]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_135 ( .clk (clk), .D ({signal_1541, signal_875}), .Q ({Ciphertext_s1[28], Ciphertext_s0[28]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_137 ( .clk (clk), .D ({signal_1539, signal_876}), .Q ({Ciphertext_s1[27], Ciphertext_s0[27]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_139 ( .clk (clk), .D ({signal_1537, signal_877}), .Q ({Ciphertext_s1[26], Ciphertext_s0[26]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_141 ( .clk (clk), .D ({signal_1535, signal_878}), .Q ({Ciphertext_s1[25], Ciphertext_s0[25]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_143 ( .clk (clk), .D ({signal_1533, signal_879}), .Q ({Ciphertext_s1[24], Ciphertext_s0[24]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_145 ( .clk (clk), .D ({signal_1531, signal_880}), .Q ({Ciphertext_s1[23], Ciphertext_s0[23]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_147 ( .clk (clk), .D ({signal_1529, signal_881}), .Q ({Ciphertext_s1[22], Ciphertext_s0[22]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_149 ( .clk (clk), .D ({signal_1527, signal_882}), .Q ({Ciphertext_s1[21], Ciphertext_s0[21]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_151 ( .clk (clk), .D ({signal_1525, signal_883}), .Q ({Ciphertext_s1[20], Ciphertext_s0[20]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_153 ( .clk (clk), .D ({signal_1523, signal_884}), .Q ({Ciphertext_s1[19], Ciphertext_s0[19]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_155 ( .clk (clk), .D ({signal_1521, signal_885}), .Q ({Ciphertext_s1[18], Ciphertext_s0[18]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_157 ( .clk (clk), .D ({signal_1519, signal_886}), .Q ({Ciphertext_s1[17], Ciphertext_s0[17]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_159 ( .clk (clk), .D ({signal_1517, signal_887}), .Q ({Ciphertext_s1[16], Ciphertext_s0[16]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_161 ( .clk (clk), .D ({signal_1515, signal_888}), .Q ({Ciphertext_s1[15], Ciphertext_s0[15]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_163 ( .clk (clk), .D ({signal_1513, signal_889}), .Q ({Ciphertext_s1[14], Ciphertext_s0[14]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_165 ( .clk (clk), .D ({signal_1511, signal_890}), .Q ({Ciphertext_s1[13], Ciphertext_s0[13]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_167 ( .clk (clk), .D ({signal_1509, signal_891}), .Q ({Ciphertext_s1[12], Ciphertext_s0[12]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_169 ( .clk (clk), .D ({signal_1507, signal_892}), .Q ({Ciphertext_s1[11], Ciphertext_s0[11]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_171 ( .clk (clk), .D ({signal_1505, signal_893}), .Q ({Ciphertext_s1[10], Ciphertext_s0[10]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_173 ( .clk (clk), .D ({signal_1503, signal_894}), .Q ({Ciphertext_s1[9], Ciphertext_s0[9]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_175 ( .clk (clk), .D ({signal_1501, signal_895}), .Q ({Ciphertext_s1[8], Ciphertext_s0[8]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_177 ( .clk (clk), .D ({signal_1499, signal_896}), .Q ({Ciphertext_s1[7], Ciphertext_s0[7]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_179 ( .clk (clk), .D ({signal_1497, signal_897}), .Q ({Ciphertext_s1[6], Ciphertext_s0[6]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_181 ( .clk (clk), .D ({signal_1495, signal_898}), .Q ({Ciphertext_s1[5], Ciphertext_s0[5]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_183 ( .clk (clk), .D ({signal_1493, signal_899}), .Q ({Ciphertext_s1[4], Ciphertext_s0[4]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_185 ( .clk (clk), .D ({signal_1491, signal_900}), .Q ({Ciphertext_s1[3], Ciphertext_s0[3]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_187 ( .clk (clk), .D ({signal_1489, signal_901}), .Q ({Ciphertext_s1[2], Ciphertext_s0[2]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_189 ( .clk (clk), .D ({signal_1487, signal_902}), .Q ({Ciphertext_s1[1], Ciphertext_s0[1]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_191 ( .clk (clk), .D ({signal_1485, signal_903}), .Q ({Ciphertext_s1[0], Ciphertext_s0[0]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_834 ( .clk (clk), .D ({signal_1937, signal_1935}), .Q ({signal_1257, signal_1132}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_836 ( .clk (clk), .D ({signal_1941, signal_1939}), .Q ({signal_1254, signal_1133}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_838 ( .clk (clk), .D ({signal_1945, signal_1943}), .Q ({signal_1251, signal_1134}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_840 ( .clk (clk), .D ({signal_1949, signal_1947}), .Q ({signal_1248, signal_1135}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_842 ( .clk (clk), .D ({signal_1953, signal_1951}), .Q ({signal_1245, signal_1136}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_844 ( .clk (clk), .D ({signal_1957, signal_1955}), .Q ({signal_1242, signal_1137}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_846 ( .clk (clk), .D ({signal_1961, signal_1959}), .Q ({signal_1239, signal_1138}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_848 ( .clk (clk), .D ({signal_1965, signal_1963}), .Q ({signal_1236, signal_1139}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_850 ( .clk (clk), .D ({signal_1969, signal_1967}), .Q ({signal_1233, signal_1140}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_852 ( .clk (clk), .D ({signal_1973, signal_1971}), .Q ({signal_1230, signal_1141}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_854 ( .clk (clk), .D ({signal_1977, signal_1975}), .Q ({signal_1227, signal_1142}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_856 ( .clk (clk), .D ({signal_1981, signal_1979}), .Q ({signal_1224, signal_1143}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_858 ( .clk (clk), .D ({signal_1985, signal_1983}), .Q ({signal_1221, signal_1144}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_860 ( .clk (clk), .D ({signal_1989, signal_1987}), .Q ({signal_1218, signal_1145}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_862 ( .clk (clk), .D ({signal_1993, signal_1991}), .Q ({signal_1215, signal_1146}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_864 ( .clk (clk), .D ({signal_1997, signal_1995}), .Q ({signal_1212, signal_1147}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_866 ( .clk (clk), .D ({signal_2001, signal_1999}), .Q ({signal_1209, signal_1148}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_868 ( .clk (clk), .D ({signal_2005, signal_2003}), .Q ({signal_1206, signal_1149}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_870 ( .clk (clk), .D ({signal_2009, signal_2007}), .Q ({signal_1203, signal_1150}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_872 ( .clk (clk), .D ({signal_2013, signal_2011}), .Q ({signal_1200, signal_1151}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_874 ( .clk (clk), .D ({signal_2017, signal_2015}), .Q ({signal_1197, signal_1152}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_876 ( .clk (clk), .D ({signal_2021, signal_2019}), .Q ({signal_1194, signal_1153}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_878 ( .clk (clk), .D ({signal_2025, signal_2023}), .Q ({signal_1191, signal_1154}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_880 ( .clk (clk), .D ({signal_2029, signal_2027}), .Q ({signal_1188, signal_1155}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_882 ( .clk (clk), .D ({signal_2033, signal_2031}), .Q ({signal_1185, signal_1156}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_884 ( .clk (clk), .D ({signal_2037, signal_2035}), .Q ({signal_1182, signal_1157}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_886 ( .clk (clk), .D ({signal_2041, signal_2039}), .Q ({signal_1179, signal_1158}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_888 ( .clk (clk), .D ({signal_2045, signal_2043}), .Q ({signal_1176, signal_1159}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_890 ( .clk (clk), .D ({signal_2049, signal_2047}), .Q ({signal_1173, signal_1160}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_892 ( .clk (clk), .D ({signal_2053, signal_2051}), .Q ({signal_1170, signal_1161}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_894 ( .clk (clk), .D ({signal_2057, signal_2055}), .Q ({signal_1167, signal_1162}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_896 ( .clk (clk), .D ({signal_2061, signal_2059}), .Q ({signal_1164, signal_1163}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_898 ( .clk (clk), .D ({signal_2065, signal_2063}), .Q ({signal_1329, signal_1108}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_900 ( .clk (clk), .D ({signal_2069, signal_2067}), .Q ({signal_1326, signal_1109}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_902 ( .clk (clk), .D ({signal_2073, signal_2071}), .Q ({signal_1323, signal_1110}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_904 ( .clk (clk), .D ({signal_2077, signal_2075}), .Q ({signal_1320, signal_1111}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_906 ( .clk (clk), .D ({signal_2081, signal_2079}), .Q ({signal_1353, signal_1100}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_908 ( .clk (clk), .D ({signal_2085, signal_2083}), .Q ({signal_1350, signal_1101}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_910 ( .clk (clk), .D ({signal_2089, signal_2087}), .Q ({signal_1347, signal_1102}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_912 ( .clk (clk), .D ({signal_2093, signal_2091}), .Q ({signal_1344, signal_1103}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_914 ( .clk (clk), .D ({signal_2097, signal_2095}), .Q ({signal_1305, signal_1116}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_916 ( .clk (clk), .D ({signal_2101, signal_2099}), .Q ({signal_1302, signal_1117}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_918 ( .clk (clk), .D ({signal_2105, signal_2103}), .Q ({signal_1299, signal_1118}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_920 ( .clk (clk), .D ({signal_2109, signal_2107}), .Q ({signal_1296, signal_1119}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_922 ( .clk (clk), .D ({signal_2113, signal_2111}), .Q ({signal_1269, signal_1128}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_924 ( .clk (clk), .D ({signal_2117, signal_2115}), .Q ({signal_1266, signal_1129}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_926 ( .clk (clk), .D ({signal_2121, signal_2119}), .Q ({signal_1263, signal_1130}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_928 ( .clk (clk), .D ({signal_2125, signal_2123}), .Q ({signal_1260, signal_1131}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_930 ( .clk (clk), .D ({signal_2129, signal_2127}), .Q ({signal_1281, signal_1124}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_932 ( .clk (clk), .D ({signal_2133, signal_2131}), .Q ({signal_1278, signal_1125}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_934 ( .clk (clk), .D ({signal_2137, signal_2135}), .Q ({signal_1275, signal_1126}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_936 ( .clk (clk), .D ({signal_2141, signal_2139}), .Q ({signal_1272, signal_1127}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_938 ( .clk (clk), .D ({signal_2145, signal_2143}), .Q ({signal_1317, signal_1112}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_940 ( .clk (clk), .D ({signal_2149, signal_2147}), .Q ({signal_1314, signal_1113}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_942 ( .clk (clk), .D ({signal_2153, signal_2151}), .Q ({signal_1311, signal_1114}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_944 ( .clk (clk), .D ({signal_2157, signal_2155}), .Q ({signal_1308, signal_1115}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_946 ( .clk (clk), .D ({signal_2161, signal_2159}), .Q ({signal_1293, signal_1120}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_948 ( .clk (clk), .D ({signal_2165, signal_2163}), .Q ({signal_1290, signal_1121}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_950 ( .clk (clk), .D ({signal_2169, signal_2167}), .Q ({signal_1287, signal_1122}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_952 ( .clk (clk), .D ({signal_2173, signal_2171}), .Q ({signal_1284, signal_1123}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_954 ( .clk (clk), .D ({signal_2177, signal_2175}), .Q ({signal_1341, signal_1104}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_956 ( .clk (clk), .D ({signal_2181, signal_2179}), .Q ({signal_1338, signal_1105}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_958 ( .clk (clk), .D ({signal_2185, signal_2183}), .Q ({signal_1335, signal_1106}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_960 ( .clk (clk), .D ({signal_2189, signal_2187}), .Q ({signal_1332, signal_1107}) ) ;
    DFF_X1 cell_968 ( .CK (clk), .D (signal_2191), .Q (signal_939), .QN () ) ;
    DFF_X1 cell_970 ( .CK (clk), .D (signal_2193), .Q (signal_940), .QN () ) ;
    DFF_X1 cell_972 ( .CK (clk), .D (signal_2195), .Q (signal_1025), .QN () ) ;
    DFF_X1 cell_974 ( .CK (clk), .D (signal_2197), .Q (signal_1026), .QN () ) ;
    DFF_X1 cell_976 ( .CK (clk), .D (signal_2199), .Q (signal_943), .QN () ) ;
    DFF_X1 cell_978 ( .CK (clk), .D (signal_2201), .Q (signal_1028), .QN () ) ;
endmodule
