/* modified netlist. Source: module LED in file /LED_round-based/AGEMA/LED.v */
/* clock gating is added to the circuit, the latency increased 16 time(s)  */

module LED_HPC2_BDDsylvan_ClockGating_d1 (IN_plaintext_s0, IN_key_s0, IN_reset, CLK, IN_key_s1, IN_plaintext_s1, Fresh, OUT_ciphertext_s0, OUT_done, OUT_ciphertext_s1, Synch);
    input [63:0] IN_plaintext_s0 ;
    input [127:0] IN_key_s0 ;
    input IN_reset ;
    input CLK ;
    input [127:0] IN_key_s1 ;
    input [63:0] IN_plaintext_s1 ;
    input [597:0] Fresh ;
    output [63:0] OUT_ciphertext_s0 ;
    output OUT_done ;
    output [63:0] OUT_ciphertext_s1 ;
    output Synch ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_285 ;
    wire signal_286 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_295 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_356 ;
    wire signal_375 ;
    wire signal_394 ;
    wire signal_413 ;
    wire signal_432 ;
    wire signal_451 ;
    wire signal_470 ;
    wire signal_489 ;
    wire signal_508 ;
    wire signal_527 ;
    wire signal_546 ;
    wire signal_565 ;
    wire signal_584 ;
    wire signal_603 ;
    wire signal_622 ;
    wire signal_641 ;
    wire signal_656 ;
    wire signal_657 ;
    wire signal_658 ;
    wire signal_659 ;
    wire signal_660 ;
    wire signal_661 ;
    wire signal_662 ;
    wire signal_663 ;
    wire signal_664 ;
    wire signal_665 ;
    wire signal_666 ;
    wire signal_667 ;
    wire signal_668 ;
    wire signal_669 ;
    wire signal_670 ;
    wire signal_671 ;
    wire signal_672 ;
    wire signal_673 ;
    wire signal_674 ;
    wire signal_675 ;
    wire signal_676 ;
    wire signal_677 ;
    wire signal_678 ;
    wire signal_679 ;
    wire signal_680 ;
    wire signal_681 ;
    wire signal_682 ;
    wire signal_683 ;
    wire signal_684 ;
    wire signal_685 ;
    wire signal_686 ;
    wire signal_687 ;
    wire signal_688 ;
    wire signal_689 ;
    wire signal_690 ;
    wire signal_691 ;
    wire signal_692 ;
    wire signal_693 ;
    wire signal_694 ;
    wire signal_695 ;
    wire signal_696 ;
    wire signal_697 ;
    wire signal_698 ;
    wire signal_699 ;
    wire signal_700 ;
    wire signal_701 ;
    wire signal_702 ;
    wire signal_703 ;
    wire signal_704 ;
    wire signal_705 ;
    wire signal_706 ;
    wire signal_707 ;
    wire signal_708 ;
    wire signal_709 ;
    wire signal_710 ;
    wire signal_711 ;
    wire signal_712 ;
    wire signal_713 ;
    wire signal_714 ;
    wire signal_715 ;
    wire signal_716 ;
    wire signal_717 ;
    wire signal_718 ;
    wire signal_719 ;
    wire signal_720 ;
    wire signal_721 ;
    wire signal_722 ;
    wire signal_723 ;
    wire signal_724 ;
    wire signal_725 ;
    wire signal_726 ;
    wire signal_727 ;
    wire signal_728 ;
    wire signal_729 ;
    wire signal_730 ;
    wire signal_731 ;
    wire signal_732 ;
    wire signal_733 ;
    wire signal_734 ;
    wire signal_735 ;
    wire signal_736 ;
    wire signal_737 ;
    wire signal_738 ;
    wire signal_739 ;
    wire signal_740 ;
    wire signal_741 ;
    wire signal_742 ;
    wire signal_743 ;
    wire signal_744 ;
    wire signal_745 ;
    wire signal_746 ;
    wire signal_747 ;
    wire signal_748 ;
    wire signal_749 ;
    wire signal_750 ;
    wire signal_751 ;
    wire signal_752 ;
    wire signal_753 ;
    wire signal_754 ;
    wire signal_755 ;
    wire signal_756 ;
    wire signal_757 ;
    wire signal_758 ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_768 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_771 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_774 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_777 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_780 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_783 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_786 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_789 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_792 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_879 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_885 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_888 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_891 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_894 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_897 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_900 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_903 ;
    wire signal_904 ;
    wire signal_905 ;
    wire signal_906 ;
    wire signal_907 ;
    wire signal_908 ;
    wire signal_909 ;
    wire signal_910 ;
    wire signal_911 ;
    wire signal_912 ;
    wire signal_914 ;
    wire signal_915 ;
    wire signal_916 ;
    wire signal_918 ;
    wire signal_919 ;
    wire signal_920 ;
    wire signal_922 ;
    wire signal_923 ;
    wire signal_924 ;
    wire signal_926 ;
    wire signal_927 ;
    wire signal_928 ;
    wire signal_929 ;
    wire signal_930 ;
    wire signal_932 ;
    wire signal_933 ;
    wire signal_934 ;
    wire signal_936 ;
    wire signal_937 ;
    wire signal_938 ;
    wire signal_940 ;
    wire signal_941 ;
    wire signal_942 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1020 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1023 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1276 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1279 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1282 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1285 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1288 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1294 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1297 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1300 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1303 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1309 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1494 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1499 ;
    wire signal_1500 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1503 ;
    wire signal_1504 ;
    wire signal_1505 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1509 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1512 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1518 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1521 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1527 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1530 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1536 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1539 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1564 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1623 ;
    wire signal_1624 ;
    wire signal_1625 ;
    wire signal_1626 ;
    wire signal_1627 ;
    wire signal_1628 ;
    wire signal_1629 ;
    wire signal_1630 ;
    wire signal_1631 ;
    wire signal_1632 ;
    wire signal_1633 ;
    wire signal_1634 ;
    wire signal_1635 ;
    wire signal_1636 ;
    wire signal_1637 ;
    wire signal_1638 ;
    wire signal_1639 ;
    wire signal_1640 ;
    wire signal_1641 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1657 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1660 ;
    wire signal_1661 ;
    wire signal_1662 ;
    wire signal_1663 ;
    wire signal_1664 ;
    wire signal_1665 ;
    wire signal_1666 ;
    wire signal_1667 ;
    wire signal_1668 ;
    wire signal_1669 ;
    wire signal_1670 ;
    wire signal_1671 ;
    wire signal_1672 ;
    wire signal_1673 ;
    wire signal_1674 ;
    wire signal_1675 ;
    wire signal_1676 ;
    wire signal_1677 ;
    wire signal_1678 ;
    wire signal_1679 ;
    wire signal_1680 ;
    wire signal_1681 ;
    wire signal_1682 ;
    wire signal_1683 ;
    wire signal_1684 ;
    wire signal_1685 ;
    wire signal_1686 ;
    wire signal_1687 ;
    wire signal_1688 ;
    wire signal_1689 ;
    wire signal_1690 ;
    wire signal_1691 ;
    wire signal_1692 ;
    wire signal_1693 ;
    wire signal_1694 ;
    wire signal_1695 ;
    wire signal_1696 ;
    wire signal_1697 ;
    wire signal_1698 ;
    wire signal_1699 ;
    wire signal_1700 ;
    wire signal_1701 ;
    wire signal_1702 ;
    wire signal_1703 ;
    wire signal_1704 ;
    wire signal_1705 ;
    wire signal_1706 ;
    wire signal_1707 ;
    wire signal_1708 ;
    wire signal_1709 ;
    wire signal_1710 ;
    wire signal_1711 ;
    wire signal_1712 ;
    wire signal_1713 ;
    wire signal_1714 ;
    wire signal_1715 ;
    wire signal_1716 ;
    wire signal_1717 ;
    wire signal_1718 ;
    wire signal_1719 ;
    wire signal_1720 ;
    wire signal_1721 ;
    wire signal_1722 ;
    wire signal_1723 ;
    wire signal_1724 ;
    wire signal_1725 ;
    wire signal_1726 ;
    wire signal_1727 ;
    wire signal_1728 ;
    wire signal_1729 ;
    wire signal_1730 ;
    wire signal_1731 ;
    wire signal_1732 ;
    wire signal_1733 ;
    wire signal_1734 ;
    wire signal_1735 ;
    wire signal_1736 ;
    wire signal_1737 ;
    wire signal_1738 ;
    wire signal_1739 ;
    wire signal_1740 ;
    wire signal_1741 ;
    wire signal_1742 ;
    wire signal_1743 ;
    wire signal_1744 ;
    wire signal_1745 ;
    wire signal_1746 ;
    wire signal_1747 ;
    wire signal_1748 ;
    wire signal_1749 ;
    wire signal_1750 ;
    wire signal_1751 ;
    wire signal_1752 ;
    wire signal_1753 ;
    wire signal_1754 ;
    wire signal_1755 ;
    wire signal_1756 ;
    wire signal_1757 ;
    wire signal_1758 ;
    wire signal_1759 ;
    wire signal_1760 ;
    wire signal_1761 ;
    wire signal_1762 ;
    wire signal_1763 ;
    wire signal_1764 ;
    wire signal_1765 ;
    wire signal_1766 ;
    wire signal_1767 ;
    wire signal_1768 ;
    wire signal_1769 ;
    wire signal_1770 ;
    wire signal_1771 ;
    wire signal_1772 ;
    wire signal_1773 ;
    wire signal_1774 ;
    wire signal_1775 ;
    wire signal_1776 ;
    wire signal_1777 ;
    wire signal_1778 ;
    wire signal_1779 ;
    wire signal_1780 ;
    wire signal_1781 ;
    wire signal_1782 ;
    wire signal_1783 ;
    wire signal_1784 ;
    wire signal_1785 ;
    wire signal_1786 ;
    wire signal_1787 ;
    wire signal_1788 ;
    wire signal_1789 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1792 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1795 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1813 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1844 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1856 ;
    wire signal_1859 ;
    wire signal_1862 ;
    wire signal_1865 ;
    wire signal_1868 ;
    wire signal_1871 ;
    wire signal_1874 ;
    wire signal_1877 ;
    wire signal_1880 ;
    wire signal_1883 ;
    wire signal_1886 ;
    wire signal_1889 ;
    wire signal_1892 ;
    wire signal_1894 ;
    wire signal_1896 ;
    wire signal_1898 ;
    wire signal_1900 ;
    wire signal_1902 ;
    wire signal_1904 ;
    wire signal_1906 ;
    wire signal_1908 ;
    wire signal_1910 ;
    wire signal_1912 ;
    wire signal_1914 ;
    wire signal_1916 ;
    wire signal_1918 ;
    wire signal_1921 ;
    wire signal_1924 ;
    wire signal_1927 ;
    wire signal_1930 ;
    wire signal_1933 ;
    wire signal_1936 ;
    wire signal_1939 ;
    wire signal_1942 ;
    wire signal_1945 ;
    wire signal_1948 ;
    wire signal_1951 ;
    wire signal_1954 ;
    wire signal_1957 ;
    wire signal_1960 ;
    wire signal_1963 ;
    wire signal_1966 ;
    wire signal_1969 ;
    wire signal_1972 ;
    wire signal_1975 ;
    wire signal_1978 ;
    wire signal_1981 ;
    wire signal_1984 ;
    wire signal_1987 ;
    wire signal_1990 ;
    wire signal_1993 ;
    wire signal_1996 ;
    wire signal_1999 ;
    wire signal_2002 ;
    wire signal_2005 ;
    wire signal_2008 ;
    wire signal_2011 ;
    wire signal_2014 ;
    wire signal_2017 ;
    wire signal_2020 ;
    wire signal_2023 ;
    wire signal_2026 ;
    wire signal_2029 ;
    wire signal_2032 ;
    wire signal_2035 ;
    wire signal_2038 ;
    wire signal_2041 ;
    wire signal_2044 ;
    wire signal_2047 ;
    wire signal_2050 ;
    wire signal_2053 ;
    wire signal_2056 ;
    wire signal_2059 ;
    wire signal_2062 ;
    wire signal_2065 ;
    wire signal_2068 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2080 ;
    wire signal_2082 ;
    wire signal_2084 ;
    wire signal_2086 ;
    wire signal_2088 ;
    wire signal_2090 ;
    wire signal_2092 ;
    wire signal_2094 ;
    wire signal_2096 ;
    wire signal_2098 ;
    wire signal_2100 ;
    wire signal_2102 ;
    wire signal_2104 ;
    wire signal_2106 ;
    wire signal_2108 ;
    wire signal_2110 ;
    wire signal_2112 ;
    wire signal_2114 ;
    wire signal_2116 ;
    wire signal_2118 ;
    wire signal_2120 ;
    wire signal_2122 ;
    wire signal_2124 ;
    wire signal_2126 ;
    wire signal_2128 ;
    wire signal_2130 ;
    wire signal_2132 ;
    wire signal_2134 ;
    wire signal_2136 ;
    wire signal_2138 ;
    wire signal_2140 ;
    wire signal_2142 ;
    wire signal_2144 ;
    wire signal_2146 ;
    wire signal_2148 ;
    wire signal_2150 ;
    wire signal_2152 ;
    wire signal_2154 ;
    wire signal_2156 ;
    wire signal_2158 ;
    wire signal_2160 ;
    wire signal_2162 ;
    wire signal_2164 ;
    wire signal_2166 ;
    wire signal_2168 ;
    wire signal_2170 ;
    wire signal_2172 ;
    wire signal_2174 ;
    wire signal_2176 ;
    wire signal_2178 ;
    wire signal_2180 ;
    wire signal_2181 ;
    wire signal_2182 ;
    wire signal_2183 ;
    wire signal_2184 ;
    wire signal_2185 ;
    wire signal_2186 ;
    wire signal_2187 ;
    wire signal_2188 ;
    wire signal_2189 ;
    wire signal_2190 ;
    wire signal_2191 ;
    wire signal_2192 ;
    wire signal_2193 ;
    wire signal_2194 ;
    wire signal_2195 ;
    wire signal_2196 ;
    wire signal_2197 ;
    wire signal_2198 ;
    wire signal_2199 ;
    wire signal_2200 ;
    wire signal_2201 ;
    wire signal_2202 ;
    wire signal_2203 ;
    wire signal_2204 ;
    wire signal_2205 ;
    wire signal_2206 ;
    wire signal_2207 ;
    wire signal_2208 ;
    wire signal_2209 ;
    wire signal_2210 ;
    wire signal_2211 ;
    wire signal_2212 ;
    wire signal_2213 ;
    wire signal_2214 ;
    wire signal_2215 ;
    wire signal_2216 ;
    wire signal_2217 ;
    wire signal_2218 ;
    wire signal_2219 ;
    wire signal_2220 ;
    wire signal_2221 ;
    wire signal_2222 ;
    wire signal_2223 ;
    wire signal_2224 ;
    wire signal_2225 ;
    wire signal_2226 ;
    wire signal_2227 ;
    wire signal_2228 ;
    wire signal_2229 ;
    wire signal_2230 ;
    wire signal_2231 ;
    wire signal_2232 ;
    wire signal_2233 ;
    wire signal_2234 ;
    wire signal_2235 ;
    wire signal_2236 ;
    wire signal_2237 ;
    wire signal_2238 ;
    wire signal_2239 ;
    wire signal_2240 ;
    wire signal_2241 ;
    wire signal_2242 ;
    wire signal_2243 ;
    wire signal_2244 ;
    wire signal_2245 ;
    wire signal_2246 ;
    wire signal_2247 ;
    wire signal_2248 ;
    wire signal_2249 ;
    wire signal_2250 ;
    wire signal_2251 ;
    wire signal_2252 ;
    wire signal_2253 ;
    wire signal_2254 ;
    wire signal_2255 ;
    wire signal_2256 ;
    wire signal_2257 ;
    wire signal_2258 ;
    wire signal_2259 ;
    wire signal_2260 ;
    wire signal_2261 ;
    wire signal_2262 ;
    wire signal_2263 ;
    wire signal_2264 ;
    wire signal_2265 ;
    wire signal_2266 ;
    wire signal_2267 ;
    wire signal_2268 ;
    wire signal_2269 ;
    wire signal_2270 ;
    wire signal_2271 ;
    wire signal_2272 ;
    wire signal_2273 ;
    wire signal_2274 ;
    wire signal_2275 ;
    wire signal_2276 ;
    wire signal_2277 ;
    wire signal_2278 ;
    wire signal_2279 ;
    wire signal_2280 ;
    wire signal_2281 ;
    wire signal_2282 ;
    wire signal_2283 ;
    wire signal_2284 ;
    wire signal_2285 ;
    wire signal_2286 ;
    wire signal_2287 ;
    wire signal_2288 ;
    wire signal_2289 ;
    wire signal_2290 ;
    wire signal_2291 ;
    wire signal_2292 ;
    wire signal_2293 ;
    wire signal_2294 ;
    wire signal_2295 ;
    wire signal_2296 ;
    wire signal_2297 ;
    wire signal_2298 ;
    wire signal_2299 ;
    wire signal_2300 ;
    wire signal_2301 ;
    wire signal_2302 ;
    wire signal_2303 ;
    wire signal_2304 ;
    wire signal_2305 ;
    wire signal_2306 ;
    wire signal_2307 ;
    wire signal_2308 ;
    wire signal_2309 ;
    wire signal_2310 ;
    wire signal_2311 ;
    wire signal_2312 ;
    wire signal_2313 ;
    wire signal_2314 ;
    wire signal_2315 ;
    wire signal_2316 ;
    wire signal_2317 ;
    wire signal_2318 ;
    wire signal_2319 ;
    wire signal_2320 ;
    wire signal_2321 ;
    wire signal_2322 ;
    wire signal_2323 ;
    wire signal_2324 ;
    wire signal_2325 ;
    wire signal_2326 ;
    wire signal_2327 ;
    wire signal_2328 ;
    wire signal_2329 ;
    wire signal_2330 ;
    wire signal_2331 ;
    wire signal_2332 ;
    wire signal_2333 ;
    wire signal_2334 ;
    wire signal_2335 ;
    wire signal_2336 ;
    wire signal_2337 ;
    wire signal_2338 ;
    wire signal_2339 ;
    wire signal_2340 ;
    wire signal_2341 ;
    wire signal_2342 ;
    wire signal_2343 ;
    wire signal_2344 ;
    wire signal_2345 ;
    wire signal_2346 ;
    wire signal_2347 ;
    wire signal_2348 ;
    wire signal_2349 ;
    wire signal_2350 ;
    wire signal_2351 ;
    wire signal_2352 ;
    wire signal_2353 ;
    wire signal_2354 ;
    wire signal_2355 ;
    wire signal_2356 ;
    wire signal_2357 ;
    wire signal_2358 ;
    wire signal_2359 ;
    wire signal_2360 ;
    wire signal_2361 ;
    wire signal_2362 ;
    wire signal_2363 ;
    wire signal_2364 ;
    wire signal_2365 ;
    wire signal_2366 ;
    wire signal_2367 ;
    wire signal_2368 ;
    wire signal_2369 ;
    wire signal_2370 ;
    wire signal_2371 ;
    wire signal_2372 ;
    wire signal_2373 ;
    wire signal_2374 ;
    wire signal_2375 ;
    wire signal_2376 ;
    wire signal_2377 ;
    wire signal_2378 ;
    wire signal_2379 ;
    wire signal_2380 ;
    wire signal_2381 ;
    wire signal_2382 ;
    wire signal_2383 ;
    wire signal_2384 ;
    wire signal_2385 ;
    wire signal_2386 ;
    wire signal_2387 ;
    wire signal_2388 ;
    wire signal_2389 ;
    wire signal_2390 ;
    wire signal_2391 ;
    wire signal_2392 ;
    wire signal_2393 ;
    wire signal_2394 ;
    wire signal_2395 ;
    wire signal_2396 ;
    wire signal_2397 ;
    wire signal_2398 ;
    wire signal_2399 ;
    wire signal_2400 ;
    wire signal_2401 ;
    wire signal_2402 ;
    wire signal_2403 ;
    wire signal_2404 ;
    wire signal_2405 ;
    wire signal_2406 ;
    wire signal_2407 ;
    wire signal_2408 ;
    wire signal_2409 ;
    wire signal_2410 ;
    wire signal_2411 ;
    wire signal_2412 ;
    wire signal_2413 ;
    wire signal_2414 ;
    wire signal_2415 ;
    wire signal_2416 ;
    wire signal_2417 ;
    wire signal_2418 ;
    wire signal_2419 ;
    wire signal_2420 ;
    wire signal_2421 ;
    wire signal_2422 ;
    wire signal_2423 ;
    wire signal_2424 ;
    wire signal_2425 ;
    wire signal_2426 ;
    wire signal_2427 ;
    wire signal_2428 ;
    wire signal_2429 ;
    wire signal_2430 ;
    wire signal_2431 ;
    wire signal_2432 ;
    wire signal_2433 ;
    wire signal_2434 ;
    wire signal_2435 ;
    wire signal_2436 ;
    wire signal_2437 ;
    wire signal_2438 ;
    wire signal_2439 ;
    wire signal_2440 ;
    wire signal_2441 ;
    wire signal_2442 ;
    wire signal_2443 ;
    wire signal_2444 ;
    wire signal_2445 ;
    wire signal_2446 ;
    wire signal_2447 ;
    wire signal_2448 ;
    wire signal_2449 ;
    wire signal_2450 ;
    wire signal_2451 ;
    wire signal_2452 ;
    wire signal_2453 ;
    wire signal_2454 ;
    wire signal_2455 ;
    wire signal_2456 ;
    wire signal_2457 ;
    wire signal_2458 ;
    wire signal_2459 ;
    wire signal_2460 ;
    wire signal_2461 ;
    wire signal_2462 ;
    wire signal_2463 ;
    wire signal_2464 ;
    wire signal_2465 ;
    wire signal_2466 ;
    wire signal_2467 ;
    wire signal_2468 ;
    wire signal_2469 ;
    wire signal_2470 ;
    wire signal_2471 ;
    wire signal_2472 ;
    wire signal_2473 ;
    wire signal_2474 ;
    wire signal_2475 ;
    wire signal_2476 ;
    wire signal_2477 ;
    wire signal_2478 ;
    wire signal_2479 ;
    wire signal_2480 ;
    wire signal_2481 ;
    wire signal_2482 ;
    wire signal_2483 ;
    wire signal_2484 ;
    wire signal_2485 ;
    wire signal_2486 ;
    wire signal_2487 ;
    wire signal_2488 ;
    wire signal_2489 ;
    wire signal_2490 ;
    wire signal_2491 ;
    wire signal_2492 ;
    wire signal_2493 ;
    wire signal_2494 ;
    wire signal_2495 ;
    wire signal_2496 ;
    wire signal_2497 ;
    wire signal_2498 ;
    wire signal_2499 ;
    wire signal_2500 ;
    wire signal_2501 ;
    wire signal_2502 ;
    wire signal_2503 ;
    wire signal_2504 ;
    wire signal_2505 ;
    wire signal_2506 ;
    wire signal_2507 ;
    wire signal_2508 ;
    wire signal_2509 ;
    wire signal_2510 ;
    wire signal_2511 ;
    wire signal_2512 ;
    wire signal_2513 ;
    wire signal_2514 ;
    wire signal_2515 ;
    wire signal_2516 ;
    wire signal_2517 ;
    wire signal_2518 ;
    wire signal_2519 ;
    wire signal_2520 ;
    wire signal_2521 ;
    wire signal_2522 ;
    wire signal_2523 ;
    wire signal_2524 ;
    wire signal_2525 ;
    wire signal_2526 ;
    wire signal_2527 ;
    wire signal_2528 ;
    wire signal_2529 ;
    wire signal_2530 ;
    wire signal_2531 ;
    wire signal_2532 ;
    wire signal_2533 ;
    wire signal_2534 ;
    wire signal_2535 ;
    wire signal_2536 ;
    wire signal_2537 ;
    wire signal_2538 ;
    wire signal_2539 ;
    wire signal_2540 ;
    wire signal_2541 ;
    wire signal_2542 ;
    wire signal_2543 ;
    wire signal_2544 ;
    wire signal_2545 ;
    wire signal_2546 ;
    wire signal_2547 ;
    wire signal_2548 ;
    wire signal_2549 ;
    wire signal_2550 ;
    wire signal_2551 ;
    wire signal_2552 ;
    wire signal_2553 ;
    wire signal_2554 ;
    wire signal_2555 ;
    wire signal_2556 ;
    wire signal_2557 ;
    wire signal_2558 ;
    wire signal_2559 ;
    wire signal_2560 ;
    wire signal_2561 ;
    wire signal_2562 ;
    wire signal_2563 ;
    wire signal_2564 ;
    wire signal_2565 ;
    wire signal_2566 ;
    wire signal_2567 ;
    wire signal_2568 ;
    wire signal_2569 ;
    wire signal_2570 ;
    wire signal_2571 ;
    wire signal_2572 ;
    wire signal_2573 ;
    wire signal_2574 ;
    wire signal_2575 ;
    wire signal_2576 ;
    wire signal_2577 ;
    wire signal_2578 ;
    wire signal_2579 ;
    wire signal_2580 ;
    wire signal_2581 ;
    wire signal_2582 ;
    wire signal_2583 ;
    wire signal_2584 ;
    wire signal_2585 ;
    wire signal_2586 ;
    wire signal_2587 ;
    wire signal_2588 ;
    wire signal_2589 ;
    wire signal_2590 ;
    wire signal_2591 ;
    wire signal_2592 ;
    wire signal_2593 ;
    wire signal_2594 ;
    wire signal_2595 ;
    wire signal_2596 ;
    wire signal_2597 ;
    wire signal_2598 ;
    wire signal_2599 ;
    wire signal_2600 ;
    wire signal_2601 ;
    wire signal_2602 ;
    wire signal_2603 ;
    wire signal_2604 ;
    wire signal_2605 ;
    wire signal_2606 ;
    wire signal_2607 ;
    wire signal_2608 ;
    wire signal_2609 ;
    wire signal_2610 ;
    wire signal_2611 ;
    wire signal_2612 ;
    wire signal_2613 ;
    wire signal_2614 ;
    wire signal_2615 ;
    wire signal_2616 ;
    wire signal_2617 ;
    wire signal_2618 ;
    wire signal_2619 ;
    wire signal_2620 ;
    wire signal_2621 ;
    wire signal_2622 ;
    wire signal_2623 ;
    wire signal_2624 ;
    wire signal_2625 ;
    wire signal_2626 ;
    wire signal_2627 ;
    wire signal_2628 ;
    wire signal_2629 ;
    wire signal_2630 ;
    wire signal_2631 ;
    wire signal_2632 ;
    wire signal_2633 ;
    wire signal_2634 ;
    wire signal_2635 ;
    wire signal_2636 ;
    wire signal_2637 ;
    wire signal_2638 ;
    wire signal_2639 ;
    wire signal_2640 ;
    wire signal_2641 ;
    wire signal_2642 ;
    wire signal_2643 ;
    wire signal_2644 ;
    wire signal_2645 ;
    wire signal_2646 ;
    wire signal_2647 ;
    wire signal_2648 ;
    wire signal_2649 ;
    wire signal_2650 ;
    wire signal_2651 ;
    wire signal_2652 ;
    wire signal_2653 ;
    wire signal_2654 ;
    wire signal_2655 ;
    wire signal_2656 ;
    wire signal_2657 ;
    wire signal_2658 ;
    wire signal_2659 ;
    wire signal_2660 ;
    wire signal_2661 ;
    wire signal_2662 ;
    wire signal_2663 ;
    wire signal_2664 ;
    wire signal_2665 ;
    wire signal_2666 ;
    wire signal_2667 ;
    wire signal_2668 ;
    wire signal_2669 ;
    wire signal_2670 ;
    wire signal_2671 ;
    wire signal_2672 ;
    wire signal_2673 ;
    wire signal_2674 ;
    wire signal_2675 ;
    wire signal_2676 ;
    wire signal_2677 ;
    wire signal_2678 ;
    wire signal_2679 ;
    wire signal_2680 ;
    wire signal_2681 ;
    wire signal_2682 ;
    wire signal_2683 ;
    wire signal_2684 ;
    wire signal_2685 ;
    wire signal_2686 ;
    wire signal_2687 ;
    wire signal_2688 ;
    wire signal_2689 ;
    wire signal_2690 ;
    wire signal_2691 ;
    wire signal_2692 ;
    wire signal_2693 ;
    wire signal_2694 ;
    wire signal_2695 ;
    wire signal_2696 ;
    wire signal_2697 ;
    wire signal_2698 ;
    wire signal_2699 ;
    wire signal_2700 ;
    wire signal_2701 ;
    wire signal_2702 ;
    wire signal_2703 ;
    wire signal_2704 ;
    wire signal_2705 ;
    wire signal_2706 ;
    wire signal_2707 ;
    wire signal_2708 ;
    wire signal_2709 ;
    wire signal_2710 ;
    wire signal_2711 ;
    wire signal_2712 ;
    wire signal_2713 ;
    wire signal_2714 ;
    wire signal_2715 ;
    wire signal_2716 ;
    wire signal_2717 ;
    wire signal_2718 ;
    wire signal_2719 ;
    wire signal_2720 ;
    wire signal_2721 ;
    wire signal_2722 ;
    wire signal_2723 ;
    wire signal_2724 ;
    wire signal_2725 ;
    wire signal_2726 ;
    wire signal_2727 ;
    wire signal_2728 ;
    wire signal_2729 ;
    wire signal_2730 ;
    wire signal_2731 ;
    wire signal_2732 ;
    wire signal_2733 ;
    wire signal_2734 ;
    wire signal_2735 ;
    wire signal_2736 ;
    wire signal_2737 ;
    wire signal_2738 ;
    wire signal_2739 ;
    wire signal_2740 ;
    wire signal_2741 ;
    wire signal_2742 ;
    wire signal_2743 ;
    wire signal_2744 ;
    wire signal_2745 ;
    wire signal_2746 ;
    wire signal_2747 ;
    wire signal_2748 ;
    wire signal_2749 ;
    wire signal_2750 ;
    wire signal_2751 ;
    wire signal_2752 ;
    wire signal_2753 ;
    wire signal_2754 ;
    wire signal_2755 ;
    wire signal_2756 ;
    wire signal_2757 ;
    wire signal_2758 ;
    wire signal_2759 ;
    wire signal_2760 ;
    wire signal_2761 ;
    wire signal_2762 ;
    wire signal_2763 ;
    wire signal_2764 ;
    wire signal_2765 ;
    wire signal_2766 ;
    wire signal_2767 ;
    wire signal_2768 ;
    wire signal_2769 ;
    wire signal_2770 ;
    wire signal_2771 ;
    wire signal_2772 ;
    wire signal_2773 ;
    wire signal_2774 ;
    wire signal_2775 ;
    wire signal_2776 ;
    wire signal_2777 ;
    wire signal_2778 ;
    wire signal_2779 ;
    wire signal_2780 ;
    wire signal_2781 ;
    wire signal_2782 ;
    wire signal_2783 ;
    wire signal_2784 ;
    wire signal_2785 ;
    wire signal_2786 ;
    wire signal_2787 ;
    wire signal_2788 ;
    wire signal_2789 ;
    wire signal_2790 ;
    wire signal_2791 ;
    wire signal_2792 ;
    wire signal_2793 ;
    wire signal_2794 ;
    wire signal_2795 ;
    wire signal_2796 ;
    wire signal_2797 ;
    wire signal_2798 ;
    wire signal_2799 ;
    wire signal_2800 ;
    wire signal_2801 ;
    wire signal_2802 ;
    wire signal_2803 ;
    wire signal_2804 ;
    wire signal_2805 ;
    wire signal_2806 ;
    wire signal_2807 ;
    wire signal_2808 ;
    wire signal_2809 ;
    wire signal_2810 ;
    wire signal_2811 ;
    wire signal_2812 ;
    wire signal_2813 ;
    wire signal_2814 ;
    wire signal_2815 ;
    wire signal_2816 ;
    wire signal_2817 ;
    wire signal_2818 ;
    wire signal_2819 ;
    wire signal_2820 ;
    wire signal_2821 ;
    wire signal_2822 ;
    wire signal_2823 ;
    wire signal_2824 ;
    wire signal_2825 ;
    wire signal_2826 ;
    wire signal_2827 ;
    wire signal_2828 ;
    wire signal_2829 ;
    wire signal_2830 ;
    wire signal_2831 ;
    wire signal_2832 ;
    wire signal_2833 ;
    wire signal_2834 ;
    wire signal_2835 ;
    wire signal_2836 ;
    wire signal_2837 ;
    wire signal_2838 ;
    wire signal_2839 ;
    wire signal_2840 ;
    wire signal_2841 ;
    wire signal_2842 ;
    wire signal_2843 ;
    wire signal_2844 ;
    wire signal_2845 ;
    wire signal_2846 ;
    wire signal_2847 ;
    wire signal_2848 ;
    wire signal_2849 ;
    wire signal_2850 ;
    wire signal_2851 ;
    wire signal_2852 ;
    wire signal_2853 ;
    wire signal_2854 ;
    wire signal_2855 ;
    wire signal_2856 ;
    wire signal_2857 ;
    wire signal_2858 ;
    wire signal_2859 ;
    wire signal_2860 ;
    wire signal_2861 ;
    wire signal_2862 ;
    wire signal_2863 ;
    wire signal_2864 ;
    wire signal_2865 ;
    wire signal_2866 ;
    wire signal_2867 ;
    wire signal_2868 ;
    wire signal_2869 ;
    wire signal_2870 ;
    wire signal_2871 ;
    wire signal_2872 ;
    wire signal_2873 ;
    wire signal_2874 ;
    wire signal_2875 ;
    wire signal_2876 ;
    wire signal_2877 ;
    wire signal_2878 ;
    wire signal_2879 ;
    wire signal_2880 ;
    wire signal_2881 ;
    wire signal_2882 ;
    wire signal_2883 ;
    wire signal_2884 ;
    wire signal_2885 ;
    wire signal_2886 ;
    wire signal_2887 ;
    wire signal_2888 ;
    wire signal_2889 ;
    wire signal_2890 ;
    wire signal_2891 ;
    wire signal_2892 ;
    wire signal_2893 ;
    wire signal_2894 ;
    wire signal_2895 ;
    wire signal_2896 ;
    wire signal_2897 ;
    wire signal_2898 ;
    wire signal_2899 ;
    wire signal_2900 ;
    wire signal_2901 ;
    wire signal_2902 ;
    wire signal_2903 ;
    wire signal_2904 ;
    wire signal_2905 ;
    wire signal_2906 ;
    wire signal_2907 ;
    wire signal_2908 ;
    wire signal_2909 ;
    wire signal_2910 ;
    wire signal_2911 ;
    wire signal_2912 ;
    wire signal_2913 ;
    wire signal_2914 ;
    wire signal_2915 ;
    wire signal_2916 ;
    wire signal_2917 ;
    wire signal_2918 ;
    wire signal_2919 ;
    wire signal_2920 ;
    wire signal_2921 ;
    wire signal_2922 ;
    wire signal_2923 ;
    wire signal_2924 ;
    wire signal_2925 ;
    wire signal_2926 ;
    wire signal_2927 ;
    wire signal_2928 ;
    wire signal_2929 ;
    wire signal_2930 ;
    wire signal_2931 ;
    wire signal_2932 ;
    wire signal_2933 ;
    wire signal_2934 ;
    wire signal_2935 ;
    wire signal_2936 ;
    wire signal_2937 ;
    wire signal_2938 ;
    wire signal_2939 ;
    wire signal_2940 ;
    wire signal_2941 ;
    wire signal_2942 ;
    wire signal_2943 ;
    wire signal_2944 ;
    wire signal_2945 ;
    wire signal_2946 ;
    wire signal_2947 ;
    wire signal_2948 ;
    wire signal_2949 ;
    wire signal_2950 ;
    wire signal_2951 ;
    wire signal_2952 ;
    wire signal_2953 ;
    wire signal_2955 ;
    wire signal_2957 ;
    wire signal_2958 ;
    wire signal_2959 ;
    wire signal_2960 ;
    wire signal_2961 ;
    wire signal_2962 ;
    wire signal_2963 ;
    wire signal_2964 ;
    wire signal_2965 ;
    wire signal_2966 ;
    wire signal_2967 ;
    wire signal_2968 ;
    wire signal_2969 ;
    wire signal_2970 ;
    wire signal_2971 ;
    wire signal_2972 ;
    wire signal_2973 ;
    wire signal_2974 ;
    wire signal_2975 ;
    wire signal_2976 ;
    wire signal_2977 ;
    wire signal_2978 ;
    wire signal_2979 ;
    wire signal_2980 ;
    wire signal_2981 ;
    wire signal_2982 ;
    wire signal_2983 ;
    wire signal_2984 ;
    wire signal_2985 ;
    wire signal_2986 ;
    wire signal_2987 ;
    wire signal_2988 ;
    wire signal_2989 ;
    wire signal_2990 ;
    wire signal_2992 ;
    wire signal_2994 ;
    wire signal_2996 ;
    wire signal_2998 ;
    wire signal_3000 ;
    wire signal_3001 ;
    wire signal_3002 ;
    wire signal_3003 ;
    wire signal_3004 ;
    wire signal_3005 ;
    wire signal_3006 ;
    wire signal_3007 ;
    wire signal_3008 ;
    wire signal_3009 ;
    wire signal_3010 ;
    wire signal_3011 ;
    wire signal_3012 ;
    wire signal_3013 ;
    wire signal_3014 ;
    wire signal_3015 ;
    wire signal_3016 ;
    wire signal_3017 ;
    wire signal_3018 ;
    wire signal_3019 ;
    wire signal_3020 ;
    wire signal_3021 ;
    wire signal_3022 ;
    wire signal_3023 ;
    wire signal_3024 ;
    wire signal_3026 ;
    wire signal_3028 ;
    wire signal_3030 ;
    wire signal_3032 ;
    wire signal_3034 ;
    wire signal_3036 ;
    wire signal_3038 ;
    wire signal_3040 ;
    wire signal_3041 ;
    wire signal_3042 ;
    wire signal_3043 ;
    wire signal_3044 ;
    wire signal_3045 ;
    wire signal_3046 ;
    wire signal_3047 ;
    wire signal_3048 ;
    wire signal_3049 ;
    wire signal_3050 ;
    wire signal_3051 ;
    wire signal_3052 ;
    wire signal_3053 ;
    wire signal_3054 ;
    wire signal_3055 ;
    wire signal_3056 ;
    wire signal_3057 ;
    wire signal_3058 ;
    wire signal_3059 ;
    wire signal_3060 ;
    wire signal_3061 ;
    wire signal_3062 ;
    wire signal_3063 ;
    wire signal_3065 ;
    wire signal_3067 ;
    wire signal_3069 ;
    wire signal_3071 ;
    wire signal_3073 ;
    wire signal_3075 ;
    wire signal_3077 ;
    wire signal_3078 ;
    wire signal_3079 ;
    wire signal_3080 ;
    wire signal_3081 ;
    wire signal_3082 ;
    wire signal_3083 ;
    wire signal_3084 ;
    wire signal_3085 ;
    wire signal_3086 ;
    wire signal_3087 ;
    wire signal_3088 ;
    wire signal_3089 ;
    wire signal_3090 ;
    wire signal_3091 ;
    wire signal_3092 ;
    wire signal_3093 ;
    wire signal_3094 ;
    wire signal_3095 ;
    wire signal_3096 ;
    wire signal_3097 ;
    wire signal_3098 ;
    wire signal_3099 ;
    wire signal_3100 ;
    wire signal_3101 ;
    wire signal_3102 ;
    wire signal_3103 ;
    wire signal_3104 ;
    wire signal_3105 ;
    wire signal_3106 ;
    wire signal_3107 ;
    wire signal_3108 ;
    wire signal_3109 ;
    wire signal_3110 ;
    wire signal_3112 ;
    wire signal_3114 ;
    wire signal_3116 ;
    wire signal_3118 ;
    wire signal_3120 ;
    wire signal_3121 ;
    wire signal_3122 ;
    wire signal_3123 ;
    wire signal_3124 ;
    wire signal_3125 ;
    wire signal_3126 ;
    wire signal_3127 ;
    wire signal_3128 ;
    wire signal_3129 ;
    wire signal_3130 ;
    wire signal_3131 ;
    wire signal_3132 ;
    wire signal_3133 ;
    wire signal_3134 ;
    wire signal_3135 ;
    wire signal_3136 ;
    wire signal_3137 ;
    wire signal_3138 ;
    wire signal_3139 ;
    wire signal_3140 ;
    wire signal_3141 ;
    wire signal_3143 ;
    wire signal_3145 ;
    wire signal_3147 ;
    wire signal_3149 ;
    wire signal_3151 ;
    wire signal_3153 ;
    wire signal_3155 ;
    wire signal_3157 ;
    wire signal_3159 ;
    wire signal_3161 ;
    wire signal_3163 ;
    wire signal_3164 ;
    wire signal_3165 ;
    wire signal_3166 ;
    wire signal_3167 ;
    wire signal_3168 ;
    wire signal_3169 ;
    wire signal_3170 ;
    wire signal_3171 ;
    wire signal_3172 ;
    wire signal_3173 ;
    wire signal_3174 ;
    wire signal_3175 ;
    wire signal_3176 ;
    wire signal_3177 ;
    wire signal_3178 ;
    wire signal_3179 ;
    wire signal_3180 ;
    wire signal_3181 ;
    wire signal_3182 ;
    wire signal_3183 ;
    wire signal_3184 ;
    wire signal_3185 ;
    wire signal_3186 ;
    wire signal_3187 ;
    wire signal_3189 ;
    wire signal_3191 ;
    wire signal_3193 ;
    wire signal_3195 ;
    wire signal_3197 ;
    wire signal_3198 ;
    wire signal_3199 ;
    wire signal_3200 ;
    wire signal_3201 ;
    wire signal_3202 ;
    wire signal_3203 ;
    wire signal_3204 ;
    wire signal_3205 ;
    wire signal_3206 ;
    wire signal_3207 ;
    wire signal_3208 ;
    wire signal_3209 ;
    wire signal_3210 ;
    wire signal_3211 ;
    wire signal_3212 ;
    wire signal_3213 ;
    wire signal_3215 ;
    wire signal_3217 ;
    wire signal_3219 ;
    wire signal_3221 ;
    wire signal_3223 ;
    wire signal_3225 ;
    wire signal_3227 ;
    wire signal_3229 ;
    wire signal_3231 ;
    wire signal_3233 ;
    wire signal_3234 ;
    wire signal_3235 ;
    wire signal_3236 ;
    wire signal_3237 ;
    wire signal_3238 ;
    wire signal_3239 ;
    wire signal_3240 ;
    wire signal_3241 ;
    wire signal_3243 ;
    wire signal_3245 ;
    wire signal_3247 ;
    wire signal_3249 ;
    wire signal_3251 ;
    wire signal_3252 ;
    wire signal_3253 ;
    wire signal_3254 ;
    wire signal_3255 ;
    wire signal_3256 ;
    wire signal_3257 ;
    wire signal_3258 ;
    wire signal_3259 ;
    wire signal_3261 ;
    wire signal_3263 ;
    wire signal_3265 ;
    wire signal_3267 ;
    wire signal_3269 ;
    wire signal_3271 ;
    wire signal_3870 ;

    /* cells in depth 0 */
    NOR2_X1 cell_0 ( .A1 (signal_875), .A2 (signal_878), .ZN (signal_266) ) ;
    NAND2_X1 cell_1 ( .A1 (signal_879), .A2 (signal_266), .ZN (signal_267) ) ;
    NOR2_X1 cell_2 ( .A1 (signal_874), .A2 (signal_267), .ZN (signal_268) ) ;
    NAND2_X1 cell_3 ( .A1 (signal_876), .A2 (signal_268), .ZN (signal_269) ) ;
    NOR2_X1 cell_4 ( .A1 (signal_877), .A2 (signal_269), .ZN (signal_270) ) ;
    NOR2_X1 cell_5 ( .A1 (OUT_done), .A2 (signal_270), .ZN (signal_271) ) ;
    NOR2_X1 cell_6 ( .A1 (IN_reset), .A2 (signal_271), .ZN (signal_265) ) ;
    NAND2_X1 cell_7 ( .A1 (signal_273), .A2 (signal_274), .ZN (signal_272) ) ;
    XNOR2_X1 cell_8 ( .A (signal_304), .B (signal_275), .ZN (signal_274) ) ;
    XOR2_X1 cell_9 ( .A (signal_309), .B (signal_307), .Z (signal_275) ) ;
    NAND2_X1 cell_10 ( .A1 (signal_276), .A2 (signal_277), .ZN (signal_273) ) ;
    NAND2_X1 cell_11 ( .A1 (signal_278), .A2 (signal_279), .ZN (signal_277) ) ;
    NOR2_X1 cell_12 ( .A1 (signal_302), .A2 (signal_289), .ZN (signal_279) ) ;
    NOR2_X1 cell_13 ( .A1 (signal_306), .A2 (signal_309), .ZN (signal_278) ) ;
    NAND2_X1 cell_14 ( .A1 (signal_289), .A2 (signal_280), .ZN (signal_276) ) ;
    AND2_X1 cell_15 ( .A1 (signal_306), .A2 (signal_309), .ZN (signal_280) ) ;
    NAND2_X1 cell_16 ( .A1 (signal_298), .A2 (signal_283), .ZN (signal_282) ) ;
    NOR2_X1 cell_17 ( .A1 (signal_300), .A2 (signal_284), .ZN (signal_283) ) ;
    NAND2_X1 cell_18 ( .A1 (signal_296), .A2 (signal_876), .ZN (signal_284) ) ;
    NAND2_X1 cell_19 ( .A1 (signal_292), .A2 (signal_290), .ZN (signal_281) ) ;
    NOR2_X1 cell_20 ( .A1 (signal_292), .A2 (IN_reset), .ZN (signal_291) ) ;
    NOR2_X1 cell_21 ( .A1 (IN_reset), .A2 (signal_294), .ZN (signal_293) ) ;
    NOR2_X1 cell_22 ( .A1 (IN_reset), .A2 (signal_296), .ZN (signal_295) ) ;
    NOR2_X1 cell_23 ( .A1 (IN_reset), .A2 (signal_298), .ZN (signal_297) ) ;
    NOR2_X1 cell_24 ( .A1 (IN_reset), .A2 (signal_300), .ZN (signal_299) ) ;
    NOR2_X1 cell_25 ( .A1 (signal_289), .A2 (IN_reset), .ZN (signal_303) ) ;
    NOR2_X1 cell_26 ( .A1 (signal_306), .A2 (IN_reset), .ZN (signal_305) ) ;
    NOR2_X1 cell_27 ( .A1 (signal_309), .A2 (IN_reset), .ZN (signal_308) ) ;
    NOR2_X1 cell_28 ( .A1 (signal_288), .A2 (IN_reset), .ZN (signal_310) ) ;
    OR2_X1 cell_29 ( .A1 (signal_288), .A2 (signal_276), .ZN (signal_286) ) ;
    NAND2_X1 cell_30 ( .A1 (signal_272), .A2 (signal_286), .ZN (signal_311) ) ;
    NOR2_X1 cell_31 ( .A1 (signal_281), .A2 (signal_282), .ZN (signal_340) ) ;
    INV_X1 cell_32 ( .A (signal_286), .ZN (signal_285) ) ;
    OR2_X1 cell_33 ( .A1 (IN_reset), .A2 (signal_287), .ZN (signal_301) ) ;
    XNOR2_X1 cell_34 ( .A (signal_292), .B (signal_290), .ZN (signal_287) ) ;
    INV_X1 cell_35 ( .A (signal_340), .ZN (signal_341) ) ;
    INV_X1 cell_36 ( .A (signal_341), .ZN (signal_344) ) ;
    INV_X1 cell_37 ( .A (signal_341), .ZN (signal_342) ) ;
    INV_X1 cell_38 ( .A (signal_341), .ZN (signal_343) ) ;
    INV_X1 cell_167 ( .A (signal_345), .ZN (signal_346) ) ;
    INV_X1 cell_168 ( .A (signal_285), .ZN (signal_345) ) ;
    INV_X1 cell_169 ( .A (signal_345), .ZN (signal_348) ) ;
    INV_X1 cell_170 ( .A (signal_345), .ZN (signal_347) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_171 ( .s (signal_285), .b ({IN_key_s1[64], IN_key_s0[64]}), .a ({IN_key_s1[0], IN_key_s0[0]}), .c ({signal_1856, signal_1135}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_172 ( .s (signal_346), .b ({IN_key_s1[65], IN_key_s0[65]}), .a ({IN_key_s1[1], IN_key_s0[1]}), .c ({signal_1921, signal_1134}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_173 ( .s (signal_346), .b ({IN_key_s1[66], IN_key_s0[66]}), .a ({IN_key_s1[2], IN_key_s0[2]}), .c ({signal_1924, signal_1133}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_174 ( .s (signal_285), .b ({IN_key_s1[67], IN_key_s0[67]}), .a ({IN_key_s1[3], IN_key_s0[3]}), .c ({signal_1859, signal_1132}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_175 ( .s (signal_346), .b ({IN_key_s1[68], IN_key_s0[68]}), .a ({IN_key_s1[4], IN_key_s0[4]}), .c ({signal_1927, signal_1131}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_176 ( .s (signal_346), .b ({IN_key_s1[69], IN_key_s0[69]}), .a ({IN_key_s1[5], IN_key_s0[5]}), .c ({signal_1930, signal_1130}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_177 ( .s (signal_346), .b ({IN_key_s1[70], IN_key_s0[70]}), .a ({IN_key_s1[6], IN_key_s0[6]}), .c ({signal_1933, signal_1129}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_178 ( .s (signal_346), .b ({IN_key_s1[71], IN_key_s0[71]}), .a ({IN_key_s1[7], IN_key_s0[7]}), .c ({signal_1936, signal_1128}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_179 ( .s (signal_346), .b ({IN_key_s1[72], IN_key_s0[72]}), .a ({IN_key_s1[8], IN_key_s0[8]}), .c ({signal_1939, signal_1127}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_180 ( .s (signal_346), .b ({IN_key_s1[73], IN_key_s0[73]}), .a ({IN_key_s1[9], IN_key_s0[9]}), .c ({signal_1942, signal_1126}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_181 ( .s (signal_346), .b ({IN_key_s1[74], IN_key_s0[74]}), .a ({IN_key_s1[10], IN_key_s0[10]}), .c ({signal_1945, signal_1125}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_182 ( .s (signal_346), .b ({IN_key_s1[75], IN_key_s0[75]}), .a ({IN_key_s1[11], IN_key_s0[11]}), .c ({signal_1948, signal_1124}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_183 ( .s (signal_346), .b ({IN_key_s1[76], IN_key_s0[76]}), .a ({IN_key_s1[12], IN_key_s0[12]}), .c ({signal_1951, signal_1123}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_184 ( .s (signal_346), .b ({IN_key_s1[77], IN_key_s0[77]}), .a ({IN_key_s1[13], IN_key_s0[13]}), .c ({signal_1954, signal_1122}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_185 ( .s (signal_346), .b ({IN_key_s1[78], IN_key_s0[78]}), .a ({IN_key_s1[14], IN_key_s0[14]}), .c ({signal_1957, signal_1121}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_186 ( .s (signal_346), .b ({IN_key_s1[79], IN_key_s0[79]}), .a ({IN_key_s1[15], IN_key_s0[15]}), .c ({signal_1960, signal_1120}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_187 ( .s (signal_285), .b ({IN_key_s1[80], IN_key_s0[80]}), .a ({IN_key_s1[16], IN_key_s0[16]}), .c ({signal_1862, signal_1119}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_188 ( .s (signal_347), .b ({IN_key_s1[81], IN_key_s0[81]}), .a ({IN_key_s1[17], IN_key_s0[17]}), .c ({signal_1963, signal_1118}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_189 ( .s (signal_348), .b ({IN_key_s1[82], IN_key_s0[82]}), .a ({IN_key_s1[18], IN_key_s0[18]}), .c ({signal_1966, signal_1117}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_190 ( .s (signal_285), .b ({IN_key_s1[83], IN_key_s0[83]}), .a ({IN_key_s1[19], IN_key_s0[19]}), .c ({signal_1865, signal_1116}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_191 ( .s (signal_346), .b ({IN_key_s1[84], IN_key_s0[84]}), .a ({IN_key_s1[20], IN_key_s0[20]}), .c ({signal_1969, signal_1115}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_192 ( .s (signal_348), .b ({IN_key_s1[85], IN_key_s0[85]}), .a ({IN_key_s1[21], IN_key_s0[21]}), .c ({signal_1972, signal_1114}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_193 ( .s (signal_285), .b ({IN_key_s1[86], IN_key_s0[86]}), .a ({IN_key_s1[22], IN_key_s0[22]}), .c ({signal_1868, signal_1113}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_194 ( .s (signal_348), .b ({IN_key_s1[87], IN_key_s0[87]}), .a ({IN_key_s1[23], IN_key_s0[23]}), .c ({signal_1975, signal_1112}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_195 ( .s (signal_285), .b ({IN_key_s1[88], IN_key_s0[88]}), .a ({IN_key_s1[24], IN_key_s0[24]}), .c ({signal_1871, signal_1111}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_196 ( .s (signal_348), .b ({IN_key_s1[89], IN_key_s0[89]}), .a ({IN_key_s1[25], IN_key_s0[25]}), .c ({signal_1978, signal_1110}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_197 ( .s (signal_285), .b ({IN_key_s1[90], IN_key_s0[90]}), .a ({IN_key_s1[26], IN_key_s0[26]}), .c ({signal_1874, signal_1109}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_198 ( .s (signal_348), .b ({IN_key_s1[91], IN_key_s0[91]}), .a ({IN_key_s1[27], IN_key_s0[27]}), .c ({signal_1981, signal_1108}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_199 ( .s (signal_285), .b ({IN_key_s1[92], IN_key_s0[92]}), .a ({IN_key_s1[28], IN_key_s0[28]}), .c ({signal_1877, signal_1107}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_200 ( .s (signal_347), .b ({IN_key_s1[93], IN_key_s0[93]}), .a ({IN_key_s1[29], IN_key_s0[29]}), .c ({signal_1984, signal_1106}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_201 ( .s (signal_347), .b ({IN_key_s1[94], IN_key_s0[94]}), .a ({IN_key_s1[30], IN_key_s0[30]}), .c ({signal_1987, signal_1105}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_202 ( .s (signal_347), .b ({IN_key_s1[95], IN_key_s0[95]}), .a ({IN_key_s1[31], IN_key_s0[31]}), .c ({signal_1990, signal_1104}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_203 ( .s (signal_285), .b ({IN_key_s1[96], IN_key_s0[96]}), .a ({IN_key_s1[32], IN_key_s0[32]}), .c ({signal_1880, signal_1103}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_204 ( .s (signal_348), .b ({IN_key_s1[97], IN_key_s0[97]}), .a ({IN_key_s1[33], IN_key_s0[33]}), .c ({signal_1993, signal_1102}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_205 ( .s (signal_285), .b ({IN_key_s1[98], IN_key_s0[98]}), .a ({IN_key_s1[34], IN_key_s0[34]}), .c ({signal_1883, signal_1101}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_206 ( .s (signal_285), .b ({IN_key_s1[99], IN_key_s0[99]}), .a ({IN_key_s1[35], IN_key_s0[35]}), .c ({signal_1886, signal_1100}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_207 ( .s (signal_285), .b ({IN_key_s1[100], IN_key_s0[100]}), .a ({IN_key_s1[36], IN_key_s0[36]}), .c ({signal_1889, signal_1099}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_208 ( .s (signal_347), .b ({IN_key_s1[101], IN_key_s0[101]}), .a ({IN_key_s1[37], IN_key_s0[37]}), .c ({signal_1996, signal_1098}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_209 ( .s (signal_347), .b ({IN_key_s1[102], IN_key_s0[102]}), .a ({IN_key_s1[38], IN_key_s0[38]}), .c ({signal_1999, signal_1097}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_210 ( .s (signal_285), .b ({IN_key_s1[103], IN_key_s0[103]}), .a ({IN_key_s1[39], IN_key_s0[39]}), .c ({signal_1892, signal_1096}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_211 ( .s (signal_347), .b ({IN_key_s1[104], IN_key_s0[104]}), .a ({IN_key_s1[40], IN_key_s0[40]}), .c ({signal_2002, signal_1095}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_212 ( .s (signal_347), .b ({IN_key_s1[105], IN_key_s0[105]}), .a ({IN_key_s1[41], IN_key_s0[41]}), .c ({signal_2005, signal_1094}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_213 ( .s (signal_347), .b ({IN_key_s1[106], IN_key_s0[106]}), .a ({IN_key_s1[42], IN_key_s0[42]}), .c ({signal_2008, signal_1093}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_214 ( .s (signal_347), .b ({IN_key_s1[107], IN_key_s0[107]}), .a ({IN_key_s1[43], IN_key_s0[43]}), .c ({signal_2011, signal_1092}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_215 ( .s (signal_347), .b ({IN_key_s1[108], IN_key_s0[108]}), .a ({IN_key_s1[44], IN_key_s0[44]}), .c ({signal_2014, signal_1091}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_216 ( .s (signal_347), .b ({IN_key_s1[109], IN_key_s0[109]}), .a ({IN_key_s1[45], IN_key_s0[45]}), .c ({signal_2017, signal_1090}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_217 ( .s (signal_347), .b ({IN_key_s1[110], IN_key_s0[110]}), .a ({IN_key_s1[46], IN_key_s0[46]}), .c ({signal_2020, signal_1089}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_218 ( .s (signal_347), .b ({IN_key_s1[111], IN_key_s0[111]}), .a ({IN_key_s1[47], IN_key_s0[47]}), .c ({signal_2023, signal_1088}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_219 ( .s (signal_347), .b ({IN_key_s1[112], IN_key_s0[112]}), .a ({IN_key_s1[48], IN_key_s0[48]}), .c ({signal_2026, signal_1087}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_220 ( .s (signal_347), .b ({IN_key_s1[113], IN_key_s0[113]}), .a ({IN_key_s1[49], IN_key_s0[49]}), .c ({signal_2029, signal_1086}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_221 ( .s (signal_347), .b ({IN_key_s1[114], IN_key_s0[114]}), .a ({IN_key_s1[50], IN_key_s0[50]}), .c ({signal_2032, signal_1085}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_222 ( .s (signal_347), .b ({IN_key_s1[115], IN_key_s0[115]}), .a ({IN_key_s1[51], IN_key_s0[51]}), .c ({signal_2035, signal_1084}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_223 ( .s (signal_348), .b ({IN_key_s1[116], IN_key_s0[116]}), .a ({IN_key_s1[52], IN_key_s0[52]}), .c ({signal_2038, signal_1083}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_224 ( .s (signal_348), .b ({IN_key_s1[117], IN_key_s0[117]}), .a ({IN_key_s1[53], IN_key_s0[53]}), .c ({signal_2041, signal_1082}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_225 ( .s (signal_348), .b ({IN_key_s1[118], IN_key_s0[118]}), .a ({IN_key_s1[54], IN_key_s0[54]}), .c ({signal_2044, signal_1081}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_226 ( .s (signal_348), .b ({IN_key_s1[119], IN_key_s0[119]}), .a ({IN_key_s1[55], IN_key_s0[55]}), .c ({signal_2047, signal_1080}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_227 ( .s (signal_348), .b ({IN_key_s1[120], IN_key_s0[120]}), .a ({IN_key_s1[56], IN_key_s0[56]}), .c ({signal_2050, signal_1079}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_228 ( .s (signal_348), .b ({IN_key_s1[121], IN_key_s0[121]}), .a ({IN_key_s1[57], IN_key_s0[57]}), .c ({signal_2053, signal_1078}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_229 ( .s (signal_348), .b ({IN_key_s1[122], IN_key_s0[122]}), .a ({IN_key_s1[58], IN_key_s0[58]}), .c ({signal_2056, signal_1077}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_230 ( .s (signal_348), .b ({IN_key_s1[123], IN_key_s0[123]}), .a ({IN_key_s1[59], IN_key_s0[59]}), .c ({signal_2059, signal_1076}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_231 ( .s (signal_348), .b ({IN_key_s1[124], IN_key_s0[124]}), .a ({IN_key_s1[60], IN_key_s0[60]}), .c ({signal_2062, signal_1075}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_232 ( .s (signal_348), .b ({IN_key_s1[125], IN_key_s0[125]}), .a ({IN_key_s1[61], IN_key_s0[61]}), .c ({signal_2065, signal_1074}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_233 ( .s (signal_348), .b ({IN_key_s1[126], IN_key_s0[126]}), .a ({IN_key_s1[62], IN_key_s0[62]}), .c ({signal_2068, signal_1073}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_234 ( .s (signal_348), .b ({IN_key_s1[127], IN_key_s0[127]}), .a ({IN_key_s1[63], IN_key_s0[63]}), .c ({signal_2071, signal_1072}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_235 ( .a ({OUT_ciphertext_s1[9], OUT_ciphertext_s0[9]}), .b ({signal_1942, signal_1126}), .c ({signal_2080, signal_1062}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_236 ( .a ({OUT_ciphertext_s1[8], OUT_ciphertext_s0[8]}), .b ({signal_1939, signal_1127}), .c ({signal_2082, signal_1063}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_237 ( .a ({OUT_ciphertext_s1[7], OUT_ciphertext_s0[7]}), .b ({signal_1936, signal_1128}), .c ({signal_2084, signal_1064}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_238 ( .a ({OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}), .b ({signal_1933, signal_1129}), .c ({signal_2086, signal_1065}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_239 ( .a ({OUT_ciphertext_s1[63], OUT_ciphertext_s0[63]}), .b ({signal_2071, signal_1072}), .c ({signal_2088, signal_1008}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_240 ( .a ({OUT_ciphertext_s1[62], OUT_ciphertext_s0[62]}), .b ({signal_2068, signal_1073}), .c ({signal_2090, signal_1009}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_241 ( .a ({OUT_ciphertext_s1[61], OUT_ciphertext_s0[61]}), .b ({signal_2065, signal_1074}), .c ({signal_2092, signal_1010}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_242 ( .a ({OUT_ciphertext_s1[60], OUT_ciphertext_s0[60]}), .b ({signal_2062, signal_1075}), .c ({signal_2094, signal_1011}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_243 ( .a ({OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}), .b ({signal_1930, signal_1130}), .c ({signal_2096, signal_1066}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_244 ( .a ({OUT_ciphertext_s1[59], OUT_ciphertext_s0[59]}), .b ({signal_2059, signal_1076}), .c ({signal_2098, signal_1012}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_245 ( .a ({OUT_ciphertext_s1[58], OUT_ciphertext_s0[58]}), .b ({signal_2056, signal_1077}), .c ({signal_2100, signal_1013}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_246 ( .a ({OUT_ciphertext_s1[57], OUT_ciphertext_s0[57]}), .b ({signal_2053, signal_1078}), .c ({signal_2102, signal_1014}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_247 ( .a ({OUT_ciphertext_s1[56], OUT_ciphertext_s0[56]}), .b ({signal_2050, signal_1079}), .c ({signal_2104, signal_1015}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_248 ( .a ({OUT_ciphertext_s1[55], OUT_ciphertext_s0[55]}), .b ({signal_2047, signal_1080}), .c ({signal_2106, signal_1016}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_249 ( .a ({OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}), .b ({signal_2044, signal_1081}), .c ({signal_2108, signal_1017}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_250 ( .a ({OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}), .b ({signal_2041, signal_1082}), .c ({signal_2110, signal_1018}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_251 ( .a ({OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}), .b ({signal_2038, signal_1083}), .c ({signal_2112, signal_1019}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_252 ( .a ({OUT_ciphertext_s1[51], OUT_ciphertext_s0[51]}), .b ({signal_2035, signal_1084}), .c ({signal_2114, signal_1020}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_253 ( .a ({OUT_ciphertext_s1[50], OUT_ciphertext_s0[50]}), .b ({signal_2032, signal_1085}), .c ({signal_2116, signal_1021}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_254 ( .a ({OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}), .b ({signal_1927, signal_1131}), .c ({signal_2118, signal_1067}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_255 ( .a ({OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}), .b ({signal_2029, signal_1086}), .c ({signal_2120, signal_1022}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_256 ( .a ({OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}), .b ({signal_2026, signal_1087}), .c ({signal_2122, signal_1023}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_257 ( .a ({OUT_ciphertext_s1[47], OUT_ciphertext_s0[47]}), .b ({signal_2023, signal_1088}), .c ({signal_2124, signal_1024}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_258 ( .a ({OUT_ciphertext_s1[46], OUT_ciphertext_s0[46]}), .b ({signal_2020, signal_1089}), .c ({signal_2126, signal_1025}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_259 ( .a ({OUT_ciphertext_s1[45], OUT_ciphertext_s0[45]}), .b ({signal_2017, signal_1090}), .c ({signal_2128, signal_1026}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_260 ( .a ({OUT_ciphertext_s1[44], OUT_ciphertext_s0[44]}), .b ({signal_2014, signal_1091}), .c ({signal_2130, signal_1027}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_261 ( .a ({OUT_ciphertext_s1[43], OUT_ciphertext_s0[43]}), .b ({signal_2011, signal_1092}), .c ({signal_2132, signal_1028}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_262 ( .a ({OUT_ciphertext_s1[42], OUT_ciphertext_s0[42]}), .b ({signal_2008, signal_1093}), .c ({signal_2134, signal_1029}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_263 ( .a ({OUT_ciphertext_s1[41], OUT_ciphertext_s0[41]}), .b ({signal_2005, signal_1094}), .c ({signal_2136, signal_1030}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_264 ( .a ({OUT_ciphertext_s1[40], OUT_ciphertext_s0[40]}), .b ({signal_2002, signal_1095}), .c ({signal_2138, signal_1031}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_265 ( .a ({OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}), .b ({signal_1859, signal_1132}), .c ({signal_1894, signal_1068}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_266 ( .a ({OUT_ciphertext_s1[39], OUT_ciphertext_s0[39]}), .b ({signal_1892, signal_1096}), .c ({signal_1896, signal_1032}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_267 ( .a ({OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}), .b ({signal_1999, signal_1097}), .c ({signal_2140, signal_1033}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_268 ( .a ({OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}), .b ({signal_1996, signal_1098}), .c ({signal_2142, signal_1034}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_269 ( .a ({OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}), .b ({signal_1889, signal_1099}), .c ({signal_1898, signal_1035}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_270 ( .a ({OUT_ciphertext_s1[35], OUT_ciphertext_s0[35]}), .b ({signal_1886, signal_1100}), .c ({signal_1900, signal_1036}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_271 ( .a ({OUT_ciphertext_s1[34], OUT_ciphertext_s0[34]}), .b ({signal_1883, signal_1101}), .c ({signal_1902, signal_1037}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_272 ( .a ({OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}), .b ({signal_1993, signal_1102}), .c ({signal_2144, signal_1038}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_273 ( .a ({OUT_ciphertext_s1[32], OUT_ciphertext_s0[32]}), .b ({signal_1880, signal_1103}), .c ({signal_1904, signal_1039}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_274 ( .a ({OUT_ciphertext_s1[31], OUT_ciphertext_s0[31]}), .b ({signal_1990, signal_1104}), .c ({signal_2146, signal_1040}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_275 ( .a ({OUT_ciphertext_s1[30], OUT_ciphertext_s0[30]}), .b ({signal_1987, signal_1105}), .c ({signal_2148, signal_1041}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_276 ( .a ({OUT_ciphertext_s1[2], OUT_ciphertext_s0[2]}), .b ({signal_1924, signal_1133}), .c ({signal_2150, signal_1069}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_277 ( .a ({OUT_ciphertext_s1[29], OUT_ciphertext_s0[29]}), .b ({signal_1984, signal_1106}), .c ({signal_2152, signal_1042}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_278 ( .a ({OUT_ciphertext_s1[28], OUT_ciphertext_s0[28]}), .b ({signal_1877, signal_1107}), .c ({signal_1906, signal_1043}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_279 ( .a ({OUT_ciphertext_s1[27], OUT_ciphertext_s0[27]}), .b ({signal_1981, signal_1108}), .c ({signal_2154, signal_1044}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_280 ( .a ({OUT_ciphertext_s1[26], OUT_ciphertext_s0[26]}), .b ({signal_1874, signal_1109}), .c ({signal_1908, signal_1045}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_281 ( .a ({OUT_ciphertext_s1[25], OUT_ciphertext_s0[25]}), .b ({signal_1978, signal_1110}), .c ({signal_2156, signal_1046}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_282 ( .a ({OUT_ciphertext_s1[24], OUT_ciphertext_s0[24]}), .b ({signal_1871, signal_1111}), .c ({signal_1910, signal_1047}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_283 ( .a ({OUT_ciphertext_s1[23], OUT_ciphertext_s0[23]}), .b ({signal_1975, signal_1112}), .c ({signal_2158, signal_1048}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_284 ( .a ({OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}), .b ({signal_1868, signal_1113}), .c ({signal_1912, signal_1049}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_285 ( .a ({OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}), .b ({signal_1972, signal_1114}), .c ({signal_2160, signal_1050}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_286 ( .a ({OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}), .b ({signal_1969, signal_1115}), .c ({signal_2162, signal_1051}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_287 ( .a ({OUT_ciphertext_s1[1], OUT_ciphertext_s0[1]}), .b ({signal_1921, signal_1134}), .c ({signal_2164, signal_1070}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_288 ( .a ({OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}), .b ({signal_1865, signal_1116}), .c ({signal_1914, signal_1052}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_289 ( .a ({OUT_ciphertext_s1[18], OUT_ciphertext_s0[18]}), .b ({signal_1966, signal_1117}), .c ({signal_2166, signal_1053}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_290 ( .a ({OUT_ciphertext_s1[17], OUT_ciphertext_s0[17]}), .b ({signal_1963, signal_1118}), .c ({signal_2168, signal_1054}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_291 ( .a ({OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}), .b ({signal_1862, signal_1119}), .c ({signal_1916, signal_1055}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_292 ( .a ({OUT_ciphertext_s1[15], OUT_ciphertext_s0[15]}), .b ({signal_1960, signal_1120}), .c ({signal_2170, signal_1056}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_293 ( .a ({OUT_ciphertext_s1[14], OUT_ciphertext_s0[14]}), .b ({signal_1957, signal_1121}), .c ({signal_2172, signal_1057}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_294 ( .a ({OUT_ciphertext_s1[13], OUT_ciphertext_s0[13]}), .b ({signal_1954, signal_1122}), .c ({signal_2174, signal_1058}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_295 ( .a ({OUT_ciphertext_s1[12], OUT_ciphertext_s0[12]}), .b ({signal_1951, signal_1123}), .c ({signal_2176, signal_1059}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_296 ( .a ({OUT_ciphertext_s1[11], OUT_ciphertext_s0[11]}), .b ({signal_1948, signal_1124}), .c ({signal_2178, signal_1060}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_297 ( .a ({OUT_ciphertext_s1[10], OUT_ciphertext_s0[10]}), .b ({signal_1945, signal_1125}), .c ({signal_2180, signal_1061}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_298 ( .a ({OUT_ciphertext_s1[0], OUT_ciphertext_s0[0]}), .b ({signal_1856, signal_1135}), .c ({signal_1918, signal_1071}) ) ;
    INV_X1 cell_299 ( .A (signal_349), .ZN (signal_351) ) ;
    INV_X1 cell_300 ( .A (signal_311), .ZN (signal_349) ) ;
    INV_X1 cell_301 ( .A (signal_349), .ZN (signal_350) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_302 ( .s (signal_311), .b ({OUT_ciphertext_s1[0], OUT_ciphertext_s0[0]}), .a ({signal_1918, signal_1071}), .c ({signal_2072, signal_312}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_303 ( .s (signal_311), .b ({OUT_ciphertext_s1[1], OUT_ciphertext_s0[1]}), .a ({signal_2164, signal_1070}), .c ({signal_2192, signal_313}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_304 ( .s (signal_311), .b ({OUT_ciphertext_s1[2], OUT_ciphertext_s0[2]}), .a ({signal_2150, signal_1069}), .c ({signal_2193, signal_314}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_305 ( .s (signal_311), .b ({OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}), .a ({signal_1894, signal_1068}), .c ({signal_2073, signal_315}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_306 ( .s (signal_350), .b ({OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}), .a ({signal_2118, signal_1067}), .c ({signal_2194, signal_316}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_307 ( .s (signal_350), .b ({OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}), .a ({signal_2096, signal_1066}), .c ({signal_2195, signal_317}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_308 ( .s (signal_350), .b ({OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}), .a ({signal_2086, signal_1065}), .c ({signal_2196, signal_318}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_309 ( .s (signal_350), .b ({OUT_ciphertext_s1[7], OUT_ciphertext_s0[7]}), .a ({signal_2084, signal_1064}), .c ({signal_2197, signal_1000}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_310 ( .s (signal_350), .b ({OUT_ciphertext_s1[8], OUT_ciphertext_s0[8]}), .a ({signal_2082, signal_1063}), .c ({signal_2198, signal_999}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_311 ( .s (signal_350), .b ({OUT_ciphertext_s1[9], OUT_ciphertext_s0[9]}), .a ({signal_2080, signal_1062}), .c ({signal_2199, signal_998}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_312 ( .s (signal_350), .b ({OUT_ciphertext_s1[10], OUT_ciphertext_s0[10]}), .a ({signal_2180, signal_1061}), .c ({signal_2200, signal_997}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_313 ( .s (signal_350), .b ({OUT_ciphertext_s1[11], OUT_ciphertext_s0[11]}), .a ({signal_2178, signal_1060}), .c ({signal_2201, signal_996}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_314 ( .s (signal_350), .b ({OUT_ciphertext_s1[12], OUT_ciphertext_s0[12]}), .a ({signal_2176, signal_1059}), .c ({signal_2202, signal_995}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_315 ( .s (signal_350), .b ({OUT_ciphertext_s1[13], OUT_ciphertext_s0[13]}), .a ({signal_2174, signal_1058}), .c ({signal_2203, signal_994}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_316 ( .s (signal_350), .b ({OUT_ciphertext_s1[14], OUT_ciphertext_s0[14]}), .a ({signal_2172, signal_1057}), .c ({signal_2204, signal_993}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_317 ( .s (signal_350), .b ({OUT_ciphertext_s1[15], OUT_ciphertext_s0[15]}), .a ({signal_2170, signal_1056}), .c ({signal_2205, signal_992}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_318 ( .s (signal_311), .b ({OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}), .a ({signal_1916, signal_1055}), .c ({signal_2074, signal_319}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_319 ( .s (signal_311), .b ({OUT_ciphertext_s1[17], OUT_ciphertext_s0[17]}), .a ({signal_2168, signal_1054}), .c ({signal_2206, signal_320}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_320 ( .s (signal_311), .b ({OUT_ciphertext_s1[18], OUT_ciphertext_s0[18]}), .a ({signal_2166, signal_1053}), .c ({signal_2207, signal_321}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_321 ( .s (signal_311), .b ({OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}), .a ({signal_1914, signal_1052}), .c ({signal_2075, signal_322}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_322 ( .s (signal_350), .b ({OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}), .a ({signal_2162, signal_1051}), .c ({signal_2208, signal_323}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_323 ( .s (signal_311), .b ({OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}), .a ({signal_2160, signal_1050}), .c ({signal_2209, signal_324}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_324 ( .s (signal_311), .b ({OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}), .a ({signal_1912, signal_1049}), .c ({signal_2076, signal_325}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_325 ( .s (signal_311), .b ({OUT_ciphertext_s1[23], OUT_ciphertext_s0[23]}), .a ({signal_2158, signal_1048}), .c ({signal_2210, signal_984}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_326 ( .s (signal_311), .b ({OUT_ciphertext_s1[24], OUT_ciphertext_s0[24]}), .a ({signal_1910, signal_1047}), .c ({signal_2077, signal_983}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_327 ( .s (signal_311), .b ({OUT_ciphertext_s1[25], OUT_ciphertext_s0[25]}), .a ({signal_2156, signal_1046}), .c ({signal_2211, signal_982}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_328 ( .s (signal_311), .b ({OUT_ciphertext_s1[26], OUT_ciphertext_s0[26]}), .a ({signal_1908, signal_1045}), .c ({signal_2078, signal_981}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_329 ( .s (signal_311), .b ({OUT_ciphertext_s1[27], OUT_ciphertext_s0[27]}), .a ({signal_2154, signal_1044}), .c ({signal_2212, signal_980}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_330 ( .s (signal_351), .b ({OUT_ciphertext_s1[28], OUT_ciphertext_s0[28]}), .a ({signal_1906, signal_1043}), .c ({signal_2181, signal_979}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_331 ( .s (signal_351), .b ({OUT_ciphertext_s1[29], OUT_ciphertext_s0[29]}), .a ({signal_2152, signal_1042}), .c ({signal_2213, signal_978}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_332 ( .s (signal_351), .b ({OUT_ciphertext_s1[30], OUT_ciphertext_s0[30]}), .a ({signal_2148, signal_1041}), .c ({signal_2214, signal_977}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_333 ( .s (signal_351), .b ({OUT_ciphertext_s1[31], OUT_ciphertext_s0[31]}), .a ({signal_2146, signal_1040}), .c ({signal_2215, signal_976}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_334 ( .s (signal_351), .b ({OUT_ciphertext_s1[32], OUT_ciphertext_s0[32]}), .a ({signal_1904, signal_1039}), .c ({signal_2182, signal_326}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_335 ( .s (signal_351), .b ({OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}), .a ({signal_2144, signal_1038}), .c ({signal_2216, signal_327}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_336 ( .s (signal_351), .b ({OUT_ciphertext_s1[34], OUT_ciphertext_s0[34]}), .a ({signal_1902, signal_1037}), .c ({signal_2183, signal_328}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_337 ( .s (signal_351), .b ({OUT_ciphertext_s1[35], OUT_ciphertext_s0[35]}), .a ({signal_1900, signal_1036}), .c ({signal_2184, signal_329}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_338 ( .s (signal_351), .b ({OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}), .a ({signal_1898, signal_1035}), .c ({signal_2185, signal_330}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_339 ( .s (signal_311), .b ({OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}), .a ({signal_2142, signal_1034}), .c ({signal_2217, signal_331}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_340 ( .s (signal_351), .b ({OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}), .a ({signal_2140, signal_1033}), .c ({signal_2218, signal_332}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_341 ( .s (signal_351), .b ({OUT_ciphertext_s1[39], OUT_ciphertext_s0[39]}), .a ({signal_1896, signal_1032}), .c ({signal_2186, signal_968}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_342 ( .s (signal_351), .b ({OUT_ciphertext_s1[40], OUT_ciphertext_s0[40]}), .a ({signal_2138, signal_1031}), .c ({signal_2219, signal_967}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_343 ( .s (signal_351), .b ({OUT_ciphertext_s1[41], OUT_ciphertext_s0[41]}), .a ({signal_2136, signal_1030}), .c ({signal_2220, signal_966}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_344 ( .s (signal_351), .b ({OUT_ciphertext_s1[42], OUT_ciphertext_s0[42]}), .a ({signal_2134, signal_1029}), .c ({signal_2221, signal_965}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_345 ( .s (signal_351), .b ({OUT_ciphertext_s1[43], OUT_ciphertext_s0[43]}), .a ({signal_2132, signal_1028}), .c ({signal_2222, signal_964}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_346 ( .s (signal_351), .b ({OUT_ciphertext_s1[44], OUT_ciphertext_s0[44]}), .a ({signal_2130, signal_1027}), .c ({signal_2223, signal_963}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_347 ( .s (signal_351), .b ({OUT_ciphertext_s1[45], OUT_ciphertext_s0[45]}), .a ({signal_2128, signal_1026}), .c ({signal_2224, signal_962}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_348 ( .s (signal_351), .b ({OUT_ciphertext_s1[46], OUT_ciphertext_s0[46]}), .a ({signal_2126, signal_1025}), .c ({signal_2225, signal_961}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_349 ( .s (signal_351), .b ({OUT_ciphertext_s1[47], OUT_ciphertext_s0[47]}), .a ({signal_2124, signal_1024}), .c ({signal_2226, signal_960}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_350 ( .s (signal_351), .b ({OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}), .a ({signal_2122, signal_1023}), .c ({signal_2227, signal_333}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_351 ( .s (signal_351), .b ({OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}), .a ({signal_2120, signal_1022}), .c ({signal_2228, signal_334}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_352 ( .s (signal_311), .b ({OUT_ciphertext_s1[50], OUT_ciphertext_s0[50]}), .a ({signal_2116, signal_1021}), .c ({signal_2229, signal_335}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_353 ( .s (signal_351), .b ({OUT_ciphertext_s1[51], OUT_ciphertext_s0[51]}), .a ({signal_2114, signal_1020}), .c ({signal_2230, signal_336}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_354 ( .s (signal_351), .b ({OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}), .a ({signal_2112, signal_1019}), .c ({signal_2231, signal_337}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_355 ( .s (signal_351), .b ({OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}), .a ({signal_2110, signal_1018}), .c ({signal_2232, signal_338}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_356 ( .s (signal_351), .b ({OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}), .a ({signal_2108, signal_1017}), .c ({signal_2233, signal_339}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_357 ( .s (signal_351), .b ({OUT_ciphertext_s1[55], OUT_ciphertext_s0[55]}), .a ({signal_2106, signal_1016}), .c ({signal_2234, signal_952}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_358 ( .s (signal_351), .b ({OUT_ciphertext_s1[56], OUT_ciphertext_s0[56]}), .a ({signal_2104, signal_1015}), .c ({signal_2235, signal_951}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_359 ( .s (signal_351), .b ({OUT_ciphertext_s1[57], OUT_ciphertext_s0[57]}), .a ({signal_2102, signal_1014}), .c ({signal_2236, signal_950}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_360 ( .s (signal_351), .b ({OUT_ciphertext_s1[58], OUT_ciphertext_s0[58]}), .a ({signal_2100, signal_1013}), .c ({signal_2237, signal_949}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_361 ( .s (signal_351), .b ({OUT_ciphertext_s1[59], OUT_ciphertext_s0[59]}), .a ({signal_2098, signal_1012}), .c ({signal_2238, signal_948}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_362 ( .s (signal_351), .b ({OUT_ciphertext_s1[60], OUT_ciphertext_s0[60]}), .a ({signal_2094, signal_1011}), .c ({signal_2239, signal_947}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_363 ( .s (signal_351), .b ({OUT_ciphertext_s1[61], OUT_ciphertext_s0[61]}), .a ({signal_2092, signal_1010}), .c ({signal_2240, signal_946}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_364 ( .s (signal_351), .b ({OUT_ciphertext_s1[62], OUT_ciphertext_s0[62]}), .a ({signal_2090, signal_1009}), .c ({signal_2241, signal_945}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_365 ( .s (signal_351), .b ({OUT_ciphertext_s1[63], OUT_ciphertext_s0[63]}), .a ({signal_2088, signal_1008}), .c ({signal_2242, signal_944}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_366 ( .a ({1'b0, signal_874}), .b ({signal_2196, signal_318}), .c ({signal_2247, signal_1001}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_367 ( .a ({1'b0, signal_875}), .b ({signal_2195, signal_317}), .c ({signal_2248, signal_1002}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_368 ( .a ({1'b0, signal_877}), .b ({signal_2233, signal_339}), .c ({signal_2249, signal_953}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_369 ( .a ({1'b0, signal_878}), .b ({signal_2232, signal_338}), .c ({signal_2250, signal_954}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_370 ( .a ({1'b0, signal_879}), .b ({signal_2231, signal_337}), .c ({signal_2251, signal_955}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_371 ( .a ({1'b0, 1'b0}), .b ({signal_2230, signal_336}), .c ({signal_2252, signal_956}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_372 ( .a ({1'b0, 1'b0}), .b ({signal_2229, signal_335}), .c ({signal_2253, signal_957}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_373 ( .a ({1'b0, signal_876}), .b ({signal_2194, signal_316}), .c ({signal_2254, signal_1003}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_374 ( .a ({1'b0, 1'b0}), .b ({signal_2228, signal_334}), .c ({signal_2255, signal_958}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_375 ( .a ({1'b0, 1'b0}), .b ({signal_2227, signal_333}), .c ({signal_2256, signal_959}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_376 ( .a ({1'b0, 1'b1}), .b ({signal_2073, signal_315}), .c ({signal_2187, signal_1004}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_377 ( .a ({1'b0, signal_874}), .b ({signal_2218, signal_332}), .c ({signal_2257, signal_969}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_378 ( .a ({1'b0, signal_875}), .b ({signal_2217, signal_331}), .c ({signal_2258, signal_970}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_379 ( .a ({1'b0, signal_876}), .b ({signal_2185, signal_330}), .c ({signal_2243, signal_971}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_380 ( .a ({1'b0, 1'b0}), .b ({signal_2184, signal_329}), .c ({signal_2244, signal_972}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_381 ( .a ({1'b0, 1'b0}), .b ({signal_2183, signal_328}), .c ({signal_2245, signal_973}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_382 ( .a ({1'b0, 1'b0}), .b ({signal_2216, signal_327}), .c ({signal_2259, signal_974}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_383 ( .a ({1'b0, 1'b0}), .b ({signal_2182, signal_326}), .c ({signal_2246, signal_975}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_384 ( .a ({1'b0, 1'b0}), .b ({signal_2193, signal_314}), .c ({signal_2260, signal_1005}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_385 ( .a ({1'b0, signal_877}), .b ({signal_2076, signal_325}), .c ({signal_2188, signal_985}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_386 ( .a ({1'b0, signal_878}), .b ({signal_2209, signal_324}), .c ({signal_2261, signal_986}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_387 ( .a ({1'b0, signal_879}), .b ({signal_2208, signal_323}), .c ({signal_2262, signal_987}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_388 ( .a ({1'b0, 1'b0}), .b ({signal_2192, signal_313}), .c ({signal_2263, signal_1006}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_389 ( .a ({1'b0, 1'b1}), .b ({signal_2075, signal_322}), .c ({signal_2189, signal_988}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_390 ( .a ({1'b0, 1'b0}), .b ({signal_2207, signal_321}), .c ({signal_2264, signal_989}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_391 ( .a ({1'b0, 1'b0}), .b ({signal_2206, signal_320}), .c ({signal_2265, signal_990}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_392 ( .a ({1'b0, 1'b0}), .b ({signal_2074, signal_319}), .c ({signal_2190, signal_991}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_393 ( .a ({1'b0, 1'b0}), .b ({signal_2072, signal_312}), .c ({signal_2191, signal_1007}) ) ;
    INV_X1 cell_978 ( .A (signal_808), .ZN (signal_309) ) ;
    INV_X1 cell_980 ( .A (signal_307), .ZN (signal_306) ) ;
    INV_X1 cell_982 ( .A (signal_304), .ZN (signal_289) ) ;
    INV_X1 cell_984 ( .A (signal_288), .ZN (signal_302) ) ;
    INV_X1 cell_986 ( .A (signal_879), .ZN (signal_300) ) ;
    INV_X1 cell_988 ( .A (signal_878), .ZN (signal_298) ) ;
    INV_X1 cell_990 ( .A (signal_877), .ZN (signal_296) ) ;
    INV_X1 cell_992 ( .A (signal_876), .ZN (signal_294) ) ;
    INV_X1 cell_994 ( .A (signal_875), .ZN (signal_292) ) ;
    INV_X1 cell_996 ( .A (signal_874), .ZN (signal_290) ) ;
    ClockGatingController #(17) cell_1726 ( .clk (CLK), .rst (IN_reset), .GatedClk (signal_3870), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1128 ( .s ({signal_2201, signal_996}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[0]), .c ({signal_2266, signal_1328}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1129 ( .s ({signal_2201, signal_996}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[1]), .c ({signal_2267, signal_1329}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1130 ( .s ({signal_2205, signal_992}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[2]), .c ({signal_2268, signal_1330}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1131 ( .s ({signal_2205, signal_992}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[3]), .c ({signal_2269, signal_1331}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1132 ( .s ({signal_2212, signal_980}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[4]), .c ({signal_2270, signal_1332}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1133 ( .s ({signal_2212, signal_980}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[5]), .c ({signal_2271, signal_1333}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1134 ( .s ({signal_2215, signal_976}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[6]), .c ({signal_2272, signal_1334}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1135 ( .s ({signal_2215, signal_976}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[7]), .c ({signal_2273, signal_1335}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1136 ( .s ({signal_2222, signal_964}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[8]), .c ({signal_2274, signal_1336}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1137 ( .s ({signal_2222, signal_964}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[9]), .c ({signal_2275, signal_1337}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1138 ( .s ({signal_2226, signal_960}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[10]), .c ({signal_2276, signal_1338}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1139 ( .s ({signal_2226, signal_960}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[11]), .c ({signal_2277, signal_1339}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1140 ( .s ({signal_2238, signal_948}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[12]), .c ({signal_2278, signal_1340}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1141 ( .s ({signal_2238, signal_948}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[13]), .c ({signal_2279, signal_1341}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1142 ( .s ({signal_2242, signal_944}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[14]), .c ({signal_2280, signal_1342}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1143 ( .s ({signal_2242, signal_944}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[15]), .c ({signal_2281, signal_1343}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1144 ( .s ({signal_2260, signal_1005}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[16]), .c ({signal_2290, signal_1344}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1145 ( .s ({signal_2263, signal_1006}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[17]), .c ({signal_2291, signal_1345}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1146 ( .s ({signal_2263, signal_1006}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[18]), .c ({signal_2292, signal_1346}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1147 ( .s ({signal_2254, signal_1003}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[19]), .c ({signal_2293, signal_1347}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1148 ( .s ({signal_2254, signal_1003}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[20]), .c ({signal_2294, signal_1348}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1149 ( .s ({signal_2248, signal_1002}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[21]), .c ({signal_2295, signal_1349}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1150 ( .s ({signal_2264, signal_989}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[22]), .c ({signal_2296, signal_1350}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1151 ( .s ({signal_2265, signal_990}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[23]), .c ({signal_2297, signal_1351}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1152 ( .s ({signal_2265, signal_990}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[24]), .c ({signal_2298, signal_1352}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1153 ( .s ({signal_2262, signal_987}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[25]), .c ({signal_2299, signal_1353}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1154 ( .s ({signal_2262, signal_987}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[26]), .c ({signal_2300, signal_1354}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1155 ( .s ({signal_2261, signal_986}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[27]), .c ({signal_2301, signal_1355}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1156 ( .s ({signal_2246, signal_975}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[28]), .c ({signal_2282, signal_1356}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1157 ( .s ({signal_2259, signal_974}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[29]), .c ({signal_2302, signal_1357}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1158 ( .s ({signal_2259, signal_974}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[30]), .c ({signal_2303, signal_1358}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1159 ( .s ({signal_2257, signal_969}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[31]), .c ({signal_2304, signal_1359}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1160 ( .s ({signal_2258, signal_970}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[32]), .c ({signal_2305, signal_1360}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1161 ( .s ({signal_2258, signal_970}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[33]), .c ({signal_2306, signal_1361}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1162 ( .s ({signal_2256, signal_959}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[34]), .c ({signal_2307, signal_1362}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1163 ( .s ({signal_2256, signal_959}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[35]), .c ({signal_2308, signal_1363}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1164 ( .s ({signal_2255, signal_958}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[36]), .c ({signal_2309, signal_1364}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1165 ( .s ({signal_2251, signal_955}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[37]), .c ({signal_2310, signal_1365}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1166 ( .s ({signal_2251, signal_955}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[38]), .c ({signal_2311, signal_1366}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1167 ( .s ({signal_2250, signal_954}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[39]), .c ({signal_2312, signal_1367}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1168 ( .s ({signal_2221, signal_965}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[40]), .c ({signal_2283, signal_1368}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1169 ( .s ({signal_2241, signal_945}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[41]), .c ({signal_2284, signal_1369}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1170 ( .s ({signal_2225, signal_961}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[42]), .c ({signal_2285, signal_1370}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1171 ( .s ({signal_2257, signal_969}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[43]), .c ({signal_2313, signal_1371}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1172 ( .s ({signal_2264, signal_989}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[44]), .c ({signal_2314, signal_1372}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1173 ( .s ({signal_2261, signal_986}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[45]), .c ({signal_2315, signal_1373}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1174 ( .s ({signal_2255, signal_958}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[46]), .c ({signal_2316, signal_1374}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1175 ( .s ({signal_2248, signal_1002}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[47]), .c ({signal_2317, signal_1375}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1176 ( .s ({signal_2250, signal_954}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[48]), .c ({signal_2318, signal_1376}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1177 ( .s ({signal_2246, signal_975}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[49]), .c ({signal_2286, signal_1377}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1178 ( .s ({signal_2200, signal_997}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[50]), .c ({signal_2287, signal_1378}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1179 ( .s ({signal_2204, signal_993}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[51]), .c ({signal_2288, signal_1379}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1180 ( .s ({signal_2237, signal_949}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[52]), .c ({signal_2289, signal_1380}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1181 ( .s ({signal_2260, signal_1005}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[53]), .c ({signal_2319, signal_1381}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1182 ( .s ({signal_2200, signal_997}), .b ({1'b0, 1'b0}), .a ({signal_2266, signal_1328}), .clk (CLK), .r (Fresh[54]), .c ({signal_2320, signal_1382}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1183 ( .s ({signal_2200, signal_997}), .b ({signal_2267, signal_1329}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[55]), .c ({signal_2321, signal_1383}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1184 ( .s ({signal_2200, signal_997}), .b ({signal_2266, signal_1328}), .a ({signal_2267, signal_1329}), .clk (CLK), .r (Fresh[56]), .c ({signal_2322, signal_1384}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1185 ( .s ({signal_2204, signal_993}), .b ({1'b0, 1'b0}), .a ({signal_2268, signal_1330}), .clk (CLK), .r (Fresh[57]), .c ({signal_2323, signal_1385}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1186 ( .s ({signal_2204, signal_993}), .b ({signal_2269, signal_1331}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[58]), .c ({signal_2324, signal_1386}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1187 ( .s ({signal_2204, signal_993}), .b ({signal_2268, signal_1330}), .a ({signal_2269, signal_1331}), .clk (CLK), .r (Fresh[59]), .c ({signal_2325, signal_1387}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1188 ( .s ({signal_2211, signal_982}), .b ({1'b0, 1'b1}), .a ({signal_2270, signal_1332}), .clk (CLK), .r (Fresh[60]), .c ({signal_2326, signal_1388}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1189 ( .s ({signal_2211, signal_982}), .b ({signal_2271, signal_1333}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[61]), .c ({signal_2327, signal_1389}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1190 ( .s ({signal_2211, signal_982}), .b ({signal_2271, signal_1333}), .a ({signal_2270, signal_1332}), .clk (CLK), .r (Fresh[62]), .c ({signal_2328, signal_1390}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1191 ( .s ({signal_2214, signal_977}), .b ({1'b0, 1'b0}), .a ({signal_2272, signal_1334}), .clk (CLK), .r (Fresh[63]), .c ({signal_2329, signal_1391}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1192 ( .s ({signal_2214, signal_977}), .b ({signal_2273, signal_1335}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[64]), .c ({signal_2330, signal_1392}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1193 ( .s ({signal_2214, signal_977}), .b ({signal_2272, signal_1334}), .a ({signal_2273, signal_1335}), .clk (CLK), .r (Fresh[65]), .c ({signal_2331, signal_1393}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1194 ( .s ({signal_2221, signal_965}), .b ({1'b0, 1'b0}), .a ({signal_2274, signal_1336}), .clk (CLK), .r (Fresh[66]), .c ({signal_2332, signal_1394}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1195 ( .s ({signal_2221, signal_965}), .b ({signal_2275, signal_1337}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[67]), .c ({signal_2333, signal_1395}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1196 ( .s ({signal_2221, signal_965}), .b ({signal_2274, signal_1336}), .a ({signal_2275, signal_1337}), .clk (CLK), .r (Fresh[68]), .c ({signal_2334, signal_1396}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1197 ( .s ({signal_2225, signal_961}), .b ({1'b0, 1'b0}), .a ({signal_2276, signal_1338}), .clk (CLK), .r (Fresh[69]), .c ({signal_2335, signal_1397}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1198 ( .s ({signal_2225, signal_961}), .b ({signal_2277, signal_1339}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[70]), .c ({signal_2336, signal_1398}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1199 ( .s ({signal_2225, signal_961}), .b ({signal_2276, signal_1338}), .a ({signal_2277, signal_1339}), .clk (CLK), .r (Fresh[71]), .c ({signal_2337, signal_1399}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1200 ( .s ({signal_2237, signal_949}), .b ({1'b0, 1'b0}), .a ({signal_2278, signal_1340}), .clk (CLK), .r (Fresh[72]), .c ({signal_2338, signal_1400}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1201 ( .s ({signal_2237, signal_949}), .b ({signal_2279, signal_1341}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[73]), .c ({signal_2339, signal_1401}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1202 ( .s ({signal_2237, signal_949}), .b ({signal_2278, signal_1340}), .a ({signal_2279, signal_1341}), .clk (CLK), .r (Fresh[74]), .c ({signal_2340, signal_1402}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1203 ( .s ({signal_2241, signal_945}), .b ({1'b0, 1'b0}), .a ({signal_2280, signal_1342}), .clk (CLK), .r (Fresh[75]), .c ({signal_2341, signal_1403}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1204 ( .s ({signal_2241, signal_945}), .b ({signal_2281, signal_1343}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[76]), .c ({signal_2342, signal_1404}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1205 ( .s ({signal_2241, signal_945}), .b ({signal_2280, signal_1342}), .a ({signal_2281, signal_1343}), .clk (CLK), .r (Fresh[77]), .c ({signal_2343, signal_1405}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1206 ( .s ({signal_2260, signal_1005}), .b ({signal_2291, signal_1345}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[78]), .c ({signal_2380, signal_1406}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1207 ( .s ({signal_2260, signal_1005}), .b ({signal_2292, signal_1346}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[79]), .c ({signal_2381, signal_1407}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1208 ( .s ({signal_2248, signal_1002}), .b ({1'b0, 1'b0}), .a ({signal_2294, signal_1348}), .clk (CLK), .r (Fresh[80]), .c ({signal_2382, signal_1408}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1209 ( .s ({signal_2248, signal_1002}), .b ({1'b0, 1'b1}), .a ({signal_2294, signal_1348}), .clk (CLK), .r (Fresh[81]), .c ({signal_2383, signal_1409}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1210 ( .s ({signal_2264, signal_989}), .b ({signal_2297, signal_1351}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[82]), .c ({signal_2384, signal_1410}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1211 ( .s ({signal_2264, signal_989}), .b ({signal_2298, signal_1352}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[83]), .c ({signal_2385, signal_1411}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1212 ( .s ({signal_2261, signal_986}), .b ({1'b0, 1'b1}), .a ({signal_2300, signal_1354}), .clk (CLK), .r (Fresh[84]), .c ({signal_2386, signal_1412}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1213 ( .s ({signal_2261, signal_986}), .b ({1'b0, 1'b0}), .a ({signal_2300, signal_1354}), .clk (CLK), .r (Fresh[85]), .c ({signal_2387, signal_1413}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1214 ( .s ({signal_2246, signal_975}), .b ({signal_2302, signal_1357}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[86]), .c ({signal_2388, signal_1414}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1215 ( .s ({signal_2246, signal_975}), .b ({1'b0, 1'b1}), .a ({signal_2303, signal_1358}), .clk (CLK), .r (Fresh[87]), .c ({signal_2389, signal_1415}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1216 ( .s ({signal_2257, signal_969}), .b ({signal_2305, signal_1360}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[88]), .c ({signal_2390, signal_1416}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1217 ( .s ({signal_2257, signal_969}), .b ({signal_2306, signal_1361}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[89]), .c ({signal_2391, signal_1417}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1218 ( .s ({signal_2255, signal_958}), .b ({1'b0, 1'b0}), .a ({signal_2308, signal_1363}), .clk (CLK), .r (Fresh[90]), .c ({signal_2392, signal_1418}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1219 ( .s ({signal_2255, signal_958}), .b ({1'b0, 1'b1}), .a ({signal_2308, signal_1363}), .clk (CLK), .r (Fresh[91]), .c ({signal_2393, signal_1419}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1220 ( .s ({signal_2250, signal_954}), .b ({1'b0, 1'b0}), .a ({signal_2311, signal_1366}), .clk (CLK), .r (Fresh[92]), .c ({signal_2394, signal_1420}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1221 ( .s ({signal_2250, signal_954}), .b ({1'b0, 1'b1}), .a ({signal_2311, signal_1366}), .clk (CLK), .r (Fresh[93]), .c ({signal_2395, signal_1421}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1222 ( .s ({signal_2221, signal_965}), .b ({signal_2275, signal_1337}), .a ({signal_2274, signal_1336}), .clk (CLK), .r (Fresh[94]), .c ({signal_2344, signal_1422}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1223 ( .s ({signal_2221, signal_965}), .b ({1'b0, 1'b1}), .a ({signal_2275, signal_1337}), .clk (CLK), .r (Fresh[95]), .c ({signal_2345, signal_1423}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1224 ( .s ({signal_2221, signal_965}), .b ({signal_2274, signal_1336}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[96]), .c ({signal_2346, signal_1424}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1225 ( .s ({signal_2221, signal_965}), .b ({1'b0, 1'b0}), .a ({signal_2275, signal_1337}), .clk (CLK), .r (Fresh[97]), .c ({signal_2347, signal_1425}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1226 ( .s ({signal_2221, signal_965}), .b ({1'b0, 1'b1}), .a ({signal_2274, signal_1336}), .clk (CLK), .r (Fresh[98]), .c ({signal_2348, signal_1426}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1227 ( .s ({signal_2241, signal_945}), .b ({1'b0, 1'b0}), .a ({signal_2281, signal_1343}), .clk (CLK), .r (Fresh[99]), .c ({signal_2349, signal_1427}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1228 ( .s ({signal_2241, signal_945}), .b ({1'b0, 1'b1}), .a ({signal_2280, signal_1342}), .clk (CLK), .r (Fresh[100]), .c ({signal_2350, signal_1428}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1229 ( .s ({signal_2241, signal_945}), .b ({signal_2281, signal_1343}), .a ({signal_2280, signal_1342}), .clk (CLK), .r (Fresh[101]), .c ({signal_2351, signal_1429}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1230 ( .s ({signal_2225, signal_961}), .b ({signal_2277, signal_1339}), .a ({signal_2276, signal_1338}), .clk (CLK), .r (Fresh[102]), .c ({signal_2352, signal_1430}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1231 ( .s ({signal_2225, signal_961}), .b ({1'b0, 1'b0}), .a ({signal_2277, signal_1339}), .clk (CLK), .r (Fresh[103]), .c ({signal_2353, signal_1431}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1232 ( .s ({signal_2225, signal_961}), .b ({1'b0, 1'b1}), .a ({signal_2276, signal_1338}), .clk (CLK), .r (Fresh[104]), .c ({signal_2354, signal_1432}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1233 ( .s ({signal_2255, signal_958}), .b ({signal_2307, signal_1362}), .a ({signal_2308, signal_1363}), .clk (CLK), .r (Fresh[105]), .c ({signal_2396, signal_1433}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1234 ( .s ({signal_2255, signal_958}), .b ({1'b0, 1'b0}), .a ({signal_2307, signal_1362}), .clk (CLK), .r (Fresh[106]), .c ({signal_2397, signal_1434}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1235 ( .s ({signal_2225, signal_961}), .b ({1'b0, 1'b1}), .a ({signal_2277, signal_1339}), .clk (CLK), .r (Fresh[107]), .c ({signal_2355, signal_1435}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1236 ( .s ({signal_2225, signal_961}), .b ({signal_2276, signal_1338}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[108]), .c ({signal_2356, signal_1436}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1237 ( .s ({signal_2214, signal_977}), .b ({signal_2273, signal_1335}), .a ({signal_2272, signal_1334}), .clk (CLK), .r (Fresh[109]), .c ({signal_2357, signal_1437}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1238 ( .s ({signal_2214, signal_977}), .b ({1'b0, 1'b1}), .a ({signal_2273, signal_1335}), .clk (CLK), .r (Fresh[110]), .c ({signal_2358, signal_1438}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1239 ( .s ({signal_2214, signal_977}), .b ({signal_2272, signal_1334}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[111]), .c ({signal_2359, signal_1439}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1240 ( .s ({signal_2246, signal_975}), .b ({signal_2302, signal_1357}), .a ({signal_2303, signal_1358}), .clk (CLK), .r (Fresh[112]), .c ({signal_2398, signal_1440}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1241 ( .s ({signal_2246, signal_975}), .b ({1'b0, 1'b0}), .a ({signal_2302, signal_1357}), .clk (CLK), .r (Fresh[113]), .c ({signal_2399, signal_1441}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1242 ( .s ({signal_2237, signal_949}), .b ({signal_2279, signal_1341}), .a ({signal_2278, signal_1340}), .clk (CLK), .r (Fresh[114]), .c ({signal_2360, signal_1442}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1243 ( .s ({signal_2222, signal_964}), .b ({signal_2301, signal_1355}), .a ({signal_2315, signal_1373}), .clk (CLK), .r (Fresh[115]), .c ({signal_2400, signal_1443}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1244 ( .s ({signal_2222, signal_964}), .b ({signal_2315, signal_1373}), .a ({signal_2301, signal_1355}), .clk (CLK), .r (Fresh[116]), .c ({signal_2401, signal_1444}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1245 ( .s ({signal_2261, signal_986}), .b ({1'b0, 1'b0}), .a ({signal_2299, signal_1353}), .clk (CLK), .r (Fresh[117]), .c ({signal_2402, signal_1445}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1246 ( .s ({signal_2261, signal_986}), .b ({signal_2300, signal_1354}), .a ({signal_2299, signal_1353}), .clk (CLK), .r (Fresh[118]), .c ({signal_2403, signal_1446}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1247 ( .s ({signal_2261, signal_986}), .b ({signal_2299, signal_1353}), .a ({signal_2300, signal_1354}), .clk (CLK), .r (Fresh[119]), .c ({signal_2404, signal_1447}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1248 ( .s ({signal_2262, signal_987}), .b ({signal_2291, signal_1345}), .a ({signal_2292, signal_1346}), .clk (CLK), .r (Fresh[120]), .c ({signal_2405, signal_1448}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1249 ( .s ({signal_2262, signal_987}), .b ({signal_2292, signal_1346}), .a ({signal_2291, signal_1345}), .clk (CLK), .r (Fresh[121]), .c ({signal_2406, signal_1449}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1250 ( .s ({signal_2260, signal_1005}), .b ({signal_2299, signal_1353}), .a ({signal_2300, signal_1354}), .clk (CLK), .r (Fresh[122]), .c ({signal_2407, signal_1450}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1251 ( .s ({signal_2260, signal_1005}), .b ({signal_2300, signal_1354}), .a ({signal_2299, signal_1353}), .clk (CLK), .r (Fresh[123]), .c ({signal_2408, signal_1451}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1252 ( .s ({signal_2211, signal_982}), .b ({signal_2270, signal_1332}), .a ({signal_2271, signal_1333}), .clk (CLK), .r (Fresh[124]), .c ({signal_2361, signal_1452}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1253 ( .s ({signal_2211, signal_982}), .b ({1'b0, 1'b0}), .a ({signal_2271, signal_1333}), .clk (CLK), .r (Fresh[125]), .c ({signal_2362, signal_1453}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1254 ( .s ({signal_2211, signal_982}), .b ({signal_2270, signal_1332}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[126]), .c ({signal_2363, signal_1454}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1255 ( .s ({signal_2255, signal_958}), .b ({signal_2308, signal_1363}), .a ({signal_2307, signal_1362}), .clk (CLK), .r (Fresh[127]), .c ({signal_2409, signal_1455}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1256 ( .s ({signal_2246, signal_975}), .b ({signal_2303, signal_1358}), .a ({signal_2302, signal_1357}), .clk (CLK), .r (Fresh[128]), .c ({signal_2410, signal_1456}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1257 ( .s ({signal_2200, signal_997}), .b ({1'b0, 1'b0}), .a ({signal_2267, signal_1329}), .clk (CLK), .r (Fresh[129]), .c ({signal_2364, signal_1457}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1258 ( .s ({signal_2200, signal_997}), .b ({1'b0, 1'b1}), .a ({signal_2266, signal_1328}), .clk (CLK), .r (Fresh[130]), .c ({signal_2365, signal_1458}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1259 ( .s ({signal_2200, signal_997}), .b ({signal_2267, signal_1329}), .a ({signal_2266, signal_1328}), .clk (CLK), .r (Fresh[131]), .c ({signal_2366, signal_1459}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1260 ( .s ({signal_2250, signal_954}), .b ({signal_2310, signal_1365}), .a ({signal_2311, signal_1366}), .clk (CLK), .r (Fresh[132]), .c ({signal_2411, signal_1460}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1261 ( .s ({signal_2250, signal_954}), .b ({1'b0, 1'b0}), .a ({signal_2310, signal_1365}), .clk (CLK), .r (Fresh[133]), .c ({signal_2412, signal_1461}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1262 ( .s ({signal_2246, signal_975}), .b ({signal_2303, signal_1358}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[134]), .c ({signal_2413, signal_1462}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1263 ( .s ({signal_2250, signal_954}), .b ({signal_2311, signal_1366}), .a ({signal_2310, signal_1365}), .clk (CLK), .r (Fresh[135]), .c ({signal_2414, signal_1463}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1264 ( .s ({signal_2200, signal_997}), .b ({1'b0, 1'b1}), .a ({signal_2267, signal_1329}), .clk (CLK), .r (Fresh[136]), .c ({signal_2367, signal_1464}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1265 ( .s ({signal_2200, signal_997}), .b ({signal_2266, signal_1328}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[137]), .c ({signal_2368, signal_1465}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1266 ( .s ({signal_2257, signal_969}), .b ({1'b0, 1'b0}), .a ({signal_2306, signal_1361}), .clk (CLK), .r (Fresh[138]), .c ({signal_2415, signal_1466}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1267 ( .s ({signal_2257, signal_969}), .b ({1'b0, 1'b1}), .a ({signal_2305, signal_1360}), .clk (CLK), .r (Fresh[139]), .c ({signal_2416, signal_1467}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1268 ( .s ({signal_2204, signal_993}), .b ({1'b0, 1'b0}), .a ({signal_2269, signal_1331}), .clk (CLK), .r (Fresh[140]), .c ({signal_2369, signal_1468}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1269 ( .s ({signal_2204, signal_993}), .b ({1'b0, 1'b1}), .a ({signal_2268, signal_1330}), .clk (CLK), .r (Fresh[141]), .c ({signal_2370, signal_1469}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1270 ( .s ({signal_2204, signal_993}), .b ({signal_2269, signal_1331}), .a ({signal_2268, signal_1330}), .clk (CLK), .r (Fresh[142]), .c ({signal_2371, signal_1470}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1271 ( .s ({signal_2257, signal_969}), .b ({signal_2305, signal_1360}), .a ({signal_2306, signal_1361}), .clk (CLK), .r (Fresh[143]), .c ({signal_2417, signal_1471}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1272 ( .s ({signal_2257, signal_969}), .b ({signal_2306, signal_1361}), .a ({signal_2305, signal_1360}), .clk (CLK), .r (Fresh[144]), .c ({signal_2418, signal_1472}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1273 ( .s ({signal_2237, signal_949}), .b ({1'b0, 1'b0}), .a ({signal_2279, signal_1341}), .clk (CLK), .r (Fresh[145]), .c ({signal_2372, signal_1473}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1274 ( .s ({signal_2237, signal_949}), .b ({1'b0, 1'b1}), .a ({signal_2278, signal_1340}), .clk (CLK), .r (Fresh[146]), .c ({signal_2373, signal_1474}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1275 ( .s ({signal_2258, signal_970}), .b ({signal_2297, signal_1351}), .a ({signal_2298, signal_1352}), .clk (CLK), .r (Fresh[147]), .c ({signal_2419, signal_1475}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1276 ( .s ({signal_2257, signal_969}), .b ({signal_2297, signal_1351}), .a ({signal_2298, signal_1352}), .clk (CLK), .r (Fresh[148]), .c ({signal_2420, signal_1476}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1277 ( .s ({signal_2264, signal_989}), .b ({signal_2298, signal_1352}), .a ({signal_2297, signal_1351}), .clk (CLK), .r (Fresh[149]), .c ({signal_2421, signal_1477}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1278 ( .s ({signal_2264, signal_989}), .b ({signal_2297, signal_1351}), .a ({signal_2298, signal_1352}), .clk (CLK), .r (Fresh[150]), .c ({signal_2422, signal_1478}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1279 ( .s ({signal_2258, signal_970}), .b ({signal_2296, signal_1350}), .a ({signal_2314, signal_1372}), .clk (CLK), .r (Fresh[151]), .c ({signal_2423, signal_1479}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1280 ( .s ({signal_2257, signal_969}), .b ({signal_2296, signal_1350}), .a ({signal_2314, signal_1372}), .clk (CLK), .r (Fresh[152]), .c ({signal_2424, signal_1480}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1281 ( .s ({signal_2258, signal_970}), .b ({signal_2298, signal_1352}), .a ({signal_2297, signal_1351}), .clk (CLK), .r (Fresh[153]), .c ({signal_2425, signal_1481}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1282 ( .s ({signal_2258, signal_970}), .b ({signal_2314, signal_1372}), .a ({signal_2296, signal_1350}), .clk (CLK), .r (Fresh[154]), .c ({signal_2426, signal_1482}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1283 ( .s ({signal_2241, signal_945}), .b ({1'b0, 1'b1}), .a ({signal_2281, signal_1343}), .clk (CLK), .r (Fresh[155]), .c ({signal_2374, signal_1483}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1284 ( .s ({signal_2241, signal_945}), .b ({signal_2280, signal_1342}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[156]), .c ({signal_2375, signal_1484}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1285 ( .s ({signal_2260, signal_1005}), .b ({signal_2291, signal_1345}), .a ({signal_2292, signal_1346}), .clk (CLK), .r (Fresh[157]), .c ({signal_2427, signal_1485}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1286 ( .s ({signal_2260, signal_1005}), .b ({signal_2292, signal_1346}), .a ({signal_2291, signal_1345}), .clk (CLK), .r (Fresh[158]), .c ({signal_2428, signal_1486}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1287 ( .s ({signal_2260, signal_1005}), .b ({1'b0, 1'b1}), .a ({signal_2291, signal_1345}), .clk (CLK), .r (Fresh[159]), .c ({signal_2429, signal_1487}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1288 ( .s ({signal_2260, signal_1005}), .b ({1'b0, 1'b0}), .a ({signal_2292, signal_1346}), .clk (CLK), .r (Fresh[160]), .c ({signal_2430, signal_1488}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1289 ( .s ({signal_2248, signal_1002}), .b ({signal_2293, signal_1347}), .a ({signal_2294, signal_1348}), .clk (CLK), .r (Fresh[161]), .c ({signal_2431, signal_1489}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1290 ( .s ({signal_2248, signal_1002}), .b ({1'b0, 1'b0}), .a ({signal_2293, signal_1347}), .clk (CLK), .r (Fresh[162]), .c ({signal_2432, signal_1490}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1291 ( .s ({signal_2254, signal_1003}), .b ({signal_2308, signal_1363}), .a ({signal_2307, signal_1362}), .clk (CLK), .r (Fresh[163]), .c ({signal_2433, signal_1491}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1292 ( .s ({signal_2255, signal_958}), .b ({1'b0, 1'b1}), .a ({signal_2307, signal_1362}), .clk (CLK), .r (Fresh[164]), .c ({signal_2434, signal_1492}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1293 ( .s ({signal_2254, signal_1003}), .b ({signal_2309, signal_1364}), .a ({signal_2316, signal_1374}), .clk (CLK), .r (Fresh[165]), .c ({signal_2435, signal_1493}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1294 ( .s ({signal_2254, signal_1003}), .b ({signal_2307, signal_1362}), .a ({signal_2308, signal_1363}), .clk (CLK), .r (Fresh[166]), .c ({signal_2436, signal_1494}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1295 ( .s ({signal_2254, signal_1003}), .b ({signal_2316, signal_1374}), .a ({signal_2309, signal_1364}), .clk (CLK), .r (Fresh[167]), .c ({signal_2437, signal_1495}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1296 ( .s ({signal_2248, signal_1002}), .b ({signal_2294, signal_1348}), .a ({signal_2293, signal_1347}), .clk (CLK), .r (Fresh[168]), .c ({signal_2438, signal_1496}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1297 ( .s ({signal_2250, signal_954}), .b ({1'b0, 1'b1}), .a ({signal_2310, signal_1365}), .clk (CLK), .r (Fresh[169]), .c ({signal_2439, signal_1497}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1298 ( .s ({signal_2237, signal_949}), .b ({1'b0, 1'b1}), .a ({signal_2279, signal_1341}), .clk (CLK), .r (Fresh[170]), .c ({signal_2376, signal_1498}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1299 ( .s ({signal_2237, signal_949}), .b ({signal_2278, signal_1340}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[171]), .c ({signal_2377, signal_1499}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1300 ( .s ({signal_2264, signal_989}), .b ({1'b0, 1'b0}), .a ({signal_2298, signal_1352}), .clk (CLK), .r (Fresh[172]), .c ({signal_2440, signal_1500}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1301 ( .s ({signal_2264, signal_989}), .b ({1'b0, 1'b1}), .a ({signal_2297, signal_1351}), .clk (CLK), .r (Fresh[173]), .c ({signal_2441, signal_1501}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1302 ( .s ({signal_2204, signal_993}), .b ({1'b0, 1'b1}), .a ({signal_2269, signal_1331}), .clk (CLK), .r (Fresh[174]), .c ({signal_2378, signal_1502}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1303 ( .s ({signal_2204, signal_993}), .b ({signal_2268, signal_1330}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[175]), .c ({signal_2379, signal_1503}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1304 ( .s ({signal_2210, signal_984}), .b ({signal_2299, signal_1353}), .a ({signal_2300, signal_1354}), .clk (CLK), .r (Fresh[176]), .c ({signal_2442, signal_1504}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1305 ( .s ({signal_2199, signal_998}), .b ({signal_2321, signal_1383}), .a ({signal_2320, signal_1382}), .clk (CLK), .r (Fresh[177]), .c ({signal_2443, signal_1505}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1306 ( .s ({signal_2199, signal_998}), .b ({signal_2267, signal_1329}), .a ({signal_2322, signal_1384}), .clk (CLK), .r (Fresh[178]), .c ({signal_2444, signal_1506}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1307 ( .s ({signal_2203, signal_994}), .b ({signal_2324, signal_1386}), .a ({signal_2323, signal_1385}), .clk (CLK), .r (Fresh[179]), .c ({signal_2445, signal_1507}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1308 ( .s ({signal_2203, signal_994}), .b ({signal_2269, signal_1331}), .a ({signal_2325, signal_1387}), .clk (CLK), .r (Fresh[180]), .c ({signal_2446, signal_1508}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1309 ( .s ({signal_2078, signal_981}), .b ({signal_2327, signal_1389}), .a ({signal_2326, signal_1388}), .clk (CLK), .r (Fresh[181]), .c ({signal_2447, signal_1509}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1310 ( .s ({signal_2078, signal_981}), .b ({signal_2328, signal_1390}), .a ({signal_2271, signal_1333}), .clk (CLK), .r (Fresh[182]), .c ({signal_2448, signal_1510}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1311 ( .s ({signal_2213, signal_978}), .b ({signal_2330, signal_1392}), .a ({signal_2329, signal_1391}), .clk (CLK), .r (Fresh[183]), .c ({signal_2449, signal_1511}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1312 ( .s ({signal_2213, signal_978}), .b ({signal_2273, signal_1335}), .a ({signal_2331, signal_1393}), .clk (CLK), .r (Fresh[184]), .c ({signal_2450, signal_1512}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1313 ( .s ({signal_2220, signal_966}), .b ({signal_2333, signal_1395}), .a ({signal_2332, signal_1394}), .clk (CLK), .r (Fresh[185]), .c ({signal_2451, signal_1513}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1314 ( .s ({signal_2220, signal_966}), .b ({signal_2275, signal_1337}), .a ({signal_2334, signal_1396}), .clk (CLK), .r (Fresh[186]), .c ({signal_2452, signal_1514}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1315 ( .s ({signal_2224, signal_962}), .b ({signal_2336, signal_1398}), .a ({signal_2335, signal_1397}), .clk (CLK), .r (Fresh[187]), .c ({signal_2453, signal_1515}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1316 ( .s ({signal_2224, signal_962}), .b ({signal_2277, signal_1339}), .a ({signal_2337, signal_1399}), .clk (CLK), .r (Fresh[188]), .c ({signal_2454, signal_1516}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1317 ( .s ({signal_2236, signal_950}), .b ({signal_2339, signal_1401}), .a ({signal_2338, signal_1400}), .clk (CLK), .r (Fresh[189]), .c ({signal_2455, signal_1517}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1318 ( .s ({signal_2236, signal_950}), .b ({signal_2279, signal_1341}), .a ({signal_2340, signal_1402}), .clk (CLK), .r (Fresh[190]), .c ({signal_2456, signal_1518}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1319 ( .s ({signal_2240, signal_946}), .b ({signal_2342, signal_1404}), .a ({signal_2341, signal_1403}), .clk (CLK), .r (Fresh[191]), .c ({signal_2457, signal_1519}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1320 ( .s ({signal_2240, signal_946}), .b ({signal_2281, signal_1343}), .a ({signal_2343, signal_1405}), .clk (CLK), .r (Fresh[192]), .c ({signal_2458, signal_1520}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1321 ( .s ({signal_2191, signal_1007}), .b ({signal_2380, signal_1406}), .a ({signal_2290, signal_1344}), .clk (CLK), .r (Fresh[193]), .c ({signal_2499, signal_1521}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1322 ( .s ({signal_2191, signal_1007}), .b ({signal_2381, signal_1407}), .a ({signal_2292, signal_1346}), .clk (CLK), .r (Fresh[194]), .c ({signal_2500, signal_1522}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1323 ( .s ({signal_2247, signal_1001}), .b ({signal_2382, signal_1408}), .a ({signal_2293, signal_1347}), .clk (CLK), .r (Fresh[195]), .c ({signal_2501, signal_1523}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1324 ( .s ({signal_2247, signal_1001}), .b ({signal_2295, signal_1349}), .a ({signal_2383, signal_1409}), .clk (CLK), .r (Fresh[196]), .c ({signal_2502, signal_1524}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1325 ( .s ({signal_2190, signal_991}), .b ({signal_2384, signal_1410}), .a ({signal_2296, signal_1350}), .clk (CLK), .r (Fresh[197]), .c ({signal_2503, signal_1525}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1326 ( .s ({signal_2190, signal_991}), .b ({signal_2385, signal_1411}), .a ({signal_2298, signal_1352}), .clk (CLK), .r (Fresh[198]), .c ({signal_2504, signal_1526}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1327 ( .s ({signal_2210, signal_984}), .b ({signal_2386, signal_1412}), .a ({signal_2299, signal_1353}), .clk (CLK), .r (Fresh[199]), .c ({signal_2505, signal_1527}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1328 ( .s ({signal_2210, signal_984}), .b ({signal_2301, signal_1355}), .a ({signal_2387, signal_1413}), .clk (CLK), .r (Fresh[200]), .c ({signal_2506, signal_1528}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1329 ( .s ({signal_2245, signal_973}), .b ({signal_2388, signal_1414}), .a ({signal_2282, signal_1356}), .clk (CLK), .r (Fresh[201]), .c ({signal_2507, signal_1529}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1330 ( .s ({signal_2245, signal_973}), .b ({signal_2303, signal_1358}), .a ({signal_2389, signal_1415}), .clk (CLK), .r (Fresh[202]), .c ({signal_2508, signal_1530}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1331 ( .s ({signal_2243, signal_971}), .b ({signal_2390, signal_1416}), .a ({signal_2304, signal_1359}), .clk (CLK), .r (Fresh[203]), .c ({signal_2509, signal_1531}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1332 ( .s ({signal_2243, signal_971}), .b ({signal_2391, signal_1417}), .a ({signal_2306, signal_1361}), .clk (CLK), .r (Fresh[204]), .c ({signal_2510, signal_1532}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1333 ( .s ({signal_2253, signal_957}), .b ({signal_2392, signal_1418}), .a ({signal_2307, signal_1362}), .clk (CLK), .r (Fresh[205]), .c ({signal_2511, signal_1533}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1334 ( .s ({signal_2253, signal_957}), .b ({signal_2309, signal_1364}), .a ({signal_2393, signal_1419}), .clk (CLK), .r (Fresh[206]), .c ({signal_2512, signal_1534}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1335 ( .s ({signal_2249, signal_953}), .b ({signal_2394, signal_1420}), .a ({signal_2310, signal_1365}), .clk (CLK), .r (Fresh[207]), .c ({signal_2513, signal_1535}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1336 ( .s ({signal_2249, signal_953}), .b ({signal_2312, signal_1367}), .a ({signal_2395, signal_1421}), .clk (CLK), .r (Fresh[208]), .c ({signal_2514, signal_1536}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1337 ( .s ({signal_2220, signal_966}), .b ({signal_2274, signal_1336}), .a ({signal_2344, signal_1422}), .clk (CLK), .r (Fresh[209]), .c ({signal_2459, signal_1537}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1338 ( .s ({signal_2220, signal_966}), .b ({signal_2346, signal_1424}), .a ({signal_2345, signal_1423}), .clk (CLK), .r (Fresh[210]), .c ({signal_2460, signal_1538}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1339 ( .s ({signal_2220, signal_966}), .b ({signal_2344, signal_1422}), .a ({signal_2275, signal_1337}), .clk (CLK), .r (Fresh[211]), .c ({signal_2461, signal_1539}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1340 ( .s ({signal_2220, signal_966}), .b ({signal_2334, signal_1396}), .a ({signal_2274, signal_1336}), .clk (CLK), .r (Fresh[212]), .c ({signal_2462, signal_1540}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1341 ( .s ({signal_2220, signal_966}), .b ({signal_2348, signal_1426}), .a ({signal_2347, signal_1425}), .clk (CLK), .r (Fresh[213]), .c ({signal_2463, signal_1541}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1342 ( .s ({signal_2220, signal_966}), .b ({signal_2344, signal_1422}), .a ({signal_2283, signal_1368}), .clk (CLK), .r (Fresh[214]), .c ({signal_2464, signal_1542}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1343 ( .s ({signal_2240, signal_946}), .b ({signal_2350, signal_1428}), .a ({signal_2349, signal_1427}), .clk (CLK), .r (Fresh[215]), .c ({signal_2465, signal_1543}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1344 ( .s ({signal_2240, signal_946}), .b ({signal_2351, signal_1429}), .a ({signal_2284, signal_1369}), .clk (CLK), .r (Fresh[216]), .c ({signal_2466, signal_1544}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1345 ( .s ({signal_2240, signal_946}), .b ({signal_2351, signal_1429}), .a ({signal_2281, signal_1343}), .clk (CLK), .r (Fresh[217]), .c ({signal_2467, signal_1545}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1346 ( .s ({signal_2240, signal_946}), .b ({signal_2343, signal_1405}), .a ({signal_2280, signal_1342}), .clk (CLK), .r (Fresh[218]), .c ({signal_2468, signal_1546}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1347 ( .s ({signal_2224, signal_962}), .b ({signal_2352, signal_1430}), .a ({signal_2277, signal_1339}), .clk (CLK), .r (Fresh[219]), .c ({signal_2469, signal_1547}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1348 ( .s ({signal_2224, signal_962}), .b ({signal_2337, signal_1399}), .a ({signal_2276, signal_1338}), .clk (CLK), .r (Fresh[220]), .c ({signal_2470, signal_1548}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1349 ( .s ({signal_2224, signal_962}), .b ({signal_2354, signal_1432}), .a ({signal_2353, signal_1431}), .clk (CLK), .r (Fresh[221]), .c ({signal_2471, signal_1549}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1350 ( .s ({signal_2224, signal_962}), .b ({signal_2352, signal_1430}), .a ({signal_2285, signal_1370}), .clk (CLK), .r (Fresh[222]), .c ({signal_2472, signal_1550}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1351 ( .s ({signal_2253, signal_957}), .b ({signal_2396, signal_1433}), .a ({signal_2309, signal_1364}), .clk (CLK), .r (Fresh[223]), .c ({signal_2515, signal_1551}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1352 ( .s ({signal_2253, signal_957}), .b ({signal_2393, signal_1419}), .a ({signal_2397, signal_1434}), .clk (CLK), .r (Fresh[224]), .c ({signal_2516, signal_1552}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1353 ( .s ({signal_2224, signal_962}), .b ({signal_2276, signal_1338}), .a ({signal_2352, signal_1430}), .clk (CLK), .r (Fresh[225]), .c ({signal_2473, signal_1553}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1354 ( .s ({signal_2224, signal_962}), .b ({signal_2356, signal_1436}), .a ({signal_2355, signal_1435}), .clk (CLK), .r (Fresh[226]), .c ({signal_2474, signal_1554}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1355 ( .s ({signal_2213, signal_978}), .b ({signal_2272, signal_1334}), .a ({signal_2357, signal_1437}), .clk (CLK), .r (Fresh[227]), .c ({signal_2475, signal_1555}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1356 ( .s ({signal_2213, signal_978}), .b ({signal_2359, signal_1439}), .a ({signal_2358, signal_1438}), .clk (CLK), .r (Fresh[228]), .c ({signal_2476, signal_1556}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1357 ( .s ({signal_2245, signal_973}), .b ({signal_2398, signal_1440}), .a ({signal_2303, signal_1358}), .clk (CLK), .r (Fresh[229]), .c ({signal_2517, signal_1557}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1358 ( .s ({signal_2245, signal_973}), .b ({signal_2389, signal_1415}), .a ({signal_2399, signal_1441}), .clk (CLK), .r (Fresh[230]), .c ({signal_2518, signal_1558}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1359 ( .s ({signal_2243, signal_971}), .b ({signal_2313, signal_1371}), .a ({signal_2391, signal_1417}), .clk (CLK), .r (Fresh[231]), .c ({signal_2519, signal_1559}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1360 ( .s ({signal_2243, signal_971}), .b ({signal_2305, signal_1360}), .a ({signal_2390, signal_1416}), .clk (CLK), .r (Fresh[232]), .c ({signal_2520, signal_1560}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1361 ( .s ({signal_2190, signal_991}), .b ({signal_2314, signal_1372}), .a ({signal_2385, signal_1411}), .clk (CLK), .r (Fresh[233]), .c ({signal_2521, signal_1561}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1362 ( .s ({signal_2190, signal_991}), .b ({signal_2297, signal_1351}), .a ({signal_2384, signal_1410}), .clk (CLK), .r (Fresh[234]), .c ({signal_2522, signal_1562}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1363 ( .s ({signal_2236, signal_950}), .b ({signal_2360, signal_1442}), .a ({signal_2279, signal_1341}), .clk (CLK), .r (Fresh[235]), .c ({signal_2477, signal_1563}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1364 ( .s ({signal_2236, signal_950}), .b ({signal_2340, signal_1402}), .a ({signal_2278, signal_1340}), .clk (CLK), .r (Fresh[236]), .c ({signal_2478, signal_1564}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1365 ( .s ({signal_2210, signal_984}), .b ({signal_2387, signal_1413}), .a ({signal_2299, signal_1353}), .clk (CLK), .r (Fresh[237]), .c ({signal_2523, signal_1565}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1366 ( .s ({signal_2210, signal_984}), .b ({signal_2315, signal_1373}), .a ({signal_2386, signal_1412}), .clk (CLK), .r (Fresh[238]), .c ({signal_2524, signal_1566}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1367 ( .s ({signal_2221, signal_965}), .b ({signal_2401, signal_1444}), .a ({signal_2400, signal_1443}), .clk (CLK), .r (Fresh[239]), .c ({signal_2525, signal_1567}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1368 ( .s ({signal_2221, signal_965}), .b ({signal_2315, signal_1373}), .a ({signal_2401, signal_1444}), .clk (CLK), .r (Fresh[240]), .c ({signal_2526, signal_1568}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1369 ( .s ({signal_2221, signal_965}), .b ({signal_2400, signal_1443}), .a ({signal_2301, signal_1355}), .clk (CLK), .r (Fresh[241]), .c ({signal_2527, signal_1569}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1370 ( .s ({signal_2222, signal_964}), .b ({signal_2402, signal_1445}), .a ({signal_2386, signal_1412}), .clk (CLK), .r (Fresh[242]), .c ({signal_2528, signal_1570}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1371 ( .s ({signal_2222, signal_964}), .b ({signal_2386, signal_1412}), .a ({signal_2402, signal_1445}), .clk (CLK), .r (Fresh[243]), .c ({signal_2529, signal_1571}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1372 ( .s ({signal_2222, signal_964}), .b ({signal_2404, signal_1447}), .a ({signal_2403, signal_1446}), .clk (CLK), .r (Fresh[244]), .c ({signal_2530, signal_1572}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1373 ( .s ({signal_2222, signal_964}), .b ({signal_2403, signal_1446}), .a ({signal_2404, signal_1447}), .clk (CLK), .r (Fresh[245]), .c ({signal_2531, signal_1573}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1374 ( .s ({signal_2261, signal_986}), .b ({signal_2406, signal_1449}), .a ({signal_2405, signal_1448}), .clk (CLK), .r (Fresh[246]), .c ({signal_2532, signal_1574}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1375 ( .s ({signal_2261, signal_986}), .b ({signal_2405, signal_1448}), .a ({signal_2406, signal_1449}), .clk (CLK), .r (Fresh[247]), .c ({signal_2533, signal_1575}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1376 ( .s ({signal_2210, signal_984}), .b ({signal_2406, signal_1449}), .a ({signal_2405, signal_1448}), .clk (CLK), .r (Fresh[248]), .c ({signal_2534, signal_1576}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1377 ( .s ({signal_2260, signal_1005}), .b ({signal_2406, signal_1449}), .a ({signal_2405, signal_1448}), .clk (CLK), .r (Fresh[249]), .c ({signal_2535, signal_1577}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1378 ( .s ({signal_2260, signal_1005}), .b ({signal_2405, signal_1448}), .a ({signal_2406, signal_1449}), .clk (CLK), .r (Fresh[250]), .c ({signal_2536, signal_1578}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1379 ( .s ({signal_2260, signal_1005}), .b ({signal_2403, signal_1446}), .a ({signal_2404, signal_1447}), .clk (CLK), .r (Fresh[251]), .c ({signal_2537, signal_1579}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1380 ( .s ({signal_2260, signal_1005}), .b ({signal_2404, signal_1447}), .a ({signal_2403, signal_1446}), .clk (CLK), .r (Fresh[252]), .c ({signal_2538, signal_1580}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1381 ( .s ({signal_2210, signal_984}), .b ({signal_2408, signal_1451}), .a ({signal_2407, signal_1450}), .clk (CLK), .r (Fresh[253]), .c ({signal_2539, signal_1581}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1382 ( .s ({signal_2253, signal_957}), .b ({signal_2393, signal_1419}), .a ({signal_2307, signal_1362}), .clk (CLK), .r (Fresh[254]), .c ({signal_2540, signal_1582}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1383 ( .s ({signal_2253, signal_957}), .b ({signal_2316, signal_1374}), .a ({signal_2392, signal_1418}), .clk (CLK), .r (Fresh[255]), .c ({signal_2541, signal_1583}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1384 ( .s ({signal_2078, signal_981}), .b ({signal_2361, signal_1452}), .a ({signal_2270, signal_1332}), .clk (CLK), .r (Fresh[256]), .c ({signal_2479, signal_1584}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1385 ( .s ({signal_2078, signal_981}), .b ({signal_2363, signal_1454}), .a ({signal_2362, signal_1453}), .clk (CLK), .r (Fresh[257]), .c ({signal_2480, signal_1585}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1386 ( .s ({signal_2253, signal_957}), .b ({signal_2308, signal_1363}), .a ({signal_2396, signal_1433}), .clk (CLK), .r (Fresh[258]), .c ({signal_2542, signal_1586}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1387 ( .s ({signal_2253, signal_957}), .b ({signal_2307, signal_1362}), .a ({signal_2409, signal_1455}), .clk (CLK), .r (Fresh[259]), .c ({signal_2543, signal_1587}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1388 ( .s ({signal_2247, signal_1001}), .b ({signal_2383, signal_1409}), .a ({signal_2293, signal_1347}), .clk (CLK), .r (Fresh[260]), .c ({signal_2544, signal_1588}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1389 ( .s ({signal_2247, signal_1001}), .b ({signal_2317, signal_1375}), .a ({signal_2382, signal_1408}), .clk (CLK), .r (Fresh[261]), .c ({signal_2545, signal_1589}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1390 ( .s ({signal_2245, signal_973}), .b ({signal_2389, signal_1415}), .a ({signal_2282, signal_1356}), .clk (CLK), .r (Fresh[262]), .c ({signal_2546, signal_1590}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1391 ( .s ({signal_2245, signal_973}), .b ({signal_2302, signal_1357}), .a ({signal_2388, signal_1414}), .clk (CLK), .r (Fresh[263]), .c ({signal_2547, signal_1591}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1392 ( .s ({signal_2249, signal_953}), .b ({signal_2395, signal_1421}), .a ({signal_2310, signal_1365}), .clk (CLK), .r (Fresh[264]), .c ({signal_2548, signal_1592}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1393 ( .s ({signal_2249, signal_953}), .b ({signal_2318, signal_1376}), .a ({signal_2394, signal_1420}), .clk (CLK), .r (Fresh[265]), .c ({signal_2549, signal_1593}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1394 ( .s ({signal_2245, signal_973}), .b ({signal_2286, signal_1377}), .a ({signal_2398, signal_1440}), .clk (CLK), .r (Fresh[266]), .c ({signal_2550, signal_1594}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1395 ( .s ({signal_2245, signal_973}), .b ({signal_2282, signal_1356}), .a ({signal_2410, signal_1456}), .clk (CLK), .r (Fresh[267]), .c ({signal_2551, signal_1595}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1396 ( .s ({signal_2199, signal_998}), .b ({signal_2365, signal_1458}), .a ({signal_2364, signal_1457}), .clk (CLK), .r (Fresh[268]), .c ({signal_2481, signal_1596}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1397 ( .s ({signal_2199, signal_998}), .b ({signal_2366, signal_1459}), .a ({signal_2287, signal_1378}), .clk (CLK), .r (Fresh[269]), .c ({signal_2482, signal_1597}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1398 ( .s ({signal_2249, signal_953}), .b ({signal_2411, signal_1460}), .a ({signal_2312, signal_1367}), .clk (CLK), .r (Fresh[270]), .c ({signal_2552, signal_1598}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1399 ( .s ({signal_2249, signal_953}), .b ({signal_2395, signal_1421}), .a ({signal_2412, signal_1461}), .clk (CLK), .r (Fresh[271]), .c ({signal_2553, signal_1599}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1400 ( .s ({signal_2245, signal_973}), .b ({signal_2399, signal_1441}), .a ({signal_2286, signal_1377}), .clk (CLK), .r (Fresh[272]), .c ({signal_2554, signal_1600}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1401 ( .s ({signal_2245, signal_973}), .b ({signal_2303, signal_1358}), .a ({signal_2413, signal_1462}), .clk (CLK), .r (Fresh[273]), .c ({signal_2555, signal_1601}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1402 ( .s ({signal_2249, signal_953}), .b ({signal_2311, signal_1366}), .a ({signal_2411, signal_1460}), .clk (CLK), .r (Fresh[274]), .c ({signal_2556, signal_1602}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1403 ( .s ({signal_2249, signal_953}), .b ({signal_2310, signal_1365}), .a ({signal_2414, signal_1463}), .clk (CLK), .r (Fresh[275]), .c ({signal_2557, signal_1603}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1404 ( .s ({signal_2199, signal_998}), .b ({signal_2266, signal_1328}), .a ({signal_2366, signal_1459}), .clk (CLK), .r (Fresh[276]), .c ({signal_2483, signal_1604}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1405 ( .s ({signal_2199, signal_998}), .b ({signal_2368, signal_1465}), .a ({signal_2367, signal_1464}), .clk (CLK), .r (Fresh[277]), .c ({signal_2484, signal_1605}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1406 ( .s ({signal_2243, signal_971}), .b ({signal_2416, signal_1467}), .a ({signal_2415, signal_1466}), .clk (CLK), .r (Fresh[278]), .c ({signal_2558, signal_1606}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1407 ( .s ({signal_2243, signal_971}), .b ({signal_2415, signal_1466}), .a ({signal_2416, signal_1467}), .clk (CLK), .r (Fresh[279]), .c ({signal_2559, signal_1607}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1408 ( .s ({signal_2203, signal_994}), .b ({signal_2370, signal_1469}), .a ({signal_2369, signal_1468}), .clk (CLK), .r (Fresh[280]), .c ({signal_2485, signal_1608}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1409 ( .s ({signal_2203, signal_994}), .b ({signal_2371, signal_1470}), .a ({signal_2288, signal_1379}), .clk (CLK), .r (Fresh[281]), .c ({signal_2486, signal_1609}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1410 ( .s ({signal_2243, signal_971}), .b ({signal_2417, signal_1471}), .a ({signal_2306, signal_1361}), .clk (CLK), .r (Fresh[282]), .c ({signal_2560, signal_1610}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1411 ( .s ({signal_2243, signal_971}), .b ({signal_2313, signal_1371}), .a ({signal_2418, signal_1472}), .clk (CLK), .r (Fresh[283]), .c ({signal_2561, signal_1611}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1412 ( .s ({signal_2236, signal_950}), .b ({signal_2373, signal_1474}), .a ({signal_2372, signal_1473}), .clk (CLK), .r (Fresh[284]), .c ({signal_2487, signal_1612}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1413 ( .s ({signal_2236, signal_950}), .b ({signal_2360, signal_1442}), .a ({signal_2289, signal_1380}), .clk (CLK), .r (Fresh[285]), .c ({signal_2488, signal_1613}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1414 ( .s ({signal_2257, signal_969}), .b ({signal_2419, signal_1475}), .a ({signal_2297, signal_1351}), .clk (CLK), .r (Fresh[286]), .c ({signal_2562, signal_1614}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1415 ( .s ({signal_2258, signal_970}), .b ({signal_2421, signal_1477}), .a ({signal_2422, signal_1478}), .clk (CLK), .r (Fresh[287]), .c ({signal_2563, signal_1615}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1416 ( .s ({signal_2257, signal_969}), .b ({signal_2421, signal_1477}), .a ({signal_2422, signal_1478}), .clk (CLK), .r (Fresh[288]), .c ({signal_2564, signal_1616}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1417 ( .s ({signal_2258, signal_970}), .b ({signal_2422, signal_1478}), .a ({signal_2421, signal_1477}), .clk (CLK), .r (Fresh[289]), .c ({signal_2565, signal_1617}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1418 ( .s ({signal_2257, signal_969}), .b ({signal_2422, signal_1478}), .a ({signal_2421, signal_1477}), .clk (CLK), .r (Fresh[290]), .c ({signal_2566, signal_1618}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1419 ( .s ({signal_2257, signal_969}), .b ({signal_2423, signal_1479}), .a ({signal_2296, signal_1350}), .clk (CLK), .r (Fresh[291]), .c ({signal_2567, signal_1619}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1420 ( .s ({signal_2257, signal_969}), .b ({signal_2425, signal_1481}), .a ({signal_2298, signal_1352}), .clk (CLK), .r (Fresh[292]), .c ({signal_2568, signal_1620}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1421 ( .s ({signal_2257, signal_969}), .b ({signal_2426, signal_1482}), .a ({signal_2314, signal_1372}), .clk (CLK), .r (Fresh[293]), .c ({signal_2569, signal_1621}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1422 ( .s ({signal_2240, signal_946}), .b ({signal_2280, signal_1342}), .a ({signal_2351, signal_1429}), .clk (CLK), .r (Fresh[294]), .c ({signal_2489, signal_1622}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1423 ( .s ({signal_2240, signal_946}), .b ({signal_2375, signal_1484}), .a ({signal_2374, signal_1483}), .clk (CLK), .r (Fresh[295]), .c ({signal_2490, signal_1623}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1424 ( .s ({signal_2191, signal_1007}), .b ({signal_2427, signal_1485}), .a ({signal_2292, signal_1346}), .clk (CLK), .r (Fresh[296]), .c ({signal_2570, signal_1624}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1425 ( .s ({signal_2191, signal_1007}), .b ({signal_2319, signal_1381}), .a ({signal_2428, signal_1486}), .clk (CLK), .r (Fresh[297]), .c ({signal_2571, signal_1625}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1426 ( .s ({signal_2242, signal_944}), .b ({signal_2430, signal_1488}), .a ({signal_2429, signal_1487}), .clk (CLK), .r (Fresh[298]), .c ({signal_2572, signal_1626}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1427 ( .s ({signal_2242, signal_944}), .b ({signal_2429, signal_1487}), .a ({signal_2430, signal_1488}), .clk (CLK), .r (Fresh[299]), .c ({signal_2573, signal_1627}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1428 ( .s ({signal_2191, signal_1007}), .b ({signal_2319, signal_1381}), .a ({signal_2381, signal_1407}), .clk (CLK), .r (Fresh[300]), .c ({signal_2574, signal_1628}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1429 ( .s ({signal_2191, signal_1007}), .b ({signal_2291, signal_1345}), .a ({signal_2380, signal_1406}), .clk (CLK), .r (Fresh[301]), .c ({signal_2575, signal_1629}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1430 ( .s ({signal_2247, signal_1001}), .b ({signal_2431, signal_1489}), .a ({signal_2295, signal_1349}), .clk (CLK), .r (Fresh[302]), .c ({signal_2576, signal_1630}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1431 ( .s ({signal_2247, signal_1001}), .b ({signal_2383, signal_1409}), .a ({signal_2432, signal_1490}), .clk (CLK), .r (Fresh[303]), .c ({signal_2577, signal_1631}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1432 ( .s ({signal_2254, signal_1003}), .b ({signal_2397, signal_1434}), .a ({signal_2393, signal_1419}), .clk (CLK), .r (Fresh[304]), .c ({signal_2578, signal_1632}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1433 ( .s ({signal_2254, signal_1003}), .b ({signal_2434, signal_1492}), .a ({signal_2392, signal_1418}), .clk (CLK), .r (Fresh[305]), .c ({signal_2579, signal_1633}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1434 ( .s ({signal_2254, signal_1003}), .b ({signal_2393, signal_1419}), .a ({signal_2397, signal_1434}), .clk (CLK), .r (Fresh[306]), .c ({signal_2580, signal_1634}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1435 ( .s ({signal_2254, signal_1003}), .b ({signal_2392, signal_1418}), .a ({signal_2434, signal_1492}), .clk (CLK), .r (Fresh[307]), .c ({signal_2581, signal_1635}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1436 ( .s ({signal_2247, signal_1001}), .b ({signal_2438, signal_1496}), .a ({signal_2317, signal_1375}), .clk (CLK), .r (Fresh[308]), .c ({signal_2582, signal_1636}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1437 ( .s ({signal_2247, signal_1001}), .b ({signal_2432, signal_1490}), .a ({signal_2383, signal_1409}), .clk (CLK), .r (Fresh[309]), .c ({signal_2583, signal_1637}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1438 ( .s ({signal_2249, signal_953}), .b ({signal_2412, signal_1461}), .a ({signal_2311, signal_1366}), .clk (CLK), .r (Fresh[310]), .c ({signal_2584, signal_1638}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1439 ( .s ({signal_2249, signal_953}), .b ({signal_2312, signal_1367}), .a ({signal_2439, signal_1497}), .clk (CLK), .r (Fresh[311]), .c ({signal_2585, signal_1639}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1440 ( .s ({signal_2213, signal_978}), .b ({signal_2357, signal_1437}), .a ({signal_2273, signal_1335}), .clk (CLK), .r (Fresh[312]), .c ({signal_2491, signal_1640}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1441 ( .s ({signal_2213, signal_978}), .b ({signal_2331, signal_1393}), .a ({signal_2272, signal_1334}), .clk (CLK), .r (Fresh[313]), .c ({signal_2492, signal_1641}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1442 ( .s ({signal_2236, signal_950}), .b ({signal_2278, signal_1340}), .a ({signal_2360, signal_1442}), .clk (CLK), .r (Fresh[314]), .c ({signal_2493, signal_1642}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1443 ( .s ({signal_2236, signal_950}), .b ({signal_2377, signal_1499}), .a ({signal_2376, signal_1498}), .clk (CLK), .r (Fresh[315]), .c ({signal_2494, signal_1643}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1444 ( .s ({signal_2205, signal_992}), .b ({signal_2441, signal_1501}), .a ({signal_2440, signal_1500}), .clk (CLK), .r (Fresh[316]), .c ({signal_2586, signal_1644}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1445 ( .s ({signal_2205, signal_992}), .b ({signal_2440, signal_1500}), .a ({signal_2441, signal_1501}), .clk (CLK), .r (Fresh[317]), .c ({signal_2587, signal_1645}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1446 ( .s ({signal_2204, signal_993}), .b ({signal_2441, signal_1501}), .a ({signal_2440, signal_1500}), .clk (CLK), .r (Fresh[318]), .c ({signal_2588, signal_1646}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1447 ( .s ({signal_2204, signal_993}), .b ({signal_2440, signal_1500}), .a ({signal_2441, signal_1501}), .clk (CLK), .r (Fresh[319]), .c ({signal_2589, signal_1647}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1448 ( .s ({signal_2203, signal_994}), .b ({signal_2268, signal_1330}), .a ({signal_2371, signal_1470}), .clk (CLK), .r (Fresh[320]), .c ({signal_2495, signal_1648}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1449 ( .s ({signal_2203, signal_994}), .b ({signal_2379, signal_1503}), .a ({signal_2378, signal_1502}), .clk (CLK), .r (Fresh[321]), .c ({signal_2496, signal_1649}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1450 ( .s ({signal_2190, signal_991}), .b ({signal_2441, signal_1501}), .a ({signal_2440, signal_1500}), .clk (CLK), .r (Fresh[322]), .c ({signal_2590, signal_1650}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1451 ( .s ({signal_2190, signal_991}), .b ({signal_2440, signal_1500}), .a ({signal_2441, signal_1501}), .clk (CLK), .r (Fresh[323]), .c ({signal_2591, signal_1651}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1452 ( .s ({signal_2210, signal_984}), .b ({signal_2403, signal_1446}), .a ({signal_2404, signal_1447}), .clk (CLK), .r (Fresh[324]), .c ({signal_2592, signal_1652}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1453 ( .s ({signal_2221, signal_965}), .b ({signal_2400, signal_1443}), .a ({signal_2401, signal_1444}), .clk (CLK), .r (Fresh[325]), .c ({signal_2593, signal_1653}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1454 ( .s ({signal_2078, signal_981}), .b ({signal_2271, signal_1333}), .a ({signal_2361, signal_1452}), .clk (CLK), .r (Fresh[326]), .c ({signal_2497, signal_1654}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1455 ( .s ({signal_2078, signal_981}), .b ({signal_2270, signal_1332}), .a ({signal_2328, signal_1390}), .clk (CLK), .r (Fresh[327]), .c ({signal_2498, signal_1655}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1456 ( .s ({signal_2257, signal_969}), .b ({signal_2298, signal_1352}), .a ({signal_2419, signal_1475}), .clk (CLK), .r (Fresh[328]), .c ({signal_2594, signal_1656}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1457 ( .s ({signal_2257, signal_969}), .b ({signal_2297, signal_1351}), .a ({signal_2425, signal_1481}), .clk (CLK), .r (Fresh[329]), .c ({signal_2595, signal_1657}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1458 ( .s ({signal_2257, signal_969}), .b ({signal_2314, signal_1372}), .a ({signal_2423, signal_1479}), .clk (CLK), .r (Fresh[330]), .c ({signal_2596, signal_1658}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1459 ( .s ({signal_2257, signal_969}), .b ({signal_2296, signal_1350}), .a ({signal_2426, signal_1482}), .clk (CLK), .r (Fresh[331]), .c ({signal_2597, signal_1659}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    mux2_masked #(.security_order(1), .pipeline(0)) cell_40 ( .s (signal_343), .b ({signal_2960, signal_1326}), .a ({signal_2192, signal_313}), .c ({signal_2984, signal_1262}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_42 ( .s (signal_342), .b ({signal_2922, signal_1324}), .a ({signal_2073, signal_315}), .c ({signal_2949, signal_1260}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_44 ( .s (signal_342), .b ({signal_2965, signal_1322}), .a ({signal_2195, signal_317}), .c ({signal_2986, signal_1258}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_46 ( .s (signal_342), .b ({signal_2882, signal_1320}), .a ({signal_2197, signal_1000}), .c ({signal_2918, signal_1256}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_48 ( .s (signal_342), .b ({signal_2932, signal_1318}), .a ({signal_2199, signal_998}), .c ({signal_2951, signal_1254}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_50 ( .s (signal_342), .b ({signal_2885, signal_1316}), .a ({signal_2201, signal_996}), .c ({signal_2919, signal_1252}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_52 ( .s (signal_342), .b ({signal_2935, signal_1314}), .a ({signal_2203, signal_994}), .c ({signal_2952, signal_1250}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_54 ( .s (signal_342), .b ({signal_2936, signal_1312}), .a ({signal_2205, signal_992}), .c ({signal_2953, signal_1248}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_57 ( .s (signal_343), .b ({signal_3041, signal_1309}), .a ({signal_2207, signal_321}), .c ({signal_3059, signal_1245}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_61 ( .s (signal_343), .b ({signal_3045, signal_1305}), .a ({signal_2076, signal_325}), .c ({signal_3060, signal_1241}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_65 ( .s (signal_343), .b ({signal_3010, signal_1301}), .a ({signal_2078, signal_981}), .c ({signal_3022, signal_1237}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_69 ( .s (signal_344), .b ({signal_3014, signal_1297}), .a ({signal_2214, signal_977}), .c ({signal_3024, signal_1233}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_104 ( .s (IN_reset), .b ({signal_2984, signal_1262}), .a ({IN_plaintext_s1[1], IN_plaintext_s0[1]}), .c ({signal_3028, signal_1198}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_106 ( .s (IN_reset), .b ({signal_2949, signal_1260}), .a ({IN_plaintext_s1[3], IN_plaintext_s0[3]}), .c ({signal_2992, signal_1196}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_108 ( .s (IN_reset), .b ({signal_2986, signal_1258}), .a ({IN_plaintext_s1[5], IN_plaintext_s0[5]}), .c ({signal_3032, signal_1194}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_110 ( .s (IN_reset), .b ({signal_2918, signal_1256}), .a ({IN_plaintext_s1[7], IN_plaintext_s0[7]}), .c ({signal_2955, signal_1192}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_112 ( .s (IN_reset), .b ({signal_2951, signal_1254}), .a ({IN_plaintext_s1[9], IN_plaintext_s0[9]}), .c ({signal_2996, signal_1190}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_114 ( .s (IN_reset), .b ({signal_2919, signal_1252}), .a ({IN_plaintext_s1[11], IN_plaintext_s0[11]}), .c ({signal_2957, signal_1188}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_116 ( .s (IN_reset), .b ({signal_2952, signal_1250}), .a ({IN_plaintext_s1[13], IN_plaintext_s0[13]}), .c ({signal_2998, signal_1186}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_118 ( .s (IN_reset), .b ({signal_2953, signal_1248}), .a ({IN_plaintext_s1[15], IN_plaintext_s0[15]}), .c ({signal_3000, signal_1184}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_121 ( .s (IN_reset), .b ({signal_3059, signal_1245}), .a ({IN_plaintext_s1[18], IN_plaintext_s0[18]}), .c ({signal_3112, signal_1181}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_125 ( .s (IN_reset), .b ({signal_3060, signal_1241}), .a ({IN_plaintext_s1[22], IN_plaintext_s0[22]}), .c ({signal_3114, signal_1177}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_129 ( .s (IN_reset), .b ({signal_3022, signal_1237}), .a ({IN_plaintext_s1[26], IN_plaintext_s0[26]}), .c ({signal_3073, signal_1173}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_133 ( .s (IN_reset), .b ({signal_3024, signal_1233}), .a ({IN_plaintext_s1[30], IN_plaintext_s0[30]}), .c ({signal_3077, signal_1169}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_412 ( .a ({signal_2191, signal_1007}), .b ({signal_2641, signal_356}), .c ({signal_2734, signal_940}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_435 ( .a ({signal_2254, signal_1003}), .b ({signal_2642, signal_375}), .c ({signal_2735, signal_936}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_458 ( .a ({signal_2198, signal_999}), .b ({signal_2598, signal_394}), .c ({signal_2633, signal_932}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_481 ( .a ({signal_2202, signal_995}), .b ({signal_2599, signal_413}), .c ({signal_2634, signal_928}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_504 ( .a ({signal_2190, signal_991}), .b ({signal_2643, signal_432}), .c ({signal_2736, signal_924}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_527 ( .a ({signal_2262, signal_987}), .b ({signal_2644, signal_451}), .c ({signal_2737, signal_920}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_550 ( .a ({signal_2077, signal_983}), .b ({signal_2600, signal_470}), .c ({signal_2635, signal_916}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_573 ( .a ({signal_2181, signal_979}), .b ({signal_2601, signal_489}), .c ({signal_2636, signal_912}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_596 ( .a ({signal_2246, signal_975}), .b ({signal_2645, signal_508}), .c ({signal_2738, signal_908}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_619 ( .a ({signal_2243, signal_971}), .b ({signal_2646, signal_527}), .c ({signal_2739, signal_904}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_642 ( .a ({signal_2219, signal_967}), .b ({signal_2602, signal_546}), .c ({signal_2637, signal_900}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_665 ( .a ({signal_2223, signal_963}), .b ({signal_2603, signal_565}), .c ({signal_2638, signal_896}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_688 ( .a ({signal_2256, signal_959}), .b ({signal_2647, signal_584}), .c ({signal_2740, signal_892}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_711 ( .a ({signal_2251, signal_955}), .b ({signal_2648, signal_603}), .c ({signal_2741, signal_888}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_734 ( .a ({signal_2235, signal_951}), .b ({signal_2604, signal_622}), .c ({signal_2639, signal_884}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_757 ( .a ({signal_2239, signal_947}), .b ({signal_2605, signal_641}), .c ({signal_2640, signal_880}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_763 ( .a ({signal_2922, signal_1324}), .b ({signal_2622, signal_882}), .c ({signal_2958, signal_657}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_766 ( .a ({signal_2609, signal_881}), .b ({signal_2879, signal_660}), .c ({signal_2920, signal_658}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_771 ( .a ({signal_2640, signal_880}), .b ({signal_2960, signal_1326}), .c ({signal_3001, signal_665}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_774 ( .a ({signal_2608, signal_901}), .b ({signal_2922, signal_1324}), .c ({signal_2959, signal_668}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_780 ( .a ({signal_2640, signal_880}), .b ({signal_2606, signal_902}), .c ({signal_2742, signal_671}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_782 ( .a ({signal_3002, signal_672}), .b ({signal_2878, signal_673}), .c ({signal_3041, signal_1309}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_783 ( .a ({signal_2816, signal_674}), .b ({signal_2622, signal_882}), .c ({signal_2878, signal_673}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_784 ( .a ({signal_2960, signal_1326}), .b ({signal_2712, signal_923}), .c ({signal_3002, signal_672}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_785 ( .a ({signal_2921, signal_675}), .b ({signal_2743, signal_676}), .c ({signal_2960, signal_1326}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_786 ( .a ({signal_2607, signal_903}), .b ({signal_2637, signal_900}), .c ({signal_2743, signal_676}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_787 ( .a ({signal_2746, signal_677}), .b ({signal_2879, signal_660}), .c ({signal_2921, signal_675}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_788 ( .a ({signal_2815, signal_678}), .b ({signal_2688, signal_941}), .c ({signal_2879, signal_660}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_789 ( .a ({signal_2653, signal_922}), .b ({signal_2734, signal_940}), .c ({signal_2815, signal_678}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_793 ( .a ({signal_2608, signal_901}), .b ({signal_2637, signal_900}), .c ({signal_2744, signal_681}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_796 ( .a ({signal_2922, signal_1324}), .b ({signal_2640, signal_880}), .c ({signal_2961, signal_684}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_799 ( .a ({signal_2609, signal_881}), .b ({signal_2637, signal_900}), .c ({signal_2745, signal_686}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_809 ( .a ({signal_2640, signal_880}), .b ({signal_2610, signal_883}), .c ({signal_2746, signal_677}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_811 ( .a ({signal_2640, signal_880}), .b ({signal_2637, signal_900}), .c ({signal_2747, signal_692}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_813 ( .a ({signal_2880, signal_693}), .b ({signal_2609, signal_881}), .c ({signal_2922, signal_1324}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_814 ( .a ({signal_2816, signal_674}), .b ({signal_2695, signal_942}), .c ({signal_2880, signal_693}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_815 ( .a ({signal_2608, signal_901}), .b ({signal_2737, signal_920}), .c ({signal_2816, signal_674}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_817 ( .a ({signal_2882, signal_1320}), .b ({signal_2671, signal_894}), .c ({signal_2923, signal_695}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_820 ( .a ({signal_2649, signal_893}), .b ({signal_2881, signal_698}), .c ({signal_2924, signal_696}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_825 ( .a ({signal_2740, signal_892}), .b ({signal_2965, signal_1322}), .c ({signal_3006, signal_703}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_828 ( .a ({signal_2612, signal_897}), .b ({signal_2882, signal_1320}), .c ({signal_2925, signal_706}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_834 ( .a ({signal_2740, signal_892}), .b ({signal_2613, signal_898}), .c ({signal_2817, signal_709}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_836 ( .a ({signal_3007, signal_710}), .b ({signal_2818, signal_711}), .c ({signal_3045, signal_1305}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_837 ( .a ({signal_2751, signal_712}), .b ({signal_2671, signal_894}), .c ({signal_2818, signal_711}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_838 ( .a ({signal_2965, signal_1322}), .b ({signal_2632, signal_919}), .c ({signal_3007, signal_710}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_839 ( .a ({signal_2926, signal_713}), .b ({signal_2748, signal_714}), .c ({signal_2965, signal_1322}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_840 ( .a ({signal_2611, signal_899}), .b ({signal_2638, signal_896}), .c ({signal_2748, signal_714}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_841 ( .a ({signal_2820, signal_715}), .b ({signal_2881, signal_698}), .c ({signal_2926, signal_713}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_842 ( .a ({signal_2819, signal_716}), .b ({signal_2696, signal_937}), .c ({signal_2881, signal_698}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_843 ( .a ({signal_2617, signal_918}), .b ({signal_2735, signal_936}), .c ({signal_2819, signal_716}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_847 ( .a ({signal_2612, signal_897}), .b ({signal_2638, signal_896}), .c ({signal_2749, signal_719}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_850 ( .a ({signal_2882, signal_1320}), .b ({signal_2740, signal_892}), .c ({signal_2927, signal_722}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_853 ( .a ({signal_2649, signal_893}), .b ({signal_2638, signal_896}), .c ({signal_2750, signal_724}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_863 ( .a ({signal_2740, signal_892}), .b ({signal_2672, signal_895}), .c ({signal_2820, signal_715}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_865 ( .a ({signal_2740, signal_892}), .b ({signal_2638, signal_896}), .c ({signal_2821, signal_730}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_867 ( .a ({signal_2822, signal_731}), .b ({signal_2649, signal_893}), .c ({signal_2882, signal_1320}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_868 ( .a ({signal_2751, signal_712}), .b ({signal_2673, signal_938}), .c ({signal_2822, signal_731}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_869 ( .a ({signal_2612, signal_897}), .b ({signal_2635, signal_916}), .c ({signal_2751, signal_712}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_871 ( .a ({signal_2885, signal_1316}), .b ({signal_2675, signal_890}), .c ({signal_2930, signal_733}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_874 ( .a ({signal_2677, signal_889}), .b ({signal_2826, signal_736}), .c ({signal_2883, signal_734}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_879 ( .a ({signal_2741, signal_888}), .b ({signal_2932, signal_1318}), .c ({signal_2969, signal_741}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_882 ( .a ({signal_2650, signal_909}), .b ({signal_2885, signal_1316}), .c ({signal_2931, signal_744}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_888 ( .a ({signal_2741, signal_888}), .b ({signal_2674, signal_910}), .c ({signal_2823, signal_747}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_890 ( .a ({signal_2970, signal_748}), .b ({signal_2824, signal_749}), .c ({signal_3010, signal_1301}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_891 ( .a ({signal_2753, signal_750}), .b ({signal_2675, signal_890}), .c ({signal_2824, signal_749}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_892 ( .a ({signal_2932, signal_1318}), .b ({signal_2631, signal_915}), .c ({signal_2970, signal_748}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_893 ( .a ({signal_2884, signal_751}), .b ({signal_2825, signal_752}), .c ({signal_2932, signal_1318}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_894 ( .a ({signal_2676, signal_911}), .b ({signal_2738, signal_908}), .c ({signal_2825, signal_752}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_895 ( .a ({signal_2829, signal_753}), .b ({signal_2826, signal_736}), .c ({signal_2884, signal_751}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_896 ( .a ({signal_2752, signal_754}), .b ({signal_2618, signal_933}), .c ({signal_2826, signal_736}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_897 ( .a ({signal_2615, signal_914}), .b ({signal_2633, signal_932}), .c ({signal_2752, signal_754}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_901 ( .a ({signal_2650, signal_909}), .b ({signal_2738, signal_908}), .c ({signal_2827, signal_757}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_904 ( .a ({signal_2885, signal_1316}), .b ({signal_2741, signal_888}), .c ({signal_2933, signal_760}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_907 ( .a ({signal_2677, signal_889}), .b ({signal_2738, signal_908}), .c ({signal_2828, signal_762}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_917 ( .a ({signal_2741, signal_888}), .b ({signal_2679, signal_891}), .c ({signal_2829, signal_753}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_919 ( .a ({signal_2741, signal_888}), .b ({signal_2738, signal_908}), .c ({signal_2830, signal_768}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_921 ( .a ({signal_2831, signal_769}), .b ({signal_2677, signal_889}), .c ({signal_2885, signal_1316}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_922 ( .a ({signal_2753, signal_750}), .b ({signal_2619, signal_934}), .c ({signal_2831, signal_769}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_923 ( .a ({signal_2650, signal_909}), .b ({signal_2636, signal_912}), .c ({signal_2753, signal_750}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_925 ( .a ({signal_2936, signal_1312}), .b ({signal_2627, signal_886}), .c ({signal_2975, signal_771}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_928 ( .a ({signal_2621, signal_885}), .b ({signal_2833, signal_774}), .c ({signal_2886, signal_772}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_933 ( .a ({signal_2639, signal_884}), .b ({signal_2935, signal_1314}), .c ({signal_2976, signal_779}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_936 ( .a ({signal_2681, signal_905}), .b ({signal_2936, signal_1312}), .c ({signal_2977, signal_782}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_942 ( .a ({signal_2639, signal_884}), .b ({signal_2651, signal_906}), .c ({signal_2754, signal_785}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_944 ( .a ({signal_2978, signal_786}), .b ({signal_2887, signal_787}), .c ({signal_3014, signal_1297}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_945 ( .a ({signal_2837, signal_788}), .b ({signal_2627, signal_886}), .c ({signal_2887, signal_787}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_946 ( .a ({signal_2935, signal_1314}), .b ({signal_2711, signal_927}), .c ({signal_2978, signal_786}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_947 ( .a ({signal_2888, signal_789}), .b ({signal_2832, signal_790}), .c ({signal_2935, signal_1314}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_948 ( .a ({signal_2680, signal_907}), .b ({signal_2739, signal_904}), .c ({signal_2832, signal_790}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_949 ( .a ({signal_2756, signal_791}), .b ({signal_2833, signal_774}), .c ({signal_2888, signal_789}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_950 ( .a ({signal_2755, signal_792}), .b ({signal_2620, signal_929}), .c ({signal_2833, signal_774}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_951 ( .a ({signal_2652, signal_926}), .b ({signal_2634, signal_928}), .c ({signal_2755, signal_792}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_955 ( .a ({signal_2681, signal_905}), .b ({signal_2739, signal_904}), .c ({signal_2834, signal_795}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_958 ( .a ({signal_2936, signal_1312}), .b ({signal_2639, signal_884}), .c ({signal_2979, signal_798}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_961 ( .a ({signal_2621, signal_885}), .b ({signal_2739, signal_904}), .c ({signal_2835, signal_800}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_971 ( .a ({signal_2639, signal_884}), .b ({signal_2616, signal_887}), .c ({signal_2756, signal_791}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_973 ( .a ({signal_2639, signal_884}), .b ({signal_2739, signal_904}), .c ({signal_2836, signal_806}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_975 ( .a ({signal_2889, signal_807}), .b ({signal_2621, signal_885}), .c ({signal_2936, signal_1312}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_976 ( .a ({signal_2837, signal_788}), .b ({signal_2629, signal_930}), .c ({signal_2889, signal_807}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_977 ( .a ({signal_2681, signal_905}), .b ({signal_2736, signal_924}), .c ({signal_2837, signal_788}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1460 ( .s ({signal_2198, signal_999}), .b ({signal_2444, signal_1506}), .a ({signal_2443, signal_1505}), .clk (CLK), .r (Fresh[332]), .c ({signal_2598, signal_394}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1461 ( .s ({signal_2202, signal_995}), .b ({signal_2446, signal_1508}), .a ({signal_2445, signal_1507}), .clk (CLK), .r (Fresh[333]), .c ({signal_2599, signal_413}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1462 ( .s ({signal_2077, signal_983}), .b ({signal_2448, signal_1510}), .a ({signal_2447, signal_1509}), .clk (CLK), .r (Fresh[334]), .c ({signal_2600, signal_470}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1463 ( .s ({signal_2181, signal_979}), .b ({signal_2450, signal_1512}), .a ({signal_2449, signal_1511}), .clk (CLK), .r (Fresh[335]), .c ({signal_2601, signal_489}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1464 ( .s ({signal_2219, signal_967}), .b ({signal_2452, signal_1514}), .a ({signal_2451, signal_1513}), .clk (CLK), .r (Fresh[336]), .c ({signal_2602, signal_546}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1465 ( .s ({signal_2223, signal_963}), .b ({signal_2454, signal_1516}), .a ({signal_2453, signal_1515}), .clk (CLK), .r (Fresh[337]), .c ({signal_2603, signal_565}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1466 ( .s ({signal_2235, signal_951}), .b ({signal_2456, signal_1518}), .a ({signal_2455, signal_1517}), .clk (CLK), .r (Fresh[338]), .c ({signal_2604, signal_622}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1467 ( .s ({signal_2239, signal_947}), .b ({signal_2458, signal_1520}), .a ({signal_2457, signal_1519}), .clk (CLK), .r (Fresh[339]), .c ({signal_2605, signal_641}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1468 ( .s ({signal_2187, signal_1004}), .b ({signal_2500, signal_1522}), .a ({signal_2499, signal_1521}), .clk (CLK), .r (Fresh[340]), .c ({signal_2641, signal_356}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1469 ( .s ({signal_2197, signal_1000}), .b ({signal_2502, signal_1524}), .a ({signal_2501, signal_1523}), .clk (CLK), .r (Fresh[341]), .c ({signal_2642, signal_375}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1470 ( .s ({signal_2189, signal_988}), .b ({signal_2504, signal_1526}), .a ({signal_2503, signal_1525}), .clk (CLK), .r (Fresh[342]), .c ({signal_2643, signal_432}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1471 ( .s ({signal_2188, signal_985}), .b ({signal_2506, signal_1528}), .a ({signal_2505, signal_1527}), .clk (CLK), .r (Fresh[343]), .c ({signal_2644, signal_451}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1472 ( .s ({signal_2244, signal_972}), .b ({signal_2508, signal_1530}), .a ({signal_2507, signal_1529}), .clk (CLK), .r (Fresh[344]), .c ({signal_2645, signal_508}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1473 ( .s ({signal_2186, signal_968}), .b ({signal_2510, signal_1532}), .a ({signal_2509, signal_1531}), .clk (CLK), .r (Fresh[345]), .c ({signal_2646, signal_527}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1474 ( .s ({signal_2252, signal_956}), .b ({signal_2512, signal_1534}), .a ({signal_2511, signal_1533}), .clk (CLK), .r (Fresh[346]), .c ({signal_2647, signal_584}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1475 ( .s ({signal_2234, signal_952}), .b ({signal_2514, signal_1536}), .a ({signal_2513, signal_1535}), .clk (CLK), .r (Fresh[347]), .c ({signal_2648, signal_603}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1476 ( .s ({signal_2219, signal_967}), .b ({signal_2460, signal_1538}), .a ({signal_2459, signal_1537}), .clk (CLK), .r (Fresh[348]), .c ({signal_2606, signal_902}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1477 ( .s ({signal_2219, signal_967}), .b ({signal_2462, signal_1540}), .a ({signal_2461, signal_1539}), .clk (CLK), .r (Fresh[349]), .c ({signal_2607, signal_903}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1478 ( .s ({signal_2219, signal_967}), .b ({signal_2464, signal_1542}), .a ({signal_2463, signal_1541}), .clk (CLK), .r (Fresh[350]), .c ({signal_2608, signal_901}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1479 ( .s ({signal_2239, signal_947}), .b ({signal_2466, signal_1544}), .a ({signal_2465, signal_1543}), .clk (CLK), .r (Fresh[351]), .c ({signal_2609, signal_881}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1480 ( .s ({signal_2239, signal_947}), .b ({signal_2468, signal_1546}), .a ({signal_2467, signal_1545}), .clk (CLK), .r (Fresh[352]), .c ({signal_2610, signal_883}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1481 ( .s ({signal_2223, signal_963}), .b ({signal_2470, signal_1548}), .a ({signal_2469, signal_1547}), .clk (CLK), .r (Fresh[353]), .c ({signal_2611, signal_899}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1482 ( .s ({signal_2223, signal_963}), .b ({signal_2472, signal_1550}), .a ({signal_2471, signal_1549}), .clk (CLK), .r (Fresh[354]), .c ({signal_2612, signal_897}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1483 ( .s ({signal_2252, signal_956}), .b ({signal_2516, signal_1552}), .a ({signal_2515, signal_1551}), .clk (CLK), .r (Fresh[355]), .c ({signal_2649, signal_893}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1484 ( .s ({signal_2223, signal_963}), .b ({signal_2474, signal_1554}), .a ({signal_2473, signal_1553}), .clk (CLK), .r (Fresh[356]), .c ({signal_2613, signal_898}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1485 ( .s ({signal_2223, signal_963}), .b ({signal_2453, signal_1515}), .a ({signal_2454, signal_1516}), .clk (CLK), .r (Fresh[357]), .c ({signal_2614, signal_1660}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1486 ( .s ({signal_2181, signal_979}), .b ({signal_2476, signal_1556}), .a ({signal_2475, signal_1555}), .clk (CLK), .r (Fresh[358]), .c ({signal_2615, signal_914}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1487 ( .s ({signal_2244, signal_972}), .b ({signal_2518, signal_1558}), .a ({signal_2517, signal_1557}), .clk (CLK), .r (Fresh[359]), .c ({signal_2650, signal_909}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1488 ( .s ({signal_2186, signal_968}), .b ({signal_2520, signal_1560}), .a ({signal_2519, signal_1559}), .clk (CLK), .r (Fresh[360]), .c ({signal_2651, signal_906}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1489 ( .s ({signal_2189, signal_988}), .b ({signal_2522, signal_1562}), .a ({signal_2521, signal_1561}), .clk (CLK), .r (Fresh[361]), .c ({signal_2652, signal_926}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1490 ( .s ({signal_2235, signal_951}), .b ({signal_2478, signal_1564}), .a ({signal_2477, signal_1563}), .clk (CLK), .r (Fresh[362]), .c ({signal_2616, signal_887}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1491 ( .s ({signal_2188, signal_985}), .b ({signal_2524, signal_1566}), .a ({signal_2523, signal_1565}), .clk (CLK), .r (Fresh[363]), .c ({signal_2653, signal_922}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1492 ( .s ({signal_2220, signal_966}), .b ({signal_2400, signal_1443}), .a ({signal_2525, signal_1567}), .clk (CLK), .r (Fresh[364]), .c ({signal_2654, signal_1661}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1493 ( .s ({signal_2220, signal_966}), .b ({signal_2527, signal_1569}), .a ({signal_2526, signal_1568}), .clk (CLK), .r (Fresh[365]), .c ({signal_2655, signal_1662}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1494 ( .s ({signal_2221, signal_965}), .b ({signal_2529, signal_1571}), .a ({signal_2528, signal_1570}), .clk (CLK), .r (Fresh[366]), .c ({signal_2656, signal_1663}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1495 ( .s ({signal_2221, signal_965}), .b ({signal_2386, signal_1412}), .a ({signal_2529, signal_1571}), .clk (CLK), .r (Fresh[367]), .c ({signal_2657, signal_1664}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1496 ( .s ({signal_2221, signal_965}), .b ({signal_2528, signal_1570}), .a ({signal_2402, signal_1445}), .clk (CLK), .r (Fresh[368]), .c ({signal_2658, signal_1665}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1497 ( .s ({signal_2221, signal_965}), .b ({signal_2531, signal_1573}), .a ({signal_2530, signal_1572}), .clk (CLK), .r (Fresh[369]), .c ({signal_2659, signal_1666}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1498 ( .s ({signal_2221, signal_965}), .b ({signal_2403, signal_1446}), .a ({signal_2531, signal_1573}), .clk (CLK), .r (Fresh[370]), .c ({signal_2660, signal_1667}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1499 ( .s ({signal_2221, signal_965}), .b ({signal_2530, signal_1572}), .a ({signal_2404, signal_1447}), .clk (CLK), .r (Fresh[371]), .c ({signal_2661, signal_1668}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1500 ( .s ({signal_2221, signal_965}), .b ({signal_2528, signal_1570}), .a ({signal_2529, signal_1571}), .clk (CLK), .r (Fresh[372]), .c ({signal_2662, signal_1669}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1501 ( .s ({signal_2221, signal_965}), .b ({signal_2402, signal_1445}), .a ({signal_2528, signal_1570}), .clk (CLK), .r (Fresh[373]), .c ({signal_2663, signal_1670}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1502 ( .s ({signal_2221, signal_965}), .b ({signal_2529, signal_1571}), .a ({signal_2386, signal_1412}), .clk (CLK), .r (Fresh[374]), .c ({signal_2664, signal_1671}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1503 ( .s ({signal_2210, signal_984}), .b ({signal_2533, signal_1575}), .a ({signal_2532, signal_1574}), .clk (CLK), .r (Fresh[375]), .c ({signal_2665, signal_1672}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1504 ( .s ({signal_2260, signal_1005}), .b ({signal_2533, signal_1575}), .a ({signal_2532, signal_1574}), .clk (CLK), .r (Fresh[376]), .c ({signal_2666, signal_1673}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1505 ( .s ({signal_2260, signal_1005}), .b ({signal_2532, signal_1574}), .a ({signal_2533, signal_1575}), .clk (CLK), .r (Fresh[377]), .c ({signal_2667, signal_1674}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1506 ( .s ({signal_2210, signal_984}), .b ({signal_2536, signal_1578}), .a ({signal_2535, signal_1577}), .clk (CLK), .r (Fresh[378]), .c ({signal_2668, signal_1675}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1507 ( .s ({signal_2210, signal_984}), .b ({signal_2538, signal_1580}), .a ({signal_2537, signal_1579}), .clk (CLK), .r (Fresh[379]), .c ({signal_2669, signal_1676}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1508 ( .s ({signal_2210, signal_984}), .b ({signal_2535, signal_1577}), .a ({signal_2536, signal_1578}), .clk (CLK), .r (Fresh[380]), .c ({signal_2670, signal_1677}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1509 ( .s ({signal_2252, signal_956}), .b ({signal_2541, signal_1583}), .a ({signal_2540, signal_1582}), .clk (CLK), .r (Fresh[381]), .c ({signal_2671, signal_894}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1510 ( .s ({signal_2077, signal_983}), .b ({signal_2480, signal_1585}), .a ({signal_2479, signal_1584}), .clk (CLK), .r (Fresh[382]), .c ({signal_2617, signal_918}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1511 ( .s ({signal_2252, signal_956}), .b ({signal_2543, signal_1587}), .a ({signal_2542, signal_1586}), .clk (CLK), .r (Fresh[383]), .c ({signal_2672, signal_895}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1512 ( .s ({signal_2197, signal_1000}), .b ({signal_2545, signal_1589}), .a ({signal_2544, signal_1588}), .clk (CLK), .r (Fresh[384]), .c ({signal_2673, signal_938}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1513 ( .s ({signal_2244, signal_972}), .b ({signal_2547, signal_1591}), .a ({signal_2546, signal_1590}), .clk (CLK), .r (Fresh[385]), .c ({signal_2674, signal_910}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1514 ( .s ({signal_2234, signal_952}), .b ({signal_2549, signal_1593}), .a ({signal_2548, signal_1592}), .clk (CLK), .r (Fresh[386]), .c ({signal_2675, signal_890}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1515 ( .s ({signal_2244, signal_972}), .b ({signal_2551, signal_1595}), .a ({signal_2550, signal_1594}), .clk (CLK), .r (Fresh[387]), .c ({signal_2676, signal_911}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1516 ( .s ({signal_2198, signal_999}), .b ({signal_2482, signal_1597}), .a ({signal_2481, signal_1596}), .clk (CLK), .r (Fresh[388]), .c ({signal_2618, signal_933}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1517 ( .s ({signal_2234, signal_952}), .b ({signal_2553, signal_1599}), .a ({signal_2552, signal_1598}), .clk (CLK), .r (Fresh[389]), .c ({signal_2677, signal_889}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1518 ( .s ({signal_2244, signal_972}), .b ({signal_2555, signal_1601}), .a ({signal_2554, signal_1600}), .clk (CLK), .r (Fresh[390]), .c ({signal_2678, signal_1678}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1519 ( .s ({signal_2234, signal_952}), .b ({signal_2557, signal_1603}), .a ({signal_2556, signal_1602}), .clk (CLK), .r (Fresh[391]), .c ({signal_2679, signal_891}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1520 ( .s ({signal_2198, signal_999}), .b ({signal_2484, signal_1605}), .a ({signal_2483, signal_1604}), .clk (CLK), .r (Fresh[392]), .c ({signal_2619, signal_934}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1521 ( .s ({signal_2186, signal_968}), .b ({signal_2559, signal_1607}), .a ({signal_2558, signal_1606}), .clk (CLK), .r (Fresh[393]), .c ({signal_2680, signal_907}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1522 ( .s ({signal_2202, signal_995}), .b ({signal_2486, signal_1609}), .a ({signal_2485, signal_1608}), .clk (CLK), .r (Fresh[394]), .c ({signal_2620, signal_929}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1523 ( .s ({signal_2186, signal_968}), .b ({signal_2561, signal_1611}), .a ({signal_2560, signal_1610}), .clk (CLK), .r (Fresh[395]), .c ({signal_2681, signal_905}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1524 ( .s ({signal_2235, signal_951}), .b ({signal_2488, signal_1613}), .a ({signal_2487, signal_1612}), .clk (CLK), .r (Fresh[396]), .c ({signal_2621, signal_885}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1525 ( .s ({signal_2243, signal_971}), .b ({signal_2420, signal_1476}), .a ({signal_2562, signal_1614}), .clk (CLK), .r (Fresh[397]), .c ({signal_2682, signal_1679}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1526 ( .s ({signal_2257, signal_969}), .b ({signal_2563, signal_1615}), .a ({signal_2421, signal_1477}), .clk (CLK), .r (Fresh[398]), .c ({signal_2683, signal_1680}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1527 ( .s ({signal_2257, signal_969}), .b ({signal_2565, signal_1617}), .a ({signal_2422, signal_1478}), .clk (CLK), .r (Fresh[399]), .c ({signal_2684, signal_1681}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1528 ( .s ({signal_2243, signal_971}), .b ({signal_2424, signal_1480}), .a ({signal_2567, signal_1619}), .clk (CLK), .r (Fresh[400]), .c ({signal_2685, signal_1682}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1529 ( .s ({signal_2243, signal_971}), .b ({signal_2425, signal_1481}), .a ({signal_2568, signal_1620}), .clk (CLK), .r (Fresh[401]), .c ({signal_2686, signal_1683}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1530 ( .s ({signal_2243, signal_971}), .b ({signal_2426, signal_1482}), .a ({signal_2569, signal_1621}), .clk (CLK), .r (Fresh[402]), .c ({signal_2687, signal_1684}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1531 ( .s ({signal_2239, signal_947}), .b ({signal_2490, signal_1623}), .a ({signal_2489, signal_1622}), .clk (CLK), .r (Fresh[403]), .c ({signal_2622, signal_882}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1532 ( .s ({signal_2187, signal_1004}), .b ({signal_2571, signal_1625}), .a ({signal_2570, signal_1624}), .clk (CLK), .r (Fresh[404]), .c ({signal_2688, signal_941}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1533 ( .s ({signal_2241, signal_945}), .b ({signal_2573, signal_1627}), .a ({signal_2572, signal_1626}), .clk (CLK), .r (Fresh[405]), .c ({signal_2689, signal_1685}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1534 ( .s ({signal_2241, signal_945}), .b ({signal_2429, signal_1487}), .a ({signal_2573, signal_1627}), .clk (CLK), .r (Fresh[406]), .c ({signal_2690, signal_1686}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1535 ( .s ({signal_2241, signal_945}), .b ({signal_2572, signal_1626}), .a ({signal_2430, signal_1488}), .clk (CLK), .r (Fresh[407]), .c ({signal_2691, signal_1687}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1536 ( .s ({signal_2241, signal_945}), .b ({signal_2572, signal_1626}), .a ({signal_2573, signal_1627}), .clk (CLK), .r (Fresh[408]), .c ({signal_2692, signal_1688}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1537 ( .s ({signal_2241, signal_945}), .b ({signal_2430, signal_1488}), .a ({signal_2572, signal_1626}), .clk (CLK), .r (Fresh[409]), .c ({signal_2693, signal_1689}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1538 ( .s ({signal_2241, signal_945}), .b ({signal_2573, signal_1627}), .a ({signal_2429, signal_1487}), .clk (CLK), .r (Fresh[410]), .c ({signal_2694, signal_1690}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1539 ( .s ({signal_2187, signal_1004}), .b ({signal_2575, signal_1629}), .a ({signal_2574, signal_1628}), .clk (CLK), .r (Fresh[411]), .c ({signal_2695, signal_942}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1540 ( .s ({signal_2197, signal_1000}), .b ({signal_2577, signal_1631}), .a ({signal_2576, signal_1630}), .clk (CLK), .r (Fresh[412]), .c ({signal_2696, signal_937}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1541 ( .s ({signal_2253, signal_957}), .b ({signal_2578, signal_1632}), .a ({signal_2433, signal_1491}), .clk (CLK), .r (Fresh[413]), .c ({signal_2697, signal_1691}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1542 ( .s ({signal_2253, signal_957}), .b ({signal_2435, signal_1493}), .a ({signal_2579, signal_1633}), .clk (CLK), .r (Fresh[414]), .c ({signal_2698, signal_1692}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1543 ( .s ({signal_2253, signal_957}), .b ({signal_2580, signal_1634}), .a ({signal_2436, signal_1494}), .clk (CLK), .r (Fresh[415]), .c ({signal_2699, signal_1693}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1544 ( .s ({signal_2253, signal_957}), .b ({signal_2437, signal_1495}), .a ({signal_2581, signal_1635}), .clk (CLK), .r (Fresh[416]), .c ({signal_2700, signal_1694}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1545 ( .s ({signal_2212, signal_980}), .b ({signal_2582, signal_1636}), .a ({signal_2576, signal_1630}), .clk (CLK), .r (Fresh[417]), .c ({signal_2701, signal_1695}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1546 ( .s ({signal_2212, signal_980}), .b ({signal_2576, signal_1630}), .a ({signal_2582, signal_1636}), .clk (CLK), .r (Fresh[418]), .c ({signal_2702, signal_1696}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1547 ( .s ({signal_2212, signal_980}), .b ({signal_2583, signal_1637}), .a ({signal_2577, signal_1631}), .clk (CLK), .r (Fresh[419]), .c ({signal_2703, signal_1697}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1548 ( .s ({signal_2212, signal_980}), .b ({signal_2577, signal_1631}), .a ({signal_2583, signal_1637}), .clk (CLK), .r (Fresh[420]), .c ({signal_2704, signal_1698}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1549 ( .s ({signal_2234, signal_952}), .b ({signal_2585, signal_1639}), .a ({signal_2584, signal_1638}), .clk (CLK), .r (Fresh[421]), .c ({signal_2705, signal_1699}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1550 ( .s ({signal_2201, signal_996}), .b ({signal_2492, signal_1641}), .a ({signal_2491, signal_1640}), .clk (CLK), .r (Fresh[422]), .c ({signal_2623, signal_1700}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1551 ( .s ({signal_2201, signal_996}), .b ({signal_2491, signal_1640}), .a ({signal_2492, signal_1641}), .clk (CLK), .r (Fresh[423]), .c ({signal_2624, signal_1701}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1552 ( .s ({signal_2200, signal_997}), .b ({signal_2492, signal_1641}), .a ({signal_2491, signal_1640}), .clk (CLK), .r (Fresh[424]), .c ({signal_2625, signal_1702}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1553 ( .s ({signal_2200, signal_997}), .b ({signal_2491, signal_1640}), .a ({signal_2492, signal_1641}), .clk (CLK), .r (Fresh[425]), .c ({signal_2626, signal_1703}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1554 ( .s ({signal_2235, signal_951}), .b ({signal_2494, signal_1643}), .a ({signal_2493, signal_1642}), .clk (CLK), .r (Fresh[426]), .c ({signal_2627, signal_886}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1555 ( .s ({signal_2235, signal_951}), .b ({signal_2455, signal_1517}), .a ({signal_2456, signal_1518}), .clk (CLK), .r (Fresh[427]), .c ({signal_2628, signal_1704}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1556 ( .s ({signal_2204, signal_993}), .b ({signal_2440, signal_1500}), .a ({signal_2586, signal_1644}), .clk (CLK), .r (Fresh[428]), .c ({signal_2706, signal_1705}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1557 ( .s ({signal_2204, signal_993}), .b ({signal_2441, signal_1501}), .a ({signal_2587, signal_1645}), .clk (CLK), .r (Fresh[429]), .c ({signal_2707, signal_1706}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1558 ( .s ({signal_2204, signal_993}), .b ({signal_2586, signal_1644}), .a ({signal_2587, signal_1645}), .clk (CLK), .r (Fresh[430]), .c ({signal_2708, signal_1707}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1559 ( .s ({signal_2204, signal_993}), .b ({signal_2587, signal_1645}), .a ({signal_2586, signal_1644}), .clk (CLK), .r (Fresh[431]), .c ({signal_2709, signal_1708}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1560 ( .s ({signal_2202, signal_995}), .b ({signal_2496, signal_1649}), .a ({signal_2495, signal_1648}), .clk (CLK), .r (Fresh[432]), .c ({signal_2629, signal_930}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1561 ( .s ({signal_2223, signal_963}), .b ({signal_2469, signal_1547}), .a ({signal_2470, signal_1548}), .clk (CLK), .r (Fresh[433]), .c ({signal_2630, signal_1709}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1562 ( .s ({signal_2181, signal_979}), .b ({signal_2492, signal_1641}), .a ({signal_2491, signal_1640}), .clk (CLK), .r (Fresh[434]), .c ({signal_2631, signal_915}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1563 ( .s ({signal_2244, signal_972}), .b ({signal_2550, signal_1594}), .a ({signal_2551, signal_1595}), .clk (CLK), .r (Fresh[435]), .c ({signal_2710, signal_1710}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1564 ( .s ({signal_2189, signal_988}), .b ({signal_2591, signal_1651}), .a ({signal_2590, signal_1650}), .clk (CLK), .r (Fresh[436]), .c ({signal_2711, signal_927}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1565 ( .s ({signal_2188, signal_985}), .b ({signal_2442, signal_1504}), .a ({signal_2592, signal_1652}), .clk (CLK), .r (Fresh[437]), .c ({signal_2712, signal_923}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1566 ( .s ({signal_2220, signal_966}), .b ({signal_2525, signal_1567}), .a ({signal_2401, signal_1444}), .clk (CLK), .r (Fresh[438]), .c ({signal_2713, signal_1711}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1567 ( .s ({signal_2220, signal_966}), .b ({signal_2593, signal_1653}), .a ({signal_2400, signal_1443}), .clk (CLK), .r (Fresh[439]), .c ({signal_2714, signal_1712}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1568 ( .s ({signal_2221, signal_965}), .b ({signal_2530, signal_1572}), .a ({signal_2531, signal_1573}), .clk (CLK), .r (Fresh[440]), .c ({signal_2715, signal_1713}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1569 ( .s ({signal_2077, signal_983}), .b ({signal_2498, signal_1655}), .a ({signal_2497, signal_1654}), .clk (CLK), .r (Fresh[441]), .c ({signal_2632, signal_919}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1570 ( .s ({signal_2243, signal_971}), .b ({signal_2595, signal_1657}), .a ({signal_2594, signal_1656}), .clk (CLK), .r (Fresh[442]), .c ({signal_2716, signal_1714}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1571 ( .s ({signal_2257, signal_969}), .b ({signal_2422, signal_1478}), .a ({signal_2563, signal_1615}), .clk (CLK), .r (Fresh[443]), .c ({signal_2717, signal_1715}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1572 ( .s ({signal_2257, signal_969}), .b ({signal_2421, signal_1477}), .a ({signal_2565, signal_1617}), .clk (CLK), .r (Fresh[444]), .c ({signal_2718, signal_1716}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1573 ( .s ({signal_2243, signal_971}), .b ({signal_2597, signal_1659}), .a ({signal_2596, signal_1658}), .clk (CLK), .r (Fresh[445]), .c ({signal_2719, signal_1717}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1574 ( .s ({signal_2243, signal_971}), .b ({signal_2594, signal_1656}), .a ({signal_2595, signal_1657}), .clk (CLK), .r (Fresh[446]), .c ({signal_2720, signal_1718}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1575 ( .s ({signal_2243, signal_971}), .b ({signal_2596, signal_1658}), .a ({signal_2597, signal_1659}), .clk (CLK), .r (Fresh[447]), .c ({signal_2721, signal_1719}) ) ;

    /* cells in depth 9 */

    /* cells in depth 10 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1576 ( .s ({signal_2212, signal_980}), .b ({signal_2614, signal_1660}), .a ({signal_2613, signal_898}), .clk (CLK), .r (Fresh[448]), .c ({signal_2722, signal_1720}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1577 ( .s ({signal_2212, signal_980}), .b ({signal_2613, signal_898}), .a ({signal_2614, signal_1660}), .clk (CLK), .r (Fresh[449]), .c ({signal_2723, signal_1721}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1578 ( .s ({signal_2211, signal_982}), .b ({signal_2614, signal_1660}), .a ({signal_2613, signal_898}), .clk (CLK), .r (Fresh[450]), .c ({signal_2724, signal_1722}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1579 ( .s ({signal_2219, signal_967}), .b ({signal_2655, signal_1662}), .a ({signal_2654, signal_1661}), .clk (CLK), .r (Fresh[451]), .c ({signal_2757, signal_1723}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1580 ( .s ({signal_2220, signal_966}), .b ({signal_2528, signal_1570}), .a ({signal_2656, signal_1663}), .clk (CLK), .r (Fresh[452]), .c ({signal_2758, signal_1724}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1581 ( .s ({signal_2220, signal_966}), .b ({signal_2658, signal_1665}), .a ({signal_2657, signal_1664}), .clk (CLK), .r (Fresh[453]), .c ({signal_2759, signal_1725}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1582 ( .s ({signal_2220, signal_966}), .b ({signal_2530, signal_1572}), .a ({signal_2659, signal_1666}), .clk (CLK), .r (Fresh[454]), .c ({signal_2760, signal_1726}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1583 ( .s ({signal_2220, signal_966}), .b ({signal_2661, signal_1668}), .a ({signal_2660, signal_1667}), .clk (CLK), .r (Fresh[455]), .c ({signal_2761, signal_1727}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1584 ( .s ({signal_2220, signal_966}), .b ({signal_2529, signal_1571}), .a ({signal_2662, signal_1669}), .clk (CLK), .r (Fresh[456]), .c ({signal_2762, signal_1728}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1585 ( .s ({signal_2220, signal_966}), .b ({signal_2664, signal_1671}), .a ({signal_2663, signal_1670}), .clk (CLK), .r (Fresh[457]), .c ({signal_2763, signal_1729}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1586 ( .s ({signal_2210, signal_984}), .b ({signal_2667, signal_1674}), .a ({signal_2666, signal_1673}), .clk (CLK), .r (Fresh[458]), .c ({signal_2764, signal_1730}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1587 ( .s ({signal_2191, signal_1007}), .b ({signal_2668, signal_1675}), .a ({signal_2534, signal_1576}), .clk (CLK), .r (Fresh[459]), .c ({signal_2765, signal_1731}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1588 ( .s ({signal_2210, signal_984}), .b ({signal_2666, signal_1673}), .a ({signal_2667, signal_1674}), .clk (CLK), .r (Fresh[460]), .c ({signal_2766, signal_1732}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1589 ( .s ({signal_2191, signal_1007}), .b ({signal_2539, signal_1581}), .a ({signal_2670, signal_1677}), .clk (CLK), .r (Fresh[461]), .c ({signal_2767, signal_1733}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1590 ( .s ({signal_2215, signal_976}), .b ({signal_2678, signal_1678}), .a ({signal_2674, signal_910}), .clk (CLK), .r (Fresh[462]), .c ({signal_2768, signal_1734}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1591 ( .s ({signal_2215, signal_976}), .b ({signal_2674, signal_910}), .a ({signal_2678, signal_1678}), .clk (CLK), .r (Fresh[463]), .c ({signal_2769, signal_1735}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1592 ( .s ({signal_2214, signal_977}), .b ({signal_2678, signal_1678}), .a ({signal_2674, signal_910}), .clk (CLK), .r (Fresh[464]), .c ({signal_2770, signal_1736}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1593 ( .s ({signal_2243, signal_971}), .b ({signal_2564, signal_1616}), .a ({signal_2683, signal_1680}), .clk (CLK), .r (Fresh[465]), .c ({signal_2771, signal_1737}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1594 ( .s ({signal_2243, signal_971}), .b ({signal_2566, signal_1618}), .a ({signal_2684, signal_1681}), .clk (CLK), .r (Fresh[466]), .c ({signal_2772, signal_1738}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1595 ( .s ({signal_2243, signal_971}), .b ({signal_2565, signal_1617}), .a ({signal_2684, signal_1681}), .clk (CLK), .r (Fresh[467]), .c ({signal_2773, signal_1739}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1596 ( .s ({signal_2243, signal_971}), .b ({signal_2563, signal_1615}), .a ({signal_2683, signal_1680}), .clk (CLK), .r (Fresh[468]), .c ({signal_2774, signal_1740}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1597 ( .s ({signal_2240, signal_946}), .b ({signal_2572, signal_1626}), .a ({signal_2689, signal_1685}), .clk (CLK), .r (Fresh[469]), .c ({signal_2775, signal_1741}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1598 ( .s ({signal_2240, signal_946}), .b ({signal_2691, signal_1687}), .a ({signal_2690, signal_1686}), .clk (CLK), .r (Fresh[470]), .c ({signal_2776, signal_1742}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1599 ( .s ({signal_2240, signal_946}), .b ({signal_2573, signal_1627}), .a ({signal_2692, signal_1688}), .clk (CLK), .r (Fresh[471]), .c ({signal_2777, signal_1743}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1600 ( .s ({signal_2240, signal_946}), .b ({signal_2694, signal_1690}), .a ({signal_2693, signal_1689}), .clk (CLK), .r (Fresh[472]), .c ({signal_2778, signal_1744}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1601 ( .s ({signal_2252, signal_956}), .b ({signal_2698, signal_1692}), .a ({signal_2697, signal_1691}), .clk (CLK), .r (Fresh[473]), .c ({signal_2779, signal_1745}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1602 ( .s ({signal_2252, signal_956}), .b ({signal_2700, signal_1694}), .a ({signal_2699, signal_1693}), .clk (CLK), .r (Fresh[474]), .c ({signal_2780, signal_1746}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1603 ( .s ({signal_2211, signal_982}), .b ({signal_2702, signal_1696}), .a ({signal_2701, signal_1695}), .clk (CLK), .r (Fresh[475]), .c ({signal_2781, signal_1747}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1604 ( .s ({signal_2211, signal_982}), .b ({signal_2704, signal_1698}), .a ({signal_2703, signal_1697}), .clk (CLK), .r (Fresh[476]), .c ({signal_2782, signal_1748}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1605 ( .s ({signal_2197, signal_1000}), .b ({signal_2703, signal_1697}), .a ({signal_2701, signal_1695}), .clk (CLK), .r (Fresh[477]), .c ({signal_2783, signal_1749}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1606 ( .s ({signal_2211, signal_982}), .b ({signal_2701, signal_1695}), .a ({signal_2702, signal_1696}), .clk (CLK), .r (Fresh[478]), .c ({signal_2784, signal_1750}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1607 ( .s ({signal_2211, signal_982}), .b ({signal_2703, signal_1697}), .a ({signal_2704, signal_1698}), .clk (CLK), .r (Fresh[479]), .c ({signal_2785, signal_1751}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1608 ( .s ({signal_2197, signal_1000}), .b ({signal_2704, signal_1698}), .a ({signal_2702, signal_1696}), .clk (CLK), .r (Fresh[480]), .c ({signal_2786, signal_1752}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1609 ( .s ({signal_2201, signal_996}), .b ({signal_2705, signal_1699}), .a ({signal_2675, signal_890}), .clk (CLK), .r (Fresh[481]), .c ({signal_2787, signal_1753}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1610 ( .s ({signal_2201, signal_996}), .b ({signal_2675, signal_890}), .a ({signal_2705, signal_1699}), .clk (CLK), .r (Fresh[482]), .c ({signal_2788, signal_1754}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1611 ( .s ({signal_2200, signal_997}), .b ({signal_2491, signal_1640}), .a ({signal_2623, signal_1700}), .clk (CLK), .r (Fresh[483]), .c ({signal_2725, signal_1755}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1612 ( .s ({signal_2200, signal_997}), .b ({signal_2492, signal_1641}), .a ({signal_2624, signal_1701}), .clk (CLK), .r (Fresh[484]), .c ({signal_2726, signal_1756}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1613 ( .s ({signal_2200, signal_997}), .b ({signal_2623, signal_1700}), .a ({signal_2624, signal_1701}), .clk (CLK), .r (Fresh[485]), .c ({signal_2727, signal_1757}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1614 ( .s ({signal_2200, signal_997}), .b ({signal_2624, signal_1701}), .a ({signal_2623, signal_1700}), .clk (CLK), .r (Fresh[486]), .c ({signal_2728, signal_1758}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1615 ( .s ({signal_2205, signal_992}), .b ({signal_2628, signal_1704}), .a ({signal_2627, signal_886}), .clk (CLK), .r (Fresh[487]), .c ({signal_2729, signal_1759}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1616 ( .s ({signal_2205, signal_992}), .b ({signal_2627, signal_886}), .a ({signal_2628, signal_1704}), .clk (CLK), .r (Fresh[488]), .c ({signal_2730, signal_1760}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1617 ( .s ({signal_2203, signal_994}), .b ({signal_2707, signal_1706}), .a ({signal_2706, signal_1705}), .clk (CLK), .r (Fresh[489]), .c ({signal_2789, signal_1761}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1618 ( .s ({signal_2203, signal_994}), .b ({signal_2708, signal_1707}), .a ({signal_2588, signal_1646}), .clk (CLK), .r (Fresh[490]), .c ({signal_2790, signal_1762}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1619 ( .s ({signal_2203, signal_994}), .b ({signal_2706, signal_1705}), .a ({signal_2707, signal_1706}), .clk (CLK), .r (Fresh[491]), .c ({signal_2791, signal_1763}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1620 ( .s ({signal_2203, signal_994}), .b ({signal_2709, signal_1708}), .a ({signal_2589, signal_1647}), .clk (CLK), .r (Fresh[492]), .c ({signal_2792, signal_1764}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1621 ( .s ({signal_2212, signal_980}), .b ({signal_2630, signal_1709}), .a ({signal_2611, signal_899}), .clk (CLK), .r (Fresh[493]), .c ({signal_2731, signal_1765}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1622 ( .s ({signal_2212, signal_980}), .b ({signal_2611, signal_899}), .a ({signal_2630, signal_1709}), .clk (CLK), .r (Fresh[494]), .c ({signal_2732, signal_1766}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1623 ( .s ({signal_2211, signal_982}), .b ({signal_2630, signal_1709}), .a ({signal_2611, signal_899}), .clk (CLK), .r (Fresh[495]), .c ({signal_2733, signal_1767}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1624 ( .s ({signal_2215, signal_976}), .b ({signal_2710, signal_1710}), .a ({signal_2676, signal_911}), .clk (CLK), .r (Fresh[496]), .c ({signal_2793, signal_1768}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1625 ( .s ({signal_2215, signal_976}), .b ({signal_2676, signal_911}), .a ({signal_2710, signal_1710}), .clk (CLK), .r (Fresh[497]), .c ({signal_2794, signal_1769}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1626 ( .s ({signal_2214, signal_977}), .b ({signal_2710, signal_1710}), .a ({signal_2676, signal_911}), .clk (CLK), .r (Fresh[498]), .c ({signal_2795, signal_1770}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1627 ( .s ({signal_2219, signal_967}), .b ({signal_2714, signal_1712}), .a ({signal_2713, signal_1711}), .clk (CLK), .r (Fresh[499]), .c ({signal_2796, signal_1771}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1628 ( .s ({signal_2220, signal_966}), .b ({signal_2656, signal_1663}), .a ({signal_2529, signal_1571}), .clk (CLK), .r (Fresh[500]), .c ({signal_2797, signal_1772}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1629 ( .s ({signal_2220, signal_966}), .b ({signal_2662, signal_1669}), .a ({signal_2528, signal_1570}), .clk (CLK), .r (Fresh[501]), .c ({signal_2798, signal_1773}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1630 ( .s ({signal_2220, signal_966}), .b ({signal_2659, signal_1666}), .a ({signal_2531, signal_1573}), .clk (CLK), .r (Fresh[502]), .c ({signal_2799, signal_1774}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1631 ( .s ({signal_2220, signal_966}), .b ({signal_2715, signal_1713}), .a ({signal_2530, signal_1572}), .clk (CLK), .r (Fresh[503]), .c ({signal_2800, signal_1775}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1632 ( .s ({signal_2243, signal_971}), .b ({signal_2718, signal_1716}), .a ({signal_2717, signal_1715}), .clk (CLK), .r (Fresh[504]), .c ({signal_2801, signal_1776}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1633 ( .s ({signal_2243, signal_971}), .b ({signal_2717, signal_1715}), .a ({signal_2718, signal_1716}), .clk (CLK), .r (Fresh[505]), .c ({signal_2802, signal_1777}) ) ;

    /* cells in depth 11 */

    /* cells in depth 12 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1634 ( .s ({signal_2211, signal_982}), .b ({signal_2723, signal_1721}), .a ({signal_2722, signal_1720}), .clk (CLK), .r (Fresh[506]), .c ({signal_2803, signal_1778}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1635 ( .s ({signal_2211, signal_982}), .b ({signal_2723, signal_1721}), .a ({signal_2613, signal_898}), .clk (CLK), .r (Fresh[507]), .c ({signal_2804, signal_1779}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1636 ( .s ({signal_2211, signal_982}), .b ({signal_2722, signal_1720}), .a ({signal_2614, signal_1660}), .clk (CLK), .r (Fresh[508]), .c ({signal_2805, signal_1780}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1637 ( .s ({signal_2219, signal_967}), .b ({signal_2759, signal_1725}), .a ({signal_2758, signal_1724}), .clk (CLK), .r (Fresh[509]), .c ({signal_2838, signal_1781}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1638 ( .s ({signal_2219, signal_967}), .b ({signal_2761, signal_1727}), .a ({signal_2760, signal_1726}), .clk (CLK), .r (Fresh[510]), .c ({signal_2839, signal_1782}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1639 ( .s ({signal_2219, signal_967}), .b ({signal_2763, signal_1729}), .a ({signal_2762, signal_1728}), .clk (CLK), .r (Fresh[511]), .c ({signal_2840, signal_1783}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1640 ( .s ({signal_2191, signal_1007}), .b ({signal_2764, signal_1730}), .a ({signal_2665, signal_1672}), .clk (CLK), .r (Fresh[512]), .c ({signal_2841, signal_1784}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1641 ( .s ({signal_2191, signal_1007}), .b ({signal_2669, signal_1676}), .a ({signal_2766, signal_1732}), .clk (CLK), .r (Fresh[513]), .c ({signal_2842, signal_1785}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1642 ( .s ({signal_2214, signal_977}), .b ({signal_2674, signal_910}), .a ({signal_2768, signal_1734}), .clk (CLK), .r (Fresh[514]), .c ({signal_2843, signal_1786}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1643 ( .s ({signal_2214, signal_977}), .b ({signal_2678, signal_1678}), .a ({signal_2769, signal_1735}), .clk (CLK), .r (Fresh[515]), .c ({signal_2844, signal_1787}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1644 ( .s ({signal_2214, signal_977}), .b ({signal_2768, signal_1734}), .a ({signal_2769, signal_1735}), .clk (CLK), .r (Fresh[516]), .c ({signal_2845, signal_1788}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1645 ( .s ({signal_2190, signal_991}), .b ({signal_2771, signal_1737}), .a ({signal_2682, signal_1679}), .clk (CLK), .r (Fresh[517]), .c ({signal_2846, signal_1789}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1646 ( .s ({signal_2190, signal_991}), .b ({signal_2685, signal_1682}), .a ({signal_2772, signal_1738}), .clk (CLK), .r (Fresh[518]), .c ({signal_2847, signal_1790}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1647 ( .s ({signal_2190, signal_991}), .b ({signal_2773, signal_1739}), .a ({signal_2686, signal_1683}), .clk (CLK), .r (Fresh[519]), .c ({signal_2848, signal_1791}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1648 ( .s ({signal_2190, signal_991}), .b ({signal_2687, signal_1684}), .a ({signal_2774, signal_1740}), .clk (CLK), .r (Fresh[520]), .c ({signal_2849, signal_1792}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1649 ( .s ({signal_2239, signal_947}), .b ({signal_2776, signal_1742}), .a ({signal_2775, signal_1741}), .clk (CLK), .r (Fresh[521]), .c ({signal_2850, signal_1793}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1650 ( .s ({signal_2239, signal_947}), .b ({signal_2778, signal_1744}), .a ({signal_2777, signal_1743}), .clk (CLK), .r (Fresh[522]), .c ({signal_2851, signal_1794}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1651 ( .s ({signal_2248, signal_1002}), .b ({signal_2780, signal_1746}), .a ({signal_2779, signal_1745}), .clk (CLK), .r (Fresh[523]), .c ({signal_2852, signal_1795}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1652 ( .s ({signal_2248, signal_1002}), .b ({signal_2779, signal_1745}), .a ({signal_2780, signal_1746}), .clk (CLK), .r (Fresh[524]), .c ({signal_2853, signal_1796}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1653 ( .s ({signal_2197, signal_1000}), .b ({signal_2782, signal_1748}), .a ({signal_2781, signal_1747}), .clk (CLK), .r (Fresh[525]), .c ({signal_2854, signal_1797}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1654 ( .s ({signal_2197, signal_1000}), .b ({signal_2785, signal_1751}), .a ({signal_2784, signal_1750}), .clk (CLK), .r (Fresh[526]), .c ({signal_2855, signal_1798}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1655 ( .s ({signal_2200, signal_997}), .b ({signal_2787, signal_1753}), .a ({signal_2788, signal_1754}), .clk (CLK), .r (Fresh[527]), .c ({signal_2856, signal_1799}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1656 ( .s ({signal_2200, signal_997}), .b ({signal_2788, signal_1754}), .a ({signal_2787, signal_1753}), .clk (CLK), .r (Fresh[528]), .c ({signal_2857, signal_1800}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1657 ( .s ({signal_2199, signal_998}), .b ({signal_2726, signal_1756}), .a ({signal_2725, signal_1755}), .clk (CLK), .r (Fresh[529]), .c ({signal_2806, signal_1801}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1658 ( .s ({signal_2199, signal_998}), .b ({signal_2727, signal_1757}), .a ({signal_2625, signal_1702}), .clk (CLK), .r (Fresh[530]), .c ({signal_2807, signal_1802}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1659 ( .s ({signal_2199, signal_998}), .b ({signal_2725, signal_1755}), .a ({signal_2726, signal_1756}), .clk (CLK), .r (Fresh[531]), .c ({signal_2808, signal_1803}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1660 ( .s ({signal_2199, signal_998}), .b ({signal_2728, signal_1758}), .a ({signal_2626, signal_1703}), .clk (CLK), .r (Fresh[532]), .c ({signal_2809, signal_1804}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1661 ( .s ({signal_2204, signal_993}), .b ({signal_2729, signal_1759}), .a ({signal_2730, signal_1760}), .clk (CLK), .r (Fresh[533]), .c ({signal_2810, signal_1805}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1662 ( .s ({signal_2204, signal_993}), .b ({signal_2730, signal_1760}), .a ({signal_2729, signal_1759}), .clk (CLK), .r (Fresh[534]), .c ({signal_2811, signal_1806}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1663 ( .s ({signal_2202, signal_995}), .b ({signal_2790, signal_1762}), .a ({signal_2789, signal_1761}), .clk (CLK), .r (Fresh[535]), .c ({signal_2858, signal_1807}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1664 ( .s ({signal_2202, signal_995}), .b ({signal_2792, signal_1764}), .a ({signal_2791, signal_1763}), .clk (CLK), .r (Fresh[536]), .c ({signal_2859, signal_1808}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1665 ( .s ({signal_2211, signal_982}), .b ({signal_2732, signal_1766}), .a ({signal_2731, signal_1765}), .clk (CLK), .r (Fresh[537]), .c ({signal_2812, signal_1809}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1666 ( .s ({signal_2211, signal_982}), .b ({signal_2732, signal_1766}), .a ({signal_2611, signal_899}), .clk (CLK), .r (Fresh[538]), .c ({signal_2813, signal_1810}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1667 ( .s ({signal_2211, signal_982}), .b ({signal_2731, signal_1765}), .a ({signal_2630, signal_1709}), .clk (CLK), .r (Fresh[539]), .c ({signal_2814, signal_1811}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1668 ( .s ({signal_2214, signal_977}), .b ({signal_2676, signal_911}), .a ({signal_2793, signal_1768}), .clk (CLK), .r (Fresh[540]), .c ({signal_2860, signal_1812}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1669 ( .s ({signal_2214, signal_977}), .b ({signal_2710, signal_1710}), .a ({signal_2794, signal_1769}), .clk (CLK), .r (Fresh[541]), .c ({signal_2861, signal_1813}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1670 ( .s ({signal_2214, signal_977}), .b ({signal_2793, signal_1768}), .a ({signal_2794, signal_1769}), .clk (CLK), .r (Fresh[542]), .c ({signal_2862, signal_1814}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1671 ( .s ({signal_2219, signal_967}), .b ({signal_2798, signal_1773}), .a ({signal_2797, signal_1772}), .clk (CLK), .r (Fresh[543]), .c ({signal_2863, signal_1815}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1672 ( .s ({signal_2219, signal_967}), .b ({signal_2800, signal_1775}), .a ({signal_2799, signal_1774}), .clk (CLK), .r (Fresh[544]), .c ({signal_2864, signal_1816}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1673 ( .s ({signal_2219, signal_967}), .b ({signal_2797, signal_1772}), .a ({signal_2798, signal_1773}), .clk (CLK), .r (Fresh[545]), .c ({signal_2865, signal_1817}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1674 ( .s ({signal_2190, signal_991}), .b ({signal_2801, signal_1776}), .a ({signal_2716, signal_1714}), .clk (CLK), .r (Fresh[546]), .c ({signal_2866, signal_1818}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1675 ( .s ({signal_2190, signal_991}), .b ({signal_2719, signal_1717}), .a ({signal_2802, signal_1777}), .clk (CLK), .r (Fresh[547]), .c ({signal_2867, signal_1819}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1676 ( .s ({signal_2190, signal_991}), .b ({signal_2802, signal_1777}), .a ({signal_2720, signal_1718}), .clk (CLK), .r (Fresh[548]), .c ({signal_2868, signal_1820}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1677 ( .s ({signal_2190, signal_991}), .b ({signal_2721, signal_1719}), .a ({signal_2801, signal_1776}), .clk (CLK), .r (Fresh[549]), .c ({signal_2869, signal_1821}) ) ;

    /* cells in depth 13 */

    /* cells in depth 14 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1678 ( .s ({signal_2078, signal_981}), .b ({signal_2724, signal_1722}), .a ({signal_2803, signal_1778}), .clk (CLK), .r (Fresh[550]), .c ({signal_2870, signal_1822}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1679 ( .s ({signal_2078, signal_981}), .b ({signal_2805, signal_1780}), .a ({signal_2804, signal_1779}), .clk (CLK), .r (Fresh[551]), .c ({signal_2871, signal_1823}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1680 ( .s ({signal_2210, signal_984}), .b ({signal_2838, signal_1781}), .a ({signal_2757, signal_1723}), .clk (CLK), .r (Fresh[552]), .c ({signal_2890, signal_1824}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1681 ( .s ({signal_2210, signal_984}), .b ({signal_2840, signal_1783}), .a ({signal_2839, signal_1782}), .clk (CLK), .r (Fresh[553]), .c ({signal_2891, signal_1825}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1682 ( .s ({signal_2188, signal_985}), .b ({signal_2765, signal_1731}), .a ({signal_2841, signal_1784}), .clk (CLK), .r (Fresh[554]), .c ({signal_2892, signal_1826}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1683 ( .s ({signal_2188, signal_985}), .b ({signal_2767, signal_1733}), .a ({signal_2842, signal_1785}), .clk (CLK), .r (Fresh[555]), .c ({signal_2893, signal_1827}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1684 ( .s ({signal_2213, signal_978}), .b ({signal_2844, signal_1787}), .a ({signal_2843, signal_1786}), .clk (CLK), .r (Fresh[556]), .c ({signal_2894, signal_1828}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1685 ( .s ({signal_2213, signal_978}), .b ({signal_2845, signal_1788}), .a ({signal_2770, signal_1736}), .clk (CLK), .r (Fresh[557]), .c ({signal_2895, signal_1829}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1686 ( .s ({signal_2189, signal_988}), .b ({signal_2847, signal_1790}), .a ({signal_2846, signal_1789}), .clk (CLK), .r (Fresh[558]), .c ({signal_2896, signal_1830}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1687 ( .s ({signal_2189, signal_988}), .b ({signal_2849, signal_1792}), .a ({signal_2848, signal_1791}), .clk (CLK), .r (Fresh[559]), .c ({signal_2897, signal_1831}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1688 ( .s ({signal_2191, signal_1007}), .b ({signal_2851, signal_1794}), .a ({signal_2850, signal_1793}), .clk (CLK), .r (Fresh[560]), .c ({signal_2898, signal_1832}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1689 ( .s ({signal_2191, signal_1007}), .b ({signal_2850, signal_1793}), .a ({signal_2851, signal_1794}), .clk (CLK), .r (Fresh[561]), .c ({signal_2899, signal_1833}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1690 ( .s ({signal_2247, signal_1001}), .b ({signal_2779, signal_1745}), .a ({signal_2852, signal_1795}), .clk (CLK), .r (Fresh[562]), .c ({signal_2900, signal_1834}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1691 ( .s ({signal_2247, signal_1001}), .b ({signal_2780, signal_1746}), .a ({signal_2853, signal_1796}), .clk (CLK), .r (Fresh[563]), .c ({signal_2901, signal_1835}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1692 ( .s ({signal_2078, signal_981}), .b ({signal_2783, signal_1749}), .a ({signal_2854, signal_1797}), .clk (CLK), .r (Fresh[564]), .c ({signal_2902, signal_1836}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1693 ( .s ({signal_2078, signal_981}), .b ({signal_2786, signal_1752}), .a ({signal_2855, signal_1798}), .clk (CLK), .r (Fresh[565]), .c ({signal_2903, signal_1837}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1694 ( .s ({signal_2199, signal_998}), .b ({signal_2856, signal_1799}), .a ({signal_2787, signal_1753}), .clk (CLK), .r (Fresh[566]), .c ({signal_2904, signal_1838}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1695 ( .s ({signal_2199, signal_998}), .b ({signal_2857, signal_1800}), .a ({signal_2788, signal_1754}), .clk (CLK), .r (Fresh[567]), .c ({signal_2905, signal_1839}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1696 ( .s ({signal_2198, signal_999}), .b ({signal_2807, signal_1802}), .a ({signal_2806, signal_1801}), .clk (CLK), .r (Fresh[568]), .c ({signal_2872, signal_1840}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1697 ( .s ({signal_2198, signal_999}), .b ({signal_2809, signal_1804}), .a ({signal_2808, signal_1803}), .clk (CLK), .r (Fresh[569]), .c ({signal_2873, signal_1841}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1698 ( .s ({signal_2203, signal_994}), .b ({signal_2810, signal_1805}), .a ({signal_2729, signal_1759}), .clk (CLK), .r (Fresh[570]), .c ({signal_2874, signal_1842}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1699 ( .s ({signal_2203, signal_994}), .b ({signal_2811, signal_1806}), .a ({signal_2730, signal_1760}), .clk (CLK), .r (Fresh[571]), .c ({signal_2875, signal_1843}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1700 ( .s ({signal_2190, signal_991}), .b ({signal_2859, signal_1808}), .a ({signal_2858, signal_1807}), .clk (CLK), .r (Fresh[572]), .c ({signal_2906, signal_1844}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1701 ( .s ({signal_2190, signal_991}), .b ({signal_2858, signal_1807}), .a ({signal_2859, signal_1808}), .clk (CLK), .r (Fresh[573]), .c ({signal_2907, signal_1845}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1702 ( .s ({signal_2078, signal_981}), .b ({signal_2733, signal_1767}), .a ({signal_2812, signal_1809}), .clk (CLK), .r (Fresh[574]), .c ({signal_2876, signal_1846}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1703 ( .s ({signal_2078, signal_981}), .b ({signal_2814, signal_1811}), .a ({signal_2813, signal_1810}), .clk (CLK), .r (Fresh[575]), .c ({signal_2877, signal_1847}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1704 ( .s ({signal_2213, signal_978}), .b ({signal_2861, signal_1813}), .a ({signal_2860, signal_1812}), .clk (CLK), .r (Fresh[576]), .c ({signal_2908, signal_1848}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1705 ( .s ({signal_2213, signal_978}), .b ({signal_2862, signal_1814}), .a ({signal_2795, signal_1770}), .clk (CLK), .r (Fresh[577]), .c ({signal_2909, signal_1849}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1706 ( .s ({signal_2210, signal_984}), .b ({signal_2863, signal_1815}), .a ({signal_2796, signal_1771}), .clk (CLK), .r (Fresh[578]), .c ({signal_2910, signal_1850}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1707 ( .s ({signal_2210, signal_984}), .b ({signal_2865, signal_1817}), .a ({signal_2864, signal_1816}), .clk (CLK), .r (Fresh[579]), .c ({signal_2911, signal_1851}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1708 ( .s ({signal_2189, signal_988}), .b ({signal_2867, signal_1819}), .a ({signal_2866, signal_1818}), .clk (CLK), .r (Fresh[580]), .c ({signal_2912, signal_1852}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1709 ( .s ({signal_2189, signal_988}), .b ({signal_2869, signal_1821}), .a ({signal_2868, signal_1820}), .clk (CLK), .r (Fresh[581]), .c ({signal_2913, signal_1853}) ) ;

    /* cells in depth 15 */

    /* cells in depth 16 */
    mux2_masked #(.security_order(1), .pipeline(0)) cell_39 ( .s (signal_343), .b ({signal_2964, signal_1327}), .a ({signal_2072, signal_312}), .c ({signal_2983, signal_1263}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_41 ( .s (signal_344), .b ({signal_3004, signal_1325}), .a ({signal_2193, signal_314}), .c ({signal_3018, signal_1261}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_43 ( .s (signal_342), .b ({signal_2968, signal_1323}), .a ({signal_2194, signal_316}), .c ({signal_2985, signal_1259}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_45 ( .s (signal_342), .b ({signal_2967, signal_1321}), .a ({signal_2196, signal_318}), .c ({signal_2987, signal_1257}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_47 ( .s (signal_342), .b ({signal_2934, signal_1319}), .a ({signal_2198, signal_999}), .c ({signal_2950, signal_1255}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_49 ( .s (signal_342), .b ({signal_3012, signal_1317}), .a ({signal_2200, signal_997}), .c ({signal_3019, signal_1253}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_51 ( .s (signal_342), .b ({signal_2982, signal_1315}), .a ({signal_2202, signal_995}), .c ({signal_2988, signal_1251}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_53 ( .s (signal_342), .b ({signal_3016, signal_1313}), .a ({signal_2204, signal_993}), .c ({signal_3020, signal_1249}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_55 ( .s (signal_343), .b ({signal_3003, signal_1311}), .a ({signal_2074, signal_319}), .c ({signal_3021, signal_1247}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_56 ( .s (signal_343), .b ({signal_3083, signal_1310}), .a ({signal_2206, signal_320}), .c ({signal_3100, signal_1246}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_58 ( .s (signal_343), .b ({signal_3082, signal_1308}), .a ({signal_2075, signal_322}), .c ({signal_3101, signal_1244}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_59 ( .s (signal_343), .b ({signal_2966, signal_1307}), .a ({signal_2208, signal_323}), .c ({signal_2989, signal_1243}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_60 ( .s (signal_343), .b ({signal_3090, signal_1306}), .a ({signal_2209, signal_324}), .c ({signal_3102, signal_1242}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_62 ( .s (signal_343), .b ({signal_3047, signal_1304}), .a ({signal_2210, signal_984}), .c ({signal_3061, signal_1240}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_63 ( .s (signal_343), .b ({signal_2971, signal_1303}), .a ({signal_2077, signal_983}), .c ({signal_2990, signal_1239}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_64 ( .s (signal_343), .b ({signal_3054, signal_1302}), .a ({signal_2211, signal_982}), .c ({signal_3062, signal_1238}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_66 ( .s (signal_343), .b ({signal_3093, signal_1300}), .a ({signal_2212, signal_980}), .c ({signal_3103, signal_1236}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_67 ( .s (signal_344), .b ({signal_3015, signal_1299}), .a ({signal_2181, signal_979}), .c ({signal_3023, signal_1235}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_68 ( .s (signal_344), .b ({signal_3099, signal_1298}), .a ({signal_2213, signal_978}), .c ({signal_3104, signal_1234}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_70 ( .s (signal_344), .b ({signal_3098, signal_1296}), .a ({signal_2215, signal_976}), .c ({signal_3105, signal_1232}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_71 ( .s (signal_344), .b ({signal_3165, signal_1295}), .a ({signal_2182, signal_326}), .c ({signal_3178, signal_1231}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_72 ( .s (signal_344), .b ({signal_3167, signal_1294}), .a ({signal_2216, signal_327}), .c ({signal_3179, signal_1230}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_73 ( .s (signal_344), .b ({signal_3078, signal_1293}), .a ({signal_2183, signal_328}), .c ({signal_3106, signal_1229}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_74 ( .s (signal_344), .b ({signal_3123, signal_1292}), .a ({signal_2184, signal_329}), .c ({signal_3137, signal_1228}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_75 ( .s (signal_344), .b ({signal_3126, signal_1291}), .a ({signal_2185, signal_330}), .c ({signal_3138, signal_1227}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_76 ( .s (signal_344), .b ({signal_3128, signal_1290}), .a ({signal_2217, signal_331}), .c ({signal_3139, signal_1226}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_77 ( .s (signal_344), .b ({signal_3084, signal_1289}), .a ({signal_2218, signal_332}), .c ({signal_3107, signal_1225}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_78 ( .s (signal_344), .b ({signal_3127, signal_1288}), .a ({signal_2186, signal_968}), .c ({signal_3140, signal_1224}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_79 ( .s (signal_344), .b ({signal_3171, signal_1287}), .a ({signal_2219, signal_967}), .c ({signal_3180, signal_1223}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_80 ( .s (signal_343), .b ({signal_3173, signal_1286}), .a ({signal_2220, signal_966}), .c ({signal_3181, signal_1222}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_81 ( .s (signal_342), .b ({signal_3049, signal_1285}), .a ({signal_2221, signal_965}), .c ({signal_3063, signal_1221}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_82 ( .s (signal_340), .b ({signal_3092, signal_1284}), .a ({signal_2222, signal_964}), .c ({signal_3108, signal_1220}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_83 ( .s (signal_343), .b ({signal_3175, signal_1283}), .a ({signal_2223, signal_963}), .c ({signal_3182, signal_1219}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_84 ( .s (signal_342), .b ({signal_3177, signal_1282}), .a ({signal_2224, signal_962}), .c ({signal_3183, signal_1218}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_85 ( .s (signal_344), .b ({signal_3094, signal_1281}), .a ({signal_2225, signal_961}), .c ({signal_3109, signal_1217}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_86 ( .s (signal_340), .b ({signal_3096, signal_1280}), .a ({signal_2226, signal_960}), .c ({signal_3110, signal_1216}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_87 ( .s (signal_340), .b ({signal_3235, signal_1279}), .a ({signal_2227, signal_333}), .c ({signal_3240, signal_1215}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_88 ( .s (signal_340), .b ({signal_3252, signal_1278}), .a ({signal_2228, signal_334}), .c ({signal_3256, signal_1214}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_89 ( .s (signal_340), .b ({signal_3198, signal_1277}), .a ({signal_2229, signal_335}), .c ({signal_3209, signal_1213}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_90 ( .s (signal_340), .b ({signal_3164, signal_1276}), .a ({signal_2230, signal_336}), .c ({signal_3184, signal_1212}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_91 ( .s (signal_340), .b ({signal_3237, signal_1275}), .a ({signal_2231, signal_337}), .c ({signal_3241, signal_1211}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_92 ( .s (signal_340), .b ({signal_3253, signal_1274}), .a ({signal_2232, signal_338}), .c ({signal_3257, signal_1210}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_93 ( .s (signal_344), .b ({signal_3169, signal_1273}), .a ({signal_2233, signal_339}), .c ({signal_3185, signal_1209}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_94 ( .s (signal_343), .b ({signal_3168, signal_1272}), .a ({signal_2234, signal_952}), .c ({signal_3186, signal_1208}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_95 ( .s (signal_342), .b ({signal_3205, signal_1271}), .a ({signal_2235, signal_951}), .c ({signal_3210, signal_1207}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_96 ( .s (signal_344), .b ({signal_3254, signal_1270}), .a ({signal_2236, signal_950}), .c ({signal_3258, signal_1206}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_97 ( .s (signal_343), .b ({signal_3203, signal_1269}), .a ({signal_2237, signal_949}), .c ({signal_3211, signal_1205}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_98 ( .s (signal_342), .b ({signal_3129, signal_1268}), .a ({signal_2238, signal_948}), .c ({signal_3141, signal_1204}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_99 ( .s (signal_343), .b ({signal_3208, signal_1267}), .a ({signal_2239, signal_947}), .c ({signal_3212, signal_1203}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_100 ( .s (signal_342), .b ({signal_3255, signal_1266}), .a ({signal_2240, signal_946}), .c ({signal_3259, signal_1202}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_101 ( .s (signal_344), .b ({signal_3206, signal_1265}), .a ({signal_2241, signal_945}), .c ({signal_3213, signal_1201}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_102 ( .s (signal_344), .b ({signal_3174, signal_1264}), .a ({signal_2242, signal_944}), .c ({signal_3187, signal_1200}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_103 ( .s (IN_reset), .b ({signal_2983, signal_1263}), .a ({IN_plaintext_s1[0], IN_plaintext_s0[0]}), .c ({signal_3026, signal_1199}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_105 ( .s (IN_reset), .b ({signal_3018, signal_1261}), .a ({IN_plaintext_s1[2], IN_plaintext_s0[2]}), .c ({signal_3065, signal_1197}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_107 ( .s (IN_reset), .b ({signal_2985, signal_1259}), .a ({IN_plaintext_s1[4], IN_plaintext_s0[4]}), .c ({signal_3030, signal_1195}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_109 ( .s (IN_reset), .b ({signal_2987, signal_1257}), .a ({IN_plaintext_s1[6], IN_plaintext_s0[6]}), .c ({signal_3034, signal_1193}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_111 ( .s (IN_reset), .b ({signal_2950, signal_1255}), .a ({IN_plaintext_s1[8], IN_plaintext_s0[8]}), .c ({signal_2994, signal_1191}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_113 ( .s (IN_reset), .b ({signal_3019, signal_1253}), .a ({IN_plaintext_s1[10], IN_plaintext_s0[10]}), .c ({signal_3067, signal_1189}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_115 ( .s (IN_reset), .b ({signal_2988, signal_1251}), .a ({IN_plaintext_s1[12], IN_plaintext_s0[12]}), .c ({signal_3036, signal_1187}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_117 ( .s (IN_reset), .b ({signal_3020, signal_1249}), .a ({IN_plaintext_s1[14], IN_plaintext_s0[14]}), .c ({signal_3069, signal_1185}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_119 ( .s (IN_reset), .b ({signal_3021, signal_1247}), .a ({IN_plaintext_s1[16], IN_plaintext_s0[16]}), .c ({signal_3071, signal_1183}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_120 ( .s (IN_reset), .b ({signal_3100, signal_1246}), .a ({IN_plaintext_s1[17], IN_plaintext_s0[17]}), .c ({signal_3143, signal_1182}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_122 ( .s (IN_reset), .b ({signal_3101, signal_1244}), .a ({IN_plaintext_s1[19], IN_plaintext_s0[19]}), .c ({signal_3145, signal_1180}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_123 ( .s (IN_reset), .b ({signal_2989, signal_1243}), .a ({IN_plaintext_s1[20], IN_plaintext_s0[20]}), .c ({signal_3038, signal_1179}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_124 ( .s (IN_reset), .b ({signal_3102, signal_1242}), .a ({IN_plaintext_s1[21], IN_plaintext_s0[21]}), .c ({signal_3147, signal_1178}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_126 ( .s (IN_reset), .b ({signal_3061, signal_1240}), .a ({IN_plaintext_s1[23], IN_plaintext_s0[23]}), .c ({signal_3116, signal_1176}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_127 ( .s (IN_reset), .b ({signal_2990, signal_1239}), .a ({IN_plaintext_s1[24], IN_plaintext_s0[24]}), .c ({signal_3040, signal_1175}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_128 ( .s (IN_reset), .b ({signal_3062, signal_1238}), .a ({IN_plaintext_s1[25], IN_plaintext_s0[25]}), .c ({signal_3118, signal_1174}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_130 ( .s (IN_reset), .b ({signal_3103, signal_1236}), .a ({IN_plaintext_s1[27], IN_plaintext_s0[27]}), .c ({signal_3149, signal_1172}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_131 ( .s (IN_reset), .b ({signal_3023, signal_1235}), .a ({IN_plaintext_s1[28], IN_plaintext_s0[28]}), .c ({signal_3075, signal_1171}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_132 ( .s (IN_reset), .b ({signal_3104, signal_1234}), .a ({IN_plaintext_s1[29], IN_plaintext_s0[29]}), .c ({signal_3151, signal_1170}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_134 ( .s (IN_reset), .b ({signal_3105, signal_1232}), .a ({IN_plaintext_s1[31], IN_plaintext_s0[31]}), .c ({signal_3153, signal_1168}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_135 ( .s (IN_reset), .b ({signal_3178, signal_1231}), .a ({IN_plaintext_s1[32], IN_plaintext_s0[32]}), .c ({signal_3215, signal_1167}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_136 ( .s (IN_reset), .b ({signal_3179, signal_1230}), .a ({IN_plaintext_s1[33], IN_plaintext_s0[33]}), .c ({signal_3217, signal_1166}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_137 ( .s (IN_reset), .b ({signal_3106, signal_1229}), .a ({IN_plaintext_s1[34], IN_plaintext_s0[34]}), .c ({signal_3155, signal_1165}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_138 ( .s (IN_reset), .b ({signal_3137, signal_1228}), .a ({IN_plaintext_s1[35], IN_plaintext_s0[35]}), .c ({signal_3189, signal_1164}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_139 ( .s (IN_reset), .b ({signal_3138, signal_1227}), .a ({IN_plaintext_s1[36], IN_plaintext_s0[36]}), .c ({signal_3191, signal_1163}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_140 ( .s (IN_reset), .b ({signal_3139, signal_1226}), .a ({IN_plaintext_s1[37], IN_plaintext_s0[37]}), .c ({signal_3193, signal_1162}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_141 ( .s (IN_reset), .b ({signal_3107, signal_1225}), .a ({IN_plaintext_s1[38], IN_plaintext_s0[38]}), .c ({signal_3157, signal_1161}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_142 ( .s (IN_reset), .b ({signal_3140, signal_1224}), .a ({IN_plaintext_s1[39], IN_plaintext_s0[39]}), .c ({signal_3195, signal_1160}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_143 ( .s (IN_reset), .b ({signal_3180, signal_1223}), .a ({IN_plaintext_s1[40], IN_plaintext_s0[40]}), .c ({signal_3219, signal_1159}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_144 ( .s (IN_reset), .b ({signal_3181, signal_1222}), .a ({IN_plaintext_s1[41], IN_plaintext_s0[41]}), .c ({signal_3221, signal_1158}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_145 ( .s (IN_reset), .b ({signal_3063, signal_1221}), .a ({IN_plaintext_s1[42], IN_plaintext_s0[42]}), .c ({signal_3120, signal_1157}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_146 ( .s (IN_reset), .b ({signal_3108, signal_1220}), .a ({IN_plaintext_s1[43], IN_plaintext_s0[43]}), .c ({signal_3159, signal_1156}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_147 ( .s (IN_reset), .b ({signal_3182, signal_1219}), .a ({IN_plaintext_s1[44], IN_plaintext_s0[44]}), .c ({signal_3223, signal_1155}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_148 ( .s (IN_reset), .b ({signal_3183, signal_1218}), .a ({IN_plaintext_s1[45], IN_plaintext_s0[45]}), .c ({signal_3225, signal_1154}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_149 ( .s (IN_reset), .b ({signal_3109, signal_1217}), .a ({IN_plaintext_s1[46], IN_plaintext_s0[46]}), .c ({signal_3161, signal_1153}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_150 ( .s (IN_reset), .b ({signal_3110, signal_1216}), .a ({IN_plaintext_s1[47], IN_plaintext_s0[47]}), .c ({signal_3163, signal_1152}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_151 ( .s (IN_reset), .b ({signal_3240, signal_1215}), .a ({IN_plaintext_s1[48], IN_plaintext_s0[48]}), .c ({signal_3261, signal_1151}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_152 ( .s (IN_reset), .b ({signal_3256, signal_1214}), .a ({IN_plaintext_s1[49], IN_plaintext_s0[49]}), .c ({signal_3265, signal_1150}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_153 ( .s (IN_reset), .b ({signal_3209, signal_1213}), .a ({IN_plaintext_s1[50], IN_plaintext_s0[50]}), .c ({signal_3243, signal_1149}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_154 ( .s (IN_reset), .b ({signal_3184, signal_1212}), .a ({IN_plaintext_s1[51], IN_plaintext_s0[51]}), .c ({signal_3227, signal_1148}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_155 ( .s (IN_reset), .b ({signal_3241, signal_1211}), .a ({IN_plaintext_s1[52], IN_plaintext_s0[52]}), .c ({signal_3263, signal_1147}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_156 ( .s (IN_reset), .b ({signal_3257, signal_1210}), .a ({IN_plaintext_s1[53], IN_plaintext_s0[53]}), .c ({signal_3267, signal_1146}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_157 ( .s (IN_reset), .b ({signal_3185, signal_1209}), .a ({IN_plaintext_s1[54], IN_plaintext_s0[54]}), .c ({signal_3229, signal_1145}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_158 ( .s (IN_reset), .b ({signal_3186, signal_1208}), .a ({IN_plaintext_s1[55], IN_plaintext_s0[55]}), .c ({signal_3231, signal_1144}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_159 ( .s (IN_reset), .b ({signal_3210, signal_1207}), .a ({IN_plaintext_s1[56], IN_plaintext_s0[56]}), .c ({signal_3245, signal_1143}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_160 ( .s (IN_reset), .b ({signal_3258, signal_1206}), .a ({IN_plaintext_s1[57], IN_plaintext_s0[57]}), .c ({signal_3269, signal_1142}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_161 ( .s (IN_reset), .b ({signal_3211, signal_1205}), .a ({IN_plaintext_s1[58], IN_plaintext_s0[58]}), .c ({signal_3247, signal_1141}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_162 ( .s (IN_reset), .b ({signal_3141, signal_1204}), .a ({IN_plaintext_s1[59], IN_plaintext_s0[59]}), .c ({signal_3197, signal_1140}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_163 ( .s (IN_reset), .b ({signal_3212, signal_1203}), .a ({IN_plaintext_s1[60], IN_plaintext_s0[60]}), .c ({signal_3249, signal_1139}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_164 ( .s (IN_reset), .b ({signal_3259, signal_1202}), .a ({IN_plaintext_s1[61], IN_plaintext_s0[61]}), .c ({signal_3271, signal_1138}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_165 ( .s (IN_reset), .b ({signal_3213, signal_1201}), .a ({IN_plaintext_s1[62], IN_plaintext_s0[62]}), .c ({signal_3251, signal_1137}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_166 ( .s (IN_reset), .b ({signal_3187, signal_1200}), .a ({IN_plaintext_s1[63], IN_plaintext_s0[63]}), .c ({signal_3233, signal_1136}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_762 ( .a ({signal_3121, signal_656}), .b ({signal_2958, signal_657}), .c ({signal_3164, signal_1276}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_764 ( .a ({signal_3078, signal_1293}), .b ({signal_3041, signal_1309}), .c ({signal_3121, signal_656}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_765 ( .a ({signal_2920, signal_658}), .b ({signal_3044, signal_659}), .c ({signal_3078, signal_1293}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_767 ( .a ({signal_3079, signal_661}), .b ({signal_3167, signal_1294}), .c ({signal_3198, signal_1277}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_768 ( .a ({signal_3004, signal_1325}), .b ({signal_3044, signal_659}), .c ({signal_3079, signal_661}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_769 ( .a ({signal_3234, signal_662}), .b ({signal_3124, signal_663}), .c ({signal_3252, signal_1278}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_770 ( .a ({signal_3199, signal_664}), .b ({signal_3001, signal_665}), .c ({signal_3234, signal_662}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_772 ( .a ({signal_3165, signal_1295}), .b ({signal_3166, signal_666}), .c ({signal_3199, signal_664}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_773 ( .a ({signal_3122, signal_667}), .b ({signal_2959, signal_668}), .c ({signal_3165, signal_1295}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_775 ( .a ({signal_2610, signal_883}), .b ({signal_3082, signal_1308}), .c ({signal_3122, signal_667}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_776 ( .a ({signal_3200, signal_669}), .b ({signal_2964, signal_1327}), .c ({signal_3235, signal_1279}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_777 ( .a ({signal_3082, signal_1308}), .b ({signal_3166, signal_666}), .c ({signal_3200, signal_669}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_778 ( .a ({signal_2609, signal_881}), .b ({signal_3123, signal_1292}), .c ({signal_3166, signal_666}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_779 ( .a ({signal_3080, signal_670}), .b ({signal_2742, signal_671}), .c ({signal_3123, signal_1292}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_781 ( .a ({signal_3041, signal_1309}), .b ({signal_3004, signal_1325}), .c ({signal_3080, signal_670}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_790 ( .a ({signal_3081, signal_679}), .b ({signal_3124, signal_663}), .c ({signal_3167, signal_1294}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_791 ( .a ({signal_3003, signal_1311}), .b ({signal_3082, signal_1308}), .c ({signal_3124, signal_663}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_792 ( .a ({signal_3042, signal_680}), .b ({signal_2744, signal_681}), .c ({signal_3081, signal_679}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_794 ( .a ({signal_3005, signal_682}), .b ({signal_2622, signal_882}), .c ({signal_3042, signal_680}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_795 ( .a ({signal_2947, signal_683}), .b ({signal_2961, signal_684}), .c ({signal_3003, signal_1311}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_798 ( .a ({signal_3043, signal_685}), .b ({signal_2745, signal_686}), .c ({signal_3082, signal_1308}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_800 ( .a ({signal_3004, signal_1325}), .b ({signal_2653, signal_922}), .c ({signal_3043, signal_685}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_801 ( .a ({signal_2941, signal_687}), .b ({signal_2962, signal_688}), .c ({signal_3004, signal_1325}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_802 ( .a ({signal_2937, signal_689}), .b ({signal_2734, signal_940}), .c ({signal_2962, signal_688}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_804 ( .a ({signal_2746, signal_677}), .b ({signal_3044, signal_659}), .c ({signal_3083, signal_1310}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_805 ( .a ({signal_2963, signal_690}), .b ({signal_3005, signal_682}), .c ({signal_3044, signal_659}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_806 ( .a ({signal_2922, signal_1324}), .b ({signal_2964, signal_1327}), .c ({signal_3005, signal_682}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_807 ( .a ({signal_2737, signal_920}), .b ({signal_2937, signal_689}), .c ({signal_2963, signal_690}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_810 ( .a ({signal_2938, signal_691}), .b ({signal_2747, signal_692}), .c ({signal_2964, signal_1327}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_816 ( .a ({signal_3125, signal_694}), .b ({signal_2923, signal_695}), .c ({signal_3168, signal_1272}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_818 ( .a ({signal_3084, signal_1289}), .b ({signal_3045, signal_1305}), .c ({signal_3125, signal_694}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_819 ( .a ({signal_2924, signal_696}), .b ({signal_3048, signal_697}), .c ({signal_3084, signal_1289}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_821 ( .a ({signal_3085, signal_699}), .b ({signal_3128, signal_1290}), .c ({signal_3169, signal_1273}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_822 ( .a ({signal_2967, signal_1321}), .b ({signal_3048, signal_697}), .c ({signal_3085, signal_699}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_823 ( .a ({signal_3236, signal_700}), .b ({signal_3088, signal_701}), .c ({signal_3253, signal_1274}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_824 ( .a ({signal_3201, signal_702}), .b ({signal_3006, signal_703}), .c ({signal_3236, signal_700}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_826 ( .a ({signal_3126, signal_1291}), .b ({signal_3170, signal_704}), .c ({signal_3201, signal_702}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_827 ( .a ({signal_3086, signal_705}), .b ({signal_2925, signal_706}), .c ({signal_3126, signal_1291}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_829 ( .a ({signal_2672, signal_895}), .b ({signal_3047, signal_1304}), .c ({signal_3086, signal_705}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_830 ( .a ({signal_3202, signal_707}), .b ({signal_2968, signal_1323}), .c ({signal_3237, signal_1275}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_831 ( .a ({signal_3047, signal_1304}), .b ({signal_3170, signal_704}), .c ({signal_3202, signal_707}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_832 ( .a ({signal_2649, signal_893}), .b ({signal_3127, signal_1288}), .c ({signal_3170, signal_704}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_833 ( .a ({signal_3087, signal_708}), .b ({signal_2817, signal_709}), .c ({signal_3127, signal_1288}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_835 ( .a ({signal_3045, signal_1305}), .b ({signal_2967, signal_1321}), .c ({signal_3087, signal_708}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_844 ( .a ({signal_3089, signal_717}), .b ({signal_3088, signal_701}), .c ({signal_3128, signal_1290}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_845 ( .a ({signal_2966, signal_1307}), .b ({signal_3047, signal_1304}), .c ({signal_3088, signal_701}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_846 ( .a ({signal_3046, signal_718}), .b ({signal_2749, signal_719}), .c ({signal_3089, signal_717}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_848 ( .a ({signal_3009, signal_720}), .b ({signal_2671, signal_894}), .c ({signal_3046, signal_718}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_849 ( .a ({signal_2917, signal_721}), .b ({signal_2927, signal_722}), .c ({signal_2966, signal_1307}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_852 ( .a ({signal_3008, signal_723}), .b ({signal_2750, signal_724}), .c ({signal_3047, signal_1304}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_854 ( .a ({signal_2967, signal_1321}), .b ({signal_2617, signal_918}), .c ({signal_3008, signal_723}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_855 ( .a ({signal_2942, signal_725}), .b ({signal_2928, signal_726}), .c ({signal_2967, signal_1321}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_856 ( .a ({signal_2914, signal_727}), .b ({signal_2735, signal_936}), .c ({signal_2928, signal_726}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_858 ( .a ({signal_2820, signal_715}), .b ({signal_3048, signal_697}), .c ({signal_3090, signal_1306}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_859 ( .a ({signal_2929, signal_728}), .b ({signal_3009, signal_720}), .c ({signal_3048, signal_697}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_860 ( .a ({signal_2882, signal_1320}), .b ({signal_2968, signal_1323}), .c ({signal_3009, signal_720}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_861 ( .a ({signal_2635, signal_916}), .b ({signal_2914, signal_727}), .c ({signal_2929, signal_728}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_864 ( .a ({signal_2943, signal_729}), .b ({signal_2821, signal_730}), .c ({signal_2968, signal_1323}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_870 ( .a ({signal_3091, signal_732}), .b ({signal_2930, signal_733}), .c ({signal_3129, signal_1268}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_872 ( .a ({signal_3049, signal_1285}), .b ({signal_3010, signal_1301}), .c ({signal_3091, signal_732}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_873 ( .a ({signal_2883, signal_734}), .b ({signal_3013, signal_735}), .c ({signal_3049, signal_1285}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_875 ( .a ({signal_3050, signal_737}), .b ({signal_3173, signal_1286}), .c ({signal_3203, signal_1269}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_876 ( .a ({signal_3012, signal_1317}), .b ({signal_3013, signal_735}), .c ({signal_3050, signal_737}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_877 ( .a ({signal_3238, signal_738}), .b ({signal_3132, signal_739}), .c ({signal_3254, signal_1270}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_878 ( .a ({signal_3204, signal_740}), .b ({signal_2969, signal_741}), .c ({signal_3238, signal_738}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_880 ( .a ({signal_3171, signal_1287}), .b ({signal_3131, signal_742}), .c ({signal_3204, signal_740}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_881 ( .a ({signal_3130, signal_743}), .b ({signal_2931, signal_744}), .c ({signal_3171, signal_1287}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_883 ( .a ({signal_2679, signal_891}), .b ({signal_3093, signal_1300}), .c ({signal_3130, signal_743}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_884 ( .a ({signal_3172, signal_745}), .b ({signal_2934, signal_1319}), .c ({signal_3205, signal_1271}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_885 ( .a ({signal_3093, signal_1300}), .b ({signal_3131, signal_742}), .c ({signal_3172, signal_745}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_886 ( .a ({signal_2677, signal_889}), .b ({signal_3092, signal_1284}), .c ({signal_3131, signal_742}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_887 ( .a ({signal_3051, signal_746}), .b ({signal_2823, signal_747}), .c ({signal_3092, signal_1284}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_889 ( .a ({signal_3010, signal_1301}), .b ({signal_3012, signal_1317}), .c ({signal_3051, signal_746}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_898 ( .a ({signal_3052, signal_755}), .b ({signal_3132, signal_739}), .c ({signal_3173, signal_1286}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_899 ( .a ({signal_2971, signal_1303}), .b ({signal_3093, signal_1300}), .c ({signal_3132, signal_739}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_900 ( .a ({signal_3011, signal_756}), .b ({signal_2827, signal_757}), .c ({signal_3052, signal_755}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_902 ( .a ({signal_2973, signal_758}), .b ({signal_2675, signal_890}), .c ({signal_3011, signal_756}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_903 ( .a ({signal_2946, signal_759}), .b ({signal_2933, signal_760}), .c ({signal_2971, signal_1303}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_906 ( .a ({signal_3053, signal_761}), .b ({signal_2828, signal_762}), .c ({signal_3093, signal_1300}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_908 ( .a ({signal_3012, signal_1317}), .b ({signal_2615, signal_914}), .c ({signal_3053, signal_761}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_909 ( .a ({signal_2944, signal_763}), .b ({signal_2972, signal_764}), .c ({signal_3012, signal_1317}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_910 ( .a ({signal_2939, signal_765}), .b ({signal_2633, signal_932}), .c ({signal_2972, signal_764}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_912 ( .a ({signal_2829, signal_753}), .b ({signal_3013, signal_735}), .c ({signal_3054, signal_1302}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_913 ( .a ({signal_2974, signal_766}), .b ({signal_2973, signal_758}), .c ({signal_3013, signal_735}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_914 ( .a ({signal_2885, signal_1316}), .b ({signal_2934, signal_1319}), .c ({signal_2973, signal_758}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_915 ( .a ({signal_2636, signal_912}), .b ({signal_2939, signal_765}), .c ({signal_2974, signal_766}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_918 ( .a ({signal_2915, signal_767}), .b ({signal_2830, signal_768}), .c ({signal_2934, signal_1319}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_924 ( .a ({signal_3133, signal_770}), .b ({signal_2975, signal_771}), .c ({signal_3174, signal_1264}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_926 ( .a ({signal_3094, signal_1281}), .b ({signal_3014, signal_1297}), .c ({signal_3133, signal_770}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_927 ( .a ({signal_2886, signal_772}), .b ({signal_3058, signal_773}), .c ({signal_3094, signal_1281}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_929 ( .a ({signal_3095, signal_775}), .b ({signal_3177, signal_1282}), .c ({signal_3206, signal_1265}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_930 ( .a ({signal_3016, signal_1313}), .b ({signal_3058, signal_773}), .c ({signal_3095, signal_775}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_931 ( .a ({signal_3239, signal_776}), .b ({signal_3136, signal_777}), .c ({signal_3255, signal_1266}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_932 ( .a ({signal_3207, signal_778}), .b ({signal_2976, signal_779}), .c ({signal_3239, signal_776}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_934 ( .a ({signal_3175, signal_1283}), .b ({signal_3135, signal_780}), .c ({signal_3207, signal_778}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_935 ( .a ({signal_3134, signal_781}), .b ({signal_2977, signal_782}), .c ({signal_3175, signal_1283}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_937 ( .a ({signal_2616, signal_887}), .b ({signal_3098, signal_1296}), .c ({signal_3134, signal_781}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_938 ( .a ({signal_3176, signal_783}), .b ({signal_2982, signal_1315}), .c ({signal_3208, signal_1267}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_939 ( .a ({signal_3098, signal_1296}), .b ({signal_3135, signal_780}), .c ({signal_3176, signal_783}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_940 ( .a ({signal_2621, signal_885}), .b ({signal_3096, signal_1280}), .c ({signal_3135, signal_780}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_941 ( .a ({signal_3055, signal_784}), .b ({signal_2754, signal_785}), .c ({signal_3096, signal_1280}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_943 ( .a ({signal_3014, signal_1297}), .b ({signal_3016, signal_1313}), .c ({signal_3055, signal_784}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_952 ( .a ({signal_3097, signal_793}), .b ({signal_3136, signal_777}), .c ({signal_3177, signal_1282}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_953 ( .a ({signal_3015, signal_1299}), .b ({signal_3098, signal_1296}), .c ({signal_3136, signal_777}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_954 ( .a ({signal_3056, signal_794}), .b ({signal_2834, signal_795}), .c ({signal_3097, signal_793}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_956 ( .a ({signal_3017, signal_796}), .b ({signal_2627, signal_886}), .c ({signal_3056, signal_794}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_957 ( .a ({signal_2948, signal_797}), .b ({signal_2979, signal_798}), .c ({signal_3015, signal_1299}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_960 ( .a ({signal_3057, signal_799}), .b ({signal_2835, signal_800}), .c ({signal_3098, signal_1296}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_962 ( .a ({signal_3016, signal_1313}), .b ({signal_2652, signal_926}), .c ({signal_3057, signal_799}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_963 ( .a ({signal_2916, signal_801}), .b ({signal_2980, signal_802}), .c ({signal_3016, signal_1313}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_964 ( .a ({signal_2940, signal_803}), .b ({signal_2634, signal_928}), .c ({signal_2980, signal_802}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_966 ( .a ({signal_2756, signal_791}), .b ({signal_3058, signal_773}), .c ({signal_3099, signal_1298}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_967 ( .a ({signal_2981, signal_804}), .b ({signal_3017, signal_796}), .c ({signal_3058, signal_773}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_968 ( .a ({signal_2936, signal_1312}), .b ({signal_2982, signal_1315}), .c ({signal_3017, signal_796}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_969 ( .a ({signal_2736, signal_924}), .b ({signal_2940, signal_803}), .c ({signal_2981, signal_804}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_972 ( .a ({signal_2945, signal_805}), .b ({signal_2836, signal_806}), .c ({signal_2982, signal_1315}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1710 ( .s ({signal_2077, signal_983}), .b ({signal_2871, signal_1823}), .a ({signal_2870, signal_1822}), .clk (CLK), .r (Fresh[582]), .c ({signal_2914, signal_727}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1711 ( .s ({signal_2188, signal_985}), .b ({signal_2891, signal_1825}), .a ({signal_2890, signal_1824}), .clk (CLK), .r (Fresh[583]), .c ({signal_2937, signal_689}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1712 ( .s ({signal_2187, signal_1004}), .b ({signal_2893, signal_1827}), .a ({signal_2892, signal_1826}), .clk (CLK), .r (Fresh[584]), .c ({signal_2938, signal_691}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1713 ( .s ({signal_2181, signal_979}), .b ({signal_2895, signal_1829}), .a ({signal_2894, signal_1828}), .clk (CLK), .r (Fresh[585]), .c ({signal_2939, signal_765}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1714 ( .s ({signal_2186, signal_968}), .b ({signal_2897, signal_1831}), .a ({signal_2896, signal_1830}), .clk (CLK), .r (Fresh[586]), .c ({signal_2940, signal_803}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1715 ( .s ({signal_2187, signal_1004}), .b ({signal_2899, signal_1833}), .a ({signal_2898, signal_1832}), .clk (CLK), .r (Fresh[587]), .c ({signal_2941, signal_687}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1716 ( .s ({signal_2197, signal_1000}), .b ({signal_2901, signal_1835}), .a ({signal_2900, signal_1834}), .clk (CLK), .r (Fresh[588]), .c ({signal_2942, signal_725}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1717 ( .s ({signal_2077, signal_983}), .b ({signal_2903, signal_1837}), .a ({signal_2902, signal_1836}), .clk (CLK), .r (Fresh[589]), .c ({signal_2943, signal_729}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1718 ( .s ({signal_2198, signal_999}), .b ({signal_2905, signal_1839}), .a ({signal_2904, signal_1838}), .clk (CLK), .r (Fresh[590]), .c ({signal_2944, signal_763}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1719 ( .s ({signal_2181, signal_979}), .b ({signal_2873, signal_1841}), .a ({signal_2872, signal_1840}), .clk (CLK), .r (Fresh[591]), .c ({signal_2915, signal_767}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1720 ( .s ({signal_2202, signal_995}), .b ({signal_2875, signal_1843}), .a ({signal_2874, signal_1842}), .clk (CLK), .r (Fresh[592]), .c ({signal_2916, signal_801}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1721 ( .s ({signal_2189, signal_988}), .b ({signal_2907, signal_1845}), .a ({signal_2906, signal_1844}), .clk (CLK), .r (Fresh[593]), .c ({signal_2945, signal_805}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1722 ( .s ({signal_2077, signal_983}), .b ({signal_2877, signal_1847}), .a ({signal_2876, signal_1846}), .clk (CLK), .r (Fresh[594]), .c ({signal_2917, signal_721}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1723 ( .s ({signal_2181, signal_979}), .b ({signal_2909, signal_1849}), .a ({signal_2908, signal_1848}), .clk (CLK), .r (Fresh[595]), .c ({signal_2946, signal_759}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1724 ( .s ({signal_2188, signal_985}), .b ({signal_2911, signal_1851}), .a ({signal_2910, signal_1850}), .clk (CLK), .r (Fresh[596]), .c ({signal_2947, signal_683}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1725 ( .s ({signal_2186, signal_968}), .b ({signal_2913, signal_1853}), .a ({signal_2912, signal_1852}), .clk (CLK), .r (Fresh[597]), .c ({signal_2948, signal_797}) ) ;

    /* register cells */
    DFF_X1 cell_979 ( .CK (signal_3870), .D (signal_310), .Q (signal_808), .QN () ) ;
    DFF_X1 cell_981 ( .CK (signal_3870), .D (signal_308), .Q (signal_307), .QN () ) ;
    DFF_X1 cell_983 ( .CK (signal_3870), .D (signal_305), .Q (signal_304), .QN () ) ;
    DFF_X1 cell_985 ( .CK (signal_3870), .D (signal_303), .Q (signal_288), .QN () ) ;
    DFF_X1 cell_987 ( .CK (signal_3870), .D (signal_301), .Q (signal_879), .QN () ) ;
    DFF_X1 cell_989 ( .CK (signal_3870), .D (signal_299), .Q (signal_878), .QN () ) ;
    DFF_X1 cell_991 ( .CK (signal_3870), .D (signal_297), .Q (signal_877), .QN () ) ;
    DFF_X1 cell_993 ( .CK (signal_3870), .D (signal_295), .Q (signal_876), .QN () ) ;
    DFF_X1 cell_995 ( .CK (signal_3870), .D (signal_293), .Q (signal_875), .QN () ) ;
    DFF_X1 cell_997 ( .CK (signal_3870), .D (signal_291), .Q (signal_874), .QN () ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_999 ( .clk (signal_3870), .D ({signal_3026, signal_1199}), .Q ({OUT_ciphertext_s1[0], OUT_ciphertext_s0[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1001 ( .clk (signal_3870), .D ({signal_3028, signal_1198}), .Q ({OUT_ciphertext_s1[1], OUT_ciphertext_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1003 ( .clk (signal_3870), .D ({signal_3065, signal_1197}), .Q ({OUT_ciphertext_s1[2], OUT_ciphertext_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1005 ( .clk (signal_3870), .D ({signal_2992, signal_1196}), .Q ({OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1007 ( .clk (signal_3870), .D ({signal_3030, signal_1195}), .Q ({OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1009 ( .clk (signal_3870), .D ({signal_3032, signal_1194}), .Q ({OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1011 ( .clk (signal_3870), .D ({signal_3034, signal_1193}), .Q ({OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1013 ( .clk (signal_3870), .D ({signal_2955, signal_1192}), .Q ({OUT_ciphertext_s1[7], OUT_ciphertext_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1015 ( .clk (signal_3870), .D ({signal_2994, signal_1191}), .Q ({OUT_ciphertext_s1[8], OUT_ciphertext_s0[8]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1017 ( .clk (signal_3870), .D ({signal_2996, signal_1190}), .Q ({OUT_ciphertext_s1[9], OUT_ciphertext_s0[9]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1019 ( .clk (signal_3870), .D ({signal_3067, signal_1189}), .Q ({OUT_ciphertext_s1[10], OUT_ciphertext_s0[10]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1021 ( .clk (signal_3870), .D ({signal_2957, signal_1188}), .Q ({OUT_ciphertext_s1[11], OUT_ciphertext_s0[11]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1023 ( .clk (signal_3870), .D ({signal_3036, signal_1187}), .Q ({OUT_ciphertext_s1[12], OUT_ciphertext_s0[12]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1025 ( .clk (signal_3870), .D ({signal_2998, signal_1186}), .Q ({OUT_ciphertext_s1[13], OUT_ciphertext_s0[13]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1027 ( .clk (signal_3870), .D ({signal_3069, signal_1185}), .Q ({OUT_ciphertext_s1[14], OUT_ciphertext_s0[14]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1029 ( .clk (signal_3870), .D ({signal_3000, signal_1184}), .Q ({OUT_ciphertext_s1[15], OUT_ciphertext_s0[15]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1031 ( .clk (signal_3870), .D ({signal_3071, signal_1183}), .Q ({OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1033 ( .clk (signal_3870), .D ({signal_3143, signal_1182}), .Q ({OUT_ciphertext_s1[17], OUT_ciphertext_s0[17]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1035 ( .clk (signal_3870), .D ({signal_3112, signal_1181}), .Q ({OUT_ciphertext_s1[18], OUT_ciphertext_s0[18]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1037 ( .clk (signal_3870), .D ({signal_3145, signal_1180}), .Q ({OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1039 ( .clk (signal_3870), .D ({signal_3038, signal_1179}), .Q ({OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1041 ( .clk (signal_3870), .D ({signal_3147, signal_1178}), .Q ({OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1043 ( .clk (signal_3870), .D ({signal_3114, signal_1177}), .Q ({OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1045 ( .clk (signal_3870), .D ({signal_3116, signal_1176}), .Q ({OUT_ciphertext_s1[23], OUT_ciphertext_s0[23]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1047 ( .clk (signal_3870), .D ({signal_3040, signal_1175}), .Q ({OUT_ciphertext_s1[24], OUT_ciphertext_s0[24]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1049 ( .clk (signal_3870), .D ({signal_3118, signal_1174}), .Q ({OUT_ciphertext_s1[25], OUT_ciphertext_s0[25]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1051 ( .clk (signal_3870), .D ({signal_3073, signal_1173}), .Q ({OUT_ciphertext_s1[26], OUT_ciphertext_s0[26]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1053 ( .clk (signal_3870), .D ({signal_3149, signal_1172}), .Q ({OUT_ciphertext_s1[27], OUT_ciphertext_s0[27]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1055 ( .clk (signal_3870), .D ({signal_3075, signal_1171}), .Q ({OUT_ciphertext_s1[28], OUT_ciphertext_s0[28]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1057 ( .clk (signal_3870), .D ({signal_3151, signal_1170}), .Q ({OUT_ciphertext_s1[29], OUT_ciphertext_s0[29]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1059 ( .clk (signal_3870), .D ({signal_3077, signal_1169}), .Q ({OUT_ciphertext_s1[30], OUT_ciphertext_s0[30]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1061 ( .clk (signal_3870), .D ({signal_3153, signal_1168}), .Q ({OUT_ciphertext_s1[31], OUT_ciphertext_s0[31]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1063 ( .clk (signal_3870), .D ({signal_3215, signal_1167}), .Q ({OUT_ciphertext_s1[32], OUT_ciphertext_s0[32]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1065 ( .clk (signal_3870), .D ({signal_3217, signal_1166}), .Q ({OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1067 ( .clk (signal_3870), .D ({signal_3155, signal_1165}), .Q ({OUT_ciphertext_s1[34], OUT_ciphertext_s0[34]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1069 ( .clk (signal_3870), .D ({signal_3189, signal_1164}), .Q ({OUT_ciphertext_s1[35], OUT_ciphertext_s0[35]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1071 ( .clk (signal_3870), .D ({signal_3191, signal_1163}), .Q ({OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1073 ( .clk (signal_3870), .D ({signal_3193, signal_1162}), .Q ({OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1075 ( .clk (signal_3870), .D ({signal_3157, signal_1161}), .Q ({OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1077 ( .clk (signal_3870), .D ({signal_3195, signal_1160}), .Q ({OUT_ciphertext_s1[39], OUT_ciphertext_s0[39]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1079 ( .clk (signal_3870), .D ({signal_3219, signal_1159}), .Q ({OUT_ciphertext_s1[40], OUT_ciphertext_s0[40]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1081 ( .clk (signal_3870), .D ({signal_3221, signal_1158}), .Q ({OUT_ciphertext_s1[41], OUT_ciphertext_s0[41]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1083 ( .clk (signal_3870), .D ({signal_3120, signal_1157}), .Q ({OUT_ciphertext_s1[42], OUT_ciphertext_s0[42]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1085 ( .clk (signal_3870), .D ({signal_3159, signal_1156}), .Q ({OUT_ciphertext_s1[43], OUT_ciphertext_s0[43]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1087 ( .clk (signal_3870), .D ({signal_3223, signal_1155}), .Q ({OUT_ciphertext_s1[44], OUT_ciphertext_s0[44]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1089 ( .clk (signal_3870), .D ({signal_3225, signal_1154}), .Q ({OUT_ciphertext_s1[45], OUT_ciphertext_s0[45]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1091 ( .clk (signal_3870), .D ({signal_3161, signal_1153}), .Q ({OUT_ciphertext_s1[46], OUT_ciphertext_s0[46]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1093 ( .clk (signal_3870), .D ({signal_3163, signal_1152}), .Q ({OUT_ciphertext_s1[47], OUT_ciphertext_s0[47]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1095 ( .clk (signal_3870), .D ({signal_3261, signal_1151}), .Q ({OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1097 ( .clk (signal_3870), .D ({signal_3265, signal_1150}), .Q ({OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1099 ( .clk (signal_3870), .D ({signal_3243, signal_1149}), .Q ({OUT_ciphertext_s1[50], OUT_ciphertext_s0[50]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1101 ( .clk (signal_3870), .D ({signal_3227, signal_1148}), .Q ({OUT_ciphertext_s1[51], OUT_ciphertext_s0[51]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1103 ( .clk (signal_3870), .D ({signal_3263, signal_1147}), .Q ({OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1105 ( .clk (signal_3870), .D ({signal_3267, signal_1146}), .Q ({OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1107 ( .clk (signal_3870), .D ({signal_3229, signal_1145}), .Q ({OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1109 ( .clk (signal_3870), .D ({signal_3231, signal_1144}), .Q ({OUT_ciphertext_s1[55], OUT_ciphertext_s0[55]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1111 ( .clk (signal_3870), .D ({signal_3245, signal_1143}), .Q ({OUT_ciphertext_s1[56], OUT_ciphertext_s0[56]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1113 ( .clk (signal_3870), .D ({signal_3269, signal_1142}), .Q ({OUT_ciphertext_s1[57], OUT_ciphertext_s0[57]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1115 ( .clk (signal_3870), .D ({signal_3247, signal_1141}), .Q ({OUT_ciphertext_s1[58], OUT_ciphertext_s0[58]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1117 ( .clk (signal_3870), .D ({signal_3197, signal_1140}), .Q ({OUT_ciphertext_s1[59], OUT_ciphertext_s0[59]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1119 ( .clk (signal_3870), .D ({signal_3249, signal_1139}), .Q ({OUT_ciphertext_s1[60], OUT_ciphertext_s0[60]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1121 ( .clk (signal_3870), .D ({signal_3271, signal_1138}), .Q ({OUT_ciphertext_s1[61], OUT_ciphertext_s0[61]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1123 ( .clk (signal_3870), .D ({signal_3251, signal_1137}), .Q ({OUT_ciphertext_s1[62], OUT_ciphertext_s0[62]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1125 ( .clk (signal_3870), .D ({signal_3233, signal_1136}), .Q ({OUT_ciphertext_s1[63], OUT_ciphertext_s0[63]}) ) ;
    DFF_X1 cell_1127 ( .CK (signal_3870), .D (signal_265), .Q (OUT_done), .QN () ) ;
endmodule
