/* modified netlist. Source: module Midori64 in file /Midori_round_based/AGEMA/Midori64.v */
/* clock gating is added to the circuit, the latency increased 2 time(s)  */

module Midori64_GHPC_ANF_ClockGating_d1 (DataIn_s0, key_s0, clk, reset, enc_dec, key_s1, DataIn_s1, Fresh, DataOut_s0, done, DataOut_s1, Synch);
    input [63:0] DataIn_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input reset ;
    input enc_dec ;
    input [127:0] key_s1 ;
    input [63:0] DataIn_s1 ;
    input [63:0] Fresh ;
    output [63:0] DataOut_s0 ;
    output done ;
    output [63:0] DataOut_s1 ;
    output Synch ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_286 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_295 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_352 ;
    wire signal_353 ;
    wire signal_354 ;
    wire signal_355 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_359 ;
    wire signal_360 ;
    wire signal_361 ;
    wire signal_362 ;
    wire signal_363 ;
    wire signal_364 ;
    wire signal_365 ;
    wire signal_366 ;
    wire signal_367 ;
    wire signal_368 ;
    wire signal_369 ;
    wire signal_370 ;
    wire signal_371 ;
    wire signal_372 ;
    wire signal_373 ;
    wire signal_374 ;
    wire signal_375 ;
    wire signal_376 ;
    wire signal_377 ;
    wire signal_378 ;
    wire signal_379 ;
    wire signal_380 ;
    wire signal_381 ;
    wire signal_382 ;
    wire signal_383 ;
    wire signal_384 ;
    wire signal_385 ;
    wire signal_386 ;
    wire signal_387 ;
    wire signal_388 ;
    wire signal_389 ;
    wire signal_390 ;
    wire signal_391 ;
    wire signal_392 ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_415 ;
    wire signal_416 ;
    wire signal_417 ;
    wire signal_418 ;
    wire signal_419 ;
    wire signal_420 ;
    wire signal_421 ;
    wire signal_422 ;
    wire signal_423 ;
    wire signal_424 ;
    wire signal_425 ;
    wire signal_426 ;
    wire signal_427 ;
    wire signal_428 ;
    wire signal_429 ;
    wire signal_430 ;
    wire signal_431 ;
    wire signal_432 ;
    wire signal_433 ;
    wire signal_434 ;
    wire signal_435 ;
    wire signal_436 ;
    wire signal_437 ;
    wire signal_438 ;
    wire signal_439 ;
    wire signal_440 ;
    wire signal_441 ;
    wire signal_442 ;
    wire signal_443 ;
    wire signal_444 ;
    wire signal_445 ;
    wire signal_446 ;
    wire signal_447 ;
    wire signal_448 ;
    wire signal_449 ;
    wire signal_450 ;
    wire signal_451 ;
    wire signal_452 ;
    wire signal_453 ;
    wire signal_454 ;
    wire signal_455 ;
    wire signal_456 ;
    wire signal_457 ;
    wire signal_458 ;
    wire signal_459 ;
    wire signal_460 ;
    wire signal_462 ;
    wire signal_464 ;
    wire signal_466 ;
    wire signal_468 ;
    wire signal_470 ;
    wire signal_472 ;
    wire signal_474 ;
    wire signal_476 ;
    wire signal_478 ;
    wire signal_480 ;
    wire signal_482 ;
    wire signal_484 ;
    wire signal_486 ;
    wire signal_488 ;
    wire signal_490 ;
    wire signal_492 ;
    wire signal_494 ;
    wire signal_496 ;
    wire signal_498 ;
    wire signal_500 ;
    wire signal_502 ;
    wire signal_504 ;
    wire signal_506 ;
    wire signal_508 ;
    wire signal_510 ;
    wire signal_512 ;
    wire signal_514 ;
    wire signal_516 ;
    wire signal_518 ;
    wire signal_520 ;
    wire signal_522 ;
    wire signal_524 ;
    wire signal_526 ;
    wire signal_528 ;
    wire signal_530 ;
    wire signal_532 ;
    wire signal_534 ;
    wire signal_536 ;
    wire signal_538 ;
    wire signal_540 ;
    wire signal_542 ;
    wire signal_544 ;
    wire signal_546 ;
    wire signal_548 ;
    wire signal_550 ;
    wire signal_552 ;
    wire signal_554 ;
    wire signal_556 ;
    wire signal_558 ;
    wire signal_560 ;
    wire signal_562 ;
    wire signal_564 ;
    wire signal_566 ;
    wire signal_568 ;
    wire signal_570 ;
    wire signal_572 ;
    wire signal_574 ;
    wire signal_576 ;
    wire signal_578 ;
    wire signal_580 ;
    wire signal_582 ;
    wire signal_584 ;
    wire signal_586 ;
    wire signal_828 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_831 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_834 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_837 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_840 ;
    wire signal_841 ;
    wire signal_842 ;
    wire signal_843 ;
    wire signal_844 ;
    wire signal_845 ;
    wire signal_846 ;
    wire signal_847 ;
    wire signal_848 ;
    wire signal_849 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_852 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_855 ;
    wire signal_856 ;
    wire signal_857 ;
    wire signal_858 ;
    wire signal_859 ;
    wire signal_860 ;
    wire signal_861 ;
    wire signal_862 ;
    wire signal_863 ;
    wire signal_864 ;
    wire signal_865 ;
    wire signal_866 ;
    wire signal_867 ;
    wire signal_868 ;
    wire signal_869 ;
    wire signal_870 ;
    wire signal_871 ;
    wire signal_872 ;
    wire signal_873 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_879 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_885 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_888 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_891 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_894 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_897 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_900 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_903 ;
    wire signal_904 ;
    wire signal_905 ;
    wire signal_906 ;
    wire signal_907 ;
    wire signal_908 ;
    wire signal_909 ;
    wire signal_910 ;
    wire signal_911 ;
    wire signal_912 ;
    wire signal_913 ;
    wire signal_914 ;
    wire signal_915 ;
    wire signal_916 ;
    wire signal_917 ;
    wire signal_918 ;
    wire signal_919 ;
    wire signal_920 ;
    wire signal_921 ;
    wire signal_922 ;
    wire signal_923 ;
    wire signal_924 ;
    wire signal_925 ;
    wire signal_926 ;
    wire signal_927 ;
    wire signal_928 ;
    wire signal_929 ;
    wire signal_930 ;
    wire signal_931 ;
    wire signal_932 ;
    wire signal_933 ;
    wire signal_934 ;
    wire signal_935 ;
    wire signal_936 ;
    wire signal_937 ;
    wire signal_938 ;
    wire signal_939 ;
    wire signal_940 ;
    wire signal_941 ;
    wire signal_942 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1020 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1023 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1276 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1279 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1282 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1285 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1288 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1294 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1297 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1300 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1303 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1309 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1458 ;
    wire signal_1461 ;
    wire signal_1464 ;
    wire signal_1467 ;
    wire signal_1470 ;
    wire signal_1473 ;
    wire signal_1476 ;
    wire signal_1479 ;
    wire signal_1482 ;
    wire signal_1485 ;
    wire signal_1488 ;
    wire signal_1491 ;
    wire signal_1494 ;
    wire signal_1497 ;
    wire signal_1500 ;
    wire signal_1503 ;
    wire signal_1506 ;
    wire signal_1509 ;
    wire signal_1512 ;
    wire signal_1515 ;
    wire signal_1518 ;
    wire signal_1521 ;
    wire signal_1524 ;
    wire signal_1527 ;
    wire signal_1530 ;
    wire signal_1533 ;
    wire signal_1536 ;
    wire signal_1539 ;
    wire signal_1542 ;
    wire signal_1545 ;
    wire signal_1548 ;
    wire signal_1551 ;
    wire signal_1554 ;
    wire signal_1557 ;
    wire signal_1560 ;
    wire signal_1563 ;
    wire signal_1566 ;
    wire signal_1569 ;
    wire signal_1572 ;
    wire signal_1575 ;
    wire signal_1578 ;
    wire signal_1581 ;
    wire signal_1584 ;
    wire signal_1587 ;
    wire signal_1590 ;
    wire signal_1593 ;
    wire signal_1596 ;
    wire signal_1599 ;
    wire signal_1602 ;
    wire signal_1605 ;
    wire signal_1608 ;
    wire signal_1611 ;
    wire signal_1614 ;
    wire signal_1617 ;
    wire signal_1620 ;
    wire signal_1623 ;
    wire signal_1626 ;
    wire signal_1629 ;
    wire signal_1632 ;
    wire signal_1635 ;
    wire signal_1638 ;
    wire signal_1641 ;
    wire signal_1644 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1657 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1660 ;
    wire signal_1662 ;
    wire signal_1664 ;
    wire signal_1666 ;
    wire signal_1668 ;
    wire signal_1670 ;
    wire signal_1672 ;
    wire signal_1674 ;
    wire signal_1676 ;
    wire signal_1678 ;
    wire signal_1680 ;
    wire signal_1682 ;
    wire signal_1684 ;
    wire signal_1686 ;
    wire signal_1688 ;
    wire signal_1690 ;
    wire signal_1692 ;
    wire signal_1694 ;
    wire signal_1696 ;
    wire signal_1698 ;
    wire signal_1700 ;
    wire signal_1702 ;
    wire signal_1704 ;
    wire signal_1706 ;
    wire signal_1708 ;
    wire signal_1710 ;
    wire signal_1712 ;
    wire signal_1714 ;
    wire signal_1716 ;
    wire signal_1718 ;
    wire signal_1720 ;
    wire signal_1722 ;
    wire signal_1724 ;
    wire signal_1726 ;
    wire signal_1728 ;
    wire signal_1730 ;
    wire signal_1732 ;
    wire signal_1734 ;
    wire signal_1736 ;
    wire signal_1738 ;
    wire signal_1740 ;
    wire signal_1742 ;
    wire signal_1744 ;
    wire signal_1746 ;
    wire signal_1748 ;
    wire signal_1750 ;
    wire signal_1752 ;
    wire signal_1754 ;
    wire signal_1756 ;
    wire signal_1758 ;
    wire signal_1760 ;
    wire signal_1762 ;
    wire signal_1764 ;
    wire signal_1766 ;
    wire signal_1768 ;
    wire signal_1770 ;
    wire signal_1772 ;
    wire signal_1774 ;
    wire signal_1776 ;
    wire signal_1778 ;
    wire signal_1780 ;
    wire signal_1782 ;
    wire signal_1784 ;
    wire signal_1786 ;
    wire signal_1788 ;
    wire signal_1789 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1792 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1795 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1813 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1844 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1854 ;
    wire signal_1855 ;
    wire signal_1856 ;
    wire signal_1857 ;
    wire signal_1858 ;
    wire signal_1859 ;
    wire signal_1860 ;
    wire signal_1861 ;
    wire signal_1862 ;
    wire signal_1863 ;
    wire signal_1864 ;
    wire signal_1865 ;
    wire signal_1866 ;
    wire signal_1867 ;
    wire signal_1868 ;
    wire signal_1869 ;
    wire signal_1870 ;
    wire signal_1871 ;
    wire signal_1872 ;
    wire signal_1873 ;
    wire signal_1874 ;
    wire signal_1875 ;
    wire signal_1876 ;
    wire signal_1877 ;
    wire signal_1878 ;
    wire signal_1879 ;
    wire signal_1880 ;
    wire signal_1881 ;
    wire signal_1882 ;
    wire signal_1883 ;
    wire signal_1884 ;
    wire signal_1885 ;
    wire signal_1886 ;
    wire signal_1887 ;
    wire signal_1888 ;
    wire signal_1889 ;
    wire signal_1890 ;
    wire signal_1891 ;
    wire signal_1892 ;
    wire signal_1893 ;
    wire signal_1894 ;
    wire signal_1895 ;
    wire signal_1896 ;
    wire signal_1897 ;
    wire signal_1898 ;
    wire signal_1899 ;
    wire signal_1900 ;
    wire signal_1901 ;
    wire signal_1902 ;
    wire signal_1903 ;
    wire signal_1904 ;
    wire signal_1905 ;
    wire signal_1906 ;
    wire signal_1907 ;
    wire signal_1908 ;
    wire signal_1909 ;
    wire signal_1910 ;
    wire signal_1911 ;
    wire signal_1912 ;
    wire signal_1913 ;
    wire signal_1914 ;
    wire signal_1915 ;
    wire signal_1916 ;
    wire signal_1981 ;
    wire signal_1982 ;
    wire signal_1983 ;
    wire signal_1984 ;
    wire signal_1985 ;
    wire signal_1986 ;
    wire signal_1987 ;
    wire signal_1988 ;
    wire signal_1989 ;
    wire signal_1990 ;
    wire signal_1991 ;
    wire signal_1992 ;
    wire signal_1993 ;
    wire signal_1994 ;
    wire signal_1995 ;
    wire signal_1996 ;
    wire signal_1997 ;
    wire signal_1998 ;
    wire signal_1999 ;
    wire signal_2000 ;
    wire signal_2001 ;
    wire signal_2002 ;
    wire signal_2003 ;
    wire signal_2004 ;
    wire signal_2005 ;
    wire signal_2006 ;
    wire signal_2007 ;
    wire signal_2008 ;
    wire signal_2009 ;
    wire signal_2010 ;
    wire signal_2011 ;
    wire signal_2012 ;
    wire signal_2013 ;
    wire signal_2014 ;
    wire signal_2015 ;
    wire signal_2016 ;
    wire signal_2017 ;
    wire signal_2018 ;
    wire signal_2019 ;
    wire signal_2020 ;
    wire signal_2021 ;
    wire signal_2022 ;
    wire signal_2023 ;
    wire signal_2024 ;
    wire signal_2025 ;
    wire signal_2026 ;
    wire signal_2027 ;
    wire signal_2028 ;
    wire signal_2029 ;
    wire signal_2030 ;
    wire signal_2031 ;
    wire signal_2032 ;
    wire signal_2033 ;
    wire signal_2034 ;
    wire signal_2035 ;
    wire signal_2036 ;
    wire signal_2037 ;
    wire signal_2038 ;
    wire signal_2039 ;
    wire signal_2040 ;
    wire signal_2041 ;
    wire signal_2042 ;
    wire signal_2043 ;
    wire signal_2044 ;
    wire signal_2045 ;
    wire signal_2046 ;
    wire signal_2047 ;
    wire signal_2048 ;
    wire signal_2049 ;
    wire signal_2050 ;
    wire signal_2051 ;
    wire signal_2052 ;
    wire signal_2053 ;
    wire signal_2054 ;
    wire signal_2055 ;
    wire signal_2056 ;
    wire signal_2057 ;
    wire signal_2058 ;
    wire signal_2059 ;
    wire signal_2060 ;
    wire signal_2061 ;
    wire signal_2062 ;
    wire signal_2063 ;
    wire signal_2064 ;
    wire signal_2065 ;
    wire signal_2066 ;
    wire signal_2067 ;
    wire signal_2068 ;
    wire signal_2069 ;
    wire signal_2070 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2079 ;
    wire signal_2080 ;
    wire signal_2081 ;
    wire signal_2082 ;
    wire signal_2083 ;
    wire signal_2084 ;
    wire signal_2085 ;
    wire signal_2086 ;
    wire signal_2087 ;
    wire signal_2088 ;
    wire signal_2089 ;
    wire signal_2090 ;
    wire signal_2091 ;
    wire signal_2092 ;
    wire signal_2093 ;
    wire signal_2094 ;
    wire signal_2095 ;
    wire signal_2096 ;
    wire signal_2097 ;
    wire signal_2098 ;
    wire signal_2099 ;
    wire signal_2100 ;
    wire signal_2101 ;
    wire signal_2102 ;
    wire signal_2103 ;
    wire signal_2104 ;
    wire signal_2105 ;
    wire signal_2106 ;
    wire signal_2107 ;
    wire signal_2108 ;
    wire signal_2109 ;
    wire signal_2110 ;
    wire signal_2111 ;
    wire signal_2112 ;
    wire signal_2113 ;
    wire signal_2114 ;
    wire signal_2115 ;
    wire signal_2116 ;
    wire signal_2117 ;
    wire signal_2118 ;
    wire signal_2119 ;
    wire signal_2120 ;
    wire signal_2121 ;
    wire signal_2122 ;
    wire signal_2123 ;
    wire signal_2124 ;
    wire signal_2125 ;
    wire signal_2126 ;
    wire signal_2127 ;
    wire signal_2128 ;
    wire signal_2129 ;
    wire signal_2130 ;
    wire signal_2131 ;
    wire signal_2132 ;
    wire signal_2133 ;
    wire signal_2134 ;
    wire signal_2135 ;
    wire signal_2136 ;
    wire signal_2137 ;
    wire signal_2138 ;
    wire signal_2139 ;
    wire signal_2140 ;
    wire signal_2141 ;
    wire signal_2142 ;
    wire signal_2143 ;
    wire signal_2144 ;
    wire signal_2145 ;
    wire signal_2146 ;
    wire signal_2147 ;
    wire signal_2148 ;
    wire signal_2149 ;
    wire signal_2150 ;
    wire signal_2151 ;
    wire signal_2152 ;
    wire signal_2153 ;
    wire signal_2154 ;
    wire signal_2155 ;
    wire signal_2156 ;
    wire signal_2157 ;
    wire signal_2158 ;
    wire signal_2159 ;
    wire signal_2160 ;
    wire signal_2161 ;
    wire signal_2162 ;
    wire signal_2163 ;
    wire signal_2164 ;
    wire signal_2165 ;
    wire signal_2166 ;
    wire signal_2167 ;
    wire signal_2168 ;
    wire signal_2169 ;
    wire signal_2170 ;
    wire signal_2171 ;
    wire signal_2172 ;
    wire signal_2173 ;
    wire signal_2174 ;
    wire signal_2175 ;
    wire signal_2176 ;
    wire signal_2177 ;
    wire signal_2178 ;
    wire signal_2179 ;
    wire signal_2180 ;
    wire signal_2181 ;
    wire signal_2182 ;
    wire signal_2183 ;
    wire signal_2184 ;
    wire signal_2185 ;
    wire signal_2186 ;
    wire signal_2187 ;
    wire signal_2188 ;
    wire signal_2189 ;
    wire signal_2190 ;
    wire signal_2191 ;
    wire signal_2192 ;
    wire signal_2193 ;
    wire signal_2194 ;
    wire signal_2195 ;
    wire signal_2196 ;
    wire signal_2197 ;
    wire signal_2198 ;
    wire signal_2199 ;
    wire signal_2200 ;
    wire signal_2201 ;
    wire signal_2202 ;
    wire signal_2203 ;
    wire signal_2204 ;
    wire signal_2205 ;
    wire signal_2206 ;
    wire signal_2207 ;
    wire signal_2208 ;
    wire signal_2209 ;
    wire signal_2210 ;
    wire signal_2211 ;
    wire signal_2212 ;
    wire signal_2213 ;
    wire signal_2214 ;
    wire signal_2215 ;
    wire signal_2216 ;
    wire signal_2217 ;
    wire signal_2218 ;
    wire signal_2219 ;
    wire signal_2220 ;
    wire signal_2221 ;
    wire signal_2222 ;
    wire signal_2223 ;
    wire signal_2224 ;
    wire signal_2225 ;
    wire signal_2226 ;
    wire signal_2227 ;
    wire signal_2228 ;
    wire signal_2229 ;
    wire signal_2230 ;
    wire signal_2231 ;
    wire signal_2232 ;
    wire signal_2233 ;
    wire signal_2234 ;
    wire signal_2235 ;
    wire signal_2236 ;
    wire signal_2237 ;
    wire signal_2238 ;
    wire signal_2239 ;
    wire signal_2240 ;
    wire signal_2241 ;
    wire signal_2242 ;
    wire signal_2243 ;
    wire signal_2244 ;
    wire signal_2245 ;
    wire signal_2246 ;
    wire signal_2247 ;
    wire signal_2248 ;
    wire signal_2249 ;
    wire signal_2250 ;
    wire signal_2251 ;
    wire signal_2252 ;
    wire signal_2253 ;
    wire signal_2254 ;
    wire signal_2255 ;
    wire signal_2256 ;
    wire signal_2257 ;
    wire signal_2258 ;
    wire signal_2259 ;
    wire signal_2260 ;
    wire signal_2261 ;
    wire signal_2262 ;
    wire signal_2263 ;
    wire signal_2264 ;
    wire signal_2265 ;
    wire signal_2266 ;
    wire signal_2267 ;
    wire signal_2268 ;
    wire signal_2269 ;
    wire signal_2270 ;
    wire signal_2271 ;
    wire signal_2272 ;
    wire signal_2273 ;
    wire signal_2274 ;
    wire signal_2275 ;
    wire signal_2276 ;
    wire signal_2277 ;
    wire signal_2278 ;
    wire signal_2279 ;
    wire signal_2280 ;
    wire signal_2281 ;
    wire signal_2282 ;
    wire signal_2283 ;
    wire signal_2284 ;
    wire signal_2285 ;
    wire signal_2286 ;
    wire signal_2287 ;
    wire signal_2288 ;
    wire signal_2289 ;
    wire signal_2290 ;
    wire signal_2291 ;
    wire signal_2292 ;
    wire signal_2293 ;
    wire signal_2294 ;
    wire signal_2295 ;
    wire signal_2296 ;
    wire signal_2297 ;
    wire signal_2298 ;
    wire signal_2299 ;
    wire signal_2300 ;
    wire signal_2301 ;
    wire signal_2302 ;
    wire signal_2303 ;
    wire signal_2304 ;
    wire signal_2305 ;
    wire signal_2306 ;
    wire signal_2307 ;
    wire signal_2308 ;
    wire signal_2309 ;
    wire signal_2310 ;
    wire signal_2311 ;
    wire signal_2312 ;
    wire signal_2313 ;
    wire signal_2314 ;
    wire signal_2315 ;
    wire signal_2316 ;
    wire signal_2317 ;
    wire signal_2318 ;
    wire signal_2319 ;
    wire signal_2320 ;
    wire signal_2321 ;
    wire signal_2322 ;
    wire signal_2323 ;
    wire signal_2324 ;
    wire signal_2325 ;
    wire signal_2326 ;
    wire signal_2327 ;
    wire signal_2328 ;
    wire signal_2329 ;
    wire signal_2330 ;
    wire signal_2331 ;
    wire signal_2332 ;
    wire signal_2333 ;
    wire signal_2334 ;
    wire signal_2335 ;
    wire signal_2336 ;
    wire signal_2337 ;
    wire signal_2338 ;
    wire signal_2339 ;
    wire signal_2340 ;
    wire signal_2341 ;
    wire signal_2342 ;
    wire signal_2343 ;
    wire signal_2344 ;
    wire signal_2345 ;
    wire signal_2346 ;
    wire signal_2347 ;
    wire signal_2348 ;
    wire signal_2349 ;
    wire signal_2350 ;
    wire signal_2351 ;
    wire signal_2352 ;
    wire signal_2353 ;
    wire signal_2354 ;
    wire signal_2355 ;
    wire signal_2356 ;
    wire signal_2357 ;
    wire signal_2358 ;
    wire signal_2359 ;
    wire signal_2360 ;
    wire signal_2361 ;
    wire signal_2362 ;
    wire signal_2363 ;
    wire signal_2364 ;
    wire signal_2365 ;
    wire signal_2366 ;
    wire signal_2367 ;
    wire signal_2368 ;
    wire signal_2369 ;
    wire signal_2370 ;
    wire signal_2371 ;
    wire signal_2372 ;
    wire signal_2373 ;
    wire signal_2374 ;
    wire signal_2375 ;
    wire signal_2376 ;
    wire signal_2377 ;
    wire signal_2378 ;
    wire signal_2379 ;
    wire signal_2380 ;
    wire signal_2381 ;
    wire signal_2382 ;
    wire signal_2383 ;
    wire signal_2384 ;
    wire signal_2385 ;
    wire signal_2386 ;
    wire signal_2387 ;
    wire signal_2388 ;
    wire signal_2389 ;
    wire signal_2390 ;
    wire signal_2391 ;
    wire signal_2392 ;
    wire signal_2393 ;
    wire signal_2394 ;
    wire signal_2395 ;
    wire signal_2396 ;
    wire signal_2397 ;
    wire signal_2398 ;
    wire signal_2399 ;
    wire signal_2400 ;
    wire signal_2401 ;
    wire signal_2402 ;
    wire signal_2403 ;
    wire signal_2404 ;
    wire signal_2405 ;
    wire signal_2406 ;
    wire signal_2407 ;
    wire signal_2408 ;
    wire signal_2409 ;
    wire signal_2410 ;
    wire signal_2411 ;
    wire signal_2412 ;
    wire signal_2413 ;
    wire signal_2414 ;
    wire signal_2415 ;
    wire signal_2416 ;
    wire signal_2417 ;
    wire signal_2418 ;
    wire signal_2419 ;
    wire signal_2420 ;
    wire signal_2421 ;
    wire signal_2422 ;
    wire signal_2423 ;
    wire signal_2424 ;
    wire signal_2425 ;
    wire signal_2426 ;
    wire signal_2427 ;
    wire signal_2428 ;
    wire signal_2429 ;
    wire signal_2430 ;
    wire signal_2431 ;
    wire signal_2432 ;
    wire signal_2433 ;
    wire signal_2434 ;
    wire signal_2435 ;
    wire signal_2436 ;
    wire signal_2437 ;
    wire signal_2438 ;
    wire signal_2439 ;
    wire signal_2440 ;
    wire signal_2441 ;
    wire signal_2442 ;
    wire signal_2443 ;
    wire signal_2444 ;
    wire signal_2445 ;
    wire signal_2446 ;
    wire signal_2447 ;
    wire signal_2448 ;
    wire signal_2449 ;
    wire signal_2450 ;
    wire signal_2451 ;
    wire signal_2452 ;
    wire signal_2453 ;
    wire signal_2454 ;
    wire signal_2455 ;
    wire signal_2456 ;
    wire signal_2457 ;
    wire signal_2458 ;
    wire signal_2459 ;
    wire signal_2460 ;
    wire signal_2461 ;
    wire signal_2462 ;
    wire signal_2463 ;
    wire signal_2528 ;

    /* cells in depth 0 */
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_0 ( .a ({key_s1[73], key_s0[73]}), .b ({key_s1[9], key_s0[9]}), .c ({signal_1458, signal_914}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1 ( .a ({key_s1[72], key_s0[72]}), .b ({key_s1[8], key_s0[8]}), .c ({signal_1461, signal_915}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_2 ( .a ({key_s1[71], key_s0[71]}), .b ({key_s1[7], key_s0[7]}), .c ({signal_1464, signal_916}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3 ( .a ({key_s1[6], key_s0[6]}), .b ({key_s1[70], key_s0[70]}), .c ({signal_1467, signal_917}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_4 ( .a ({key_s1[127], key_s0[127]}), .b ({key_s1[63], key_s0[63]}), .c ({signal_1470, signal_860}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_5 ( .a ({key_s1[126], key_s0[126]}), .b ({key_s1[62], key_s0[62]}), .c ({signal_1473, signal_861}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_6 ( .a ({key_s1[125], key_s0[125]}), .b ({key_s1[61], key_s0[61]}), .c ({signal_1476, signal_862}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_7 ( .a ({key_s1[124], key_s0[124]}), .b ({key_s1[60], key_s0[60]}), .c ({signal_1479, signal_863}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_8 ( .a ({key_s1[5], key_s0[5]}), .b ({key_s1[69], key_s0[69]}), .c ({signal_1482, signal_918}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_9 ( .a ({key_s1[123], key_s0[123]}), .b ({key_s1[59], key_s0[59]}), .c ({signal_1485, signal_864}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_10 ( .a ({key_s1[122], key_s0[122]}), .b ({key_s1[58], key_s0[58]}), .c ({signal_1488, signal_865}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_11 ( .a ({key_s1[121], key_s0[121]}), .b ({key_s1[57], key_s0[57]}), .c ({signal_1491, signal_866}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_12 ( .a ({key_s1[120], key_s0[120]}), .b ({key_s1[56], key_s0[56]}), .c ({signal_1494, signal_867}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_13 ( .a ({key_s1[119], key_s0[119]}), .b ({key_s1[55], key_s0[55]}), .c ({signal_1497, signal_868}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_14 ( .a ({key_s1[118], key_s0[118]}), .b ({key_s1[54], key_s0[54]}), .c ({signal_1500, signal_869}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_15 ( .a ({key_s1[117], key_s0[117]}), .b ({key_s1[53], key_s0[53]}), .c ({signal_1503, signal_870}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_16 ( .a ({key_s1[116], key_s0[116]}), .b ({key_s1[52], key_s0[52]}), .c ({signal_1506, signal_871}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_17 ( .a ({key_s1[115], key_s0[115]}), .b ({key_s1[51], key_s0[51]}), .c ({signal_1509, signal_872}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_18 ( .a ({key_s1[114], key_s0[114]}), .b ({key_s1[50], key_s0[50]}), .c ({signal_1512, signal_873}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_19 ( .a ({key_s1[4], key_s0[4]}), .b ({key_s1[68], key_s0[68]}), .c ({signal_1515, signal_919}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_20 ( .a ({key_s1[113], key_s0[113]}), .b ({key_s1[49], key_s0[49]}), .c ({signal_1518, signal_874}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_21 ( .a ({key_s1[112], key_s0[112]}), .b ({key_s1[48], key_s0[48]}), .c ({signal_1521, signal_875}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_22 ( .a ({key_s1[111], key_s0[111]}), .b ({key_s1[47], key_s0[47]}), .c ({signal_1524, signal_876}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_23 ( .a ({key_s1[110], key_s0[110]}), .b ({key_s1[46], key_s0[46]}), .c ({signal_1527, signal_877}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_24 ( .a ({key_s1[109], key_s0[109]}), .b ({key_s1[45], key_s0[45]}), .c ({signal_1530, signal_878}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_25 ( .a ({key_s1[108], key_s0[108]}), .b ({key_s1[44], key_s0[44]}), .c ({signal_1533, signal_879}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_26 ( .a ({key_s1[107], key_s0[107]}), .b ({key_s1[43], key_s0[43]}), .c ({signal_1536, signal_880}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_27 ( .a ({key_s1[106], key_s0[106]}), .b ({key_s1[42], key_s0[42]}), .c ({signal_1539, signal_881}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_28 ( .a ({key_s1[105], key_s0[105]}), .b ({key_s1[41], key_s0[41]}), .c ({signal_1542, signal_882}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_29 ( .a ({key_s1[104], key_s0[104]}), .b ({key_s1[40], key_s0[40]}), .c ({signal_1545, signal_883}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_30 ( .a ({key_s1[3], key_s0[3]}), .b ({key_s1[67], key_s0[67]}), .c ({signal_1548, signal_920}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_31 ( .a ({key_s1[103], key_s0[103]}), .b ({key_s1[39], key_s0[39]}), .c ({signal_1551, signal_884}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_32 ( .a ({key_s1[102], key_s0[102]}), .b ({key_s1[38], key_s0[38]}), .c ({signal_1554, signal_885}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_33 ( .a ({key_s1[101], key_s0[101]}), .b ({key_s1[37], key_s0[37]}), .c ({signal_1557, signal_886}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_34 ( .a ({key_s1[100], key_s0[100]}), .b ({key_s1[36], key_s0[36]}), .c ({signal_1560, signal_887}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_35 ( .a ({key_s1[35], key_s0[35]}), .b ({key_s1[99], key_s0[99]}), .c ({signal_1563, signal_888}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_36 ( .a ({key_s1[34], key_s0[34]}), .b ({key_s1[98], key_s0[98]}), .c ({signal_1566, signal_889}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_37 ( .a ({key_s1[33], key_s0[33]}), .b ({key_s1[97], key_s0[97]}), .c ({signal_1569, signal_890}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_38 ( .a ({key_s1[32], key_s0[32]}), .b ({key_s1[96], key_s0[96]}), .c ({signal_1572, signal_891}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_39 ( .a ({key_s1[31], key_s0[31]}), .b ({key_s1[95], key_s0[95]}), .c ({signal_1575, signal_892}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_40 ( .a ({key_s1[30], key_s0[30]}), .b ({key_s1[94], key_s0[94]}), .c ({signal_1578, signal_893}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_41 ( .a ({key_s1[2], key_s0[2]}), .b ({key_s1[66], key_s0[66]}), .c ({signal_1581, signal_921}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_42 ( .a ({key_s1[29], key_s0[29]}), .b ({key_s1[93], key_s0[93]}), .c ({signal_1584, signal_894}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_43 ( .a ({key_s1[28], key_s0[28]}), .b ({key_s1[92], key_s0[92]}), .c ({signal_1587, signal_895}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_44 ( .a ({key_s1[27], key_s0[27]}), .b ({key_s1[91], key_s0[91]}), .c ({signal_1590, signal_896}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_45 ( .a ({key_s1[26], key_s0[26]}), .b ({key_s1[90], key_s0[90]}), .c ({signal_1593, signal_897}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_46 ( .a ({key_s1[25], key_s0[25]}), .b ({key_s1[89], key_s0[89]}), .c ({signal_1596, signal_898}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_47 ( .a ({key_s1[24], key_s0[24]}), .b ({key_s1[88], key_s0[88]}), .c ({signal_1599, signal_899}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_48 ( .a ({key_s1[23], key_s0[23]}), .b ({key_s1[87], key_s0[87]}), .c ({signal_1602, signal_900}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_49 ( .a ({key_s1[22], key_s0[22]}), .b ({key_s1[86], key_s0[86]}), .c ({signal_1605, signal_901}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_50 ( .a ({key_s1[21], key_s0[21]}), .b ({key_s1[85], key_s0[85]}), .c ({signal_1608, signal_902}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_51 ( .a ({key_s1[20], key_s0[20]}), .b ({key_s1[84], key_s0[84]}), .c ({signal_1611, signal_903}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_52 ( .a ({key_s1[1], key_s0[1]}), .b ({key_s1[65], key_s0[65]}), .c ({signal_1614, signal_922}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_53 ( .a ({key_s1[19], key_s0[19]}), .b ({key_s1[83], key_s0[83]}), .c ({signal_1617, signal_904}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_54 ( .a ({key_s1[18], key_s0[18]}), .b ({key_s1[82], key_s0[82]}), .c ({signal_1620, signal_905}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_55 ( .a ({key_s1[17], key_s0[17]}), .b ({key_s1[81], key_s0[81]}), .c ({signal_1623, signal_906}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_56 ( .a ({key_s1[16], key_s0[16]}), .b ({key_s1[80], key_s0[80]}), .c ({signal_1626, signal_907}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_57 ( .a ({key_s1[15], key_s0[15]}), .b ({key_s1[79], key_s0[79]}), .c ({signal_1629, signal_908}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_58 ( .a ({key_s1[14], key_s0[14]}), .b ({key_s1[78], key_s0[78]}), .c ({signal_1632, signal_909}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_59 ( .a ({key_s1[13], key_s0[13]}), .b ({key_s1[77], key_s0[77]}), .c ({signal_1635, signal_910}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_60 ( .a ({key_s1[12], key_s0[12]}), .b ({key_s1[76], key_s0[76]}), .c ({signal_1638, signal_911}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_61 ( .a ({key_s1[11], key_s0[11]}), .b ({key_s1[75], key_s0[75]}), .c ({signal_1641, signal_912}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_62 ( .a ({key_s1[10], key_s0[10]}), .b ({key_s1[74], key_s0[74]}), .c ({signal_1644, signal_913}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_63 ( .a ({key_s1[0], key_s0[0]}), .b ({key_s1[64], key_s0[64]}), .c ({signal_1647, signal_923}) ) ;
    NOR2_X1 cell_64 ( .A1 (signal_266), .A2 (signal_267), .ZN (done) ) ;
    NAND2_X1 cell_65 ( .A1 (signal_927), .A2 (signal_926), .ZN (signal_267) ) ;
    NAND2_X1 cell_66 ( .A1 (signal_925), .A2 (signal_924), .ZN (signal_266) ) ;
    INV_X1 cell_67 ( .A (signal_268), .ZN (signal_278) ) ;
    MUX2_X1 cell_68 ( .S (signal_281), .A (signal_269), .B (signal_270), .Z (signal_268) ) ;
    NOR2_X1 cell_69 ( .A1 (reset), .A2 (signal_271), .ZN (signal_282) ) ;
    XNOR2_X1 cell_70 ( .A (signal_927), .B (signal_926), .ZN (signal_271) ) ;
    MUX2_X1 cell_71 ( .S (signal_924), .A (signal_272), .B (signal_273), .Z (signal_280) ) ;
    NAND2_X1 cell_72 ( .A1 (signal_269), .A2 (signal_274), .ZN (signal_273) ) ;
    NAND2_X1 cell_73 ( .A1 (signal_281), .A2 (signal_277), .ZN (signal_274) ) ;
    NOR2_X1 cell_74 ( .A1 (signal_275), .A2 (signal_283), .ZN (signal_269) ) ;
    NOR2_X1 cell_75 ( .A1 (signal_926), .A2 (reset), .ZN (signal_275) ) ;
    NOR2_X1 cell_76 ( .A1 (signal_281), .A2 (signal_270), .ZN (signal_272) ) ;
    NAND2_X1 cell_77 ( .A1 (signal_926), .A2 (signal_276), .ZN (signal_270) ) ;
    NOR2_X1 cell_78 ( .A1 (reset), .A2 (signal_279), .ZN (signal_276) ) ;
    NOR2_X1 cell_79 ( .A1 (reset), .A2 (signal_927), .ZN (signal_283) ) ;
    INV_X1 cell_80 ( .A (reset), .ZN (signal_277) ) ;
    INV_X1 cell_81 ( .A (signal_927), .ZN (signal_279) ) ;
    INV_X1 cell_85 ( .A (signal_925), .ZN (signal_281) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_153 ( .a ({signal_1458, signal_914}), .b ({DataIn_s1[9], DataIn_s0[9]}), .c ({signal_1662, signal_982}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_154 ( .a ({signal_1461, signal_915}), .b ({DataIn_s1[8], DataIn_s0[8]}), .c ({signal_1664, signal_983}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_155 ( .a ({signal_1464, signal_916}), .b ({DataIn_s1[7], DataIn_s0[7]}), .c ({signal_1666, signal_984}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_156 ( .a ({signal_1467, signal_917}), .b ({DataIn_s1[6], DataIn_s0[6]}), .c ({signal_1668, signal_985}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_157 ( .a ({signal_1470, signal_860}), .b ({DataIn_s1[63], DataIn_s0[63]}), .c ({signal_1670, signal_928}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_158 ( .a ({signal_1473, signal_861}), .b ({DataIn_s1[62], DataIn_s0[62]}), .c ({signal_1672, signal_929}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_159 ( .a ({signal_1476, signal_862}), .b ({DataIn_s1[61], DataIn_s0[61]}), .c ({signal_1674, signal_930}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_160 ( .a ({signal_1479, signal_863}), .b ({DataIn_s1[60], DataIn_s0[60]}), .c ({signal_1676, signal_931}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_161 ( .a ({signal_1482, signal_918}), .b ({DataIn_s1[5], DataIn_s0[5]}), .c ({signal_1678, signal_986}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_162 ( .a ({signal_1485, signal_864}), .b ({DataIn_s1[59], DataIn_s0[59]}), .c ({signal_1680, signal_932}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_163 ( .a ({signal_1488, signal_865}), .b ({DataIn_s1[58], DataIn_s0[58]}), .c ({signal_1682, signal_933}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_164 ( .a ({signal_1491, signal_866}), .b ({DataIn_s1[57], DataIn_s0[57]}), .c ({signal_1684, signal_934}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_165 ( .a ({signal_1494, signal_867}), .b ({DataIn_s1[56], DataIn_s0[56]}), .c ({signal_1686, signal_935}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_166 ( .a ({signal_1497, signal_868}), .b ({DataIn_s1[55], DataIn_s0[55]}), .c ({signal_1688, signal_936}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_167 ( .a ({signal_1500, signal_869}), .b ({DataIn_s1[54], DataIn_s0[54]}), .c ({signal_1690, signal_937}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_168 ( .a ({signal_1503, signal_870}), .b ({DataIn_s1[53], DataIn_s0[53]}), .c ({signal_1692, signal_938}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_169 ( .a ({signal_1506, signal_871}), .b ({DataIn_s1[52], DataIn_s0[52]}), .c ({signal_1694, signal_939}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_170 ( .a ({signal_1509, signal_872}), .b ({DataIn_s1[51], DataIn_s0[51]}), .c ({signal_1696, signal_940}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_171 ( .a ({signal_1512, signal_873}), .b ({DataIn_s1[50], DataIn_s0[50]}), .c ({signal_1698, signal_941}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_172 ( .a ({signal_1515, signal_919}), .b ({DataIn_s1[4], DataIn_s0[4]}), .c ({signal_1700, signal_987}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_173 ( .a ({signal_1518, signal_874}), .b ({DataIn_s1[49], DataIn_s0[49]}), .c ({signal_1702, signal_942}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_174 ( .a ({signal_1521, signal_875}), .b ({DataIn_s1[48], DataIn_s0[48]}), .c ({signal_1704, signal_943}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_175 ( .a ({signal_1524, signal_876}), .b ({DataIn_s1[47], DataIn_s0[47]}), .c ({signal_1706, signal_944}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_176 ( .a ({signal_1527, signal_877}), .b ({DataIn_s1[46], DataIn_s0[46]}), .c ({signal_1708, signal_945}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_177 ( .a ({signal_1530, signal_878}), .b ({DataIn_s1[45], DataIn_s0[45]}), .c ({signal_1710, signal_946}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_178 ( .a ({signal_1533, signal_879}), .b ({DataIn_s1[44], DataIn_s0[44]}), .c ({signal_1712, signal_947}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_179 ( .a ({signal_1536, signal_880}), .b ({DataIn_s1[43], DataIn_s0[43]}), .c ({signal_1714, signal_948}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_180 ( .a ({signal_1539, signal_881}), .b ({DataIn_s1[42], DataIn_s0[42]}), .c ({signal_1716, signal_949}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_181 ( .a ({signal_1542, signal_882}), .b ({DataIn_s1[41], DataIn_s0[41]}), .c ({signal_1718, signal_950}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_182 ( .a ({signal_1545, signal_883}), .b ({DataIn_s1[40], DataIn_s0[40]}), .c ({signal_1720, signal_951}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_183 ( .a ({signal_1548, signal_920}), .b ({DataIn_s1[3], DataIn_s0[3]}), .c ({signal_1722, signal_988}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_184 ( .a ({signal_1551, signal_884}), .b ({DataIn_s1[39], DataIn_s0[39]}), .c ({signal_1724, signal_952}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_185 ( .a ({signal_1554, signal_885}), .b ({DataIn_s1[38], DataIn_s0[38]}), .c ({signal_1726, signal_953}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_186 ( .a ({signal_1557, signal_886}), .b ({DataIn_s1[37], DataIn_s0[37]}), .c ({signal_1728, signal_954}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_187 ( .a ({signal_1560, signal_887}), .b ({DataIn_s1[36], DataIn_s0[36]}), .c ({signal_1730, signal_955}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_188 ( .a ({signal_1563, signal_888}), .b ({DataIn_s1[35], DataIn_s0[35]}), .c ({signal_1732, signal_956}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_189 ( .a ({signal_1566, signal_889}), .b ({DataIn_s1[34], DataIn_s0[34]}), .c ({signal_1734, signal_957}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_190 ( .a ({signal_1569, signal_890}), .b ({DataIn_s1[33], DataIn_s0[33]}), .c ({signal_1736, signal_958}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_191 ( .a ({signal_1572, signal_891}), .b ({DataIn_s1[32], DataIn_s0[32]}), .c ({signal_1738, signal_959}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_192 ( .a ({signal_1575, signal_892}), .b ({DataIn_s1[31], DataIn_s0[31]}), .c ({signal_1740, signal_960}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_193 ( .a ({signal_1578, signal_893}), .b ({DataIn_s1[30], DataIn_s0[30]}), .c ({signal_1742, signal_961}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_194 ( .a ({signal_1581, signal_921}), .b ({DataIn_s1[2], DataIn_s0[2]}), .c ({signal_1744, signal_989}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_195 ( .a ({signal_1584, signal_894}), .b ({DataIn_s1[29], DataIn_s0[29]}), .c ({signal_1746, signal_962}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_196 ( .a ({signal_1587, signal_895}), .b ({DataIn_s1[28], DataIn_s0[28]}), .c ({signal_1748, signal_963}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_197 ( .a ({signal_1590, signal_896}), .b ({DataIn_s1[27], DataIn_s0[27]}), .c ({signal_1750, signal_964}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_198 ( .a ({signal_1593, signal_897}), .b ({DataIn_s1[26], DataIn_s0[26]}), .c ({signal_1752, signal_965}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_199 ( .a ({signal_1596, signal_898}), .b ({DataIn_s1[25], DataIn_s0[25]}), .c ({signal_1754, signal_966}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_200 ( .a ({signal_1599, signal_899}), .b ({DataIn_s1[24], DataIn_s0[24]}), .c ({signal_1756, signal_967}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_201 ( .a ({signal_1602, signal_900}), .b ({DataIn_s1[23], DataIn_s0[23]}), .c ({signal_1758, signal_968}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_202 ( .a ({signal_1605, signal_901}), .b ({DataIn_s1[22], DataIn_s0[22]}), .c ({signal_1760, signal_969}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_203 ( .a ({signal_1608, signal_902}), .b ({DataIn_s1[21], DataIn_s0[21]}), .c ({signal_1762, signal_970}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_204 ( .a ({signal_1611, signal_903}), .b ({DataIn_s1[20], DataIn_s0[20]}), .c ({signal_1764, signal_971}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_205 ( .a ({signal_1614, signal_922}), .b ({DataIn_s1[1], DataIn_s0[1]}), .c ({signal_1766, signal_990}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_206 ( .a ({signal_1617, signal_904}), .b ({DataIn_s1[19], DataIn_s0[19]}), .c ({signal_1768, signal_972}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_207 ( .a ({signal_1620, signal_905}), .b ({DataIn_s1[18], DataIn_s0[18]}), .c ({signal_1770, signal_973}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_208 ( .a ({signal_1623, signal_906}), .b ({DataIn_s1[17], DataIn_s0[17]}), .c ({signal_1772, signal_974}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_209 ( .a ({signal_1626, signal_907}), .b ({DataIn_s1[16], DataIn_s0[16]}), .c ({signal_1774, signal_975}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_210 ( .a ({signal_1629, signal_908}), .b ({DataIn_s1[15], DataIn_s0[15]}), .c ({signal_1776, signal_976}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_211 ( .a ({signal_1632, signal_909}), .b ({DataIn_s1[14], DataIn_s0[14]}), .c ({signal_1778, signal_977}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_212 ( .a ({signal_1635, signal_910}), .b ({DataIn_s1[13], DataIn_s0[13]}), .c ({signal_1780, signal_978}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_213 ( .a ({signal_1638, signal_911}), .b ({DataIn_s1[12], DataIn_s0[12]}), .c ({signal_1782, signal_979}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_214 ( .a ({signal_1641, signal_912}), .b ({DataIn_s1[11], DataIn_s0[11]}), .c ({signal_1784, signal_980}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_215 ( .a ({signal_1644, signal_913}), .b ({DataIn_s1[10], DataIn_s0[10]}), .c ({signal_1786, signal_981}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_216 ( .a ({signal_1647, signal_923}), .b ({DataIn_s1[0], DataIn_s0[0]}), .c ({signal_1788, signal_991}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_283 ( .a ({signal_1653, signal_310}), .b ({1'b0, signal_1453}), .c ({signal_2254, signal_286}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_290 ( .a ({signal_2038, signal_362}), .b ({1'b0, signal_1440}), .c ({signal_2310, signal_287}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_296 ( .a ({signal_2034, signal_358}), .b ({1'b0, signal_1441}), .c ({signal_2311, signal_288}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_301 ( .a ({signal_2030, signal_354}), .b ({1'b0, signal_1442}), .c ({signal_2312, signal_289}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_305 ( .a ({signal_1652, signal_306}), .b ({1'b0, signal_1454}), .c ({signal_2313, signal_290}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_308 ( .a ({signal_2026, signal_350}), .b ({1'b0, signal_1443}), .c ({signal_2378, signal_291}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_313 ( .a ({signal_2022, signal_346}), .b ({1'b0, signal_1444}), .c ({signal_2255, signal_292}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_318 ( .a ({signal_2018, signal_342}), .b ({1'b0, signal_1445}), .c ({signal_2314, signal_293}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_324 ( .a ({signal_2014, signal_338}), .b ({1'b0, signal_1446}), .c ({signal_2256, signal_294}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_329 ( .a ({signal_2010, signal_334}), .b ({1'b0, signal_1447}), .c ({signal_2315, signal_295}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_335 ( .a ({signal_2006, signal_330}), .b ({1'b0, signal_1448}), .c ({signal_2372, signal_296}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_340 ( .a ({signal_2003, signal_326}), .b ({1'b0, signal_1449}), .c ({signal_2316, signal_297}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_345 ( .a ({signal_1999, signal_322}), .b ({1'b0, signal_1450}), .c ({signal_2257, signal_298}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_351 ( .a ({signal_1995, signal_318}), .b ({1'b0, signal_1451}), .c ({signal_2317, signal_299}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_356 ( .a ({signal_1994, signal_314}), .b ({1'b0, signal_1452}), .c ({signal_2318, signal_300}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_360 ( .a ({signal_1648, signal_302}), .b ({1'b0, signal_1455}), .c ({signal_2319, signal_301}) ) ;
    NAND2_X1 cell_361 ( .A1 (signal_366), .A2 (signal_367), .ZN (signal_1446) ) ;
    NOR2_X1 cell_362 ( .A1 (signal_368), .A2 (signal_369), .ZN (signal_366) ) ;
    OR2_X1 cell_363 ( .A1 (signal_370), .A2 (signal_371), .ZN (signal_369) ) ;
    NAND2_X1 cell_364 ( .A1 (signal_372), .A2 (signal_373), .ZN (signal_1447) ) ;
    NAND2_X1 cell_365 ( .A1 (signal_374), .A2 (signal_375), .ZN (signal_1448) ) ;
    NOR2_X1 cell_366 ( .A1 (signal_1444), .A2 (signal_376), .ZN (signal_375) ) ;
    NAND2_X1 cell_367 ( .A1 (signal_377), .A2 (signal_378), .ZN (signal_376) ) ;
    NOR2_X1 cell_368 ( .A1 (signal_379), .A2 (signal_380), .ZN (signal_377) ) ;
    NAND2_X1 cell_369 ( .A1 (signal_381), .A2 (signal_382), .ZN (signal_1449) ) ;
    NOR2_X1 cell_370 ( .A1 (signal_383), .A2 (signal_384), .ZN (signal_382) ) ;
    NAND2_X1 cell_371 ( .A1 (signal_385), .A2 (signal_386), .ZN (signal_1450) ) ;
    NOR2_X1 cell_372 ( .A1 (signal_371), .A2 (signal_387), .ZN (signal_386) ) ;
    NAND2_X1 cell_373 ( .A1 (signal_388), .A2 (signal_378), .ZN (signal_387) ) ;
    NAND2_X1 cell_374 ( .A1 (signal_389), .A2 (signal_388), .ZN (signal_1451) ) ;
    NOR2_X1 cell_375 ( .A1 (signal_390), .A2 (signal_391), .ZN (signal_388) ) ;
    NAND2_X1 cell_376 ( .A1 (signal_392), .A2 (signal_393), .ZN (signal_1452) ) ;
    NOR2_X1 cell_377 ( .A1 (signal_368), .A2 (signal_394), .ZN (signal_392) ) ;
    NAND2_X1 cell_378 ( .A1 (signal_395), .A2 (signal_378), .ZN (signal_394) ) ;
    INV_X1 cell_379 ( .A (signal_396), .ZN (signal_395) ) ;
    OR2_X1 cell_380 ( .A1 (signal_368), .A2 (signal_397), .ZN (signal_1453) ) ;
    NAND2_X1 cell_381 ( .A1 (signal_381), .A2 (signal_398), .ZN (signal_397) ) ;
    NOR2_X1 cell_382 ( .A1 (signal_399), .A2 (signal_371), .ZN (signal_381) ) ;
    NAND2_X1 cell_383 ( .A1 (signal_400), .A2 (signal_373), .ZN (signal_368) ) ;
    NAND2_X1 cell_384 ( .A1 (signal_401), .A2 (signal_402), .ZN (signal_1454) ) ;
    NOR2_X1 cell_385 ( .A1 (signal_396), .A2 (signal_403), .ZN (signal_402) ) ;
    OR2_X1 cell_386 ( .A1 (signal_371), .A2 (signal_379), .ZN (signal_403) ) ;
    INV_X1 cell_387 ( .A (signal_400), .ZN (signal_379) ) ;
    NAND2_X1 cell_388 ( .A1 (signal_404), .A2 (signal_405), .ZN (signal_400) ) ;
    NAND2_X1 cell_389 ( .A1 (signal_406), .A2 (signal_407), .ZN (signal_405) ) ;
    NOR2_X1 cell_390 ( .A1 (signal_455), .A2 (signal_408), .ZN (signal_371) ) ;
    MUX2_X1 cell_391 ( .S (signal_925), .A (signal_409), .B (signal_410), .Z (signal_408) ) ;
    NAND2_X1 cell_392 ( .A1 (signal_411), .A2 (signal_412), .ZN (signal_1440) ) ;
    NOR2_X1 cell_393 ( .A1 (signal_383), .A2 (signal_396), .ZN (signal_411) ) ;
    NAND2_X1 cell_394 ( .A1 (signal_413), .A2 (signal_389), .ZN (signal_1441) ) ;
    NOR2_X1 cell_395 ( .A1 (signal_414), .A2 (signal_415), .ZN (signal_389) ) ;
    NAND2_X1 cell_396 ( .A1 (signal_367), .A2 (signal_378), .ZN (signal_415) ) ;
    OR2_X1 cell_397 ( .A1 (signal_454), .A2 (signal_416), .ZN (signal_378) ) ;
    MUX2_X1 cell_398 ( .S (signal_925), .A (signal_417), .B (signal_418), .Z (signal_416) ) ;
    NAND2_X1 cell_399 ( .A1 (signal_398), .A2 (signal_419), .ZN (signal_1442) ) ;
    NOR2_X1 cell_400 ( .A1 (signal_420), .A2 (signal_421), .ZN (signal_419) ) ;
    INV_X1 cell_401 ( .A (signal_413), .ZN (signal_421) ) ;
    NOR2_X1 cell_402 ( .A1 (signal_422), .A2 (signal_391), .ZN (signal_398) ) ;
    NAND2_X1 cell_403 ( .A1 (signal_423), .A2 (signal_393), .ZN (signal_1443) ) ;
    INV_X1 cell_404 ( .A (signal_399), .ZN (signal_393) ) ;
    NOR2_X1 cell_405 ( .A1 (signal_380), .A2 (signal_424), .ZN (signal_423) ) ;
    NAND2_X1 cell_406 ( .A1 (signal_372), .A2 (signal_413), .ZN (signal_424) ) ;
    NOR2_X1 cell_407 ( .A1 (signal_390), .A2 (signal_414), .ZN (signal_372) ) ;
    NAND2_X1 cell_408 ( .A1 (signal_385), .A2 (signal_425), .ZN (signal_414) ) ;
    NAND2_X1 cell_409 ( .A1 (signal_454), .A2 (signal_426), .ZN (signal_425) ) ;
    NAND2_X1 cell_410 ( .A1 (signal_418), .A2 (signal_406), .ZN (signal_426) ) ;
    NOR2_X1 cell_411 ( .A1 (signal_383), .A2 (signal_427), .ZN (signal_385) ) ;
    NOR2_X1 cell_412 ( .A1 (signal_455), .A2 (signal_428), .ZN (signal_427) ) ;
    MUX2_X1 cell_413 ( .S (signal_925), .A (signal_407), .B (signal_417), .Z (signal_428) ) ;
    NOR2_X1 cell_414 ( .A1 (signal_454), .A2 (signal_429), .ZN (signal_383) ) ;
    MUX2_X1 cell_415 ( .S (signal_925), .A (signal_409), .B (signal_430), .Z (signal_429) ) ;
    OR2_X1 cell_416 ( .A1 (signal_384), .A2 (signal_370), .ZN (signal_1444) ) ;
    NAND2_X1 cell_417 ( .A1 (signal_413), .A2 (signal_373), .ZN (signal_384) ) ;
    NAND2_X1 cell_418 ( .A1 (signal_431), .A2 (signal_432), .ZN (signal_373) ) ;
    AND2_X1 cell_419 ( .A1 (signal_455), .A2 (signal_925), .ZN (signal_432) ) ;
    NOR2_X1 cell_420 ( .A1 (signal_433), .A2 (signal_396), .ZN (signal_413) ) ;
    NOR2_X1 cell_421 ( .A1 (signal_454), .A2 (signal_434), .ZN (signal_396) ) ;
    MUX2_X1 cell_422 ( .S (signal_925), .A (signal_418), .B (signal_417), .Z (signal_434) ) ;
    NOR2_X1 cell_423 ( .A1 (signal_454), .A2 (signal_435), .ZN (signal_433) ) ;
    MUX2_X1 cell_424 ( .S (signal_925), .A (signal_430), .B (signal_409), .Z (signal_435) ) ;
    NAND2_X1 cell_425 ( .A1 (signal_436), .A2 (signal_412), .ZN (signal_1445) ) ;
    NOR2_X1 cell_426 ( .A1 (signal_437), .A2 (signal_370), .ZN (signal_412) ) ;
    NOR2_X1 cell_427 ( .A1 (signal_455), .A2 (signal_438), .ZN (signal_370) ) ;
    MUX2_X1 cell_428 ( .S (signal_925), .A (signal_418), .B (signal_406), .Z (signal_438) ) ;
    INV_X1 cell_429 ( .A (signal_439), .ZN (signal_437) ) ;
    INV_X1 cell_430 ( .A (signal_390), .ZN (signal_436) ) ;
    NAND2_X1 cell_431 ( .A1 (signal_401), .A2 (signal_439), .ZN (signal_1455) ) ;
    NOR2_X1 cell_432 ( .A1 (signal_380), .A2 (signal_391), .ZN (signal_439) ) ;
    NOR2_X1 cell_433 ( .A1 (signal_455), .A2 (signal_440), .ZN (signal_391) ) ;
    MUX2_X1 cell_434 ( .S (signal_925), .A (signal_410), .B (signal_409), .Z (signal_440) ) ;
    NAND2_X1 cell_435 ( .A1 (signal_441), .A2 (signal_442), .ZN (signal_409) ) ;
    NAND2_X1 cell_436 ( .A1 (signal_443), .A2 (signal_926), .ZN (signal_410) ) ;
    NOR2_X1 cell_437 ( .A1 (signal_455), .A2 (signal_444), .ZN (signal_380) ) ;
    MUX2_X1 cell_438 ( .S (signal_925), .A (signal_417), .B (signal_407), .Z (signal_444) ) ;
    NAND2_X1 cell_439 ( .A1 (enc_dec), .A2 (signal_431), .ZN (signal_407) ) ;
    NOR2_X1 cell_440 ( .A1 (signal_924), .A2 (signal_442), .ZN (signal_431) ) ;
    NAND2_X1 cell_441 ( .A1 (signal_445), .A2 (signal_442), .ZN (signal_417) ) ;
    NOR2_X1 cell_442 ( .A1 (signal_399), .A2 (signal_446), .ZN (signal_401) ) ;
    NAND2_X1 cell_443 ( .A1 (signal_374), .A2 (signal_367), .ZN (signal_446) ) ;
    NAND2_X1 cell_444 ( .A1 (signal_420), .A2 (signal_447), .ZN (signal_367) ) ;
    OR2_X1 cell_445 ( .A1 (signal_443), .A2 (signal_441), .ZN (signal_447) ) ;
    AND2_X1 cell_446 ( .A1 (signal_926), .A2 (signal_404), .ZN (signal_420) ) ;
    NOR2_X1 cell_447 ( .A1 (signal_454), .A2 (signal_925), .ZN (signal_404) ) ;
    NOR2_X1 cell_448 ( .A1 (signal_390), .A2 (signal_422), .ZN (signal_374) ) ;
    NOR2_X1 cell_449 ( .A1 (signal_455), .A2 (signal_448), .ZN (signal_422) ) ;
    MUX2_X1 cell_450 ( .S (signal_925), .A (signal_406), .B (signal_418), .Z (signal_448) ) ;
    NAND2_X1 cell_451 ( .A1 (enc_dec), .A2 (signal_449), .ZN (signal_418) ) ;
    NOR2_X1 cell_452 ( .A1 (signal_924), .A2 (signal_926), .ZN (signal_449) ) ;
    NAND2_X1 cell_453 ( .A1 (signal_926), .A2 (signal_445), .ZN (signal_406) ) ;
    NOR2_X1 cell_454 ( .A1 (enc_dec), .A2 (signal_450), .ZN (signal_445) ) ;
    INV_X1 cell_455 ( .A (signal_924), .ZN (signal_450) ) ;
    NOR2_X1 cell_456 ( .A1 (signal_455), .A2 (signal_451), .ZN (signal_390) ) ;
    MUX2_X1 cell_457 ( .S (signal_925), .A (signal_430), .B (signal_452), .Z (signal_451) ) ;
    NOR2_X1 cell_458 ( .A1 (signal_455), .A2 (signal_453), .ZN (signal_399) ) ;
    MUX2_X1 cell_459 ( .S (signal_925), .A (signal_452), .B (signal_430), .Z (signal_453) ) ;
    NAND2_X1 cell_460 ( .A1 (signal_443), .A2 (signal_442), .ZN (signal_430) ) ;
    INV_X1 cell_461 ( .A (signal_926), .ZN (signal_442) ) ;
    NOR2_X1 cell_462 ( .A1 (enc_dec), .A2 (signal_924), .ZN (signal_443) ) ;
    NAND2_X1 cell_463 ( .A1 (signal_441), .A2 (signal_926), .ZN (signal_452) ) ;
    AND2_X1 cell_464 ( .A1 (enc_dec), .A2 (signal_924), .ZN (signal_441) ) ;
    INV_X1 cell_465 ( .A (signal_454), .ZN (signal_455) ) ;
    INV_X1 cell_466 ( .A (signal_927), .ZN (signal_454) ) ;
    INV_X1 cell_467 ( .A (signal_927), .ZN (signal_456) ) ;
    INV_X1 cell_468 ( .A (signal_456), .ZN (signal_459) ) ;
    INV_X1 cell_469 ( .A (signal_456), .ZN (signal_458) ) ;
    INV_X1 cell_470 ( .A (signal_456), .ZN (signal_457) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_471 ( .s (signal_927), .b ({key_s1[64], key_s0[64]}), .a ({key_s1[0], key_s0[0]}), .c ({signal_1648, signal_302}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_472 ( .s (signal_927), .b ({key_s1[65], key_s0[65]}), .a ({key_s1[1], key_s0[1]}), .c ({signal_1649, signal_303}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_473 ( .s (signal_927), .b ({key_s1[66], key_s0[66]}), .a ({key_s1[2], key_s0[2]}), .c ({signal_1650, signal_304}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_474 ( .s (signal_927), .b ({key_s1[67], key_s0[67]}), .a ({key_s1[3], key_s0[3]}), .c ({signal_1651, signal_305}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_475 ( .s (signal_927), .b ({key_s1[68], key_s0[68]}), .a ({key_s1[4], key_s0[4]}), .c ({signal_1652, signal_306}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_476 ( .s (signal_459), .b ({key_s1[69], key_s0[69]}), .a ({key_s1[5], key_s0[5]}), .c ({signal_1991, signal_307}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_477 ( .s (signal_457), .b ({key_s1[70], key_s0[70]}), .a ({key_s1[6], key_s0[6]}), .c ({signal_1992, signal_308}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_478 ( .s (signal_458), .b ({key_s1[71], key_s0[71]}), .a ({key_s1[7], key_s0[7]}), .c ({signal_1993, signal_309}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_479 ( .s (signal_927), .b ({key_s1[72], key_s0[72]}), .a ({key_s1[8], key_s0[8]}), .c ({signal_1653, signal_310}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_480 ( .s (signal_927), .b ({key_s1[73], key_s0[73]}), .a ({key_s1[9], key_s0[9]}), .c ({signal_1654, signal_311}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_481 ( .s (signal_927), .b ({key_s1[74], key_s0[74]}), .a ({key_s1[10], key_s0[10]}), .c ({signal_1655, signal_312}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_482 ( .s (signal_927), .b ({key_s1[75], key_s0[75]}), .a ({key_s1[11], key_s0[11]}), .c ({signal_1656, signal_313}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_483 ( .s (signal_458), .b ({key_s1[76], key_s0[76]}), .a ({key_s1[12], key_s0[12]}), .c ({signal_1994, signal_314}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_484 ( .s (signal_927), .b ({key_s1[77], key_s0[77]}), .a ({key_s1[13], key_s0[13]}), .c ({signal_1657, signal_315}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_485 ( .s (signal_927), .b ({key_s1[78], key_s0[78]}), .a ({key_s1[14], key_s0[14]}), .c ({signal_1658, signal_316}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_486 ( .s (signal_927), .b ({key_s1[79], key_s0[79]}), .a ({key_s1[15], key_s0[15]}), .c ({signal_1659, signal_317}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_487 ( .s (signal_457), .b ({key_s1[80], key_s0[80]}), .a ({key_s1[16], key_s0[16]}), .c ({signal_1995, signal_318}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_488 ( .s (signal_459), .b ({key_s1[81], key_s0[81]}), .a ({key_s1[17], key_s0[17]}), .c ({signal_1996, signal_319}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_489 ( .s (signal_457), .b ({key_s1[82], key_s0[82]}), .a ({key_s1[18], key_s0[18]}), .c ({signal_1997, signal_320}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_490 ( .s (signal_457), .b ({key_s1[83], key_s0[83]}), .a ({key_s1[19], key_s0[19]}), .c ({signal_1998, signal_321}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_491 ( .s (signal_457), .b ({key_s1[84], key_s0[84]}), .a ({key_s1[20], key_s0[20]}), .c ({signal_1999, signal_322}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_492 ( .s (signal_457), .b ({key_s1[85], key_s0[85]}), .a ({key_s1[21], key_s0[21]}), .c ({signal_2000, signal_323}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_493 ( .s (signal_458), .b ({key_s1[86], key_s0[86]}), .a ({key_s1[22], key_s0[22]}), .c ({signal_2001, signal_324}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_494 ( .s (signal_459), .b ({key_s1[87], key_s0[87]}), .a ({key_s1[23], key_s0[23]}), .c ({signal_2002, signal_325}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_495 ( .s (signal_457), .b ({key_s1[88], key_s0[88]}), .a ({key_s1[24], key_s0[24]}), .c ({signal_2003, signal_326}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_496 ( .s (signal_458), .b ({key_s1[89], key_s0[89]}), .a ({key_s1[25], key_s0[25]}), .c ({signal_2004, signal_327}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_497 ( .s (signal_927), .b ({key_s1[90], key_s0[90]}), .a ({key_s1[26], key_s0[26]}), .c ({signal_1660, signal_328}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_498 ( .s (signal_457), .b ({key_s1[91], key_s0[91]}), .a ({key_s1[27], key_s0[27]}), .c ({signal_2005, signal_329}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_499 ( .s (signal_457), .b ({key_s1[92], key_s0[92]}), .a ({key_s1[28], key_s0[28]}), .c ({signal_2006, signal_330}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_500 ( .s (signal_457), .b ({key_s1[93], key_s0[93]}), .a ({key_s1[29], key_s0[29]}), .c ({signal_2007, signal_331}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_501 ( .s (signal_457), .b ({key_s1[94], key_s0[94]}), .a ({key_s1[30], key_s0[30]}), .c ({signal_2008, signal_332}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_502 ( .s (signal_457), .b ({key_s1[95], key_s0[95]}), .a ({key_s1[31], key_s0[31]}), .c ({signal_2009, signal_333}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_503 ( .s (signal_457), .b ({key_s1[96], key_s0[96]}), .a ({key_s1[32], key_s0[32]}), .c ({signal_2010, signal_334}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_504 ( .s (signal_457), .b ({key_s1[97], key_s0[97]}), .a ({key_s1[33], key_s0[33]}), .c ({signal_2011, signal_335}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_505 ( .s (signal_457), .b ({key_s1[98], key_s0[98]}), .a ({key_s1[34], key_s0[34]}), .c ({signal_2012, signal_336}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_506 ( .s (signal_457), .b ({key_s1[99], key_s0[99]}), .a ({key_s1[35], key_s0[35]}), .c ({signal_2013, signal_337}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_507 ( .s (signal_457), .b ({key_s1[100], key_s0[100]}), .a ({key_s1[36], key_s0[36]}), .c ({signal_2014, signal_338}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_508 ( .s (signal_457), .b ({key_s1[101], key_s0[101]}), .a ({key_s1[37], key_s0[37]}), .c ({signal_2015, signal_339}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_509 ( .s (signal_457), .b ({key_s1[102], key_s0[102]}), .a ({key_s1[38], key_s0[38]}), .c ({signal_2016, signal_340}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_510 ( .s (signal_457), .b ({key_s1[103], key_s0[103]}), .a ({key_s1[39], key_s0[39]}), .c ({signal_2017, signal_341}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_511 ( .s (signal_458), .b ({key_s1[104], key_s0[104]}), .a ({key_s1[40], key_s0[40]}), .c ({signal_2018, signal_342}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_512 ( .s (signal_458), .b ({key_s1[105], key_s0[105]}), .a ({key_s1[41], key_s0[41]}), .c ({signal_2019, signal_343}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_513 ( .s (signal_458), .b ({key_s1[106], key_s0[106]}), .a ({key_s1[42], key_s0[42]}), .c ({signal_2020, signal_344}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_514 ( .s (signal_458), .b ({key_s1[107], key_s0[107]}), .a ({key_s1[43], key_s0[43]}), .c ({signal_2021, signal_345}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_515 ( .s (signal_458), .b ({key_s1[108], key_s0[108]}), .a ({key_s1[44], key_s0[44]}), .c ({signal_2022, signal_346}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_516 ( .s (signal_458), .b ({key_s1[109], key_s0[109]}), .a ({key_s1[45], key_s0[45]}), .c ({signal_2023, signal_347}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_517 ( .s (signal_458), .b ({key_s1[110], key_s0[110]}), .a ({key_s1[46], key_s0[46]}), .c ({signal_2024, signal_348}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_518 ( .s (signal_458), .b ({key_s1[111], key_s0[111]}), .a ({key_s1[47], key_s0[47]}), .c ({signal_2025, signal_349}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_519 ( .s (signal_458), .b ({key_s1[112], key_s0[112]}), .a ({key_s1[48], key_s0[48]}), .c ({signal_2026, signal_350}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_520 ( .s (signal_458), .b ({key_s1[113], key_s0[113]}), .a ({key_s1[49], key_s0[49]}), .c ({signal_2027, signal_351}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_521 ( .s (signal_458), .b ({key_s1[114], key_s0[114]}), .a ({key_s1[50], key_s0[50]}), .c ({signal_2028, signal_352}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_522 ( .s (signal_458), .b ({key_s1[115], key_s0[115]}), .a ({key_s1[51], key_s0[51]}), .c ({signal_2029, signal_353}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_523 ( .s (signal_459), .b ({key_s1[116], key_s0[116]}), .a ({key_s1[52], key_s0[52]}), .c ({signal_2030, signal_354}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_524 ( .s (signal_459), .b ({key_s1[117], key_s0[117]}), .a ({key_s1[53], key_s0[53]}), .c ({signal_2031, signal_355}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_525 ( .s (signal_459), .b ({key_s1[118], key_s0[118]}), .a ({key_s1[54], key_s0[54]}), .c ({signal_2032, signal_356}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_526 ( .s (signal_459), .b ({key_s1[119], key_s0[119]}), .a ({key_s1[55], key_s0[55]}), .c ({signal_2033, signal_357}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_527 ( .s (signal_459), .b ({key_s1[120], key_s0[120]}), .a ({key_s1[56], key_s0[56]}), .c ({signal_2034, signal_358}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_528 ( .s (signal_459), .b ({key_s1[121], key_s0[121]}), .a ({key_s1[57], key_s0[57]}), .c ({signal_2035, signal_359}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_529 ( .s (signal_459), .b ({key_s1[122], key_s0[122]}), .a ({key_s1[58], key_s0[58]}), .c ({signal_2036, signal_360}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_530 ( .s (signal_459), .b ({key_s1[123], key_s0[123]}), .a ({key_s1[59], key_s0[59]}), .c ({signal_2037, signal_361}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_531 ( .s (signal_459), .b ({key_s1[124], key_s0[124]}), .a ({key_s1[60], key_s0[60]}), .c ({signal_2038, signal_362}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_532 ( .s (signal_459), .b ({key_s1[125], key_s0[125]}), .a ({key_s1[61], key_s0[61]}), .c ({signal_2039, signal_363}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_533 ( .s (signal_459), .b ({key_s1[126], key_s0[126]}), .a ({key_s1[62], key_s0[62]}), .c ({signal_2040, signal_364}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_534 ( .s (signal_459), .b ({key_s1[127], key_s0[127]}), .a ({key_s1[63], key_s0[63]}), .c ({signal_2041, signal_365}) ) ;
    ClockGatingController #(3) cell_1256 ( .clk (clk), .rst (reset), .GatedClk (signal_2528), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_89 ( .a ({signal_1458, signal_914}), .b ({signal_1907, signal_1302}), .c ({DataOut_s1[9], DataOut_s0[9]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_90 ( .a ({signal_1461, signal_915}), .b ({signal_1908, signal_1303}), .c ({DataOut_s1[8], DataOut_s0[8]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_91 ( .a ({signal_1464, signal_916}), .b ({signal_1869, signal_1264}), .c ({DataOut_s1[7], DataOut_s0[7]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_92 ( .a ({signal_1467, signal_917}), .b ({signal_1870, signal_1265}), .c ({DataOut_s1[6], DataOut_s0[6]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_93 ( .a ({signal_1470, signal_860}), .b ({signal_1853, signal_1248}), .c ({DataOut_s1[63], DataOut_s0[63]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_94 ( .a ({signal_1473, signal_861}), .b ({signal_1854, signal_1249}), .c ({DataOut_s1[62], DataOut_s0[62]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_95 ( .a ({signal_1476, signal_862}), .b ({signal_1855, signal_1250}), .c ({DataOut_s1[61], DataOut_s0[61]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_96 ( .a ({signal_1479, signal_863}), .b ({signal_1856, signal_1251}), .c ({DataOut_s1[60], DataOut_s0[60]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_97 ( .a ({signal_1482, signal_918}), .b ({signal_1871, signal_1266}), .c ({DataOut_s1[5], DataOut_s0[5]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_98 ( .a ({signal_1485, signal_864}), .b ({signal_1881, signal_1276}), .c ({DataOut_s1[59], DataOut_s0[59]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_99 ( .a ({signal_1488, signal_865}), .b ({signal_1882, signal_1277}), .c ({DataOut_s1[58], DataOut_s0[58]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_100 ( .a ({signal_1491, signal_866}), .b ({signal_1883, signal_1278}), .c ({DataOut_s1[57], DataOut_s0[57]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_101 ( .a ({signal_1494, signal_867}), .b ({signal_1884, signal_1279}), .c ({DataOut_s1[56], DataOut_s0[56]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_102 ( .a ({signal_1497, signal_868}), .b ({signal_1909, signal_1304}), .c ({DataOut_s1[55], DataOut_s0[55]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_103 ( .a ({signal_1500, signal_869}), .b ({signal_1910, signal_1305}), .c ({DataOut_s1[54], DataOut_s0[54]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_104 ( .a ({signal_1503, signal_870}), .b ({signal_1911, signal_1306}), .c ({DataOut_s1[53], DataOut_s0[53]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_105 ( .a ({signal_1506, signal_871}), .b ({signal_1912, signal_1307}), .c ({DataOut_s1[52], DataOut_s0[52]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_106 ( .a ({signal_1509, signal_872}), .b ({signal_1889, signal_1284}), .c ({DataOut_s1[51], DataOut_s0[51]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_107 ( .a ({signal_1512, signal_873}), .b ({signal_1890, signal_1285}), .c ({DataOut_s1[50], DataOut_s0[50]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_108 ( .a ({signal_1515, signal_919}), .b ({signal_1872, signal_1267}), .c ({DataOut_s1[4], DataOut_s0[4]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_109 ( .a ({signal_1518, signal_874}), .b ({signal_1891, signal_1286}), .c ({DataOut_s1[49], DataOut_s0[49]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_110 ( .a ({signal_1521, signal_875}), .b ({signal_1892, signal_1287}), .c ({DataOut_s1[48], DataOut_s0[48]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_111 ( .a ({signal_1524, signal_876}), .b ({signal_1873, signal_1268}), .c ({DataOut_s1[47], DataOut_s0[47]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_112 ( .a ({signal_1527, signal_877}), .b ({signal_1874, signal_1269}), .c ({DataOut_s1[46], DataOut_s0[46]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_113 ( .a ({signal_1530, signal_878}), .b ({signal_1875, signal_1270}), .c ({DataOut_s1[45], DataOut_s0[45]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_114 ( .a ({signal_1533, signal_879}), .b ({signal_1876, signal_1271}), .c ({DataOut_s1[44], DataOut_s0[44]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_115 ( .a ({signal_1536, signal_880}), .b ({signal_1861, signal_1256}), .c ({DataOut_s1[43], DataOut_s0[43]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_116 ( .a ({signal_1539, signal_881}), .b ({signal_1862, signal_1257}), .c ({DataOut_s1[42], DataOut_s0[42]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_117 ( .a ({signal_1542, signal_882}), .b ({signal_1863, signal_1258}), .c ({DataOut_s1[41], DataOut_s0[41]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_118 ( .a ({signal_1545, signal_883}), .b ({signal_1864, signal_1259}), .c ({DataOut_s1[40], DataOut_s0[40]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_119 ( .a ({signal_1548, signal_920}), .b ({signal_1865, signal_1260}), .c ({DataOut_s1[3], DataOut_s0[3]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_120 ( .a ({signal_1551, signal_884}), .b ({signal_1897, signal_1292}), .c ({DataOut_s1[39], DataOut_s0[39]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_121 ( .a ({signal_1554, signal_885}), .b ({signal_1898, signal_1293}), .c ({DataOut_s1[38], DataOut_s0[38]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_122 ( .a ({signal_1557, signal_886}), .b ({signal_1899, signal_1294}), .c ({DataOut_s1[37], DataOut_s0[37]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_123 ( .a ({signal_1560, signal_887}), .b ({signal_1900, signal_1295}), .c ({DataOut_s1[36], DataOut_s0[36]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_124 ( .a ({signal_1563, signal_888}), .b ({signal_1901, signal_1296}), .c ({DataOut_s1[35], DataOut_s0[35]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_125 ( .a ({signal_1566, signal_889}), .b ({signal_1902, signal_1297}), .c ({DataOut_s1[34], DataOut_s0[34]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_126 ( .a ({signal_1569, signal_890}), .b ({signal_1903, signal_1298}), .c ({DataOut_s1[33], DataOut_s0[33]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_127 ( .a ({signal_1572, signal_891}), .b ({signal_1904, signal_1299}), .c ({DataOut_s1[32], DataOut_s0[32]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_128 ( .a ({signal_1575, signal_892}), .b ({signal_1913, signal_1308}), .c ({DataOut_s1[31], DataOut_s0[31]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_129 ( .a ({signal_1578, signal_893}), .b ({signal_1914, signal_1309}), .c ({DataOut_s1[30], DataOut_s0[30]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_130 ( .a ({signal_1581, signal_921}), .b ({signal_1866, signal_1261}), .c ({DataOut_s1[2], DataOut_s0[2]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_131 ( .a ({signal_1584, signal_894}), .b ({signal_1915, signal_1310}), .c ({DataOut_s1[29], DataOut_s0[29]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_132 ( .a ({signal_1587, signal_895}), .b ({signal_1916, signal_1311}), .c ({DataOut_s1[28], DataOut_s0[28]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_133 ( .a ({signal_1590, signal_896}), .b ({signal_1885, signal_1280}), .c ({DataOut_s1[27], DataOut_s0[27]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_134 ( .a ({signal_1593, signal_897}), .b ({signal_1886, signal_1281}), .c ({DataOut_s1[26], DataOut_s0[26]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_135 ( .a ({signal_1596, signal_898}), .b ({signal_1887, signal_1282}), .c ({DataOut_s1[25], DataOut_s0[25]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_136 ( .a ({signal_1599, signal_899}), .b ({signal_1888, signal_1283}), .c ({DataOut_s1[24], DataOut_s0[24]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_137 ( .a ({signal_1602, signal_900}), .b ({signal_1857, signal_1252}), .c ({DataOut_s1[23], DataOut_s0[23]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_138 ( .a ({signal_1605, signal_901}), .b ({signal_1858, signal_1253}), .c ({DataOut_s1[22], DataOut_s0[22]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_139 ( .a ({signal_1608, signal_902}), .b ({signal_1859, signal_1254}), .c ({DataOut_s1[21], DataOut_s0[21]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_140 ( .a ({signal_1611, signal_903}), .b ({signal_1860, signal_1255}), .c ({DataOut_s1[20], DataOut_s0[20]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_141 ( .a ({signal_1614, signal_922}), .b ({signal_1867, signal_1262}), .c ({DataOut_s1[1], DataOut_s0[1]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_142 ( .a ({signal_1617, signal_904}), .b ({signal_1877, signal_1272}), .c ({DataOut_s1[19], DataOut_s0[19]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_143 ( .a ({signal_1620, signal_905}), .b ({signal_1878, signal_1273}), .c ({DataOut_s1[18], DataOut_s0[18]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_144 ( .a ({signal_1623, signal_906}), .b ({signal_1879, signal_1274}), .c ({DataOut_s1[17], DataOut_s0[17]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_145 ( .a ({signal_1626, signal_907}), .b ({signal_1880, signal_1275}), .c ({DataOut_s1[16], DataOut_s0[16]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_146 ( .a ({signal_1629, signal_908}), .b ({signal_1893, signal_1288}), .c ({DataOut_s1[15], DataOut_s0[15]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_147 ( .a ({signal_1632, signal_909}), .b ({signal_1894, signal_1289}), .c ({DataOut_s1[14], DataOut_s0[14]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_148 ( .a ({signal_1635, signal_910}), .b ({signal_1895, signal_1290}), .c ({DataOut_s1[13], DataOut_s0[13]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_149 ( .a ({signal_1638, signal_911}), .b ({signal_1896, signal_1291}), .c ({DataOut_s1[12], DataOut_s0[12]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_150 ( .a ({signal_1641, signal_912}), .b ({signal_1905, signal_1300}), .c ({DataOut_s1[11], DataOut_s0[11]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_151 ( .a ({signal_1644, signal_913}), .b ({signal_1906, signal_1301}), .c ({DataOut_s1[10], DataOut_s0[10]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_152 ( .a ({signal_1647, signal_923}), .b ({signal_1868, signal_1263}), .c ({DataOut_s1[0], DataOut_s0[0]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_217 ( .a ({signal_1654, signal_311}), .b ({signal_1907, signal_1302}), .c ({signal_1981, signal_1238}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_218 ( .a ({signal_1908, signal_1303}), .b ({signal_2254, signal_286}), .c ({signal_2306, signal_1239}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_219 ( .a ({signal_1993, signal_309}), .b ({signal_1869, signal_1264}), .c ({signal_2042, signal_1240}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_220 ( .a ({signal_1992, signal_308}), .b ({signal_1870, signal_1265}), .c ({signal_2043, signal_1241}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_221 ( .a ({signal_2041, signal_365}), .b ({signal_1853, signal_1248}), .c ({signal_2044, signal_1184}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_222 ( .a ({signal_2040, signal_364}), .b ({signal_1854, signal_1249}), .c ({signal_2045, signal_1185}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_223 ( .a ({signal_2039, signal_363}), .b ({signal_1855, signal_1250}), .c ({signal_2046, signal_1186}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_224 ( .a ({signal_1856, signal_1251}), .b ({signal_2310, signal_287}), .c ({signal_2362, signal_1187}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_225 ( .a ({signal_1991, signal_307}), .b ({signal_1871, signal_1266}), .c ({signal_2047, signal_1242}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_226 ( .a ({signal_2037, signal_361}), .b ({signal_1881, signal_1276}), .c ({signal_2048, signal_1188}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_227 ( .a ({signal_2036, signal_360}), .b ({signal_1882, signal_1277}), .c ({signal_2049, signal_1189}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_228 ( .a ({signal_2035, signal_359}), .b ({signal_1883, signal_1278}), .c ({signal_2050, signal_1190}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_229 ( .a ({signal_1884, signal_1279}), .b ({signal_2311, signal_288}), .c ({signal_2363, signal_1191}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_230 ( .a ({signal_2033, signal_357}), .b ({signal_1909, signal_1304}), .c ({signal_2051, signal_1192}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_231 ( .a ({signal_2032, signal_356}), .b ({signal_1910, signal_1305}), .c ({signal_2052, signal_1193}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_232 ( .a ({signal_2031, signal_355}), .b ({signal_1911, signal_1306}), .c ({signal_2053, signal_1194}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_233 ( .a ({signal_1912, signal_1307}), .b ({signal_2312, signal_289}), .c ({signal_2364, signal_1195}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_234 ( .a ({signal_2029, signal_353}), .b ({signal_1889, signal_1284}), .c ({signal_2054, signal_1196}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_235 ( .a ({signal_2028, signal_352}), .b ({signal_1890, signal_1285}), .c ({signal_2055, signal_1197}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_236 ( .a ({signal_1872, signal_1267}), .b ({signal_2313, signal_290}), .c ({signal_2365, signal_1243}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_237 ( .a ({signal_2027, signal_351}), .b ({signal_1891, signal_1286}), .c ({signal_2056, signal_1198}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_238 ( .a ({signal_1892, signal_1287}), .b ({signal_2378, signal_291}), .c ({signal_2389, signal_1199}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_239 ( .a ({signal_2025, signal_349}), .b ({signal_1873, signal_1268}), .c ({signal_2057, signal_1200}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_240 ( .a ({signal_2024, signal_348}), .b ({signal_1874, signal_1269}), .c ({signal_2058, signal_1201}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_241 ( .a ({signal_2023, signal_347}), .b ({signal_1875, signal_1270}), .c ({signal_2059, signal_1202}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_242 ( .a ({signal_1876, signal_1271}), .b ({signal_2255, signal_292}), .c ({signal_2307, signal_1203}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_243 ( .a ({signal_2021, signal_345}), .b ({signal_1861, signal_1256}), .c ({signal_2060, signal_1204}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_244 ( .a ({signal_2020, signal_344}), .b ({signal_1862, signal_1257}), .c ({signal_2061, signal_1205}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_245 ( .a ({signal_2019, signal_343}), .b ({signal_1863, signal_1258}), .c ({signal_2062, signal_1206}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_246 ( .a ({signal_1864, signal_1259}), .b ({signal_2314, signal_293}), .c ({signal_2366, signal_1207}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_247 ( .a ({signal_1651, signal_305}), .b ({signal_1865, signal_1260}), .c ({signal_1982, signal_1244}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_248 ( .a ({signal_2017, signal_341}), .b ({signal_1897, signal_1292}), .c ({signal_2063, signal_1208}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_249 ( .a ({signal_2016, signal_340}), .b ({signal_1898, signal_1293}), .c ({signal_2064, signal_1209}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_250 ( .a ({signal_2015, signal_339}), .b ({signal_1899, signal_1294}), .c ({signal_2065, signal_1210}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_251 ( .a ({signal_1900, signal_1295}), .b ({signal_2256, signal_294}), .c ({signal_2308, signal_1211}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_252 ( .a ({signal_2013, signal_337}), .b ({signal_1901, signal_1296}), .c ({signal_2066, signal_1212}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_253 ( .a ({signal_2012, signal_336}), .b ({signal_1902, signal_1297}), .c ({signal_2067, signal_1213}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_254 ( .a ({signal_2011, signal_335}), .b ({signal_1903, signal_1298}), .c ({signal_2068, signal_1214}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_255 ( .a ({signal_1904, signal_1299}), .b ({signal_2315, signal_295}), .c ({signal_2367, signal_1215}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_256 ( .a ({signal_2009, signal_333}), .b ({signal_1913, signal_1308}), .c ({signal_2069, signal_1216}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_257 ( .a ({signal_2008, signal_332}), .b ({signal_1914, signal_1309}), .c ({signal_2070, signal_1217}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_258 ( .a ({signal_1650, signal_304}), .b ({signal_1866, signal_1261}), .c ({signal_1983, signal_1245}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_259 ( .a ({signal_2007, signal_331}), .b ({signal_1915, signal_1310}), .c ({signal_2071, signal_1218}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_260 ( .a ({signal_1916, signal_1311}), .b ({signal_2372, signal_296}), .c ({signal_2377, signal_1219}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_261 ( .a ({signal_2005, signal_329}), .b ({signal_1885, signal_1280}), .c ({signal_2072, signal_1220}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_262 ( .a ({signal_1660, signal_328}), .b ({signal_1886, signal_1281}), .c ({signal_1984, signal_1221}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_263 ( .a ({signal_2004, signal_327}), .b ({signal_1887, signal_1282}), .c ({signal_2073, signal_1222}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_264 ( .a ({signal_1888, signal_1283}), .b ({signal_2316, signal_297}), .c ({signal_2368, signal_1223}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_265 ( .a ({signal_2002, signal_325}), .b ({signal_1857, signal_1252}), .c ({signal_2074, signal_1224}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_266 ( .a ({signal_2001, signal_324}), .b ({signal_1858, signal_1253}), .c ({signal_2075, signal_1225}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_267 ( .a ({signal_2000, signal_323}), .b ({signal_1859, signal_1254}), .c ({signal_2076, signal_1226}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_268 ( .a ({signal_1860, signal_1255}), .b ({signal_2257, signal_298}), .c ({signal_2309, signal_1227}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_269 ( .a ({signal_1649, signal_303}), .b ({signal_1867, signal_1262}), .c ({signal_1985, signal_1246}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_270 ( .a ({signal_1998, signal_321}), .b ({signal_1877, signal_1272}), .c ({signal_2077, signal_1228}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_271 ( .a ({signal_1997, signal_320}), .b ({signal_1878, signal_1273}), .c ({signal_2078, signal_1229}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_272 ( .a ({signal_1996, signal_319}), .b ({signal_1879, signal_1274}), .c ({signal_2079, signal_1230}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_273 ( .a ({signal_1880, signal_1275}), .b ({signal_2317, signal_299}), .c ({signal_2369, signal_1231}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_274 ( .a ({signal_1659, signal_317}), .b ({signal_1893, signal_1288}), .c ({signal_1986, signal_1232}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_275 ( .a ({signal_1658, signal_316}), .b ({signal_1894, signal_1289}), .c ({signal_1987, signal_1233}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_276 ( .a ({signal_1657, signal_315}), .b ({signal_1895, signal_1290}), .c ({signal_1988, signal_1234}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_277 ( .a ({signal_1896, signal_1291}), .b ({signal_2318, signal_300}), .c ({signal_2370, signal_1235}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_278 ( .a ({signal_1656, signal_313}), .b ({signal_1905, signal_1300}), .c ({signal_1989, signal_1236}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_279 ( .a ({signal_1655, signal_312}), .b ({signal_1906, signal_1301}), .c ({signal_1990, signal_1237}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_280 ( .a ({signal_1868, signal_1263}), .b ({signal_2319, signal_301}), .c ({signal_2371, signal_1247}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_281 ( .a ({signal_1654, signal_311}), .b ({signal_2200, signal_1110}), .c ({signal_2206, signal_1046}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_282 ( .a ({signal_2406, signal_1111}), .b ({signal_2254, signal_286}), .c ({signal_2410, signal_1047}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_284 ( .a ({signal_1993, signal_309}), .b ({signal_2149, signal_1064}), .c ({signal_2158, signal_1048}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_285 ( .a ({signal_1992, signal_308}), .b ({signal_2150, signal_1065}), .c ({signal_2159, signal_1049}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_286 ( .a ({signal_2041, signal_365}), .b ({signal_2171, signal_1056}), .c ({signal_2207, signal_992}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_287 ( .a ({signal_2040, signal_364}), .b ({signal_2172, signal_1057}), .c ({signal_2208, signal_993}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_288 ( .a ({signal_2039, signal_363}), .b ({signal_2173, signal_1058}), .c ({signal_2209, signal_994}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_289 ( .a ({signal_2429, signal_1059}), .b ({signal_2310, signal_287}), .c ({signal_2441, signal_995}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_291 ( .a ({signal_1991, signal_307}), .b ({signal_2151, signal_1066}), .c ({signal_2160, signal_1050}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_292 ( .a ({signal_2037, signal_361}), .b ({signal_2174, signal_1096}), .c ({signal_2210, signal_996}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_293 ( .a ({signal_2036, signal_360}), .b ({signal_2175, signal_1097}), .c ({signal_2211, signal_997}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_294 ( .a ({signal_2035, signal_359}), .b ({signal_2164, signal_1098}), .c ({signal_2212, signal_998}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_295 ( .a ({signal_2428, signal_1099}), .b ({signal_2311, signal_288}), .c ({signal_2442, signal_999}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_297 ( .a ({signal_2033, signal_357}), .b ({signal_2165, signal_1076}), .c ({signal_2213, signal_1000}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_298 ( .a ({signal_2032, signal_356}), .b ({signal_2166, signal_1077}), .c ({signal_2214, signal_1001}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_299 ( .a ({signal_2031, signal_355}), .b ({signal_2167, signal_1078}), .c ({signal_2215, signal_1002}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_300 ( .a ({signal_2421, signal_1079}), .b ({signal_2312, signal_289}), .c ({signal_2425, signal_1003}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_302 ( .a ({signal_2029, signal_353}), .b ({signal_2168, signal_1116}), .c ({signal_2216, signal_1004}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_303 ( .a ({signal_2028, signal_352}), .b ({signal_2169, signal_1117}), .c ({signal_2217, signal_1005}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_304 ( .a ({signal_2407, signal_1067}), .b ({signal_2313, signal_290}), .c ({signal_2411, signal_1051}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_306 ( .a ({signal_2027, signal_351}), .b ({signal_2170, signal_1118}), .c ({signal_2218, signal_1006}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_307 ( .a ({signal_2398, signal_1119}), .b ({signal_2378, signal_291}), .c ({signal_2412, signal_1007}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_309 ( .a ({signal_2025, signal_349}), .b ({signal_2183, signal_1112}), .c ({signal_2219, signal_1008}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_310 ( .a ({signal_2024, signal_348}), .b ({signal_2184, signal_1113}), .c ({signal_2220, signal_1009}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_311 ( .a ({signal_2023, signal_347}), .b ({signal_2185, signal_1114}), .c ({signal_2221, signal_1010}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_312 ( .a ({signal_2401, signal_1115}), .b ({signal_2255, signal_292}), .c ({signal_2413, signal_1011}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_314 ( .a ({signal_2021, signal_345}), .b ({signal_2186, signal_1072}), .c ({signal_2222, signal_1012}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_315 ( .a ({signal_2020, signal_344}), .b ({signal_2187, signal_1073}), .c ({signal_2223, signal_1013}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_316 ( .a ({signal_2019, signal_343}), .b ({signal_2176, signal_1074}), .c ({signal_2224, signal_1014}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_317 ( .a ({signal_2399, signal_1075}), .b ({signal_2314, signal_293}), .c ({signal_2414, signal_1015}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_319 ( .a ({signal_1651, signal_305}), .b ({signal_2152, signal_1088}), .c ({signal_2161, signal_1052}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_320 ( .a ({signal_2017, signal_341}), .b ({signal_2177, signal_1100}), .c ({signal_2225, signal_1016}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_321 ( .a ({signal_2016, signal_340}), .b ({signal_2178, signal_1101}), .c ({signal_2226, signal_1017}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_322 ( .a ({signal_2015, signal_339}), .b ({signal_2179, signal_1102}), .c ({signal_2227, signal_1018}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_323 ( .a ({signal_2400, signal_1103}), .b ({signal_2256, signal_294}), .c ({signal_2415, signal_1019}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_325 ( .a ({signal_2013, signal_337}), .b ({signal_2180, signal_1060}), .c ({signal_2228, signal_1020}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_326 ( .a ({signal_2012, signal_336}), .b ({signal_2181, signal_1061}), .c ({signal_2229, signal_1021}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_327 ( .a ({signal_2011, signal_335}), .b ({signal_2182, signal_1062}), .c ({signal_2230, signal_1022}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_328 ( .a ({signal_2402, signal_1063}), .b ({signal_2315, signal_295}), .c ({signal_2416, signal_1023}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_330 ( .a ({signal_2009, signal_333}), .b ({signal_2195, signal_1092}), .c ({signal_2231, signal_1024}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_331 ( .a ({signal_2008, signal_332}), .b ({signal_2196, signal_1093}), .c ({signal_2232, signal_1025}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_332 ( .a ({signal_1650, signal_304}), .b ({signal_2153, signal_1089}), .c ({signal_2162, signal_1053}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_333 ( .a ({signal_2007, signal_331}), .b ({signal_2197, signal_1094}), .c ({signal_2233, signal_1026}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_334 ( .a ({signal_2404, signal_1095}), .b ({signal_2372, signal_296}), .c ({signal_2417, signal_1027}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_336 ( .a ({signal_2005, signal_329}), .b ({signal_2198, signal_1068}), .c ({signal_2234, signal_1028}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_337 ( .a ({signal_1660, signal_328}), .b ({signal_2199, signal_1069}), .c ({signal_2235, signal_1029}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_338 ( .a ({signal_2004, signal_327}), .b ({signal_2188, signal_1070}), .c ({signal_2236, signal_1030}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_339 ( .a ({signal_2403, signal_1071}), .b ({signal_2316, signal_297}), .c ({signal_2418, signal_1031}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_341 ( .a ({signal_2002, signal_325}), .b ({signal_2189, signal_1104}), .c ({signal_2237, signal_1032}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_342 ( .a ({signal_2001, signal_324}), .b ({signal_2190, signal_1105}), .c ({signal_2238, signal_1033}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_343 ( .a ({signal_2000, signal_323}), .b ({signal_2191, signal_1106}), .c ({signal_2239, signal_1034}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_344 ( .a ({signal_2423, signal_1107}), .b ({signal_2257, signal_298}), .c ({signal_2426, signal_1035}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_346 ( .a ({signal_1649, signal_303}), .b ({signal_2154, signal_1090}), .c ({signal_2163, signal_1054}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_347 ( .a ({signal_1998, signal_321}), .b ({signal_2192, signal_1080}), .c ({signal_2240, signal_1036}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_348 ( .a ({signal_1997, signal_320}), .b ({signal_2193, signal_1081}), .c ({signal_2241, signal_1037}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_349 ( .a ({signal_1996, signal_319}), .b ({signal_2194, signal_1082}), .c ({signal_2242, signal_1038}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_350 ( .a ({signal_2424, signal_1083}), .b ({signal_2317, signal_299}), .c ({signal_2427, signal_1039}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_352 ( .a ({signal_1659, signal_317}), .b ({signal_2201, signal_1084}), .c ({signal_2243, signal_1040}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_353 ( .a ({signal_1658, signal_316}), .b ({signal_2202, signal_1085}), .c ({signal_2244, signal_1041}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_354 ( .a ({signal_1657, signal_315}), .b ({signal_2203, signal_1086}), .c ({signal_2245, signal_1042}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_355 ( .a ({signal_2408, signal_1087}), .b ({signal_2318, signal_300}), .c ({signal_2419, signal_1043}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_357 ( .a ({signal_1656, signal_313}), .b ({signal_2204, signal_1108}), .c ({signal_2246, signal_1044}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_358 ( .a ({signal_1655, signal_312}), .b ({signal_2205, signal_1109}), .c ({signal_2247, signal_1045}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_359 ( .a ({signal_2409, signal_1091}), .b ({signal_2319, signal_301}), .c ({signal_2420, signal_1055}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_535 ( .s (reset), .b ({signal_2430, signal_1439}), .a ({signal_1788, signal_991}), .c ({signal_2443, signal_460}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_538 ( .s (reset), .b ({signal_2248, signal_1438}), .a ({signal_1766, signal_990}), .c ({signal_2258, signal_462}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_541 ( .s (reset), .b ({signal_2249, signal_1437}), .a ({signal_1744, signal_989}), .c ({signal_2259, signal_464}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_544 ( .s (reset), .b ({signal_2250, signal_1436}), .a ({signal_1722, signal_988}), .c ({signal_2260, signal_466}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_547 ( .s (reset), .b ({signal_2431, signal_1435}), .a ({signal_1700, signal_987}), .c ({signal_2444, signal_468}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_550 ( .s (reset), .b ({signal_2251, signal_1434}), .a ({signal_1678, signal_986}), .c ({signal_2261, signal_470}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_553 ( .s (reset), .b ({signal_2252, signal_1433}), .a ({signal_1668, signal_985}), .c ({signal_2262, signal_472}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_556 ( .s (reset), .b ({signal_2253, signal_1432}), .a ({signal_1666, signal_984}), .c ({signal_2263, signal_474}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_559 ( .s (reset), .b ({signal_2432, signal_1431}), .a ({signal_1664, signal_983}), .c ({signal_2445, signal_476}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_562 ( .s (reset), .b ({signal_2264, signal_1430}), .a ({signal_1662, signal_982}), .c ({signal_2320, signal_478}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_565 ( .s (reset), .b ({signal_2265, signal_1429}), .a ({signal_1786, signal_981}), .c ({signal_2321, signal_480}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_568 ( .s (reset), .b ({signal_2266, signal_1428}), .a ({signal_1784, signal_980}), .c ({signal_2322, signal_482}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_571 ( .s (reset), .b ({signal_2433, signal_1427}), .a ({signal_1782, signal_979}), .c ({signal_2446, signal_484}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_574 ( .s (reset), .b ({signal_2267, signal_1426}), .a ({signal_1780, signal_978}), .c ({signal_2323, signal_486}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_577 ( .s (reset), .b ({signal_2268, signal_1425}), .a ({signal_1778, signal_977}), .c ({signal_2324, signal_488}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_580 ( .s (reset), .b ({signal_2269, signal_1424}), .a ({signal_1776, signal_976}), .c ({signal_2325, signal_490}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_583 ( .s (reset), .b ({signal_2454, signal_1423}), .a ({signal_1774, signal_975}), .c ({signal_2457, signal_492}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_586 ( .s (reset), .b ({signal_2270, signal_1422}), .a ({signal_1772, signal_974}), .c ({signal_2326, signal_494}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_589 ( .s (reset), .b ({signal_2271, signal_1421}), .a ({signal_1770, signal_973}), .c ({signal_2327, signal_496}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_592 ( .s (reset), .b ({signal_2272, signal_1420}), .a ({signal_1768, signal_972}), .c ({signal_2328, signal_498}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_595 ( .s (reset), .b ({signal_2455, signal_1419}), .a ({signal_1764, signal_971}), .c ({signal_2458, signal_500}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_598 ( .s (reset), .b ({signal_2273, signal_1418}), .a ({signal_1762, signal_970}), .c ({signal_2329, signal_502}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_601 ( .s (reset), .b ({signal_2274, signal_1417}), .a ({signal_1760, signal_969}), .c ({signal_2330, signal_504}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_604 ( .s (reset), .b ({signal_2275, signal_1416}), .a ({signal_1758, signal_968}), .c ({signal_2331, signal_506}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_607 ( .s (reset), .b ({signal_2434, signal_1415}), .a ({signal_1756, signal_967}), .c ({signal_2447, signal_508}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_610 ( .s (reset), .b ({signal_2276, signal_1414}), .a ({signal_1754, signal_966}), .c ({signal_2332, signal_510}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_613 ( .s (reset), .b ({signal_2277, signal_1413}), .a ({signal_1752, signal_965}), .c ({signal_2333, signal_512}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_616 ( .s (reset), .b ({signal_2278, signal_1412}), .a ({signal_1750, signal_964}), .c ({signal_2334, signal_514}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_619 ( .s (reset), .b ({signal_2435, signal_1411}), .a ({signal_1748, signal_963}), .c ({signal_2448, signal_516}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_622 ( .s (reset), .b ({signal_2279, signal_1410}), .a ({signal_1746, signal_962}), .c ({signal_2335, signal_518}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_625 ( .s (reset), .b ({signal_2280, signal_1409}), .a ({signal_1742, signal_961}), .c ({signal_2336, signal_520}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_628 ( .s (reset), .b ({signal_2281, signal_1408}), .a ({signal_1740, signal_960}), .c ({signal_2337, signal_522}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_631 ( .s (reset), .b ({signal_2436, signal_1407}), .a ({signal_1738, signal_959}), .c ({signal_2449, signal_524}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_634 ( .s (reset), .b ({signal_2282, signal_1406}), .a ({signal_1736, signal_958}), .c ({signal_2338, signal_526}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_637 ( .s (reset), .b ({signal_2283, signal_1405}), .a ({signal_1734, signal_957}), .c ({signal_2339, signal_528}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_640 ( .s (reset), .b ({signal_2284, signal_1404}), .a ({signal_1732, signal_956}), .c ({signal_2340, signal_530}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_643 ( .s (reset), .b ({signal_2437, signal_1403}), .a ({signal_1730, signal_955}), .c ({signal_2450, signal_532}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_646 ( .s (reset), .b ({signal_2285, signal_1402}), .a ({signal_1728, signal_954}), .c ({signal_2341, signal_534}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_649 ( .s (reset), .b ({signal_2286, signal_1401}), .a ({signal_1726, signal_953}), .c ({signal_2342, signal_536}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_652 ( .s (reset), .b ({signal_2287, signal_1400}), .a ({signal_1724, signal_952}), .c ({signal_2343, signal_538}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_655 ( .s (reset), .b ({signal_2438, signal_1399}), .a ({signal_1720, signal_951}), .c ({signal_2451, signal_540}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_658 ( .s (reset), .b ({signal_2288, signal_1398}), .a ({signal_1718, signal_950}), .c ({signal_2344, signal_542}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_661 ( .s (reset), .b ({signal_2289, signal_1397}), .a ({signal_1716, signal_949}), .c ({signal_2345, signal_544}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_664 ( .s (reset), .b ({signal_2290, signal_1396}), .a ({signal_1714, signal_948}), .c ({signal_2346, signal_546}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_667 ( .s (reset), .b ({signal_2439, signal_1395}), .a ({signal_1712, signal_947}), .c ({signal_2452, signal_548}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_670 ( .s (reset), .b ({signal_2291, signal_1394}), .a ({signal_1710, signal_946}), .c ({signal_2347, signal_550}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_673 ( .s (reset), .b ({signal_2292, signal_1393}), .a ({signal_1708, signal_945}), .c ({signal_2348, signal_552}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_676 ( .s (reset), .b ({signal_2293, signal_1392}), .a ({signal_1706, signal_944}), .c ({signal_2349, signal_554}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_679 ( .s (reset), .b ({signal_2440, signal_1391}), .a ({signal_1704, signal_943}), .c ({signal_2453, signal_556}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_682 ( .s (reset), .b ({signal_2294, signal_1390}), .a ({signal_1702, signal_942}), .c ({signal_2350, signal_558}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_685 ( .s (reset), .b ({signal_2295, signal_1389}), .a ({signal_1698, signal_941}), .c ({signal_2351, signal_560}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_688 ( .s (reset), .b ({signal_2296, signal_1388}), .a ({signal_1696, signal_940}), .c ({signal_2352, signal_562}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_691 ( .s (reset), .b ({signal_2456, signal_1387}), .a ({signal_1694, signal_939}), .c ({signal_2459, signal_564}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_694 ( .s (reset), .b ({signal_2297, signal_1386}), .a ({signal_1692, signal_938}), .c ({signal_2353, signal_566}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_697 ( .s (reset), .b ({signal_2298, signal_1385}), .a ({signal_1690, signal_937}), .c ({signal_2354, signal_568}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_700 ( .s (reset), .b ({signal_2299, signal_1384}), .a ({signal_1688, signal_936}), .c ({signal_2355, signal_570}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_703 ( .s (reset), .b ({signal_2460, signal_1383}), .a ({signal_1686, signal_935}), .c ({signal_2462, signal_572}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_706 ( .s (reset), .b ({signal_2300, signal_1382}), .a ({signal_1684, signal_934}), .c ({signal_2356, signal_574}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_709 ( .s (reset), .b ({signal_2301, signal_1381}), .a ({signal_1682, signal_933}), .c ({signal_2357, signal_576}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_712 ( .s (reset), .b ({signal_2302, signal_1380}), .a ({signal_1680, signal_932}), .c ({signal_2358, signal_578}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_715 ( .s (reset), .b ({signal_2461, signal_1379}), .a ({signal_1676, signal_931}), .c ({signal_2463, signal_580}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_718 ( .s (reset), .b ({signal_2303, signal_1378}), .a ({signal_1674, signal_930}), .c ({signal_2359, signal_582}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_721 ( .s (reset), .b ({signal_2304, signal_1377}), .a ({signal_1672, signal_929}), .c ({signal_2360, signal_584}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_724 ( .s (reset), .b ({signal_2305, signal_1376}), .a ({signal_1670, signal_928}), .c ({signal_2361, signal_586}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1031 ( .s (enc_dec), .b ({signal_1916, signal_1311}), .a ({signal_2371, signal_1247}), .c ({signal_2379, signal_1183}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1032 ( .s (enc_dec), .b ({signal_1915, signal_1310}), .a ({signal_1985, signal_1246}), .c ({signal_2080, signal_1182}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1033 ( .s (enc_dec), .b ({signal_1914, signal_1309}), .a ({signal_1983, signal_1245}), .c ({signal_2081, signal_1181}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1034 ( .s (enc_dec), .b ({signal_1913, signal_1308}), .a ({signal_1982, signal_1244}), .c ({signal_2082, signal_1180}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1035 ( .s (enc_dec), .b ({signal_1912, signal_1307}), .a ({signal_2365, signal_1243}), .c ({signal_2380, signal_1179}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1036 ( .s (enc_dec), .b ({signal_1911, signal_1306}), .a ({signal_2047, signal_1242}), .c ({signal_2090, signal_1178}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1037 ( .s (enc_dec), .b ({signal_1910, signal_1305}), .a ({signal_2043, signal_1241}), .c ({signal_2091, signal_1177}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1038 ( .s (enc_dec), .b ({signal_1909, signal_1304}), .a ({signal_2042, signal_1240}), .c ({signal_2092, signal_1176}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1039 ( .s (enc_dec), .b ({signal_1908, signal_1303}), .a ({signal_2306, signal_1239}), .c ({signal_2373, signal_1175}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1040 ( .s (enc_dec), .b ({signal_1907, signal_1302}), .a ({signal_1981, signal_1238}), .c ({signal_2083, signal_1174}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1041 ( .s (enc_dec), .b ({signal_1906, signal_1301}), .a ({signal_1990, signal_1237}), .c ({signal_2084, signal_1173}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1042 ( .s (enc_dec), .b ({signal_1905, signal_1300}), .a ({signal_1989, signal_1236}), .c ({signal_2085, signal_1172}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1043 ( .s (enc_dec), .b ({signal_1904, signal_1299}), .a ({signal_2370, signal_1235}), .c ({signal_2381, signal_1171}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1044 ( .s (enc_dec), .b ({signal_1903, signal_1298}), .a ({signal_1988, signal_1234}), .c ({signal_2086, signal_1170}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1045 ( .s (enc_dec), .b ({signal_1902, signal_1297}), .a ({signal_1987, signal_1233}), .c ({signal_2087, signal_1169}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1046 ( .s (enc_dec), .b ({signal_1901, signal_1296}), .a ({signal_1986, signal_1232}), .c ({signal_2088, signal_1168}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1047 ( .s (enc_dec), .b ({signal_1900, signal_1295}), .a ({signal_2369, signal_1231}), .c ({signal_2382, signal_1167}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1048 ( .s (enc_dec), .b ({signal_1899, signal_1294}), .a ({signal_2079, signal_1230}), .c ({signal_2093, signal_1166}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1049 ( .s (enc_dec), .b ({signal_1898, signal_1293}), .a ({signal_2078, signal_1229}), .c ({signal_2094, signal_1165}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1050 ( .s (enc_dec), .b ({signal_1897, signal_1292}), .a ({signal_2077, signal_1228}), .c ({signal_2095, signal_1164}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1051 ( .s (enc_dec), .b ({signal_1896, signal_1291}), .a ({signal_2309, signal_1227}), .c ({signal_2374, signal_1163}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1052 ( .s (enc_dec), .b ({signal_1895, signal_1290}), .a ({signal_2076, signal_1226}), .c ({signal_2096, signal_1162}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1053 ( .s (enc_dec), .b ({signal_1894, signal_1289}), .a ({signal_2075, signal_1225}), .c ({signal_2097, signal_1161}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1054 ( .s (enc_dec), .b ({signal_1893, signal_1288}), .a ({signal_2074, signal_1224}), .c ({signal_2098, signal_1160}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1055 ( .s (enc_dec), .b ({signal_1892, signal_1287}), .a ({signal_2368, signal_1223}), .c ({signal_2383, signal_1159}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1056 ( .s (enc_dec), .b ({signal_1891, signal_1286}), .a ({signal_2073, signal_1222}), .c ({signal_2099, signal_1158}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1057 ( .s (enc_dec), .b ({signal_1890, signal_1285}), .a ({signal_1984, signal_1221}), .c ({signal_2089, signal_1157}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1058 ( .s (enc_dec), .b ({signal_1889, signal_1284}), .a ({signal_2072, signal_1220}), .c ({signal_2100, signal_1156}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1059 ( .s (enc_dec), .b ({signal_1888, signal_1283}), .a ({signal_2377, signal_1219}), .c ({signal_2390, signal_1155}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1060 ( .s (enc_dec), .b ({signal_1887, signal_1282}), .a ({signal_2071, signal_1218}), .c ({signal_2101, signal_1154}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1061 ( .s (enc_dec), .b ({signal_1886, signal_1281}), .a ({signal_2070, signal_1217}), .c ({signal_2102, signal_1153}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1062 ( .s (enc_dec), .b ({signal_1885, signal_1280}), .a ({signal_2069, signal_1216}), .c ({signal_2103, signal_1152}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1063 ( .s (enc_dec), .b ({signal_1884, signal_1279}), .a ({signal_2367, signal_1215}), .c ({signal_2384, signal_1151}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1064 ( .s (enc_dec), .b ({signal_1883, signal_1278}), .a ({signal_2068, signal_1214}), .c ({signal_2104, signal_1150}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1065 ( .s (enc_dec), .b ({signal_1882, signal_1277}), .a ({signal_2067, signal_1213}), .c ({signal_2105, signal_1149}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1066 ( .s (enc_dec), .b ({signal_1881, signal_1276}), .a ({signal_2066, signal_1212}), .c ({signal_2106, signal_1148}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1067 ( .s (enc_dec), .b ({signal_1880, signal_1275}), .a ({signal_2308, signal_1211}), .c ({signal_2375, signal_1147}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1068 ( .s (enc_dec), .b ({signal_1879, signal_1274}), .a ({signal_2065, signal_1210}), .c ({signal_2107, signal_1146}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1069 ( .s (enc_dec), .b ({signal_1878, signal_1273}), .a ({signal_2064, signal_1209}), .c ({signal_2108, signal_1145}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1070 ( .s (enc_dec), .b ({signal_1877, signal_1272}), .a ({signal_2063, signal_1208}), .c ({signal_2109, signal_1144}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1071 ( .s (enc_dec), .b ({signal_1876, signal_1271}), .a ({signal_2366, signal_1207}), .c ({signal_2385, signal_1143}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1072 ( .s (enc_dec), .b ({signal_1875, signal_1270}), .a ({signal_2062, signal_1206}), .c ({signal_2110, signal_1142}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1073 ( .s (enc_dec), .b ({signal_1874, signal_1269}), .a ({signal_2061, signal_1205}), .c ({signal_2111, signal_1141}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1074 ( .s (enc_dec), .b ({signal_1873, signal_1268}), .a ({signal_2060, signal_1204}), .c ({signal_2112, signal_1140}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1075 ( .s (enc_dec), .b ({signal_1872, signal_1267}), .a ({signal_2307, signal_1203}), .c ({signal_2376, signal_1139}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1076 ( .s (enc_dec), .b ({signal_1871, signal_1266}), .a ({signal_2059, signal_1202}), .c ({signal_2113, signal_1138}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1077 ( .s (enc_dec), .b ({signal_1870, signal_1265}), .a ({signal_2058, signal_1201}), .c ({signal_2114, signal_1137}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1078 ( .s (enc_dec), .b ({signal_1869, signal_1264}), .a ({signal_2057, signal_1200}), .c ({signal_2115, signal_1136}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1079 ( .s (enc_dec), .b ({signal_1868, signal_1263}), .a ({signal_2389, signal_1199}), .c ({signal_2397, signal_1135}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1080 ( .s (enc_dec), .b ({signal_1867, signal_1262}), .a ({signal_2056, signal_1198}), .c ({signal_2116, signal_1134}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1081 ( .s (enc_dec), .b ({signal_1866, signal_1261}), .a ({signal_2055, signal_1197}), .c ({signal_2117, signal_1133}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1082 ( .s (enc_dec), .b ({signal_1865, signal_1260}), .a ({signal_2054, signal_1196}), .c ({signal_2118, signal_1132}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1083 ( .s (enc_dec), .b ({signal_1864, signal_1259}), .a ({signal_2364, signal_1195}), .c ({signal_2386, signal_1131}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1084 ( .s (enc_dec), .b ({signal_1863, signal_1258}), .a ({signal_2053, signal_1194}), .c ({signal_2119, signal_1130}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1085 ( .s (enc_dec), .b ({signal_1862, signal_1257}), .a ({signal_2052, signal_1193}), .c ({signal_2120, signal_1129}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1086 ( .s (enc_dec), .b ({signal_1861, signal_1256}), .a ({signal_2051, signal_1192}), .c ({signal_2121, signal_1128}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1087 ( .s (enc_dec), .b ({signal_1860, signal_1255}), .a ({signal_2363, signal_1191}), .c ({signal_2387, signal_1127}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1088 ( .s (enc_dec), .b ({signal_1859, signal_1254}), .a ({signal_2050, signal_1190}), .c ({signal_2122, signal_1126}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1089 ( .s (enc_dec), .b ({signal_1858, signal_1253}), .a ({signal_2049, signal_1189}), .c ({signal_2123, signal_1125}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1090 ( .s (enc_dec), .b ({signal_1857, signal_1252}), .a ({signal_2048, signal_1188}), .c ({signal_2124, signal_1124}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1091 ( .s (enc_dec), .b ({signal_1856, signal_1251}), .a ({signal_2362, signal_1187}), .c ({signal_2388, signal_1123}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1092 ( .s (enc_dec), .b ({signal_1855, signal_1250}), .a ({signal_2046, signal_1186}), .c ({signal_2125, signal_1122}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1093 ( .s (enc_dec), .b ({signal_1854, signal_1249}), .a ({signal_2045, signal_1185}), .c ({signal_2126, signal_1121}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1094 ( .s (enc_dec), .b ({signal_1853, signal_1248}), .a ({signal_2044, signal_1184}), .c ({signal_2127, signal_1120}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1095 ( .a ({signal_2125, signal_1122}), .b ({signal_2134, signal_828}), .c ({signal_2164, signal_1098}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1096 ( .a ({signal_2388, signal_1123}), .b ({signal_2422, signal_829}), .c ({signal_2428, signal_1099}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1097 ( .a ({signal_2118, signal_1132}), .b ({signal_2131, signal_830}), .c ({signal_2165, signal_1076}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1098 ( .a ({signal_2117, signal_1133}), .b ({signal_2132, signal_831}), .c ({signal_2166, signal_1077}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1099 ( .a ({signal_2116, signal_1134}), .b ({signal_2133, signal_832}), .c ({signal_2167, signal_1078}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1100 ( .a ({signal_2397, signal_1135}), .b ({signal_2391, signal_833}), .c ({signal_2421, signal_1079}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1101 ( .a ({signal_2121, signal_1128}), .b ({signal_2131, signal_830}), .c ({signal_2168, signal_1116}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1102 ( .a ({signal_2127, signal_1120}), .b ({signal_2124, signal_1124}), .c ({signal_2131, signal_830}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1103 ( .a ({signal_2120, signal_1129}), .b ({signal_2132, signal_831}), .c ({signal_2169, signal_1117}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1104 ( .a ({signal_2126, signal_1121}), .b ({signal_2123, signal_1125}), .c ({signal_2132, signal_831}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1105 ( .a ({signal_2119, signal_1130}), .b ({signal_2133, signal_832}), .c ({signal_2170, signal_1118}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1106 ( .a ({signal_2122, signal_1126}), .b ({signal_2125, signal_1122}), .c ({signal_2133, signal_832}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1107 ( .a ({signal_2124, signal_1124}), .b ({signal_2135, signal_834}), .c ({signal_2171, signal_1056}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1108 ( .a ({signal_2123, signal_1125}), .b ({signal_2136, signal_835}), .c ({signal_2172, signal_1057}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1109 ( .a ({signal_2122, signal_1126}), .b ({signal_2134, signal_828}), .c ({signal_2173, signal_1058}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1110 ( .a ({signal_2116, signal_1134}), .b ({signal_2119, signal_1130}), .c ({signal_2134, signal_828}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1111 ( .a ({signal_2387, signal_1127}), .b ({signal_2422, signal_829}), .c ({signal_2429, signal_1059}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1112 ( .a ({signal_2386, signal_1131}), .b ({signal_2397, signal_1135}), .c ({signal_2422, signal_829}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1113 ( .a ({signal_2127, signal_1120}), .b ({signal_2135, signal_834}), .c ({signal_2174, signal_1096}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1114 ( .a ({signal_2118, signal_1132}), .b ({signal_2121, signal_1128}), .c ({signal_2135, signal_834}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1115 ( .a ({signal_2126, signal_1121}), .b ({signal_2136, signal_835}), .c ({signal_2175, signal_1097}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1116 ( .a ({signal_2117, signal_1133}), .b ({signal_2120, signal_1129}), .c ({signal_2136, signal_835}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1117 ( .a ({signal_2386, signal_1131}), .b ({signal_2391, signal_833}), .c ({signal_2398, signal_1119}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1118 ( .a ({signal_2388, signal_1123}), .b ({signal_2387, signal_1127}), .c ({signal_2391, signal_833}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1119 ( .a ({signal_2113, signal_1138}), .b ({signal_2140, signal_836}), .c ({signal_2176, signal_1074}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1120 ( .a ({signal_2376, signal_1139}), .b ({signal_2392, signal_837}), .c ({signal_2399, signal_1075}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1121 ( .a ({signal_2106, signal_1148}), .b ({signal_2137, signal_838}), .c ({signal_2177, signal_1100}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1122 ( .a ({signal_2105, signal_1149}), .b ({signal_2138, signal_839}), .c ({signal_2178, signal_1101}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1123 ( .a ({signal_2104, signal_1150}), .b ({signal_2139, signal_840}), .c ({signal_2179, signal_1102}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1124 ( .a ({signal_2384, signal_1151}), .b ({signal_2393, signal_841}), .c ({signal_2400, signal_1103}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1125 ( .a ({signal_2109, signal_1144}), .b ({signal_2137, signal_838}), .c ({signal_2180, signal_1060}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1126 ( .a ({signal_2115, signal_1136}), .b ({signal_2112, signal_1140}), .c ({signal_2137, signal_838}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1127 ( .a ({signal_2108, signal_1145}), .b ({signal_2138, signal_839}), .c ({signal_2181, signal_1061}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1128 ( .a ({signal_2114, signal_1137}), .b ({signal_2111, signal_1141}), .c ({signal_2138, signal_839}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1129 ( .a ({signal_2107, signal_1146}), .b ({signal_2139, signal_840}), .c ({signal_2182, signal_1062}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1130 ( .a ({signal_2110, signal_1142}), .b ({signal_2113, signal_1138}), .c ({signal_2139, signal_840}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1131 ( .a ({signal_2112, signal_1140}), .b ({signal_2141, signal_842}), .c ({signal_2183, signal_1112}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1132 ( .a ({signal_2111, signal_1141}), .b ({signal_2142, signal_843}), .c ({signal_2184, signal_1113}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1133 ( .a ({signal_2110, signal_1142}), .b ({signal_2140, signal_836}), .c ({signal_2185, signal_1114}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1134 ( .a ({signal_2104, signal_1150}), .b ({signal_2107, signal_1146}), .c ({signal_2140, signal_836}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1135 ( .a ({signal_2385, signal_1143}), .b ({signal_2392, signal_837}), .c ({signal_2401, signal_1115}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1136 ( .a ({signal_2375, signal_1147}), .b ({signal_2384, signal_1151}), .c ({signal_2392, signal_837}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1137 ( .a ({signal_2115, signal_1136}), .b ({signal_2141, signal_842}), .c ({signal_2186, signal_1072}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1138 ( .a ({signal_2106, signal_1148}), .b ({signal_2109, signal_1144}), .c ({signal_2141, signal_842}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1139 ( .a ({signal_2114, signal_1137}), .b ({signal_2142, signal_843}), .c ({signal_2187, signal_1073}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1140 ( .a ({signal_2105, signal_1149}), .b ({signal_2108, signal_1145}), .c ({signal_2142, signal_843}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1141 ( .a ({signal_2375, signal_1147}), .b ({signal_2393, signal_841}), .c ({signal_2402, signal_1063}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1142 ( .a ({signal_2376, signal_1139}), .b ({signal_2385, signal_1143}), .c ({signal_2393, signal_841}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1143 ( .a ({signal_2101, signal_1154}), .b ({signal_2146, signal_844}), .c ({signal_2188, signal_1070}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1144 ( .a ({signal_2390, signal_1155}), .b ({signal_2394, signal_845}), .c ({signal_2403, signal_1071}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1145 ( .a ({signal_2095, signal_1164}), .b ({signal_2143, signal_846}), .c ({signal_2189, signal_1104}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1146 ( .a ({signal_2094, signal_1165}), .b ({signal_2144, signal_847}), .c ({signal_2190, signal_1105}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1147 ( .a ({signal_2093, signal_1166}), .b ({signal_2145, signal_848}), .c ({signal_2191, signal_1106}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1148 ( .a ({signal_2382, signal_1167}), .b ({signal_2405, signal_849}), .c ({signal_2423, signal_1107}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1149 ( .a ({signal_2098, signal_1160}), .b ({signal_2143, signal_846}), .c ({signal_2192, signal_1080}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1150 ( .a ({signal_2103, signal_1152}), .b ({signal_2100, signal_1156}), .c ({signal_2143, signal_846}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1151 ( .a ({signal_2097, signal_1161}), .b ({signal_2144, signal_847}), .c ({signal_2193, signal_1081}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1152 ( .a ({signal_2102, signal_1153}), .b ({signal_2089, signal_1157}), .c ({signal_2144, signal_847}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1153 ( .a ({signal_2096, signal_1162}), .b ({signal_2145, signal_848}), .c ({signal_2194, signal_1082}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1154 ( .a ({signal_2099, signal_1158}), .b ({signal_2101, signal_1154}), .c ({signal_2145, signal_848}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1155 ( .a ({signal_2100, signal_1156}), .b ({signal_2147, signal_850}), .c ({signal_2195, signal_1092}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1156 ( .a ({signal_2089, signal_1157}), .b ({signal_2148, signal_851}), .c ({signal_2196, signal_1093}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1157 ( .a ({signal_2099, signal_1158}), .b ({signal_2146, signal_844}), .c ({signal_2197, signal_1094}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1158 ( .a ({signal_2093, signal_1166}), .b ({signal_2096, signal_1162}), .c ({signal_2146, signal_844}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1159 ( .a ({signal_2383, signal_1159}), .b ({signal_2394, signal_845}), .c ({signal_2404, signal_1095}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1160 ( .a ({signal_2374, signal_1163}), .b ({signal_2382, signal_1167}), .c ({signal_2394, signal_845}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1161 ( .a ({signal_2103, signal_1152}), .b ({signal_2147, signal_850}), .c ({signal_2198, signal_1068}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1162 ( .a ({signal_2095, signal_1164}), .b ({signal_2098, signal_1160}), .c ({signal_2147, signal_850}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1163 ( .a ({signal_2102, signal_1153}), .b ({signal_2148, signal_851}), .c ({signal_2199, signal_1069}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1164 ( .a ({signal_2094, signal_1165}), .b ({signal_2097, signal_1161}), .c ({signal_2148, signal_851}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1165 ( .a ({signal_2374, signal_1163}), .b ({signal_2405, signal_849}), .c ({signal_2424, signal_1083}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1166 ( .a ({signal_2390, signal_1155}), .b ({signal_2383, signal_1159}), .c ({signal_2405, signal_849}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1167 ( .a ({signal_2086, signal_1170}), .b ({signal_2155, signal_852}), .c ({signal_2200, signal_1110}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1168 ( .a ({signal_2381, signal_1171}), .b ({signal_2395, signal_853}), .c ({signal_2406, signal_1111}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1169 ( .a ({signal_2082, signal_1180}), .b ({signal_2128, signal_854}), .c ({signal_2149, signal_1064}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1170 ( .a ({signal_2081, signal_1181}), .b ({signal_2129, signal_855}), .c ({signal_2150, signal_1065}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1171 ( .a ({signal_2080, signal_1182}), .b ({signal_2130, signal_856}), .c ({signal_2151, signal_1066}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1172 ( .a ({signal_2379, signal_1183}), .b ({signal_2396, signal_857}), .c ({signal_2407, signal_1067}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1173 ( .a ({signal_2092, signal_1176}), .b ({signal_2128, signal_854}), .c ({signal_2152, signal_1088}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1174 ( .a ({signal_2088, signal_1168}), .b ({signal_2085, signal_1172}), .c ({signal_2128, signal_854}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1175 ( .a ({signal_2091, signal_1177}), .b ({signal_2129, signal_855}), .c ({signal_2153, signal_1089}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1176 ( .a ({signal_2087, signal_1169}), .b ({signal_2084, signal_1173}), .c ({signal_2129, signal_855}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1177 ( .a ({signal_2090, signal_1178}), .b ({signal_2130, signal_856}), .c ({signal_2154, signal_1090}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1178 ( .a ({signal_2083, signal_1174}), .b ({signal_2086, signal_1170}), .c ({signal_2130, signal_856}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1179 ( .a ({signal_2085, signal_1172}), .b ({signal_2156, signal_858}), .c ({signal_2201, signal_1084}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1180 ( .a ({signal_2084, signal_1173}), .b ({signal_2157, signal_859}), .c ({signal_2202, signal_1085}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1181 ( .a ({signal_2083, signal_1174}), .b ({signal_2155, signal_852}), .c ({signal_2203, signal_1086}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1182 ( .a ({signal_2080, signal_1182}), .b ({signal_2090, signal_1178}), .c ({signal_2155, signal_852}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1183 ( .a ({signal_2373, signal_1175}), .b ({signal_2395, signal_853}), .c ({signal_2408, signal_1087}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1184 ( .a ({signal_2380, signal_1179}), .b ({signal_2379, signal_1183}), .c ({signal_2395, signal_853}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1185 ( .a ({signal_2088, signal_1168}), .b ({signal_2156, signal_858}), .c ({signal_2204, signal_1108}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1186 ( .a ({signal_2082, signal_1180}), .b ({signal_2092, signal_1176}), .c ({signal_2156, signal_858}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1187 ( .a ({signal_2087, signal_1169}), .b ({signal_2157, signal_859}), .c ({signal_2205, signal_1109}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1188 ( .a ({signal_2081, signal_1181}), .b ({signal_2091, signal_1177}), .c ({signal_2157, signal_859}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1189 ( .a ({signal_2380, signal_1179}), .b ({signal_2396, signal_857}), .c ({signal_2409, signal_1091}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1190 ( .a ({signal_2381, signal_1171}), .b ({signal_2373, signal_1175}), .c ({signal_2396, signal_857}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1191 ( .s (enc_dec), .b ({signal_2420, signal_1055}), .a ({signal_2398, signal_1119}), .c ({signal_2430, signal_1439}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1192 ( .s (enc_dec), .b ({signal_2163, signal_1054}), .a ({signal_2170, signal_1118}), .c ({signal_2248, signal_1438}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1193 ( .s (enc_dec), .b ({signal_2162, signal_1053}), .a ({signal_2169, signal_1117}), .c ({signal_2249, signal_1437}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1194 ( .s (enc_dec), .b ({signal_2161, signal_1052}), .a ({signal_2168, signal_1116}), .c ({signal_2250, signal_1436}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1195 ( .s (enc_dec), .b ({signal_2411, signal_1051}), .a ({signal_2401, signal_1115}), .c ({signal_2431, signal_1435}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1196 ( .s (enc_dec), .b ({signal_2160, signal_1050}), .a ({signal_2185, signal_1114}), .c ({signal_2251, signal_1434}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1197 ( .s (enc_dec), .b ({signal_2159, signal_1049}), .a ({signal_2184, signal_1113}), .c ({signal_2252, signal_1433}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1198 ( .s (enc_dec), .b ({signal_2158, signal_1048}), .a ({signal_2183, signal_1112}), .c ({signal_2253, signal_1432}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1199 ( .s (enc_dec), .b ({signal_2410, signal_1047}), .a ({signal_2406, signal_1111}), .c ({signal_2432, signal_1431}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1200 ( .s (enc_dec), .b ({signal_2206, signal_1046}), .a ({signal_2200, signal_1110}), .c ({signal_2264, signal_1430}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1201 ( .s (enc_dec), .b ({signal_2247, signal_1045}), .a ({signal_2205, signal_1109}), .c ({signal_2265, signal_1429}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1202 ( .s (enc_dec), .b ({signal_2246, signal_1044}), .a ({signal_2204, signal_1108}), .c ({signal_2266, signal_1428}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1203 ( .s (enc_dec), .b ({signal_2419, signal_1043}), .a ({signal_2423, signal_1107}), .c ({signal_2433, signal_1427}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1204 ( .s (enc_dec), .b ({signal_2245, signal_1042}), .a ({signal_2191, signal_1106}), .c ({signal_2267, signal_1426}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1205 ( .s (enc_dec), .b ({signal_2244, signal_1041}), .a ({signal_2190, signal_1105}), .c ({signal_2268, signal_1425}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1206 ( .s (enc_dec), .b ({signal_2243, signal_1040}), .a ({signal_2189, signal_1104}), .c ({signal_2269, signal_1424}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1207 ( .s (enc_dec), .b ({signal_2427, signal_1039}), .a ({signal_2400, signal_1103}), .c ({signal_2454, signal_1423}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1208 ( .s (enc_dec), .b ({signal_2242, signal_1038}), .a ({signal_2179, signal_1102}), .c ({signal_2270, signal_1422}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1209 ( .s (enc_dec), .b ({signal_2241, signal_1037}), .a ({signal_2178, signal_1101}), .c ({signal_2271, signal_1421}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1210 ( .s (enc_dec), .b ({signal_2240, signal_1036}), .a ({signal_2177, signal_1100}), .c ({signal_2272, signal_1420}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1211 ( .s (enc_dec), .b ({signal_2426, signal_1035}), .a ({signal_2428, signal_1099}), .c ({signal_2455, signal_1419}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1212 ( .s (enc_dec), .b ({signal_2239, signal_1034}), .a ({signal_2164, signal_1098}), .c ({signal_2273, signal_1418}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1213 ( .s (enc_dec), .b ({signal_2238, signal_1033}), .a ({signal_2175, signal_1097}), .c ({signal_2274, signal_1417}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1214 ( .s (enc_dec), .b ({signal_2237, signal_1032}), .a ({signal_2174, signal_1096}), .c ({signal_2275, signal_1416}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1215 ( .s (enc_dec), .b ({signal_2418, signal_1031}), .a ({signal_2404, signal_1095}), .c ({signal_2434, signal_1415}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1216 ( .s (enc_dec), .b ({signal_2236, signal_1030}), .a ({signal_2197, signal_1094}), .c ({signal_2276, signal_1414}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1217 ( .s (enc_dec), .b ({signal_2235, signal_1029}), .a ({signal_2196, signal_1093}), .c ({signal_2277, signal_1413}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1218 ( .s (enc_dec), .b ({signal_2234, signal_1028}), .a ({signal_2195, signal_1092}), .c ({signal_2278, signal_1412}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1219 ( .s (enc_dec), .b ({signal_2417, signal_1027}), .a ({signal_2409, signal_1091}), .c ({signal_2435, signal_1411}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1220 ( .s (enc_dec), .b ({signal_2233, signal_1026}), .a ({signal_2154, signal_1090}), .c ({signal_2279, signal_1410}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1221 ( .s (enc_dec), .b ({signal_2232, signal_1025}), .a ({signal_2153, signal_1089}), .c ({signal_2280, signal_1409}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1222 ( .s (enc_dec), .b ({signal_2231, signal_1024}), .a ({signal_2152, signal_1088}), .c ({signal_2281, signal_1408}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1223 ( .s (enc_dec), .b ({signal_2416, signal_1023}), .a ({signal_2408, signal_1087}), .c ({signal_2436, signal_1407}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1224 ( .s (enc_dec), .b ({signal_2230, signal_1022}), .a ({signal_2203, signal_1086}), .c ({signal_2282, signal_1406}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1225 ( .s (enc_dec), .b ({signal_2229, signal_1021}), .a ({signal_2202, signal_1085}), .c ({signal_2283, signal_1405}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1226 ( .s (enc_dec), .b ({signal_2228, signal_1020}), .a ({signal_2201, signal_1084}), .c ({signal_2284, signal_1404}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1227 ( .s (enc_dec), .b ({signal_2415, signal_1019}), .a ({signal_2424, signal_1083}), .c ({signal_2437, signal_1403}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1228 ( .s (enc_dec), .b ({signal_2227, signal_1018}), .a ({signal_2194, signal_1082}), .c ({signal_2285, signal_1402}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1229 ( .s (enc_dec), .b ({signal_2226, signal_1017}), .a ({signal_2193, signal_1081}), .c ({signal_2286, signal_1401}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1230 ( .s (enc_dec), .b ({signal_2225, signal_1016}), .a ({signal_2192, signal_1080}), .c ({signal_2287, signal_1400}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1231 ( .s (enc_dec), .b ({signal_2414, signal_1015}), .a ({signal_2421, signal_1079}), .c ({signal_2438, signal_1399}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1232 ( .s (enc_dec), .b ({signal_2224, signal_1014}), .a ({signal_2167, signal_1078}), .c ({signal_2288, signal_1398}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1233 ( .s (enc_dec), .b ({signal_2223, signal_1013}), .a ({signal_2166, signal_1077}), .c ({signal_2289, signal_1397}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1234 ( .s (enc_dec), .b ({signal_2222, signal_1012}), .a ({signal_2165, signal_1076}), .c ({signal_2290, signal_1396}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1235 ( .s (enc_dec), .b ({signal_2413, signal_1011}), .a ({signal_2399, signal_1075}), .c ({signal_2439, signal_1395}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1236 ( .s (enc_dec), .b ({signal_2221, signal_1010}), .a ({signal_2176, signal_1074}), .c ({signal_2291, signal_1394}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1237 ( .s (enc_dec), .b ({signal_2220, signal_1009}), .a ({signal_2187, signal_1073}), .c ({signal_2292, signal_1393}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1238 ( .s (enc_dec), .b ({signal_2219, signal_1008}), .a ({signal_2186, signal_1072}), .c ({signal_2293, signal_1392}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1239 ( .s (enc_dec), .b ({signal_2412, signal_1007}), .a ({signal_2403, signal_1071}), .c ({signal_2440, signal_1391}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1240 ( .s (enc_dec), .b ({signal_2218, signal_1006}), .a ({signal_2188, signal_1070}), .c ({signal_2294, signal_1390}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1241 ( .s (enc_dec), .b ({signal_2217, signal_1005}), .a ({signal_2199, signal_1069}), .c ({signal_2295, signal_1389}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1242 ( .s (enc_dec), .b ({signal_2216, signal_1004}), .a ({signal_2198, signal_1068}), .c ({signal_2296, signal_1388}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1243 ( .s (enc_dec), .b ({signal_2425, signal_1003}), .a ({signal_2407, signal_1067}), .c ({signal_2456, signal_1387}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1244 ( .s (enc_dec), .b ({signal_2215, signal_1002}), .a ({signal_2151, signal_1066}), .c ({signal_2297, signal_1386}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1245 ( .s (enc_dec), .b ({signal_2214, signal_1001}), .a ({signal_2150, signal_1065}), .c ({signal_2298, signal_1385}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1246 ( .s (enc_dec), .b ({signal_2213, signal_1000}), .a ({signal_2149, signal_1064}), .c ({signal_2299, signal_1384}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1247 ( .s (enc_dec), .b ({signal_2442, signal_999}), .a ({signal_2402, signal_1063}), .c ({signal_2460, signal_1383}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1248 ( .s (enc_dec), .b ({signal_2212, signal_998}), .a ({signal_2182, signal_1062}), .c ({signal_2300, signal_1382}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1249 ( .s (enc_dec), .b ({signal_2211, signal_997}), .a ({signal_2181, signal_1061}), .c ({signal_2301, signal_1381}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1250 ( .s (enc_dec), .b ({signal_2210, signal_996}), .a ({signal_2180, signal_1060}), .c ({signal_2302, signal_1380}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1251 ( .s (enc_dec), .b ({signal_2441, signal_995}), .a ({signal_2429, signal_1059}), .c ({signal_2461, signal_1379}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1252 ( .s (enc_dec), .b ({signal_2209, signal_994}), .a ({signal_2173, signal_1058}), .c ({signal_2303, signal_1378}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1253 ( .s (enc_dec), .b ({signal_2208, signal_993}), .a ({signal_2172, signal_1057}), .c ({signal_2304, signal_1377}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1254 ( .s (enc_dec), .b ({signal_2207, signal_992}), .a ({signal_2171, signal_1056}), .c ({signal_2305, signal_1376}) ) ;
    Midori64_step2_ANF #(.low_latency(0), .pipeline(0)) cell_1255 ( .in0 ({signal_1375, signal_1374, signal_1373, signal_1372, signal_1371, signal_1370, signal_1369, signal_1368, signal_1367, signal_1366, signal_1365, signal_1364, signal_1363, signal_1362, signal_1361, signal_1360, signal_1359, signal_1358, signal_1357, signal_1356, signal_1355, signal_1354, signal_1353, signal_1352, signal_1351, signal_1350, signal_1349, signal_1348, signal_1347, signal_1346, signal_1345, signal_1344, signal_1343, signal_1342, signal_1341, signal_1340, signal_1339, signal_1338, signal_1337, signal_1336, signal_1335, signal_1334, signal_1333, signal_1332, signal_1331, signal_1330, signal_1329, signal_1328, signal_1327, signal_1326, signal_1325, signal_1324, signal_1323, signal_1322, signal_1321, signal_1320, signal_1319, signal_1318, signal_1317, signal_1316, signal_1315, signal_1314, signal_1313, signal_1312}), .in1 ({signal_1852, signal_1851, signal_1850, signal_1849, signal_1848, signal_1847, signal_1846, signal_1845, signal_1844, signal_1843, signal_1842, signal_1841, signal_1840, signal_1839, signal_1838, signal_1837, signal_1836, signal_1835, signal_1834, signal_1833, signal_1832, signal_1831, signal_1830, signal_1829, signal_1828, signal_1827, signal_1826, signal_1825, signal_1824, signal_1823, signal_1822, signal_1821, signal_1820, signal_1819, signal_1818, signal_1817, signal_1816, signal_1815, signal_1814, signal_1813, signal_1812, signal_1811, signal_1810, signal_1809, signal_1808, signal_1807, signal_1806, signal_1805, signal_1804, signal_1803, signal_1802, signal_1801, signal_1800, signal_1799, signal_1798, signal_1797, signal_1796, signal_1795, signal_1794, signal_1793, signal_1792, signal_1791, signal_1790, signal_1789}), .clk (clk), .r ({Fresh[63], Fresh[62], Fresh[61], Fresh[60], Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48], Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30], Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .out0 ({signal_1311, signal_1310, signal_1309, signal_1308, signal_1307, signal_1306, signal_1305, signal_1304, signal_1303, signal_1302, signal_1301, signal_1300, signal_1299, signal_1298, signal_1297, signal_1296, signal_1295, signal_1294, signal_1293, signal_1292, signal_1291, signal_1290, signal_1289, signal_1288, signal_1287, signal_1286, signal_1285, signal_1284, signal_1283, signal_1282, signal_1281, signal_1280, signal_1279, signal_1278, signal_1277, signal_1276, signal_1275, signal_1274, signal_1273, signal_1272, signal_1271, signal_1270, signal_1269, signal_1268, signal_1267, signal_1266, signal_1265, signal_1264, signal_1263, signal_1262, signal_1261, signal_1260, signal_1259, signal_1258, signal_1257, signal_1256, signal_1255, signal_1254, signal_1253, signal_1252, signal_1251, signal_1250, signal_1249, signal_1248}), .out1 ({signal_1916, signal_1915, signal_1914, signal_1913, signal_1912, signal_1911, signal_1910, signal_1909, signal_1908, signal_1907, signal_1906, signal_1905, signal_1904, signal_1903, signal_1902, signal_1901, signal_1900, signal_1899, signal_1898, signal_1897, signal_1896, signal_1895, signal_1894, signal_1893, signal_1892, signal_1891, signal_1890, signal_1889, signal_1888, signal_1887, signal_1886, signal_1885, signal_1884, signal_1883, signal_1882, signal_1881, signal_1880, signal_1879, signal_1878, signal_1877, signal_1876, signal_1875, signal_1874, signal_1873, signal_1872, signal_1871, signal_1870, signal_1869, signal_1868, signal_1867, signal_1866, signal_1865, signal_1864, signal_1863, signal_1862, signal_1861, signal_1860, signal_1859, signal_1858, signal_1857, signal_1856, signal_1855, signal_1854, signal_1853}) ) ;

    /* register cells */
    DFF_X1 cell_82 ( .CK (signal_2528), .D (signal_283), .Q (signal_927), .QN () ) ;
    DFF_X1 cell_84 ( .CK (signal_2528), .D (signal_282), .Q (signal_926), .QN () ) ;
    DFF_X1 cell_86 ( .CK (signal_2528), .D (signal_278), .Q (signal_925), .QN () ) ;
    DFF_X1 cell_88 ( .CK (signal_2528), .D (signal_280), .Q (signal_924), .QN () ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_537 ( .clk (signal_2528), .D ({signal_2443, signal_460}), .Q ({signal_1852, signal_1375}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_540 ( .clk (signal_2528), .D ({signal_2258, signal_462}), .Q ({signal_1851, signal_1374}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_543 ( .clk (signal_2528), .D ({signal_2259, signal_464}), .Q ({signal_1850, signal_1373}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_546 ( .clk (signal_2528), .D ({signal_2260, signal_466}), .Q ({signal_1849, signal_1372}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_549 ( .clk (signal_2528), .D ({signal_2444, signal_468}), .Q ({signal_1848, signal_1371}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_552 ( .clk (signal_2528), .D ({signal_2261, signal_470}), .Q ({signal_1847, signal_1370}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_555 ( .clk (signal_2528), .D ({signal_2262, signal_472}), .Q ({signal_1846, signal_1369}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_558 ( .clk (signal_2528), .D ({signal_2263, signal_474}), .Q ({signal_1845, signal_1368}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_561 ( .clk (signal_2528), .D ({signal_2445, signal_476}), .Q ({signal_1844, signal_1367}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_564 ( .clk (signal_2528), .D ({signal_2320, signal_478}), .Q ({signal_1843, signal_1366}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_567 ( .clk (signal_2528), .D ({signal_2321, signal_480}), .Q ({signal_1842, signal_1365}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_570 ( .clk (signal_2528), .D ({signal_2322, signal_482}), .Q ({signal_1841, signal_1364}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_573 ( .clk (signal_2528), .D ({signal_2446, signal_484}), .Q ({signal_1840, signal_1363}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_576 ( .clk (signal_2528), .D ({signal_2323, signal_486}), .Q ({signal_1839, signal_1362}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_579 ( .clk (signal_2528), .D ({signal_2324, signal_488}), .Q ({signal_1838, signal_1361}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_582 ( .clk (signal_2528), .D ({signal_2325, signal_490}), .Q ({signal_1837, signal_1360}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_585 ( .clk (signal_2528), .D ({signal_2457, signal_492}), .Q ({signal_1836, signal_1359}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_588 ( .clk (signal_2528), .D ({signal_2326, signal_494}), .Q ({signal_1835, signal_1358}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_591 ( .clk (signal_2528), .D ({signal_2327, signal_496}), .Q ({signal_1834, signal_1357}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_594 ( .clk (signal_2528), .D ({signal_2328, signal_498}), .Q ({signal_1833, signal_1356}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_597 ( .clk (signal_2528), .D ({signal_2458, signal_500}), .Q ({signal_1832, signal_1355}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_600 ( .clk (signal_2528), .D ({signal_2329, signal_502}), .Q ({signal_1831, signal_1354}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_603 ( .clk (signal_2528), .D ({signal_2330, signal_504}), .Q ({signal_1830, signal_1353}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_606 ( .clk (signal_2528), .D ({signal_2331, signal_506}), .Q ({signal_1829, signal_1352}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_609 ( .clk (signal_2528), .D ({signal_2447, signal_508}), .Q ({signal_1828, signal_1351}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_612 ( .clk (signal_2528), .D ({signal_2332, signal_510}), .Q ({signal_1827, signal_1350}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_615 ( .clk (signal_2528), .D ({signal_2333, signal_512}), .Q ({signal_1826, signal_1349}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_618 ( .clk (signal_2528), .D ({signal_2334, signal_514}), .Q ({signal_1825, signal_1348}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_621 ( .clk (signal_2528), .D ({signal_2448, signal_516}), .Q ({signal_1824, signal_1347}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_624 ( .clk (signal_2528), .D ({signal_2335, signal_518}), .Q ({signal_1823, signal_1346}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_627 ( .clk (signal_2528), .D ({signal_2336, signal_520}), .Q ({signal_1822, signal_1345}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_630 ( .clk (signal_2528), .D ({signal_2337, signal_522}), .Q ({signal_1821, signal_1344}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_633 ( .clk (signal_2528), .D ({signal_2449, signal_524}), .Q ({signal_1820, signal_1343}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_636 ( .clk (signal_2528), .D ({signal_2338, signal_526}), .Q ({signal_1819, signal_1342}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_639 ( .clk (signal_2528), .D ({signal_2339, signal_528}), .Q ({signal_1818, signal_1341}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_642 ( .clk (signal_2528), .D ({signal_2340, signal_530}), .Q ({signal_1817, signal_1340}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_645 ( .clk (signal_2528), .D ({signal_2450, signal_532}), .Q ({signal_1816, signal_1339}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_648 ( .clk (signal_2528), .D ({signal_2341, signal_534}), .Q ({signal_1815, signal_1338}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_651 ( .clk (signal_2528), .D ({signal_2342, signal_536}), .Q ({signal_1814, signal_1337}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_654 ( .clk (signal_2528), .D ({signal_2343, signal_538}), .Q ({signal_1813, signal_1336}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_657 ( .clk (signal_2528), .D ({signal_2451, signal_540}), .Q ({signal_1812, signal_1335}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_660 ( .clk (signal_2528), .D ({signal_2344, signal_542}), .Q ({signal_1811, signal_1334}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_663 ( .clk (signal_2528), .D ({signal_2345, signal_544}), .Q ({signal_1810, signal_1333}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_666 ( .clk (signal_2528), .D ({signal_2346, signal_546}), .Q ({signal_1809, signal_1332}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_669 ( .clk (signal_2528), .D ({signal_2452, signal_548}), .Q ({signal_1808, signal_1331}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_672 ( .clk (signal_2528), .D ({signal_2347, signal_550}), .Q ({signal_1807, signal_1330}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_675 ( .clk (signal_2528), .D ({signal_2348, signal_552}), .Q ({signal_1806, signal_1329}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_678 ( .clk (signal_2528), .D ({signal_2349, signal_554}), .Q ({signal_1805, signal_1328}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_681 ( .clk (signal_2528), .D ({signal_2453, signal_556}), .Q ({signal_1804, signal_1327}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_684 ( .clk (signal_2528), .D ({signal_2350, signal_558}), .Q ({signal_1803, signal_1326}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_687 ( .clk (signal_2528), .D ({signal_2351, signal_560}), .Q ({signal_1802, signal_1325}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_690 ( .clk (signal_2528), .D ({signal_2352, signal_562}), .Q ({signal_1801, signal_1324}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_693 ( .clk (signal_2528), .D ({signal_2459, signal_564}), .Q ({signal_1800, signal_1323}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_696 ( .clk (signal_2528), .D ({signal_2353, signal_566}), .Q ({signal_1799, signal_1322}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_699 ( .clk (signal_2528), .D ({signal_2354, signal_568}), .Q ({signal_1798, signal_1321}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_702 ( .clk (signal_2528), .D ({signal_2355, signal_570}), .Q ({signal_1797, signal_1320}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_705 ( .clk (signal_2528), .D ({signal_2462, signal_572}), .Q ({signal_1796, signal_1319}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_708 ( .clk (signal_2528), .D ({signal_2356, signal_574}), .Q ({signal_1795, signal_1318}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_711 ( .clk (signal_2528), .D ({signal_2357, signal_576}), .Q ({signal_1794, signal_1317}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_714 ( .clk (signal_2528), .D ({signal_2358, signal_578}), .Q ({signal_1793, signal_1316}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_717 ( .clk (signal_2528), .D ({signal_2463, signal_580}), .Q ({signal_1792, signal_1315}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_720 ( .clk (signal_2528), .D ({signal_2359, signal_582}), .Q ({signal_1791, signal_1314}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_723 ( .clk (signal_2528), .D ({signal_2360, signal_584}), .Q ({signal_1790, signal_1313}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_726 ( .clk (signal_2528), .D ({signal_2361, signal_586}), .Q ({signal_1789, signal_1312}) ) ;
endmodule
