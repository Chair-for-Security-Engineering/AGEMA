/* modified netlist. Source: module sbox in file Designs/AESSbox//Canright/AGEMA/sbox.v */
/* clock gating is added to the circuit, the latency increased 16 time(s)  */

module sbox_HPC2_AIG_ClockGating_d4 (X_s0, clk, X_s1, X_s2, X_s3, X_s4, Fresh, rst, Y_s0, Y_s1, Y_s2, Y_s3, Y_s4, Synch);
    input [7:0] X_s0 ;
    input clk ;
    input [7:0] X_s1 ;
    input [7:0] X_s2 ;
    input [7:0] X_s3 ;
    input [7:0] X_s4 ;
    input rst ;
    input [879:0] Fresh ;
    output [7:0] Y_s0 ;
    output [7:0] Y_s1 ;
    output [7:0] Y_s2 ;
    output [7:0] Y_s3 ;
    output [7:0] Y_s4 ;
    output Synch ;
    wire signal_160 ;
    wire signal_161 ;
    wire signal_162 ;
    wire signal_163 ;
    wire signal_164 ;
    wire signal_165 ;
    wire signal_166 ;
    wire signal_167 ;
    wire signal_192 ;
    wire signal_193 ;
    wire signal_194 ;
    wire signal_195 ;
    wire signal_196 ;
    wire signal_197 ;
    wire signal_198 ;
    wire signal_199 ;
    wire signal_200 ;
    wire signal_201 ;
    wire signal_202 ;
    wire signal_203 ;
    wire signal_204 ;
    wire signal_205 ;
    wire signal_206 ;
    wire signal_207 ;
    wire signal_208 ;
    wire signal_209 ;
    wire signal_210 ;
    wire signal_211 ;
    wire signal_212 ;
    wire signal_213 ;
    wire signal_214 ;
    wire signal_215 ;
    wire signal_216 ;
    wire signal_217 ;
    wire signal_218 ;
    wire signal_219 ;
    wire signal_220 ;
    wire signal_221 ;
    wire signal_222 ;
    wire signal_223 ;
    wire signal_224 ;
    wire signal_225 ;
    wire signal_226 ;
    wire signal_227 ;
    wire signal_228 ;
    wire signal_229 ;
    wire signal_230 ;
    wire signal_231 ;
    wire signal_232 ;
    wire signal_233 ;
    wire signal_234 ;
    wire signal_235 ;
    wire signal_236 ;
    wire signal_237 ;
    wire signal_238 ;
    wire signal_239 ;
    wire signal_240 ;
    wire signal_241 ;
    wire signal_242 ;
    wire signal_243 ;
    wire signal_244 ;
    wire signal_245 ;
    wire signal_246 ;
    wire signal_247 ;
    wire signal_248 ;
    wire signal_249 ;
    wire signal_250 ;
    wire signal_251 ;
    wire signal_252 ;
    wire signal_253 ;
    wire signal_254 ;
    wire signal_255 ;
    wire signal_256 ;
    wire signal_257 ;
    wire signal_258 ;
    wire signal_259 ;
    wire signal_260 ;
    wire signal_261 ;
    wire signal_262 ;
    wire signal_263 ;
    wire signal_264 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_285 ;
    wire signal_286 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_295 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_352 ;
    wire signal_353 ;
    wire signal_354 ;
    wire signal_355 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_359 ;
    wire signal_360 ;
    wire signal_361 ;
    wire signal_362 ;
    wire signal_363 ;
    wire signal_364 ;
    wire signal_365 ;
    wire signal_366 ;
    wire signal_367 ;
    wire signal_368 ;
    wire signal_369 ;
    wire signal_370 ;
    wire signal_371 ;
    wire signal_372 ;
    wire signal_373 ;
    wire signal_374 ;
    wire signal_375 ;
    wire signal_376 ;
    wire signal_377 ;
    wire signal_378 ;
    wire signal_379 ;
    wire signal_380 ;
    wire signal_381 ;
    wire signal_382 ;
    wire signal_383 ;
    wire signal_384 ;
    wire signal_385 ;
    wire signal_386 ;
    wire signal_387 ;
    wire signal_388 ;
    wire signal_389 ;
    wire signal_390 ;
    wire signal_391 ;
    wire signal_392 ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_415 ;
    wire signal_416 ;
    wire signal_417 ;
    wire signal_418 ;
    wire signal_419 ;
    wire signal_420 ;
    wire signal_421 ;
    wire signal_422 ;
    wire signal_423 ;
    wire signal_424 ;
    wire signal_425 ;
    wire signal_426 ;
    wire signal_427 ;
    wire signal_428 ;
    wire signal_429 ;
    wire signal_430 ;
    wire signal_431 ;
    wire signal_432 ;
    wire signal_433 ;
    wire signal_434 ;
    wire signal_435 ;
    wire signal_436 ;
    wire signal_441 ;
    wire signal_442 ;
    wire signal_443 ;
    wire signal_444 ;
    wire signal_453 ;
    wire signal_454 ;
    wire signal_455 ;
    wire signal_456 ;
    wire signal_465 ;
    wire signal_466 ;
    wire signal_467 ;
    wire signal_468 ;
    wire signal_469 ;
    wire signal_470 ;
    wire signal_471 ;
    wire signal_472 ;
    wire signal_473 ;
    wire signal_474 ;
    wire signal_475 ;
    wire signal_476 ;
    wire signal_481 ;
    wire signal_482 ;
    wire signal_483 ;
    wire signal_484 ;
    wire signal_485 ;
    wire signal_486 ;
    wire signal_487 ;
    wire signal_488 ;
    wire signal_489 ;
    wire signal_490 ;
    wire signal_491 ;
    wire signal_492 ;
    wire signal_493 ;
    wire signal_494 ;
    wire signal_495 ;
    wire signal_496 ;
    wire signal_497 ;
    wire signal_498 ;
    wire signal_499 ;
    wire signal_500 ;
    wire signal_505 ;
    wire signal_506 ;
    wire signal_507 ;
    wire signal_508 ;
    wire signal_509 ;
    wire signal_510 ;
    wire signal_511 ;
    wire signal_512 ;
    wire signal_517 ;
    wire signal_518 ;
    wire signal_519 ;
    wire signal_520 ;
    wire signal_521 ;
    wire signal_522 ;
    wire signal_523 ;
    wire signal_524 ;
    wire signal_525 ;
    wire signal_526 ;
    wire signal_527 ;
    wire signal_528 ;
    wire signal_529 ;
    wire signal_530 ;
    wire signal_531 ;
    wire signal_532 ;
    wire signal_533 ;
    wire signal_534 ;
    wire signal_535 ;
    wire signal_536 ;
    wire signal_537 ;
    wire signal_538 ;
    wire signal_539 ;
    wire signal_540 ;
    wire signal_541 ;
    wire signal_542 ;
    wire signal_543 ;
    wire signal_544 ;
    wire signal_545 ;
    wire signal_546 ;
    wire signal_547 ;
    wire signal_548 ;
    wire signal_549 ;
    wire signal_550 ;
    wire signal_551 ;
    wire signal_552 ;
    wire signal_553 ;
    wire signal_554 ;
    wire signal_555 ;
    wire signal_556 ;
    wire signal_557 ;
    wire signal_558 ;
    wire signal_559 ;
    wire signal_560 ;
    wire signal_561 ;
    wire signal_562 ;
    wire signal_563 ;
    wire signal_564 ;
    wire signal_565 ;
    wire signal_566 ;
    wire signal_567 ;
    wire signal_568 ;
    wire signal_569 ;
    wire signal_570 ;
    wire signal_571 ;
    wire signal_572 ;
    wire signal_573 ;
    wire signal_574 ;
    wire signal_575 ;
    wire signal_576 ;
    wire signal_577 ;
    wire signal_578 ;
    wire signal_579 ;
    wire signal_580 ;
    wire signal_581 ;
    wire signal_582 ;
    wire signal_583 ;
    wire signal_584 ;
    wire signal_585 ;
    wire signal_586 ;
    wire signal_587 ;
    wire signal_588 ;
    wire signal_589 ;
    wire signal_590 ;
    wire signal_591 ;
    wire signal_592 ;
    wire signal_593 ;
    wire signal_594 ;
    wire signal_595 ;
    wire signal_596 ;
    wire signal_597 ;
    wire signal_598 ;
    wire signal_599 ;
    wire signal_600 ;
    wire signal_601 ;
    wire signal_602 ;
    wire signal_603 ;
    wire signal_604 ;
    wire signal_605 ;
    wire signal_606 ;
    wire signal_607 ;
    wire signal_608 ;
    wire signal_609 ;
    wire signal_610 ;
    wire signal_611 ;
    wire signal_612 ;
    wire signal_613 ;
    wire signal_614 ;
    wire signal_615 ;
    wire signal_616 ;
    wire signal_617 ;
    wire signal_618 ;
    wire signal_619 ;
    wire signal_620 ;
    wire signal_621 ;
    wire signal_622 ;
    wire signal_623 ;
    wire signal_624 ;
    wire signal_625 ;
    wire signal_626 ;
    wire signal_627 ;
    wire signal_628 ;
    wire signal_629 ;
    wire signal_630 ;
    wire signal_631 ;
    wire signal_632 ;
    wire signal_633 ;
    wire signal_634 ;
    wire signal_635 ;
    wire signal_636 ;
    wire signal_637 ;
    wire signal_638 ;
    wire signal_639 ;
    wire signal_640 ;
    wire signal_641 ;
    wire signal_642 ;
    wire signal_643 ;
    wire signal_644 ;
    wire signal_645 ;
    wire signal_646 ;
    wire signal_647 ;
    wire signal_648 ;
    wire signal_649 ;
    wire signal_650 ;
    wire signal_651 ;
    wire signal_652 ;
    wire signal_653 ;
    wire signal_654 ;
    wire signal_655 ;
    wire signal_656 ;
    wire signal_657 ;
    wire signal_658 ;
    wire signal_659 ;
    wire signal_660 ;
    wire signal_661 ;
    wire signal_662 ;
    wire signal_663 ;
    wire signal_664 ;
    wire signal_665 ;
    wire signal_666 ;
    wire signal_667 ;
    wire signal_668 ;
    wire signal_669 ;
    wire signal_670 ;
    wire signal_671 ;
    wire signal_672 ;
    wire signal_673 ;
    wire signal_674 ;
    wire signal_675 ;
    wire signal_676 ;
    wire signal_677 ;
    wire signal_678 ;
    wire signal_679 ;
    wire signal_680 ;
    wire signal_681 ;
    wire signal_682 ;
    wire signal_683 ;
    wire signal_684 ;
    wire signal_685 ;
    wire signal_686 ;
    wire signal_687 ;
    wire signal_688 ;
    wire signal_689 ;
    wire signal_690 ;
    wire signal_691 ;
    wire signal_692 ;
    wire signal_693 ;
    wire signal_694 ;
    wire signal_695 ;
    wire signal_696 ;
    wire signal_697 ;
    wire signal_698 ;
    wire signal_699 ;
    wire signal_700 ;
    wire signal_701 ;
    wire signal_702 ;
    wire signal_703 ;
    wire signal_704 ;
    wire signal_705 ;
    wire signal_706 ;
    wire signal_707 ;
    wire signal_708 ;
    wire signal_709 ;
    wire signal_710 ;
    wire signal_711 ;
    wire signal_712 ;
    wire signal_713 ;
    wire signal_714 ;
    wire signal_715 ;
    wire signal_716 ;
    wire signal_717 ;
    wire signal_718 ;
    wire signal_719 ;
    wire signal_720 ;
    wire signal_721 ;
    wire signal_722 ;
    wire signal_723 ;
    wire signal_724 ;
    wire signal_725 ;
    wire signal_726 ;
    wire signal_727 ;
    wire signal_728 ;
    wire signal_729 ;
    wire signal_730 ;
    wire signal_731 ;
    wire signal_732 ;
    wire signal_733 ;
    wire signal_734 ;
    wire signal_735 ;
    wire signal_736 ;
    wire signal_737 ;
    wire signal_738 ;
    wire signal_739 ;
    wire signal_740 ;
    wire signal_741 ;
    wire signal_742 ;
    wire signal_743 ;
    wire signal_744 ;
    wire signal_745 ;
    wire signal_746 ;
    wire signal_747 ;
    wire signal_748 ;
    wire signal_749 ;
    wire signal_750 ;
    wire signal_751 ;
    wire signal_752 ;
    wire signal_753 ;
    wire signal_754 ;
    wire signal_755 ;
    wire signal_756 ;
    wire signal_757 ;
    wire signal_758 ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_768 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_771 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_774 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_777 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_780 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_783 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_786 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_789 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_792 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_809 ;
    wire signal_810 ;
    wire signal_811 ;
    wire signal_812 ;
    wire signal_813 ;
    wire signal_814 ;
    wire signal_815 ;
    wire signal_816 ;
    wire signal_817 ;
    wire signal_818 ;
    wire signal_819 ;
    wire signal_820 ;
    wire signal_821 ;
    wire signal_822 ;
    wire signal_823 ;
    wire signal_824 ;
    wire signal_825 ;
    wire signal_826 ;
    wire signal_827 ;
    wire signal_828 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_831 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_834 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_837 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_840 ;
    wire signal_841 ;
    wire signal_842 ;
    wire signal_843 ;
    wire signal_844 ;
    wire signal_845 ;
    wire signal_846 ;
    wire signal_847 ;
    wire signal_848 ;
    wire signal_849 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_852 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_855 ;
    wire signal_856 ;
    wire signal_857 ;
    wire signal_858 ;
    wire signal_859 ;
    wire signal_860 ;
    wire signal_861 ;
    wire signal_862 ;
    wire signal_863 ;
    wire signal_864 ;
    wire signal_865 ;
    wire signal_866 ;
    wire signal_867 ;
    wire signal_868 ;
    wire signal_869 ;
    wire signal_870 ;
    wire signal_871 ;
    wire signal_872 ;
    wire signal_873 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_879 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_885 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_888 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_891 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_894 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_897 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_900 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_903 ;
    wire signal_904 ;
    wire signal_905 ;
    wire signal_906 ;
    wire signal_907 ;
    wire signal_908 ;
    wire signal_909 ;
    wire signal_910 ;
    wire signal_911 ;
    wire signal_912 ;
    wire signal_913 ;
    wire signal_914 ;
    wire signal_915 ;
    wire signal_916 ;
    wire signal_917 ;
    wire signal_918 ;
    wire signal_919 ;
    wire signal_920 ;
    wire signal_921 ;
    wire signal_922 ;
    wire signal_923 ;
    wire signal_924 ;
    wire signal_925 ;
    wire signal_926 ;
    wire signal_927 ;
    wire signal_928 ;
    wire signal_929 ;
    wire signal_930 ;
    wire signal_931 ;
    wire signal_932 ;
    wire signal_933 ;
    wire signal_934 ;
    wire signal_935 ;
    wire signal_936 ;
    wire signal_937 ;
    wire signal_938 ;
    wire signal_939 ;
    wire signal_940 ;
    wire signal_941 ;
    wire signal_942 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1020 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1023 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1276 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1279 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1282 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1285 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1288 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1294 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1297 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1300 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1303 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1309 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_2390 ;

    /* cells in depth 0 */
    not_masked #(.security_order(4), .pipeline(0)) cell_176 ( .a ({X_s4[0], X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({signal_444, signal_443, signal_442, signal_441, signal_192}) ) ;
    INV_X1 cell_177 ( .A ( 1'b1 ), .ZN ( signal_193 ) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_178 ( .a ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .c ({signal_456, signal_455, signal_454, signal_453, signal_194}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_179 ( .a ({X_s4[7], X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s4[5], X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .c ({signal_468, signal_467, signal_466, signal_465, signal_195}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_180 ( .a ({X_s4[7], X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .c ({signal_472, signal_471, signal_470, signal_469, signal_196}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_181 ( .a ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({X_s4[0], X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .c ({signal_476, signal_475, signal_474, signal_473, signal_197}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_182 ( .a ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({X_s4[0], X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .c ({signal_484, signal_483, signal_482, signal_481, signal_198}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_183 ( .a ({signal_472, signal_471, signal_470, signal_469, signal_196}), .b ({signal_488, signal_487, signal_486, signal_485, signal_199}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_186 ( .a ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_472, signal_471, signal_470, signal_469, signal_196}), .c ({signal_500, signal_499, signal_498, signal_497, signal_202}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_187 ( .a ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_468, signal_467, signal_466, signal_465, signal_195}), .c ({signal_508, signal_507, signal_506, signal_505, signal_203}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_188 ( .a ({signal_468, signal_467, signal_466, signal_465, signal_195}), .b ({signal_476, signal_475, signal_474, signal_473, signal_197}), .c ({signal_512, signal_511, signal_510, signal_509, signal_204}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_189 ( .a ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_476, signal_475, signal_474, signal_473, signal_197}), .c ({signal_520, signal_519, signal_518, signal_517, signal_205}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_190 ( .a ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_484, signal_483, signal_482, signal_481, signal_198}), .c ({signal_524, signal_523, signal_522, signal_521, signal_206}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_191 ( .a ({X_s4[5], X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_476, signal_475, signal_474, signal_473, signal_197}), .c ({signal_528, signal_527, signal_526, signal_525, signal_207}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_192 ( .a ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_484, signal_483, signal_482, signal_481, signal_198}), .c ({signal_532, signal_531, signal_530, signal_529, signal_208}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_193 ( .a ({signal_512, signal_511, signal_510, signal_509, signal_204}), .b ({signal_536, signal_535, signal_534, signal_533, signal_209}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_194 ( .a ({signal_528, signal_527, signal_526, signal_525, signal_207}), .b ({signal_540, signal_539, signal_538, signal_537, signal_210}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_201 ( .a ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_528, signal_527, signal_526, signal_525, signal_207}), .c ({signal_568, signal_567, signal_566, signal_565, signal_217}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_202 ( .a ({signal_508, signal_507, signal_506, signal_505, signal_203}), .b ({signal_520, signal_519, signal_518, signal_517, signal_205}), .c ({signal_572, signal_571, signal_570, signal_569, signal_218}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_203 ( .a ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_520, signal_519, signal_518, signal_517, signal_205}), .c ({signal_576, signal_575, signal_574, signal_573, signal_219}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_204 ( .a ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_520, signal_519, signal_518, signal_517, signal_205}), .c ({signal_580, signal_579, signal_578, signal_577, signal_220}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_205 ( .a ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_528, signal_527, signal_526, signal_525, signal_207}), .c ({signal_584, signal_583, signal_582, signal_581, signal_221}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_206 ( .a ({signal_472, signal_471, signal_470, signal_469, signal_196}), .b ({signal_532, signal_531, signal_530, signal_529, signal_208}), .c ({signal_588, signal_587, signal_586, signal_585, signal_222}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_208 ( .a ({signal_568, signal_567, signal_566, signal_565, signal_217}), .b ({signal_596, signal_595, signal_594, signal_593, signal_224}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_209 ( .a ({signal_572, signal_571, signal_570, signal_569, signal_218}), .b ({signal_600, signal_599, signal_598, signal_597, signal_225}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_210 ( .a ({signal_584, signal_583, signal_582, signal_581, signal_221}), .b ({signal_604, signal_603, signal_602, signal_601, signal_226}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_211 ( .a ({signal_588, signal_587, signal_586, signal_585, signal_222}), .b ({signal_608, signal_607, signal_606, signal_605, signal_227}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_219 ( .a ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_580, signal_579, signal_578, signal_577, signal_220}), .c ({signal_640, signal_639, signal_638, signal_637, signal_235}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_220 ( .a ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_584, signal_583, signal_582, signal_581, signal_221}), .c ({signal_644, signal_643, signal_642, signal_641, signal_236}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_222 ( .a ({signal_640, signal_639, signal_638, signal_637, signal_235}), .b ({signal_652, signal_651, signal_650, signal_649, signal_238}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_223 ( .a ({signal_644, signal_643, signal_642, signal_641, signal_236}), .b ({signal_656, signal_655, signal_654, signal_653, signal_239}) ) ;
    ClockGatingController #(17) cell_429 ( .clk ( clk ), .rst ( rst ), .GatedClk ( signal_2390 ), .Synch ( Synch ) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_184 ( .a ({signal_444, signal_443, signal_442, signal_441, signal_192}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({signal_492, signal_491, signal_490, signal_489, signal_200}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_185 ( .a ({1'b0, 1'b0, 1'b0, 1'b0, signal_193}), .b ({signal_456, signal_455, signal_454, signal_453, signal_194}), .clk ( clk ), .r ({Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10]}), .c ({signal_496, signal_495, signal_494, signal_493, signal_201}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_195 ( .a ({signal_492, signal_491, signal_490, signal_489, signal_200}), .b ({signal_544, signal_543, signal_542, signal_541, signal_211}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_196 ( .a ({signal_496, signal_495, signal_494, signal_493, signal_201}), .b ({signal_548, signal_547, signal_546, signal_545, signal_212}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_197 ( .a ({1'b0, 1'b0, 1'b0, 1'b0, signal_193}), .b ({signal_508, signal_507, signal_506, signal_505, signal_203}), .clk ( clk ), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20]}), .c ({signal_552, signal_551, signal_550, signal_549, signal_213}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_198 ( .a ({1'b0, 1'b0, 1'b0, 1'b0, signal_193}), .b ({signal_524, signal_523, signal_522, signal_521, signal_206}), .clk ( clk ), .r ({Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({signal_556, signal_555, signal_554, signal_553, signal_214}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_199 ( .a ({1'b0, 1'b0, 1'b0, 1'b0, signal_193}), .b ({signal_488, signal_487, signal_486, signal_485, signal_199}), .clk ( clk ), .r ({Fresh[49], Fresh[48], Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40]}), .c ({signal_560, signal_559, signal_558, signal_557, signal_215}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_200 ( .a ({1'b0, 1'b0, 1'b0, 1'b0, signal_193}), .b ({signal_500, signal_499, signal_498, signal_497, signal_202}), .clk ( clk ), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50]}), .c ({signal_564, signal_563, signal_562, signal_561, signal_216}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_207 ( .a ({signal_552, signal_551, signal_550, signal_549, signal_213}), .b ({signal_592, signal_591, signal_590, signal_589, signal_223}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_212 ( .a ({signal_556, signal_555, signal_554, signal_553, signal_214}), .b ({signal_612, signal_611, signal_610, signal_609, signal_228}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_213 ( .a ({signal_560, signal_559, signal_558, signal_557, signal_215}), .b ({signal_616, signal_615, signal_614, signal_613, signal_229}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_214 ( .a ({signal_564, signal_563, signal_562, signal_561, signal_216}), .b ({signal_620, signal_619, signal_618, signal_617, signal_230}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_215 ( .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .b ({signal_540, signal_539, signal_538, signal_537, signal_210}), .clk ( clk ), .r ({Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({signal_624, signal_623, signal_622, signal_621, signal_231}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_216 ( .a ({1'b0, 1'b0, 1'b0, 1'b0, signal_193}), .b ({signal_576, signal_575, signal_574, signal_573, signal_219}), .clk ( clk ), .r ({Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72], Fresh[71], Fresh[70]}), .c ({signal_628, signal_627, signal_626, signal_625, signal_232}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_217 ( .a ({1'b0, 1'b0, 1'b0, 1'b0, signal_193}), .b ({signal_580, signal_579, signal_578, signal_577, signal_220}), .clk ( clk ), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84], Fresh[83], Fresh[82], Fresh[81], Fresh[80]}), .c ({signal_632, signal_631, signal_630, signal_629, signal_233}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_218 ( .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .b ({signal_536, signal_535, signal_534, signal_533, signal_209}), .clk ( clk ), .r ({Fresh[99], Fresh[98], Fresh[97], Fresh[96], Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({signal_636, signal_635, signal_634, signal_633, signal_234}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_221 ( .a ({signal_624, signal_623, signal_622, signal_621, signal_231}), .b ({signal_648, signal_647, signal_646, signal_645, signal_237}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_224 ( .a ({signal_628, signal_627, signal_626, signal_625, signal_232}), .b ({signal_660, signal_659, signal_658, signal_657, signal_240}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_225 ( .a ({signal_632, signal_631, signal_630, signal_629, signal_233}), .b ({signal_664, signal_663, signal_662, signal_661, signal_241}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_226 ( .a ({signal_636, signal_635, signal_634, signal_633, signal_234}), .b ({signal_668, signal_667, signal_666, signal_665, signal_242}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_228 ( .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .b ({signal_600, signal_599, signal_598, signal_597, signal_225}), .clk ( clk ), .r ({Fresh[109], Fresh[108], Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100]}), .c ({signal_676, signal_675, signal_674, signal_673, signal_244}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_229 ( .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .b ({signal_604, signal_603, signal_602, signal_601, signal_226}), .clk ( clk ), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114], Fresh[113], Fresh[112], Fresh[111], Fresh[110]}), .c ({signal_680, signal_679, signal_678, signal_677, signal_245}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_230 ( .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .b ({signal_596, signal_595, signal_594, signal_593, signal_224}), .clk ( clk ), .r ({Fresh[129], Fresh[128], Fresh[127], Fresh[126], Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({signal_684, signal_683, signal_682, signal_681, signal_246}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_231 ( .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .b ({signal_608, signal_607, signal_606, signal_605, signal_227}), .clk ( clk ), .r ({Fresh[139], Fresh[138], Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132], Fresh[131], Fresh[130]}), .c ({signal_688, signal_687, signal_686, signal_685, signal_247}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_232 ( .a ({signal_676, signal_675, signal_674, signal_673, signal_244}), .b ({signal_692, signal_691, signal_690, signal_689, signal_248}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_233 ( .a ({signal_680, signal_679, signal_678, signal_677, signal_245}), .b ({signal_696, signal_695, signal_694, signal_693, signal_249}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_234 ( .a ({signal_684, signal_683, signal_682, signal_681, signal_246}), .b ({signal_700, signal_699, signal_698, signal_697, signal_250}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_235 ( .a ({signal_688, signal_687, signal_686, signal_685, signal_247}), .b ({signal_704, signal_703, signal_702, signal_701, signal_251}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_238 ( .a ({1'b0, 1'b0, 1'b0, 1'b0, signal_193}), .b ({signal_656, signal_655, signal_654, signal_653, signal_239}), .clk ( clk ), .r ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144], Fresh[143], Fresh[142], Fresh[141], Fresh[140]}), .c ({signal_716, signal_715, signal_714, signal_713, signal_254}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_239 ( .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .b ({signal_652, signal_651, signal_650, signal_649, signal_238}), .clk ( clk ), .r ({Fresh[159], Fresh[158], Fresh[157], Fresh[156], Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .c ({signal_720, signal_719, signal_718, signal_717, signal_255}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_241 ( .a ({signal_716, signal_715, signal_714, signal_713, signal_254}), .b ({signal_728, signal_727, signal_726, signal_725, signal_257}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_242 ( .a ({signal_720, signal_719, signal_718, signal_717, signal_255}), .b ({signal_732, signal_731, signal_730, signal_729, signal_258}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_227 ( .a ({signal_592, signal_591, signal_590, signal_589, signal_223}), .b ({signal_544, signal_543, signal_542, signal_541, signal_211}), .clk ( clk ), .r ({Fresh[169], Fresh[168], Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162], Fresh[161], Fresh[160]}), .c ({signal_672, signal_671, signal_670, signal_669, signal_243}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_236 ( .a ({signal_612, signal_611, signal_610, signal_609, signal_228}), .b ({signal_648, signal_647, signal_646, signal_645, signal_237}), .clk ( clk ), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174], Fresh[173], Fresh[172], Fresh[171], Fresh[170]}), .c ({signal_708, signal_707, signal_706, signal_705, signal_252}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_237 ( .a ({signal_664, signal_663, signal_662, signal_661, signal_241}), .b ({signal_668, signal_667, signal_666, signal_665, signal_242}), .clk ( clk ), .r ({Fresh[189], Fresh[188], Fresh[187], Fresh[186], Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({signal_712, signal_711, signal_710, signal_709, signal_253}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_240 ( .a ({signal_712, signal_711, signal_710, signal_709, signal_253}), .b ({signal_724, signal_723, signal_722, signal_721, signal_256}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_243 ( .a ({signal_616, signal_615, signal_614, signal_613, signal_229}), .b ({signal_692, signal_691, signal_690, signal_689, signal_248}), .clk ( clk ), .r ({Fresh[199], Fresh[198], Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192], Fresh[191], Fresh[190]}), .c ({signal_736, signal_735, signal_734, signal_733, signal_259}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_244 ( .a ({signal_660, signal_659, signal_658, signal_657, signal_240}), .b ({signal_696, signal_695, signal_694, signal_693, signal_249}), .clk ( clk ), .r ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204], Fresh[203], Fresh[202], Fresh[201], Fresh[200]}), .c ({signal_740, signal_739, signal_738, signal_737, signal_260}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_245 ( .a ({signal_548, signal_547, signal_546, signal_545, signal_212}), .b ({signal_700, signal_699, signal_698, signal_697, signal_250}), .clk ( clk ), .r ({Fresh[219], Fresh[218], Fresh[217], Fresh[216], Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .c ({signal_744, signal_743, signal_742, signal_741, signal_261}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_246 ( .a ({signal_620, signal_619, signal_618, signal_617, signal_230}), .b ({signal_704, signal_703, signal_702, signal_701, signal_251}), .clk ( clk ), .r ({Fresh[229], Fresh[228], Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222], Fresh[221], Fresh[220]}), .c ({signal_748, signal_747, signal_746, signal_745, signal_262}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_247 ( .a ({signal_728, signal_727, signal_726, signal_725, signal_257}), .b ({signal_732, signal_731, signal_730, signal_729, signal_258}), .clk ( clk ), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234], Fresh[233], Fresh[232], Fresh[231], Fresh[230]}), .c ({signal_752, signal_751, signal_750, signal_749, signal_263}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_251 ( .a ({signal_672, signal_671, signal_670, signal_669, signal_243}), .b ({signal_748, signal_747, signal_746, signal_745, signal_262}), .c ({signal_768, signal_767, signal_766, signal_765, signal_267}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_252 ( .a ({signal_708, signal_707, signal_706, signal_705, signal_252}), .b ({signal_748, signal_747, signal_746, signal_745, signal_262}), .c ({signal_772, signal_771, signal_770, signal_769, signal_268}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_253 ( .a ({signal_744, signal_743, signal_742, signal_741, signal_261}), .b ({signal_712, signal_711, signal_710, signal_709, signal_253}), .c ({signal_776, signal_775, signal_774, signal_773, signal_269}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_254 ( .a ({signal_736, signal_735, signal_734, signal_733, signal_259}), .b ({signal_740, signal_739, signal_738, signal_737, signal_260}), .c ({signal_780, signal_779, signal_778, signal_777, signal_270}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_255 ( .a ({signal_740, signal_739, signal_738, signal_737, signal_260}), .b ({signal_712, signal_711, signal_710, signal_709, signal_253}), .c ({signal_784, signal_783, signal_782, signal_781, signal_271}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_256 ( .a ({signal_736, signal_735, signal_734, signal_733, signal_259}), .b ({signal_744, signal_743, signal_742, signal_741, signal_261}), .c ({signal_788, signal_787, signal_786, signal_785, signal_272}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_257 ( .a ({signal_752, signal_751, signal_750, signal_749, signal_263}), .b ({signal_792, signal_791, signal_790, signal_789, signal_273}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_258 ( .a ({signal_772, signal_771, signal_770, signal_769, signal_268}), .b ({signal_796, signal_795, signal_794, signal_793, signal_274}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_259 ( .a ({signal_776, signal_775, signal_774, signal_773, signal_269}), .b ({signal_800, signal_799, signal_798, signal_797, signal_275}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_260 ( .a ({signal_784, signal_783, signal_782, signal_781, signal_271}), .b ({signal_804, signal_803, signal_802, signal_801, signal_276}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_261 ( .a ({signal_788, signal_787, signal_786, signal_785, signal_272}), .b ({signal_808, signal_807, signal_806, signal_805, signal_277}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_264 ( .a ({signal_708, signal_707, signal_706, signal_705, signal_252}), .b ({signal_752, signal_751, signal_750, signal_749, signal_263}), .c ({signal_820, signal_819, signal_818, signal_817, signal_280}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_265 ( .a ({signal_672, signal_671, signal_670, signal_669, signal_243}), .b ({signal_752, signal_751, signal_750, signal_749, signal_263}), .c ({signal_824, signal_823, signal_822, signal_821, signal_281}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_266 ( .a ({signal_784, signal_783, signal_782, signal_781, signal_271}), .b ({signal_788, signal_787, signal_786, signal_785, signal_272}), .c ({signal_828, signal_827, signal_826, signal_825, signal_282}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_267 ( .a ({signal_820, signal_819, signal_818, signal_817, signal_280}), .b ({signal_832, signal_831, signal_830, signal_829, signal_283}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_268 ( .a ({signal_824, signal_823, signal_822, signal_821, signal_281}), .b ({signal_836, signal_835, signal_834, signal_833, signal_284}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_273 ( .a ({signal_772, signal_771, signal_770, signal_769, signal_268}), .b ({signal_824, signal_823, signal_822, signal_821, signal_281}), .c ({signal_856, signal_855, signal_854, signal_853, signal_289}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_248 ( .a ({signal_736, signal_735, signal_734, signal_733, signal_259}), .b ({signal_748, signal_747, signal_746, signal_745, signal_262}), .clk ( clk ), .r ({Fresh[249], Fresh[248], Fresh[247], Fresh[246], Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .c ({signal_756, signal_755, signal_754, signal_753, signal_264}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_249 ( .a ({signal_672, signal_671, signal_670, signal_669, signal_243}), .b ({signal_740, signal_739, signal_738, signal_737, signal_260}), .clk ( clk ), .r ({Fresh[259], Fresh[258], Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252], Fresh[251], Fresh[250]}), .c ({signal_760, signal_759, signal_758, signal_757, signal_265}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_250 ( .a ({signal_708, signal_707, signal_706, signal_705, signal_252}), .b ({signal_744, signal_743, signal_742, signal_741, signal_261}), .clk ( clk ), .r ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264], Fresh[263], Fresh[262], Fresh[261], Fresh[260]}), .c ({signal_764, signal_763, signal_762, signal_761, signal_266}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_262 ( .a ({signal_768, signal_767, signal_766, signal_765, signal_267}), .b ({signal_780, signal_779, signal_778, signal_777, signal_270}), .clk ( clk ), .r ({Fresh[279], Fresh[278], Fresh[277], Fresh[276], Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .c ({signal_812, signal_811, signal_810, signal_809, signal_278}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_263 ( .a ({signal_772, signal_771, signal_770, signal_769, signal_268}), .b ({signal_788, signal_787, signal_786, signal_785, signal_272}), .clk ( clk ), .r ({Fresh[289], Fresh[288], Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282], Fresh[281], Fresh[280]}), .c ({signal_816, signal_815, signal_814, signal_813, signal_279}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_269 ( .a ({signal_796, signal_795, signal_794, signal_793, signal_274}), .b ({signal_808, signal_807, signal_806, signal_805, signal_277}), .clk ( clk ), .r ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294], Fresh[293], Fresh[292], Fresh[291], Fresh[290]}), .c ({signal_840, signal_839, signal_838, signal_837, signal_285}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_270 ( .a ({signal_724, signal_723, signal_722, signal_721, signal_256}), .b ({signal_792, signal_791, signal_790, signal_789, signal_273}), .clk ( clk ), .r ({Fresh[309], Fresh[308], Fresh[307], Fresh[306], Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .c ({signal_844, signal_843, signal_842, signal_841, signal_286}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_271 ( .a ({signal_776, signal_775, signal_774, signal_773, signal_269}), .b ({signal_820, signal_819, signal_818, signal_817, signal_280}), .clk ( clk ), .r ({Fresh[319], Fresh[318], Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312], Fresh[311], Fresh[310]}), .c ({signal_848, signal_847, signal_846, signal_845, signal_287}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_272 ( .a ({signal_784, signal_783, signal_782, signal_781, signal_271}), .b ({signal_824, signal_823, signal_822, signal_821, signal_281}), .clk ( clk ), .r ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324], Fresh[323], Fresh[322], Fresh[321], Fresh[320]}), .c ({signal_852, signal_851, signal_850, signal_849, signal_288}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_274 ( .a ({signal_804, signal_803, signal_802, signal_801, signal_276}), .b ({signal_836, signal_835, signal_834, signal_833, signal_284}), .clk ( clk ), .r ({Fresh[339], Fresh[338], Fresh[337], Fresh[336], Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .c ({signal_860, signal_859, signal_858, signal_857, signal_290}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_275 ( .a ({signal_800, signal_799, signal_798, signal_797, signal_275}), .b ({signal_832, signal_831, signal_830, signal_829, signal_283}), .clk ( clk ), .r ({Fresh[349], Fresh[348], Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342], Fresh[341], Fresh[340]}), .c ({signal_864, signal_863, signal_862, signal_861, signal_291}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_276 ( .a ({signal_828, signal_827, signal_826, signal_825, signal_282}), .b ({signal_856, signal_855, signal_854, signal_853, signal_289}), .clk ( clk ), .r ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354], Fresh[353], Fresh[352], Fresh[351], Fresh[350]}), .c ({signal_868, signal_867, signal_866, signal_865, signal_292}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_277 ( .a ({signal_760, signal_759, signal_758, signal_757, signal_265}), .b ({signal_840, signal_839, signal_838, signal_837, signal_285}), .c ({signal_872, signal_871, signal_870, signal_869, signal_293}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_278 ( .a ({signal_812, signal_811, signal_810, signal_809, signal_278}), .b ({signal_852, signal_851, signal_850, signal_849, signal_288}), .c ({signal_876, signal_875, signal_874, signal_873, signal_294}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_279 ( .a ({signal_844, signal_843, signal_842, signal_841, signal_286}), .b ({signal_848, signal_847, signal_846, signal_845, signal_287}), .c ({signal_880, signal_879, signal_878, signal_877, signal_295}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_280 ( .a ({signal_756, signal_755, signal_754, signal_753, signal_264}), .b ({signal_860, signal_859, signal_858, signal_857, signal_290}), .c ({signal_884, signal_883, signal_882, signal_881, signal_296}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_281 ( .a ({signal_764, signal_763, signal_762, signal_761, signal_266}), .b ({signal_864, signal_863, signal_862, signal_861, signal_291}), .c ({signal_888, signal_887, signal_886, signal_885, signal_297}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_282 ( .a ({signal_812, signal_811, signal_810, signal_809, signal_278}), .b ({signal_868, signal_867, signal_866, signal_865, signal_292}), .c ({signal_892, signal_891, signal_890, signal_889, signal_298}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_283 ( .a ({signal_872, signal_871, signal_870, signal_869, signal_293}), .b ({signal_876, signal_875, signal_874, signal_873, signal_294}), .c ({signal_896, signal_895, signal_894, signal_893, signal_299}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_284 ( .a ({signal_852, signal_851, signal_850, signal_849, signal_288}), .b ({signal_868, signal_867, signal_866, signal_865, signal_292}), .c ({signal_900, signal_899, signal_898, signal_897, signal_300}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_285 ( .a ({signal_816, signal_815, signal_814, signal_813, signal_279}), .b ({signal_880, signal_879, signal_878, signal_877, signal_295}), .c ({signal_904, signal_903, signal_902, signal_901, signal_301}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_286 ( .a ({signal_896, signal_895, signal_894, signal_893, signal_299}), .b ({signal_908, signal_907, signal_906, signal_905, signal_302}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_287 ( .a ({signal_884, signal_883, signal_882, signal_881, signal_296}), .b ({signal_892, signal_891, signal_890, signal_889, signal_298}), .c ({signal_912, signal_911, signal_910, signal_909, signal_303}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_288 ( .a ({signal_888, signal_887, signal_886, signal_885, signal_297}), .b ({signal_900, signal_899, signal_898, signal_897, signal_300}), .c ({signal_916, signal_915, signal_914, signal_913, signal_304}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_289 ( .a ({signal_852, signal_851, signal_850, signal_849, signal_288}), .b ({signal_904, signal_903, signal_902, signal_901, signal_301}), .c ({signal_920, signal_919, signal_918, signal_917, signal_305}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_290 ( .a ({signal_912, signal_911, signal_910, signal_909, signal_303}), .b ({signal_924, signal_923, signal_922, signal_921, signal_306}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_291 ( .a ({signal_916, signal_915, signal_914, signal_913, signal_304}), .b ({signal_928, signal_927, signal_926, signal_925, signal_307}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_292 ( .a ({signal_920, signal_919, signal_918, signal_917, signal_305}), .b ({signal_932, signal_931, signal_930, signal_929, signal_308}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_294 ( .a ({signal_896, signal_895, signal_894, signal_893, signal_299}), .b ({signal_912, signal_911, signal_910, signal_909, signal_303}), .c ({signal_940, signal_939, signal_938, signal_937, signal_310}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_295 ( .a ({signal_916, signal_915, signal_914, signal_913, signal_304}), .b ({signal_920, signal_919, signal_918, signal_917, signal_305}), .c ({signal_944, signal_943, signal_942, signal_941, signal_311}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_296 ( .a ({signal_940, signal_939, signal_938, signal_937, signal_310}), .b ({signal_948, signal_947, signal_946, signal_945, signal_312}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_297 ( .a ({signal_944, signal_943, signal_942, signal_941, signal_311}), .b ({signal_952, signal_951, signal_950, signal_949, signal_313}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_293 ( .a ({signal_912, signal_911, signal_910, signal_909, signal_303}), .b ({signal_916, signal_915, signal_914, signal_913, signal_304}), .clk ( clk ), .r ({Fresh[369], Fresh[368], Fresh[367], Fresh[366], Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .c ({signal_936, signal_935, signal_934, signal_933, signal_309}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_298 ( .a ({signal_908, signal_907, signal_906, signal_905, signal_302}), .b ({signal_932, signal_931, signal_930, signal_929, signal_308}), .clk ( clk ), .r ({Fresh[379], Fresh[378], Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372], Fresh[371], Fresh[370]}), .c ({signal_956, signal_955, signal_954, signal_953, signal_314}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_299 ( .a ({signal_940, signal_939, signal_938, signal_937, signal_310}), .b ({signal_944, signal_943, signal_942, signal_941, signal_311}), .clk ( clk ), .r ({Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384], Fresh[383], Fresh[382], Fresh[381], Fresh[380]}), .c ({signal_960, signal_959, signal_958, signal_957, signal_315}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_300 ( .a ({signal_948, signal_947, signal_946, signal_945, signal_312}), .b ({signal_952, signal_951, signal_950, signal_949, signal_313}), .clk ( clk ), .r ({Fresh[399], Fresh[398], Fresh[397], Fresh[396], Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390]}), .c ({signal_964, signal_963, signal_962, signal_961, signal_316}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_301 ( .a ({signal_936, signal_935, signal_934, signal_933, signal_309}), .b ({signal_960, signal_959, signal_958, signal_957, signal_315}), .c ({signal_968, signal_967, signal_966, signal_965, signal_317}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_302 ( .a ({signal_968, signal_967, signal_966, signal_965, signal_317}), .b ({signal_972, signal_971, signal_970, signal_969, signal_318}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_303 ( .a ({signal_956, signal_955, signal_954, signal_953, signal_314}), .b ({signal_964, signal_963, signal_962, signal_961, signal_316}), .c ({signal_976, signal_975, signal_974, signal_973, signal_319}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_304 ( .a ({signal_976, signal_975, signal_974, signal_973, signal_319}), .b ({signal_980, signal_979, signal_978, signal_977, signal_320}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_307 ( .a ({signal_968, signal_967, signal_966, signal_965, signal_317}), .b ({signal_976, signal_975, signal_974, signal_973, signal_319}), .c ({signal_992, signal_991, signal_990, signal_989, signal_323}) ) ;

    /* cells in depth 9 */

    /* cells in depth 10 */
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_305 ( .a ({signal_932, signal_931, signal_930, signal_929, signal_308}), .b ({signal_972, signal_971, signal_970, signal_969, signal_318}), .clk ( clk ), .r ({Fresh[409], Fresh[408], Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402], Fresh[401], Fresh[400]}), .c ({signal_984, signal_983, signal_982, signal_981, signal_321}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_306 ( .a ({signal_908, signal_907, signal_906, signal_905, signal_302}), .b ({signal_972, signal_971, signal_970, signal_969, signal_318}), .clk ( clk ), .r ({Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414], Fresh[413], Fresh[412], Fresh[411], Fresh[410]}), .c ({signal_988, signal_987, signal_986, signal_985, signal_322}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_308 ( .a ({signal_928, signal_927, signal_926, signal_925, signal_307}), .b ({signal_980, signal_979, signal_978, signal_977, signal_320}), .clk ( clk ), .r ({Fresh[429], Fresh[428], Fresh[427], Fresh[426], Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420]}), .c ({signal_996, signal_995, signal_994, signal_993, signal_324}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_309 ( .a ({signal_924, signal_923, signal_922, signal_921, signal_306}), .b ({signal_980, signal_979, signal_978, signal_977, signal_320}), .clk ( clk ), .r ({Fresh[439], Fresh[438], Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432], Fresh[431], Fresh[430]}), .c ({signal_1000, signal_999, signal_998, signal_997, signal_325}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_310 ( .a ({signal_944, signal_943, signal_942, signal_941, signal_311}), .b ({signal_992, signal_991, signal_990, signal_989, signal_323}), .clk ( clk ), .r ({Fresh[449], Fresh[448], Fresh[447], Fresh[446], Fresh[445], Fresh[444], Fresh[443], Fresh[442], Fresh[441], Fresh[440]}), .c ({signal_1004, signal_1003, signal_1002, signal_1001, signal_326}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_311 ( .a ({signal_940, signal_939, signal_938, signal_937, signal_310}), .b ({signal_992, signal_991, signal_990, signal_989, signal_323}), .clk ( clk ), .r ({Fresh[459], Fresh[458], Fresh[457], Fresh[456], Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450]}), .c ({signal_1008, signal_1007, signal_1006, signal_1005, signal_327}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_312 ( .a ({signal_996, signal_995, signal_994, signal_993, signal_324}), .b ({signal_1004, signal_1003, signal_1002, signal_1001, signal_326}), .c ({signal_1012, signal_1011, signal_1010, signal_1009, signal_328}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_313 ( .a ({signal_984, signal_983, signal_982, signal_981, signal_321}), .b ({signal_1004, signal_1003, signal_1002, signal_1001, signal_326}), .c ({signal_1016, signal_1015, signal_1014, signal_1013, signal_329}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_314 ( .a ({signal_1000, signal_999, signal_998, signal_997, signal_325}), .b ({signal_1008, signal_1007, signal_1006, signal_1005, signal_327}), .c ({signal_1020, signal_1019, signal_1018, signal_1017, signal_330}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_315 ( .a ({signal_988, signal_987, signal_986, signal_985, signal_322}), .b ({signal_1008, signal_1007, signal_1006, signal_1005, signal_327}), .c ({signal_1024, signal_1023, signal_1022, signal_1021, signal_331}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_324 ( .a ({signal_1020, signal_1019, signal_1018, signal_1017, signal_330}), .b ({signal_1024, signal_1023, signal_1022, signal_1021, signal_331}), .c ({signal_1060, signal_1059, signal_1058, signal_1057, signal_340}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_325 ( .a ({signal_1012, signal_1011, signal_1010, signal_1009, signal_328}), .b ({signal_1016, signal_1015, signal_1014, signal_1013, signal_329}), .c ({signal_1064, signal_1063, signal_1062, signal_1061, signal_341}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_326 ( .a ({signal_1016, signal_1015, signal_1014, signal_1013, signal_329}), .b ({signal_1024, signal_1023, signal_1022, signal_1021, signal_331}), .c ({signal_1068, signal_1067, signal_1066, signal_1065, signal_342}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_327 ( .a ({signal_1012, signal_1011, signal_1010, signal_1009, signal_328}), .b ({signal_1020, signal_1019, signal_1018, signal_1017, signal_330}), .c ({signal_1072, signal_1071, signal_1070, signal_1069, signal_343}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_336 ( .a ({signal_1068, signal_1067, signal_1066, signal_1065, signal_342}), .b ({signal_1072, signal_1071, signal_1070, signal_1069, signal_343}), .c ({signal_1108, signal_1107, signal_1106, signal_1105, signal_352}) ) ;

    /* cells in depth 11 */

    /* cells in depth 12 */
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_316 ( .a ({signal_748, signal_747, signal_746, signal_745, signal_262}), .b ({signal_1012, signal_1011, signal_1010, signal_1009, signal_328}), .clk ( clk ), .r ({Fresh[469], Fresh[468], Fresh[467], Fresh[466], Fresh[465], Fresh[464], Fresh[463], Fresh[462], Fresh[461], Fresh[460]}), .c ({signal_1028, signal_1027, signal_1026, signal_1025, signal_332}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_317 ( .a ({signal_672, signal_671, signal_670, signal_669, signal_243}), .b ({signal_1016, signal_1015, signal_1014, signal_1013, signal_329}), .clk ( clk ), .r ({Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474], Fresh[473], Fresh[472], Fresh[471], Fresh[470]}), .c ({signal_1032, signal_1031, signal_1030, signal_1029, signal_333}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_318 ( .a ({signal_708, signal_707, signal_706, signal_705, signal_252}), .b ({signal_1020, signal_1019, signal_1018, signal_1017, signal_330}), .clk ( clk ), .r ({Fresh[489], Fresh[488], Fresh[487], Fresh[486], Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .c ({signal_1036, signal_1035, signal_1034, signal_1033, signal_334}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_319 ( .a ({signal_752, signal_751, signal_750, signal_749, signal_263}), .b ({signal_1024, signal_1023, signal_1022, signal_1021, signal_331}), .clk ( clk ), .r ({Fresh[499], Fresh[498], Fresh[497], Fresh[496], Fresh[495], Fresh[494], Fresh[493], Fresh[492], Fresh[491], Fresh[490]}), .c ({signal_1040, signal_1039, signal_1038, signal_1037, signal_335}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_320 ( .a ({signal_736, signal_735, signal_734, signal_733, signal_259}), .b ({signal_1012, signal_1011, signal_1010, signal_1009, signal_328}), .clk ( clk ), .r ({Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504], Fresh[503], Fresh[502], Fresh[501], Fresh[500]}), .c ({signal_1044, signal_1043, signal_1042, signal_1041, signal_336}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_321 ( .a ({signal_740, signal_739, signal_738, signal_737, signal_260}), .b ({signal_1016, signal_1015, signal_1014, signal_1013, signal_329}), .clk ( clk ), .r ({Fresh[519], Fresh[518], Fresh[517], Fresh[516], Fresh[515], Fresh[514], Fresh[513], Fresh[512], Fresh[511], Fresh[510]}), .c ({signal_1048, signal_1047, signal_1046, signal_1045, signal_337}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_322 ( .a ({signal_744, signal_743, signal_742, signal_741, signal_261}), .b ({signal_1020, signal_1019, signal_1018, signal_1017, signal_330}), .clk ( clk ), .r ({Fresh[529], Fresh[528], Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522], Fresh[521], Fresh[520]}), .c ({signal_1052, signal_1051, signal_1050, signal_1049, signal_338}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_323 ( .a ({signal_712, signal_711, signal_710, signal_709, signal_253}), .b ({signal_1024, signal_1023, signal_1022, signal_1021, signal_331}), .clk ( clk ), .r ({Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534], Fresh[533], Fresh[532], Fresh[531], Fresh[530]}), .c ({signal_1056, signal_1055, signal_1054, signal_1053, signal_339}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_328 ( .a ({signal_768, signal_767, signal_766, signal_765, signal_267}), .b ({signal_1064, signal_1063, signal_1062, signal_1061, signal_341}), .clk ( clk ), .r ({Fresh[549], Fresh[548], Fresh[547], Fresh[546], Fresh[545], Fresh[544], Fresh[543], Fresh[542], Fresh[541], Fresh[540]}), .c ({signal_1076, signal_1075, signal_1074, signal_1073, signal_344}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_329 ( .a ({signal_820, signal_819, signal_818, signal_817, signal_280}), .b ({signal_1060, signal_1059, signal_1058, signal_1057, signal_340}), .clk ( clk ), .r ({Fresh[559], Fresh[558], Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552], Fresh[551], Fresh[550]}), .c ({signal_1080, signal_1079, signal_1078, signal_1077, signal_345}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_330 ( .a ({signal_772, signal_771, signal_770, signal_769, signal_268}), .b ({signal_1072, signal_1071, signal_1070, signal_1069, signal_343}), .clk ( clk ), .r ({Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564], Fresh[563], Fresh[562], Fresh[561], Fresh[560]}), .c ({signal_1084, signal_1083, signal_1082, signal_1081, signal_346}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_331 ( .a ({signal_824, signal_823, signal_822, signal_821, signal_281}), .b ({signal_1068, signal_1067, signal_1066, signal_1065, signal_342}), .clk ( clk ), .r ({Fresh[579], Fresh[578], Fresh[577], Fresh[576], Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570]}), .c ({signal_1088, signal_1087, signal_1086, signal_1085, signal_347}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_332 ( .a ({signal_780, signal_779, signal_778, signal_777, signal_270}), .b ({signal_1064, signal_1063, signal_1062, signal_1061, signal_341}), .clk ( clk ), .r ({Fresh[589], Fresh[588], Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582], Fresh[581], Fresh[580]}), .c ({signal_1092, signal_1091, signal_1090, signal_1089, signal_348}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_333 ( .a ({signal_776, signal_775, signal_774, signal_773, signal_269}), .b ({signal_1060, signal_1059, signal_1058, signal_1057, signal_340}), .clk ( clk ), .r ({Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594], Fresh[593], Fresh[592], Fresh[591], Fresh[590]}), .c ({signal_1096, signal_1095, signal_1094, signal_1093, signal_349}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_334 ( .a ({signal_788, signal_787, signal_786, signal_785, signal_272}), .b ({signal_1072, signal_1071, signal_1070, signal_1069, signal_343}), .clk ( clk ), .r ({Fresh[609], Fresh[608], Fresh[607], Fresh[606], Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600]}), .c ({signal_1100, signal_1099, signal_1098, signal_1097, signal_350}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_335 ( .a ({signal_784, signal_783, signal_782, signal_781, signal_271}), .b ({signal_1068, signal_1067, signal_1066, signal_1065, signal_342}), .clk ( clk ), .r ({Fresh[619], Fresh[618], Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612], Fresh[611], Fresh[610]}), .c ({signal_1104, signal_1103, signal_1102, signal_1101, signal_351}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_337 ( .a ({signal_856, signal_855, signal_854, signal_853, signal_289}), .b ({signal_1108, signal_1107, signal_1106, signal_1105, signal_352}), .clk ( clk ), .r ({Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624], Fresh[623], Fresh[622], Fresh[621], Fresh[620]}), .c ({signal_1112, signal_1111, signal_1110, signal_1109, signal_353}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_338 ( .a ({signal_828, signal_827, signal_826, signal_825, signal_282}), .b ({signal_1108, signal_1107, signal_1106, signal_1105, signal_352}), .clk ( clk ), .r ({Fresh[639], Fresh[638], Fresh[637], Fresh[636], Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630]}), .c ({signal_1116, signal_1115, signal_1114, signal_1113, signal_354}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_339 ( .a ({signal_1028, signal_1027, signal_1026, signal_1025, signal_332}), .b ({signal_1076, signal_1075, signal_1074, signal_1073, signal_344}), .c ({signal_1120, signal_1119, signal_1118, signal_1117, signal_355}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_340 ( .a ({signal_1032, signal_1031, signal_1030, signal_1029, signal_333}), .b ({signal_1076, signal_1075, signal_1074, signal_1073, signal_344}), .c ({signal_1124, signal_1123, signal_1122, signal_1121, signal_356}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_341 ( .a ({signal_1036, signal_1035, signal_1034, signal_1033, signal_334}), .b ({signal_1080, signal_1079, signal_1078, signal_1077, signal_345}), .c ({signal_1128, signal_1127, signal_1126, signal_1125, signal_357}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_342 ( .a ({signal_1040, signal_1039, signal_1038, signal_1037, signal_335}), .b ({signal_1080, signal_1079, signal_1078, signal_1077, signal_345}), .c ({signal_1132, signal_1131, signal_1130, signal_1129, signal_358}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_343 ( .a ({signal_1084, signal_1083, signal_1082, signal_1081, signal_346}), .b ({signal_1088, signal_1087, signal_1086, signal_1085, signal_347}), .c ({signal_1136, signal_1135, signal_1134, signal_1133, signal_359}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_344 ( .a ({signal_1044, signal_1043, signal_1042, signal_1041, signal_336}), .b ({signal_1092, signal_1091, signal_1090, signal_1089, signal_348}), .c ({signal_1140, signal_1139, signal_1138, signal_1137, signal_360}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_345 ( .a ({signal_1048, signal_1047, signal_1046, signal_1045, signal_337}), .b ({signal_1092, signal_1091, signal_1090, signal_1089, signal_348}), .c ({signal_1144, signal_1143, signal_1142, signal_1141, signal_361}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_346 ( .a ({signal_1052, signal_1051, signal_1050, signal_1049, signal_338}), .b ({signal_1096, signal_1095, signal_1094, signal_1093, signal_349}), .c ({signal_1148, signal_1147, signal_1146, signal_1145, signal_362}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_347 ( .a ({signal_1056, signal_1055, signal_1054, signal_1053, signal_339}), .b ({signal_1096, signal_1095, signal_1094, signal_1093, signal_349}), .c ({signal_1152, signal_1151, signal_1150, signal_1149, signal_363}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_348 ( .a ({signal_1100, signal_1099, signal_1098, signal_1097, signal_350}), .b ({signal_1104, signal_1103, signal_1102, signal_1101, signal_351}), .c ({signal_1156, signal_1155, signal_1154, signal_1153, signal_364}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_349 ( .a ({signal_1124, signal_1123, signal_1122, signal_1121, signal_356}), .b ({signal_1136, signal_1135, signal_1134, signal_1133, signal_359}), .c ({signal_1160, signal_1159, signal_1158, signal_1157, signal_365}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_350 ( .a ({signal_1132, signal_1131, signal_1130, signal_1129, signal_358}), .b ({signal_1136, signal_1135, signal_1134, signal_1133, signal_359}), .c ({signal_1164, signal_1163, signal_1162, signal_1161, signal_366}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_351 ( .a ({signal_1088, signal_1087, signal_1086, signal_1085, signal_347}), .b ({signal_1112, signal_1111, signal_1110, signal_1109, signal_353}), .c ({signal_1168, signal_1167, signal_1166, signal_1165, signal_367}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_352 ( .a ({signal_1144, signal_1143, signal_1142, signal_1141, signal_361}), .b ({signal_1156, signal_1155, signal_1154, signal_1153, signal_364}), .c ({signal_1172, signal_1171, signal_1170, signal_1169, signal_368}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_353 ( .a ({signal_1152, signal_1151, signal_1150, signal_1149, signal_363}), .b ({signal_1156, signal_1155, signal_1154, signal_1153, signal_364}), .c ({signal_1176, signal_1175, signal_1174, signal_1173, signal_369}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_354 ( .a ({signal_1104, signal_1103, signal_1102, signal_1101, signal_351}), .b ({signal_1116, signal_1115, signal_1114, signal_1113, signal_354}), .c ({signal_1180, signal_1179, signal_1178, signal_1177, signal_370}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_355 ( .a ({signal_1172, signal_1171, signal_1170, signal_1169, signal_368}), .b ({signal_1184, signal_1183, signal_1182, signal_1181, signal_371}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_356 ( .a ({signal_1160, signal_1159, signal_1158, signal_1157, signal_365}), .b ({signal_1176, signal_1175, signal_1174, signal_1173, signal_369}), .c ({signal_1188, signal_1187, signal_1186, signal_1185, signal_372}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_357 ( .a ({signal_1160, signal_1159, signal_1158, signal_1157, signal_365}), .b ({signal_1164, signal_1163, signal_1162, signal_1161, signal_366}), .c ({signal_1192, signal_1191, signal_1190, signal_1189, signal_373}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_358 ( .a ({signal_1120, signal_1119, signal_1118, signal_1117, signal_355}), .b ({signal_1168, signal_1167, signal_1166, signal_1165, signal_367}), .c ({signal_1196, signal_1195, signal_1194, signal_1193, signal_374}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_359 ( .a ({signal_1128, signal_1127, signal_1126, signal_1125, signal_357}), .b ({signal_1168, signal_1167, signal_1166, signal_1165, signal_367}), .c ({signal_1200, signal_1199, signal_1198, signal_1197, signal_375}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_360 ( .a ({signal_1140, signal_1139, signal_1138, signal_1137, signal_360}), .b ({signal_1180, signal_1179, signal_1178, signal_1177, signal_370}), .c ({signal_1204, signal_1203, signal_1202, signal_1201, signal_376}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_361 ( .a ({signal_1148, signal_1147, signal_1146, signal_1145, signal_362}), .b ({signal_1180, signal_1179, signal_1178, signal_1177, signal_370}), .c ({signal_1208, signal_1207, signal_1206, signal_1205, signal_377}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_364 ( .a ({signal_1200, signal_1199, signal_1198, signal_1197, signal_375}), .b ({signal_1208, signal_1207, signal_1206, signal_1205, signal_377}), .c ({signal_1220, signal_1219, signal_1218, signal_1217, signal_380}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_365 ( .a ({signal_1164, signal_1163, signal_1162, signal_1161, signal_366}), .b ({signal_1208, signal_1207, signal_1206, signal_1205, signal_377}), .c ({signal_1224, signal_1223, signal_1222, signal_1221, signal_381}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_366 ( .a ({signal_1160, signal_1159, signal_1158, signal_1157, signal_365}), .b ({signal_1208, signal_1207, signal_1206, signal_1205, signal_377}), .c ({signal_1228, signal_1227, signal_1226, signal_1225, signal_382}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_367 ( .a ({signal_1196, signal_1195, signal_1194, signal_1193, signal_374}), .b ({signal_1204, signal_1203, signal_1202, signal_1201, signal_376}), .c ({signal_1232, signal_1231, signal_1230, signal_1229, signal_383}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_368 ( .a ({signal_1200, signal_1199, signal_1198, signal_1197, signal_375}), .b ({signal_1204, signal_1203, signal_1202, signal_1201, signal_376}), .c ({signal_1236, signal_1235, signal_1234, signal_1233, signal_384}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_369 ( .a ({signal_1192, signal_1191, signal_1190, signal_1189, signal_373}), .b ({signal_1208, signal_1207, signal_1206, signal_1205, signal_377}), .c ({signal_1240, signal_1239, signal_1238, signal_1237, signal_385}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_370 ( .a ({signal_1220, signal_1219, signal_1218, signal_1217, signal_380}), .b ({signal_1244, signal_1243, signal_1242, signal_1241, signal_386}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_371 ( .a ({signal_1224, signal_1223, signal_1222, signal_1221, signal_381}), .b ({signal_1248, signal_1247, signal_1246, signal_1245, signal_387}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_372 ( .a ({signal_1228, signal_1227, signal_1226, signal_1225, signal_382}), .b ({signal_1252, signal_1251, signal_1250, signal_1249, signal_388}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_373 ( .a ({signal_1236, signal_1235, signal_1234, signal_1233, signal_384}), .b ({signal_1256, signal_1255, signal_1254, signal_1253, signal_389}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_378 ( .a ({signal_1164, signal_1163, signal_1162, signal_1161, signal_366}), .b ({signal_1220, signal_1219, signal_1218, signal_1217, signal_380}), .c ({signal_1276, signal_1275, signal_1274, signal_1273, signal_394}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_379 ( .a ({signal_1200, signal_1199, signal_1198, signal_1197, signal_375}), .b ({signal_1232, signal_1231, signal_1230, signal_1229, signal_383}), .c ({signal_1280, signal_1279, signal_1278, signal_1277, signal_395}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_380 ( .a ({signal_1172, signal_1171, signal_1170, signal_1169, signal_368}), .b ({signal_1236, signal_1235, signal_1234, signal_1233, signal_384}), .c ({signal_1284, signal_1283, signal_1282, signal_1281, signal_396}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_381 ( .a ({signal_1280, signal_1279, signal_1278, signal_1277, signal_395}), .b ({signal_1288, signal_1287, signal_1286, signal_1285, signal_397}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_389 ( .a ({signal_1196, signal_1195, signal_1194, signal_1193, signal_374}), .b ({signal_1276, signal_1275, signal_1274, signal_1273, signal_394}), .c ({signal_1320, signal_1319, signal_1318, signal_1317, signal_405}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_390 ( .a ({signal_1188, signal_1187, signal_1186, signal_1185, signal_372}), .b ({signal_1280, signal_1279, signal_1278, signal_1277, signal_395}), .c ({signal_1324, signal_1323, signal_1322, signal_1321, signal_406}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_391 ( .a ({signal_1240, signal_1239, signal_1238, signal_1237, signal_385}), .b ({signal_1284, signal_1283, signal_1282, signal_1281, signal_396}), .c ({signal_1328, signal_1327, signal_1326, signal_1325, signal_407}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_392 ( .a ({signal_1192, signal_1191, signal_1190, signal_1189, signal_373}), .b ({signal_1280, signal_1279, signal_1278, signal_1277, signal_395}), .c ({signal_1332, signal_1331, signal_1330, signal_1329, signal_408}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_393 ( .a ({signal_1188, signal_1187, signal_1186, signal_1185, signal_372}), .b ({signal_1284, signal_1283, signal_1282, signal_1281, signal_396}), .c ({signal_1336, signal_1335, signal_1334, signal_1333, signal_409}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_396 ( .a ({signal_1320, signal_1319, signal_1318, signal_1317, signal_405}), .b ({signal_1348, signal_1347, signal_1346, signal_1345, signal_412}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_397 ( .a ({signal_1328, signal_1327, signal_1326, signal_1325, signal_407}), .b ({signal_1352, signal_1351, signal_1350, signal_1349, signal_413}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_398 ( .a ({signal_1332, signal_1331, signal_1330, signal_1329, signal_408}), .b ({signal_1356, signal_1355, signal_1354, signal_1353, signal_414}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_399 ( .a ({signal_1336, signal_1335, signal_1334, signal_1333, signal_409}), .b ({signal_1360, signal_1359, signal_1358, signal_1357, signal_415}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_405 ( .a ({signal_1208, signal_1207, signal_1206, signal_1205, signal_377}), .b ({signal_1324, signal_1323, signal_1322, signal_1321, signal_406}), .c ({signal_1384, signal_1383, signal_1382, signal_1381, signal_420}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(0)) cell_406 ( .a ({signal_1172, signal_1171, signal_1170, signal_1169, signal_368}), .b ({signal_1324, signal_1323, signal_1322, signal_1321, signal_406}), .c ({signal_1388, signal_1387, signal_1386, signal_1385, signal_421}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_408 ( .a ({signal_1384, signal_1383, signal_1382, signal_1381, signal_420}), .b ({signal_1396, signal_1395, signal_1394, signal_1393, signal_423}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_409 ( .a ({signal_1388, signal_1387, signal_1386, signal_1385, signal_421}), .b ({signal_1400, signal_1399, signal_1398, signal_1397, signal_424}) ) ;

    /* cells in depth 13 */

    /* cells in depth 14 */
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_362 ( .a ({1'b0, 1'b0, 1'b0, 1'b0, signal_193}), .b ({signal_1184, signal_1183, signal_1182, signal_1181, signal_371}), .clk ( clk ), .r ({Fresh[649], Fresh[648], Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642], Fresh[641], Fresh[640]}), .c ({signal_1212, signal_1211, signal_1210, signal_1209, signal_378}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_363 ( .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .b ({signal_1188, signal_1187, signal_1186, signal_1185, signal_372}), .clk ( clk ), .r ({Fresh[659], Fresh[658], Fresh[657], Fresh[656], Fresh[655], Fresh[654], Fresh[653], Fresh[652], Fresh[651], Fresh[650]}), .c ({signal_1216, signal_1215, signal_1214, signal_1213, signal_379}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_374 ( .a ({signal_1212, signal_1211, signal_1210, signal_1209, signal_378}), .b ({signal_1260, signal_1259, signal_1258, signal_1257, signal_390}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_375 ( .a ({signal_1216, signal_1215, signal_1214, signal_1213, signal_379}), .b ({signal_1264, signal_1263, signal_1262, signal_1261, signal_391}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_376 ( .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .b ({signal_1240, signal_1239, signal_1238, signal_1237, signal_385}), .clk ( clk ), .r ({Fresh[669], Fresh[668], Fresh[667], Fresh[666], Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660]}), .c ({signal_1268, signal_1267, signal_1266, signal_1265, signal_392}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_377 ( .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .b ({signal_1232, signal_1231, signal_1230, signal_1229, signal_383}), .clk ( clk ), .r ({Fresh[679], Fresh[678], Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672], Fresh[671], Fresh[670]}), .c ({signal_1272, signal_1271, signal_1270, signal_1269, signal_393}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_382 ( .a ({signal_1268, signal_1267, signal_1266, signal_1265, signal_392}), .b ({signal_1292, signal_1291, signal_1290, signal_1289, signal_398}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_383 ( .a ({signal_1272, signal_1271, signal_1270, signal_1269, signal_393}), .b ({signal_1296, signal_1295, signal_1294, signal_1293, signal_399}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_384 ( .a ({1'b0, 1'b0, 1'b0, 1'b0, signal_193}), .b ({signal_1248, signal_1247, signal_1246, signal_1245, signal_387}), .clk ( clk ), .r ({Fresh[689], Fresh[688], Fresh[687], Fresh[686], Fresh[685], Fresh[684], Fresh[683], Fresh[682], Fresh[681], Fresh[680]}), .c ({signal_1300, signal_1299, signal_1298, signal_1297, signal_400}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_385 ( .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .b ({signal_1256, signal_1255, signal_1254, signal_1253, signal_389}), .clk ( clk ), .r ({Fresh[699], Fresh[698], Fresh[697], Fresh[696], Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690]}), .c ({signal_1304, signal_1303, signal_1302, signal_1301, signal_401}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_386 ( .a ({1'b0, 1'b0, 1'b0, 1'b0, signal_193}), .b ({signal_1252, signal_1251, signal_1250, signal_1249, signal_388}), .clk ( clk ), .r ({Fresh[709], Fresh[708], Fresh[707], Fresh[706], Fresh[705], Fresh[704], Fresh[703], Fresh[702], Fresh[701], Fresh[700]}), .c ({signal_1308, signal_1307, signal_1306, signal_1305, signal_402}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_387 ( .a ({1'b0, 1'b0, 1'b0, 1'b0, signal_193}), .b ({signal_1244, signal_1243, signal_1242, signal_1241, signal_386}), .clk ( clk ), .r ({Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714], Fresh[713], Fresh[712], Fresh[711], Fresh[710]}), .c ({signal_1312, signal_1311, signal_1310, signal_1309, signal_403}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_388 ( .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .b ({signal_1276, signal_1275, signal_1274, signal_1273, signal_394}), .clk ( clk ), .r ({Fresh[729], Fresh[728], Fresh[727], Fresh[726], Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720]}), .c ({signal_1316, signal_1315, signal_1314, signal_1313, signal_404}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_394 ( .a ({signal_1300, signal_1299, signal_1298, signal_1297, signal_400}), .b ({signal_1340, signal_1339, signal_1338, signal_1337, signal_410}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_395 ( .a ({signal_1304, signal_1303, signal_1302, signal_1301, signal_401}), .b ({signal_1344, signal_1343, signal_1342, signal_1341, signal_411}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_400 ( .a ({signal_1308, signal_1307, signal_1306, signal_1305, signal_402}), .b ({signal_1364, signal_1363, signal_1362, signal_1361, signal_416}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_401 ( .a ({signal_1312, signal_1311, signal_1310, signal_1309, signal_403}), .b ({signal_1368, signal_1367, signal_1366, signal_1365, signal_417}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_402 ( .a ({signal_1316, signal_1315, signal_1314, signal_1313, signal_404}), .b ({signal_1372, signal_1371, signal_1370, signal_1369, signal_418}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_404 ( .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .b ({signal_1288, signal_1287, signal_1286, signal_1285, signal_397}), .clk ( clk ), .r ({Fresh[739], Fresh[738], Fresh[737], Fresh[736], Fresh[735], Fresh[734], Fresh[733], Fresh[732], Fresh[731], Fresh[730]}), .c ({signal_1380, signal_1379, signal_1378, signal_1377, signal_419}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_407 ( .a ({signal_1380, signal_1379, signal_1378, signal_1377, signal_419}), .b ({signal_1392, signal_1391, signal_1390, signal_1389, signal_422}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_412 ( .a ({1'b0, 1'b0, 1'b0, 1'b0, signal_193}), .b ({signal_1352, signal_1351, signal_1350, signal_1349, signal_413}), .clk ( clk ), .r ({Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744], Fresh[743], Fresh[742], Fresh[741], Fresh[740]}), .c ({signal_1412, signal_1411, signal_1410, signal_1409, signal_425}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_413 ( .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .b ({signal_1356, signal_1355, signal_1354, signal_1353, signal_414}), .clk ( clk ), .r ({Fresh[759], Fresh[758], Fresh[757], Fresh[756], Fresh[755], Fresh[754], Fresh[753], Fresh[752], Fresh[751], Fresh[750]}), .c ({signal_1416, signal_1415, signal_1414, signal_1413, signal_426}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_414 ( .a ({1'b0, 1'b0, 1'b0, 1'b0, signal_193}), .b ({signal_1348, signal_1347, signal_1346, signal_1345, signal_412}), .clk ( clk ), .r ({Fresh[769], Fresh[768], Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762], Fresh[761], Fresh[760]}), .c ({signal_1420, signal_1419, signal_1418, signal_1417, signal_427}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_415 ( .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .b ({signal_1360, signal_1359, signal_1358, signal_1357, signal_415}), .clk ( clk ), .r ({Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774], Fresh[773], Fresh[772], Fresh[771], Fresh[770]}), .c ({signal_1424, signal_1423, signal_1422, signal_1421, signal_428}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_416 ( .a ({signal_1412, signal_1411, signal_1410, signal_1409, signal_425}), .b ({signal_1428, signal_1427, signal_1426, signal_1425, signal_429}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_417 ( .a ({signal_1416, signal_1415, signal_1414, signal_1413, signal_426}), .b ({signal_1432, signal_1431, signal_1430, signal_1429, signal_430}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_418 ( .a ({signal_1420, signal_1419, signal_1418, signal_1417, signal_427}), .b ({signal_1436, signal_1435, signal_1434, signal_1433, signal_431}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_419 ( .a ({signal_1424, signal_1423, signal_1422, signal_1421, signal_428}), .b ({signal_1440, signal_1439, signal_1438, signal_1437, signal_432}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_421 ( .a ({1'b0, 1'b0, 1'b0, 1'b0, signal_193}), .b ({signal_1396, signal_1395, signal_1394, signal_1393, signal_423}), .clk ( clk ), .r ({Fresh[789], Fresh[788], Fresh[787], Fresh[786], Fresh[785], Fresh[784], Fresh[783], Fresh[782], Fresh[781], Fresh[780]}), .c ({signal_1448, signal_1447, signal_1446, signal_1445, signal_433}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_422 ( .a ({1'b0, 1'b0, 1'b0, 1'b0, signal_193}), .b ({signal_1400, signal_1399, signal_1398, signal_1397, signal_424}), .clk ( clk ), .r ({Fresh[799], Fresh[798], Fresh[797], Fresh[796], Fresh[795], Fresh[794], Fresh[793], Fresh[792], Fresh[791], Fresh[790]}), .c ({signal_1452, signal_1451, signal_1450, signal_1449, signal_434}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_423 ( .a ({signal_1448, signal_1447, signal_1446, signal_1445, signal_433}), .b ({signal_1456, signal_1455, signal_1454, signal_1453, signal_435}) ) ;
    not_masked #(.security_order(4), .pipeline(0)) cell_424 ( .a ({signal_1452, signal_1451, signal_1450, signal_1449, signal_434}), .b ({signal_1460, signal_1459, signal_1458, signal_1457, signal_436}) ) ;

    /* cells in depth 15 */

    /* cells in depth 16 */
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_403 ( .a ({signal_1260, signal_1259, signal_1258, signal_1257, signal_390}), .b ({signal_1292, signal_1291, signal_1290, signal_1289, signal_398}), .clk ( clk ), .r ({Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804], Fresh[803], Fresh[802], Fresh[801], Fresh[800]}), .c ({signal_1376, signal_1375, signal_1374, signal_1373, signal_167}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_410 ( .a ({signal_1340, signal_1339, signal_1338, signal_1337, signal_410}), .b ({signal_1344, signal_1343, signal_1342, signal_1341, signal_411}), .clk ( clk ), .r ({Fresh[819], Fresh[818], Fresh[817], Fresh[816], Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810]}), .c ({signal_1404, signal_1403, signal_1402, signal_1401, signal_160}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_411 ( .a ({signal_1368, signal_1367, signal_1366, signal_1365, signal_417}), .b ({signal_1372, signal_1371, signal_1370, signal_1369, signal_418}), .clk ( clk ), .r ({Fresh[829], Fresh[828], Fresh[827], Fresh[826], Fresh[825], Fresh[824], Fresh[823], Fresh[822], Fresh[821], Fresh[820]}), .c ({signal_1408, signal_1407, signal_1406, signal_1405, signal_166}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_420 ( .a ({signal_1364, signal_1363, signal_1362, signal_1361, signal_416}), .b ({signal_1392, signal_1391, signal_1390, signal_1389, signal_422}), .clk ( clk ), .r ({Fresh[839], Fresh[838], Fresh[837], Fresh[836], Fresh[835], Fresh[834], Fresh[833], Fresh[832], Fresh[831], Fresh[830]}), .c ({signal_1444, signal_1443, signal_1442, signal_1441, signal_163}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_425 ( .a ({signal_1428, signal_1427, signal_1426, signal_1425, signal_429}), .b ({signal_1432, signal_1431, signal_1430, signal_1429, signal_430}), .clk ( clk ), .r ({Fresh[849], Fresh[848], Fresh[847], Fresh[846], Fresh[845], Fresh[844], Fresh[843], Fresh[842], Fresh[841], Fresh[840]}), .c ({signal_1464, signal_1463, signal_1462, signal_1461, signal_164}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_426 ( .a ({signal_1436, signal_1435, signal_1434, signal_1433, signal_431}), .b ({signal_1440, signal_1439, signal_1438, signal_1437, signal_432}), .clk ( clk ), .r ({Fresh[859], Fresh[858], Fresh[857], Fresh[856], Fresh[855], Fresh[854], Fresh[853], Fresh[852], Fresh[851], Fresh[850]}), .c ({signal_1468, signal_1467, signal_1466, signal_1465, signal_165}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_427 ( .a ({signal_1456, signal_1455, signal_1454, signal_1453, signal_435}), .b ({signal_1296, signal_1295, signal_1294, signal_1293, signal_399}), .clk ( clk ), .r ({Fresh[869], Fresh[868], Fresh[867], Fresh[866], Fresh[865], Fresh[864], Fresh[863], Fresh[862], Fresh[861], Fresh[860]}), .c ({signal_1472, signal_1471, signal_1470, signal_1469, signal_161}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(0)) cell_428 ( .a ({signal_1460, signal_1459, signal_1458, signal_1457, signal_436}), .b ({signal_1264, signal_1263, signal_1262, signal_1261, signal_391}), .clk ( clk ), .r ({Fresh[879], Fresh[878], Fresh[877], Fresh[876], Fresh[875], Fresh[874], Fresh[873], Fresh[872], Fresh[871], Fresh[870]}), .c ({signal_1476, signal_1475, signal_1474, signal_1473, signal_162}) ) ;

    /* register cells */
    reg_masked #(.security_order(4), .pipeline(0)) cell_0 ( .clk ( signal_2390 ), .D ({signal_1404, signal_1403, signal_1402, signal_1401, signal_160}), .Q ({Y_s4[7], Y_s3[7], Y_s2[7], Y_s1[7], Y_s0[7]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) cell_1 ( .clk ( signal_2390 ), .D ({signal_1472, signal_1471, signal_1470, signal_1469, signal_161}), .Q ({Y_s4[6], Y_s3[6], Y_s2[6], Y_s1[6], Y_s0[6]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) cell_2 ( .clk ( signal_2390 ), .D ({signal_1476, signal_1475, signal_1474, signal_1473, signal_162}), .Q ({Y_s4[5], Y_s3[5], Y_s2[5], Y_s1[5], Y_s0[5]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) cell_3 ( .clk ( signal_2390 ), .D ({signal_1444, signal_1443, signal_1442, signal_1441, signal_163}), .Q ({Y_s4[4], Y_s3[4], Y_s2[4], Y_s1[4], Y_s0[4]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) cell_4 ( .clk ( signal_2390 ), .D ({signal_1464, signal_1463, signal_1462, signal_1461, signal_164}), .Q ({Y_s4[3], Y_s3[3], Y_s2[3], Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) cell_5 ( .clk ( signal_2390 ), .D ({signal_1468, signal_1467, signal_1466, signal_1465, signal_165}), .Q ({Y_s4[2], Y_s3[2], Y_s2[2], Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) cell_6 ( .clk ( signal_2390 ), .D ({signal_1408, signal_1407, signal_1406, signal_1405, signal_166}), .Q ({Y_s4[1], Y_s3[1], Y_s2[1], Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) cell_7 ( .clk ( signal_2390 ), .D ({signal_1376, signal_1375, signal_1374, signal_1373, signal_167}), .Q ({Y_s4[0], Y_s3[0], Y_s2[0], Y_s1[0], Y_s0[0]}) ) ;
endmodule
