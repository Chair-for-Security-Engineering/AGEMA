module Reg1(x, y);
 input [203:0] x;
 output [202:0] y;

  assign y[10] = x[203];
  assign y[75] = x[71];
  assign y[76] = x[82];
  assign y[77] = x[93];
  assign y[78] = x[104];
  assign y[79] = x[115];
  assign y[80] = x[126];
  assign y[81] = x[131];
  assign y[82] = x[132];
  assign y[83] = x[133];
  assign y[84] = x[134];
  assign y[85] = x[72];
  assign y[86] = x[73];
  assign y[87] = x[74];
  assign y[88] = x[75];
  assign y[89] = x[76];
  assign y[90] = x[77];
  assign y[91] = x[78];
  assign y[92] = x[79];
  assign y[93] = x[80];
  assign y[94] = x[81];
  assign y[95] = x[83];
  assign y[96] = x[84];
  assign y[97] = x[85];
  assign y[98] = x[86];
  assign y[99] = x[87];
  assign y[100] = x[88];
  assign y[101] = x[89];
  assign y[102] = x[90];
  assign y[103] = x[91];
  assign y[104] = x[92];
  assign y[105] = x[94];
  assign y[106] = x[95];
  assign y[107] = x[96];
  assign y[108] = x[97];
  assign y[109] = x[98];
  assign y[110] = x[99];
  assign y[111] = x[100];
  assign y[112] = x[101];
  assign y[113] = x[102];
  assign y[114] = x[103];
  assign y[115] = x[105];
  assign y[116] = x[106];
  assign y[117] = x[107];
  assign y[118] = x[108];
  assign y[119] = x[109];
  assign y[120] = x[110];
  assign y[121] = x[111];
  assign y[122] = x[112];
  assign y[123] = x[113];
  assign y[124] = x[114];
  assign y[125] = x[116];
  assign y[126] = x[117];
  assign y[127] = x[118];
  assign y[128] = x[119];
  assign y[129] = x[120];
  assign y[130] = x[121];
  assign y[131] = x[122];
  assign y[132] = x[123];
  assign y[133] = x[124];
  assign y[134] = x[125];
  assign y[135] = x[127];
  assign y[136] = x[128];
  assign y[137] = x[129];
  assign y[138] = x[130];
  assign y[139] = x[135];
  assign y[140] = x[146];
  assign y[141] = x[157];
  assign y[142] = x[168];
  assign y[143] = x[179];
  assign y[144] = x[190];
  assign y[145] = x[195];
  assign y[146] = x[196];
  assign y[147] = x[197];
  assign y[148] = x[198];
  assign y[149] = x[136];
  assign y[150] = x[137];
  assign y[151] = x[138];
  assign y[152] = x[139];
  assign y[153] = x[140];
  assign y[154] = x[141];
  assign y[155] = x[142];
  assign y[156] = x[143];
  assign y[157] = x[144];
  assign y[158] = x[145];
  assign y[159] = x[147];
  assign y[160] = x[148];
  assign y[161] = x[149];
  assign y[162] = x[150];
  assign y[163] = x[151];
  assign y[164] = x[152];
  assign y[165] = x[153];
  assign y[166] = x[154];
  assign y[167] = x[155];
  assign y[168] = x[156];
  assign y[169] = x[158];
  assign y[170] = x[159];
  assign y[171] = x[160];
  assign y[172] = x[161];
  assign y[173] = x[162];
  assign y[174] = x[163];
  assign y[175] = x[164];
  assign y[176] = x[165];
  assign y[177] = x[166];
  assign y[178] = x[167];
  assign y[179] = x[169];
  assign y[180] = x[170];
  assign y[181] = x[171];
  assign y[182] = x[172];
  assign y[183] = x[173];
  assign y[184] = x[174];
  assign y[185] = x[175];
  assign y[186] = x[176];
  assign y[187] = x[177];
  assign y[188] = x[178];
  assign y[189] = x[180];
  assign y[190] = x[181];
  assign y[191] = x[182];
  assign y[192] = x[183];
  assign y[193] = x[184];
  assign y[194] = x[185];
  assign y[195] = x[186];
  assign y[196] = x[187];
  assign y[197] = x[188];
  assign y[198] = x[189];
  assign y[199] = x[191];
  assign y[200] = x[192];
  assign y[201] = x[193];
  assign y[202] = x[194];
  register_stage #(.WIDTH(74)) inst_0(.clk(x[199]), .D({x[200],x[64],x[65],x[66],x[67],x[68],x[69],x[70],x[201],x[202],x[0],x[11],x[22],x[33],x[44],x[55],x[60],x[61],x[62],x[63],x[1],x[2],x[3],x[4],x[5],x[6],x[7],x[8],x[9],x[10],x[12],x[13],x[14],x[15],x[16],x[17],x[18],x[19],x[20],x[21],x[23],x[24],x[25],x[26],x[27],x[28],x[29],x[30],x[31],x[32],x[34],x[35],x[36],x[37],x[38],x[39],x[40],x[41],x[42],x[43],x[45],x[46],x[47],x[48],x[49],x[50],x[51],x[52],x[53],x[54],x[56],x[57],x[58],x[59]}), .Q({y[0],y[1],y[2],y[3],y[4],y[5],y[6],y[7],y[8],y[9],y[11],y[12],y[13],y[14],y[15],y[16],y[17],y[18],y[19],y[20],y[21],y[22],y[23],y[24],y[25],y[26],y[27],y[28],y[29],y[30],y[31],y[32],y[33],y[34],y[35],y[36],y[37],y[38],y[39],y[40],y[41],y[42],y[43],y[44],y[45],y[46],y[47],y[48],y[49],y[50],y[51],y[52],y[53],y[54],y[55],y[56],y[57],y[58],y[59],y[60],y[61],y[62],y[63],y[64],y[65],y[66],y[67],y[68],y[69],y[70],y[71],y[72],y[73],y[74]}));
endmodule

module Reg2(x, y);
 input [406:0] x;
 output [405:0] y;

  assign y[20] = x[405];
  assign y[21] = x[406];
  assign y[150] = x[142];
  assign y[151] = x[143];
  assign y[152] = x[164];
  assign y[153] = x[165];
  assign y[154] = x[186];
  assign y[155] = x[187];
  assign y[156] = x[208];
  assign y[157] = x[209];
  assign y[158] = x[230];
  assign y[159] = x[231];
  assign y[160] = x[252];
  assign y[161] = x[253];
  assign y[162] = x[262];
  assign y[163] = x[263];
  assign y[164] = x[264];
  assign y[165] = x[265];
  assign y[166] = x[266];
  assign y[167] = x[267];
  assign y[168] = x[268];
  assign y[169] = x[269];
  assign y[170] = x[144];
  assign y[171] = x[145];
  assign y[172] = x[146];
  assign y[173] = x[147];
  assign y[174] = x[148];
  assign y[175] = x[149];
  assign y[176] = x[150];
  assign y[177] = x[151];
  assign y[178] = x[152];
  assign y[179] = x[153];
  assign y[180] = x[154];
  assign y[181] = x[155];
  assign y[182] = x[156];
  assign y[183] = x[157];
  assign y[184] = x[158];
  assign y[185] = x[159];
  assign y[186] = x[160];
  assign y[187] = x[161];
  assign y[188] = x[162];
  assign y[189] = x[163];
  assign y[190] = x[166];
  assign y[191] = x[167];
  assign y[192] = x[168];
  assign y[193] = x[169];
  assign y[194] = x[170];
  assign y[195] = x[171];
  assign y[196] = x[172];
  assign y[197] = x[173];
  assign y[198] = x[174];
  assign y[199] = x[175];
  assign y[200] = x[176];
  assign y[201] = x[177];
  assign y[202] = x[178];
  assign y[203] = x[179];
  assign y[204] = x[180];
  assign y[205] = x[181];
  assign y[206] = x[182];
  assign y[207] = x[183];
  assign y[208] = x[184];
  assign y[209] = x[185];
  assign y[210] = x[188];
  assign y[211] = x[189];
  assign y[212] = x[190];
  assign y[213] = x[191];
  assign y[214] = x[192];
  assign y[215] = x[193];
  assign y[216] = x[194];
  assign y[217] = x[195];
  assign y[218] = x[196];
  assign y[219] = x[197];
  assign y[220] = x[198];
  assign y[221] = x[199];
  assign y[222] = x[200];
  assign y[223] = x[201];
  assign y[224] = x[202];
  assign y[225] = x[203];
  assign y[226] = x[204];
  assign y[227] = x[205];
  assign y[228] = x[206];
  assign y[229] = x[207];
  assign y[230] = x[210];
  assign y[231] = x[211];
  assign y[232] = x[212];
  assign y[233] = x[213];
  assign y[234] = x[214];
  assign y[235] = x[215];
  assign y[236] = x[216];
  assign y[237] = x[217];
  assign y[238] = x[218];
  assign y[239] = x[219];
  assign y[240] = x[220];
  assign y[241] = x[221];
  assign y[242] = x[222];
  assign y[243] = x[223];
  assign y[244] = x[224];
  assign y[245] = x[225];
  assign y[246] = x[226];
  assign y[247] = x[227];
  assign y[248] = x[228];
  assign y[249] = x[229];
  assign y[250] = x[232];
  assign y[251] = x[233];
  assign y[252] = x[234];
  assign y[253] = x[235];
  assign y[254] = x[236];
  assign y[255] = x[237];
  assign y[256] = x[238];
  assign y[257] = x[239];
  assign y[258] = x[240];
  assign y[259] = x[241];
  assign y[260] = x[242];
  assign y[261] = x[243];
  assign y[262] = x[244];
  assign y[263] = x[245];
  assign y[264] = x[246];
  assign y[265] = x[247];
  assign y[266] = x[248];
  assign y[267] = x[249];
  assign y[268] = x[250];
  assign y[269] = x[251];
  assign y[270] = x[254];
  assign y[271] = x[255];
  assign y[272] = x[256];
  assign y[273] = x[257];
  assign y[274] = x[258];
  assign y[275] = x[259];
  assign y[276] = x[260];
  assign y[277] = x[261];
  assign y[278] = x[270];
  assign y[279] = x[271];
  assign y[280] = x[292];
  assign y[281] = x[293];
  assign y[282] = x[314];
  assign y[283] = x[315];
  assign y[284] = x[336];
  assign y[285] = x[337];
  assign y[286] = x[358];
  assign y[287] = x[359];
  assign y[288] = x[380];
  assign y[289] = x[381];
  assign y[290] = x[390];
  assign y[291] = x[391];
  assign y[292] = x[392];
  assign y[293] = x[393];
  assign y[294] = x[394];
  assign y[295] = x[395];
  assign y[296] = x[396];
  assign y[297] = x[397];
  assign y[298] = x[272];
  assign y[299] = x[273];
  assign y[300] = x[274];
  assign y[301] = x[275];
  assign y[302] = x[276];
  assign y[303] = x[277];
  assign y[304] = x[278];
  assign y[305] = x[279];
  assign y[306] = x[280];
  assign y[307] = x[281];
  assign y[308] = x[282];
  assign y[309] = x[283];
  assign y[310] = x[284];
  assign y[311] = x[285];
  assign y[312] = x[286];
  assign y[313] = x[287];
  assign y[314] = x[288];
  assign y[315] = x[289];
  assign y[316] = x[290];
  assign y[317] = x[291];
  assign y[318] = x[294];
  assign y[319] = x[295];
  assign y[320] = x[296];
  assign y[321] = x[297];
  assign y[322] = x[298];
  assign y[323] = x[299];
  assign y[324] = x[300];
  assign y[325] = x[301];
  assign y[326] = x[302];
  assign y[327] = x[303];
  assign y[328] = x[304];
  assign y[329] = x[305];
  assign y[330] = x[306];
  assign y[331] = x[307];
  assign y[332] = x[308];
  assign y[333] = x[309];
  assign y[334] = x[310];
  assign y[335] = x[311];
  assign y[336] = x[312];
  assign y[337] = x[313];
  assign y[338] = x[316];
  assign y[339] = x[317];
  assign y[340] = x[318];
  assign y[341] = x[319];
  assign y[342] = x[320];
  assign y[343] = x[321];
  assign y[344] = x[322];
  assign y[345] = x[323];
  assign y[346] = x[324];
  assign y[347] = x[325];
  assign y[348] = x[326];
  assign y[349] = x[327];
  assign y[350] = x[328];
  assign y[351] = x[329];
  assign y[352] = x[330];
  assign y[353] = x[331];
  assign y[354] = x[332];
  assign y[355] = x[333];
  assign y[356] = x[334];
  assign y[357] = x[335];
  assign y[358] = x[338];
  assign y[359] = x[339];
  assign y[360] = x[340];
  assign y[361] = x[341];
  assign y[362] = x[342];
  assign y[363] = x[343];
  assign y[364] = x[344];
  assign y[365] = x[345];
  assign y[366] = x[346];
  assign y[367] = x[347];
  assign y[368] = x[348];
  assign y[369] = x[349];
  assign y[370] = x[350];
  assign y[371] = x[351];
  assign y[372] = x[352];
  assign y[373] = x[353];
  assign y[374] = x[354];
  assign y[375] = x[355];
  assign y[376] = x[356];
  assign y[377] = x[357];
  assign y[378] = x[360];
  assign y[379] = x[361];
  assign y[380] = x[362];
  assign y[381] = x[363];
  assign y[382] = x[364];
  assign y[383] = x[365];
  assign y[384] = x[366];
  assign y[385] = x[367];
  assign y[386] = x[368];
  assign y[387] = x[369];
  assign y[388] = x[370];
  assign y[389] = x[371];
  assign y[390] = x[372];
  assign y[391] = x[373];
  assign y[392] = x[374];
  assign y[393] = x[375];
  assign y[394] = x[376];
  assign y[395] = x[377];
  assign y[396] = x[378];
  assign y[397] = x[379];
  assign y[398] = x[382];
  assign y[399] = x[383];
  assign y[400] = x[384];
  assign y[401] = x[385];
  assign y[402] = x[386];
  assign y[403] = x[387];
  assign y[404] = x[388];
  assign y[405] = x[389];
  register_stage #(.WIDTH(148)) inst_0(.clk(x[398]), .D({x[399],x[400],x[128],x[129],x[130],x[131],x[132],x[133],x[134],x[135],x[136],x[137],x[138],x[139],x[140],x[141],x[401],x[402],x[403],x[404],x[0],x[1],x[22],x[23],x[44],x[45],x[66],x[67],x[88],x[89],x[110],x[111],x[120],x[121],x[122],x[123],x[124],x[125],x[126],x[127],x[2],x[3],x[4],x[5],x[6],x[7],x[8],x[9],x[10],x[11],x[12],x[13],x[14],x[15],x[16],x[17],x[18],x[19],x[20],x[21],x[24],x[25],x[26],x[27],x[28],x[29],x[30],x[31],x[32],x[33],x[34],x[35],x[36],x[37],x[38],x[39],x[40],x[41],x[42],x[43],x[46],x[47],x[48],x[49],x[50],x[51],x[52],x[53],x[54],x[55],x[56],x[57],x[58],x[59],x[60],x[61],x[62],x[63],x[64],x[65],x[68],x[69],x[70],x[71],x[72],x[73],x[74],x[75],x[76],x[77],x[78],x[79],x[80],x[81],x[82],x[83],x[84],x[85],x[86],x[87],x[90],x[91],x[92],x[93],x[94],x[95],x[96],x[97],x[98],x[99],x[100],x[101],x[102],x[103],x[104],x[105],x[106],x[107],x[108],x[109],x[112],x[113],x[114],x[115],x[116],x[117],x[118],x[119]}), .Q({y[0],y[1],y[2],y[3],y[4],y[5],y[6],y[7],y[8],y[9],y[10],y[11],y[12],y[13],y[14],y[15],y[16],y[17],y[18],y[19],y[22],y[23],y[24],y[25],y[26],y[27],y[28],y[29],y[30],y[31],y[32],y[33],y[34],y[35],y[36],y[37],y[38],y[39],y[40],y[41],y[42],y[43],y[44],y[45],y[46],y[47],y[48],y[49],y[50],y[51],y[52],y[53],y[54],y[55],y[56],y[57],y[58],y[59],y[60],y[61],y[62],y[63],y[64],y[65],y[66],y[67],y[68],y[69],y[70],y[71],y[72],y[73],y[74],y[75],y[76],y[77],y[78],y[79],y[80],y[81],y[82],y[83],y[84],y[85],y[86],y[87],y[88],y[89],y[90],y[91],y[92],y[93],y[94],y[95],y[96],y[97],y[98],y[99],y[100],y[101],y[102],y[103],y[104],y[105],y[106],y[107],y[108],y[109],y[110],y[111],y[112],y[113],y[114],y[115],y[116],y[117],y[118],y[119],y[120],y[121],y[122],y[123],y[124],y[125],y[126],y[127],y[128],y[129],y[130],y[131],y[132],y[133],y[134],y[135],y[136],y[137],y[138],y[139],y[140],y[141],y[142],y[143],y[144],y[145],y[146],y[147],y[148],y[149]}));
endmodule

module InF(x, y);
 input [192:0] x;
 output [385:0] y;

  assign y[0] = (x[0]);
  assign y[1] = (x[0]);
  assign y[2] = (x[1]);
  assign y[3] = (x[1]);
  assign y[4] = (x[2]);
  assign y[5] = (x[2]);
  assign y[6] = (x[3]);
  assign y[7] = (x[3]);
  assign y[8] = (x[4]);
  assign y[9] = (x[4]);
  assign y[10] = (x[5]);
  assign y[11] = (x[5]);
  assign y[12] = (x[6]);
  assign y[13] = (x[6]);
  assign y[14] = (x[7]);
  assign y[15] = (x[7]);
  assign y[16] = (x[8]);
  assign y[17] = (x[8]);
  assign y[18] = (x[9]);
  assign y[19] = (x[9]);
  assign y[20] = (x[10]);
  assign y[21] = (x[10]);
  assign y[22] = (x[11]);
  assign y[23] = (x[11]);
  assign y[24] = (x[12]);
  assign y[25] = (x[12]);
  assign y[26] = (x[13]);
  assign y[27] = (x[13]);
  assign y[28] = (x[14]);
  assign y[29] = (x[14]);
  assign y[30] = (x[15]);
  assign y[31] = (x[15]);
  assign y[32] = (x[16]);
  assign y[33] = (x[16]);
  assign y[34] = (x[17]);
  assign y[35] = (x[17]);
  assign y[36] = (x[18]);
  assign y[37] = (x[18]);
  assign y[38] = (x[19]);
  assign y[39] = (x[19]);
  assign y[40] = (x[20]);
  assign y[41] = (x[20]);
  assign y[42] = (x[21]);
  assign y[43] = (x[21]);
  assign y[44] = (x[22]);
  assign y[45] = (x[22]);
  assign y[46] = (x[23]);
  assign y[47] = (x[23]);
  assign y[48] = (x[24]);
  assign y[49] = (x[24]);
  assign y[50] = (x[25]);
  assign y[51] = (x[25]);
  assign y[52] = (x[26]);
  assign y[53] = (x[26]);
  assign y[54] = (x[27]);
  assign y[55] = (x[27]);
  assign y[56] = (x[28]);
  assign y[57] = (x[28]);
  assign y[58] = (x[29]);
  assign y[59] = (x[29]);
  assign y[60] = (x[30]);
  assign y[61] = (x[30]);
  assign y[62] = (x[31]);
  assign y[63] = (x[31]);
  assign y[64] = (x[32]);
  assign y[65] = (x[32]);
  assign y[66] = (x[33]);
  assign y[67] = (x[33]);
  assign y[68] = (x[34]);
  assign y[69] = (x[34]);
  assign y[70] = (x[35]);
  assign y[71] = (x[35]);
  assign y[72] = (x[36]);
  assign y[73] = (x[36]);
  assign y[74] = (x[37]);
  assign y[75] = (x[37]);
  assign y[76] = (x[38]);
  assign y[77] = (x[38]);
  assign y[78] = (x[39]);
  assign y[79] = (x[39]);
  assign y[80] = (x[40]);
  assign y[81] = (x[40]);
  assign y[82] = (x[41]);
  assign y[83] = (x[41]);
  assign y[84] = (x[42]);
  assign y[85] = (x[42]);
  assign y[86] = (x[43]);
  assign y[87] = (x[43]);
  assign y[88] = (x[44]);
  assign y[89] = (x[44]);
  assign y[90] = (x[45]);
  assign y[91] = (x[45]);
  assign y[92] = (x[46]);
  assign y[93] = (x[46]);
  assign y[94] = (x[47]);
  assign y[95] = (x[47]);
  assign y[96] = (x[48]);
  assign y[97] = (x[48]);
  assign y[98] = (x[49]);
  assign y[99] = (x[49]);
  assign y[100] = (x[50]);
  assign y[101] = (x[50]);
  assign y[102] = (x[51]);
  assign y[103] = (x[51]);
  assign y[104] = (x[52]);
  assign y[105] = (x[52]);
  assign y[106] = (x[53]);
  assign y[107] = (x[53]);
  assign y[108] = (x[54]);
  assign y[109] = (x[54]);
  assign y[110] = (x[55]);
  assign y[111] = (x[55]);
  assign y[112] = (x[56]);
  assign y[113] = (x[56]);
  assign y[114] = (x[57]);
  assign y[115] = (x[57]);
  assign y[116] = (x[58]);
  assign y[117] = (x[58]);
  assign y[118] = (x[59]);
  assign y[119] = (x[59]);
  assign y[120] = (x[60]);
  assign y[121] = (x[60]);
  assign y[122] = (x[61]);
  assign y[123] = (x[61]);
  assign y[124] = (x[62]);
  assign y[125] = (x[62]);
  assign y[126] = (x[63]);
  assign y[127] = (x[63]);
  assign y[128] = (x[64]);
  assign y[129] = (x[64]);
  assign y[130] = (x[65]);
  assign y[131] = (x[65]);
  assign y[132] = (x[66]);
  assign y[133] = (x[66]);
  assign y[134] = (x[67]);
  assign y[135] = (x[67]);
  assign y[136] = (x[68]);
  assign y[137] = (x[68]);
  assign y[138] = (x[69]);
  assign y[139] = (x[69]);
  assign y[140] = (x[70]);
  assign y[141] = (x[70]);
  assign y[142] = (x[71]);
  assign y[143] = (x[71]);
  assign y[144] = (x[72]);
  assign y[145] = (x[72]);
  assign y[146] = (x[73]);
  assign y[147] = (x[73]);
  assign y[148] = (x[74]);
  assign y[149] = (x[74]);
  assign y[150] = (x[75]);
  assign y[151] = (x[75]);
  assign y[152] = (x[76]);
  assign y[153] = (x[76]);
  assign y[154] = (x[77]);
  assign y[155] = (x[77]);
  assign y[156] = (x[78]);
  assign y[157] = (x[78]);
  assign y[158] = (x[79]);
  assign y[159] = (x[79]);
  assign y[160] = (x[80]);
  assign y[161] = (x[80]);
  assign y[162] = (x[81]);
  assign y[163] = (x[81]);
  assign y[164] = (x[82]);
  assign y[165] = (x[82]);
  assign y[166] = (x[83]);
  assign y[167] = (x[83]);
  assign y[168] = (x[84]);
  assign y[169] = (x[84]);
  assign y[170] = (x[85]);
  assign y[171] = (x[85]);
  assign y[172] = (x[86]);
  assign y[173] = (x[86]);
  assign y[174] = (x[87]);
  assign y[175] = (x[87]);
  assign y[176] = (x[88]);
  assign y[177] = (x[88]);
  assign y[178] = (x[89]);
  assign y[179] = (x[89]);
  assign y[180] = (x[90]);
  assign y[181] = (x[90]);
  assign y[182] = (x[91]);
  assign y[183] = (x[91]);
  assign y[184] = (x[92]);
  assign y[185] = (x[92]);
  assign y[186] = (x[93]);
  assign y[187] = (x[93]);
  assign y[188] = (x[94]);
  assign y[189] = (x[94]);
  assign y[190] = (x[95]);
  assign y[191] = (x[95]);
  assign y[192] = (x[96]);
  assign y[193] = (x[96]);
  assign y[194] = (x[97]);
  assign y[195] = (x[97]);
  assign y[196] = (x[98]);
  assign y[197] = (x[98]);
  assign y[198] = (x[99]);
  assign y[199] = (x[99]);
  assign y[200] = (x[100]);
  assign y[201] = (x[100]);
  assign y[202] = (x[101]);
  assign y[203] = (x[101]);
  assign y[204] = (x[102]);
  assign y[205] = (x[102]);
  assign y[206] = (x[103]);
  assign y[207] = (x[103]);
  assign y[208] = (x[104]);
  assign y[209] = (x[104]);
  assign y[210] = (x[105]);
  assign y[211] = (x[105]);
  assign y[212] = (x[106]);
  assign y[213] = (x[106]);
  assign y[214] = (x[107]);
  assign y[215] = (x[107]);
  assign y[216] = (x[108]);
  assign y[217] = (x[108]);
  assign y[218] = (x[109]);
  assign y[219] = (x[109]);
  assign y[220] = (x[110]);
  assign y[221] = (x[110]);
  assign y[222] = (x[111]);
  assign y[223] = (x[111]);
  assign y[224] = (x[112]);
  assign y[225] = (x[112]);
  assign y[226] = (x[113]);
  assign y[227] = (x[113]);
  assign y[228] = (x[114]);
  assign y[229] = (x[114]);
  assign y[230] = (x[115]);
  assign y[231] = (x[115]);
  assign y[232] = (x[116]);
  assign y[233] = (x[116]);
  assign y[234] = (x[117]);
  assign y[235] = (x[117]);
  assign y[236] = (x[118]);
  assign y[237] = (x[118]);
  assign y[238] = (x[119]);
  assign y[239] = (x[119]);
  assign y[240] = (x[120]);
  assign y[241] = (x[120]);
  assign y[242] = (x[121]);
  assign y[243] = (x[121]);
  assign y[244] = (x[122]);
  assign y[245] = (x[122]);
  assign y[246] = (x[123]);
  assign y[247] = (x[123]);
  assign y[248] = (x[124]);
  assign y[249] = (x[124]);
  assign y[250] = (x[125]);
  assign y[251] = (x[125]);
  assign y[252] = (x[126]);
  assign y[253] = (x[126]);
  assign y[254] = (x[127]);
  assign y[255] = (x[127]);
  assign y[256] = (x[128]);
  assign y[257] = (x[128]);
  assign y[258] = (x[129]);
  assign y[259] = (x[129]);
  assign y[260] = (x[130]);
  assign y[261] = (x[130]);
  assign y[262] = (x[131]);
  assign y[263] = (x[131]);
  assign y[264] = (x[132]);
  assign y[265] = (x[132]);
  assign y[266] = (x[133]);
  assign y[267] = (x[133]);
  assign y[268] = (x[134]);
  assign y[269] = (x[134]);
  assign y[270] = (x[135]);
  assign y[271] = (x[135]);
  assign y[272] = (x[136]);
  assign y[273] = (x[136]);
  assign y[274] = (x[137]);
  assign y[275] = (x[137]);
  assign y[276] = (x[138]);
  assign y[277] = (x[138]);
  assign y[278] = (x[139]);
  assign y[279] = (x[139]);
  assign y[280] = (x[140]);
  assign y[281] = (x[140]);
  assign y[282] = (x[141]);
  assign y[283] = (x[141]);
  assign y[284] = (x[142]);
  assign y[285] = (x[142]);
  assign y[286] = (x[143]);
  assign y[287] = (x[143]);
  assign y[288] = (x[144]);
  assign y[289] = (x[144]);
  assign y[290] = (x[145]);
  assign y[291] = (x[145]);
  assign y[292] = (x[146]);
  assign y[293] = (x[146]);
  assign y[294] = (x[147]);
  assign y[295] = (x[147]);
  assign y[296] = (x[148]);
  assign y[297] = (x[148]);
  assign y[298] = (x[149]);
  assign y[299] = (x[149]);
  assign y[300] = (x[150]);
  assign y[301] = (x[150]);
  assign y[302] = (x[151]);
  assign y[303] = (x[151]);
  assign y[304] = (x[152]);
  assign y[305] = (x[152]);
  assign y[306] = (x[153]);
  assign y[307] = (x[153]);
  assign y[308] = (x[154]);
  assign y[309] = (x[154]);
  assign y[310] = (x[155]);
  assign y[311] = (x[155]);
  assign y[312] = (x[156]);
  assign y[313] = (x[156]);
  assign y[314] = (x[157]);
  assign y[315] = (x[157]);
  assign y[316] = (x[158]);
  assign y[317] = (x[158]);
  assign y[318] = (x[159]);
  assign y[319] = (x[159]);
  assign y[320] = (x[160]);
  assign y[321] = (x[160]);
  assign y[322] = (x[161]);
  assign y[323] = (x[161]);
  assign y[324] = (x[162]);
  assign y[325] = (x[162]);
  assign y[326] = (x[163]);
  assign y[327] = (x[163]);
  assign y[328] = (x[164]);
  assign y[329] = (x[164]);
  assign y[330] = (x[165]);
  assign y[331] = (x[165]);
  assign y[332] = (x[166]);
  assign y[333] = (x[166]);
  assign y[334] = (x[167]);
  assign y[335] = (x[167]);
  assign y[336] = (x[168]);
  assign y[337] = (x[168]);
  assign y[338] = (x[169]);
  assign y[339] = (x[169]);
  assign y[340] = (x[170]);
  assign y[341] = (x[170]);
  assign y[342] = (x[171]);
  assign y[343] = (x[171]);
  assign y[344] = (x[172]);
  assign y[345] = (x[172]);
  assign y[346] = (x[173]);
  assign y[347] = (x[173]);
  assign y[348] = (x[174]);
  assign y[349] = (x[174]);
  assign y[350] = (x[175]);
  assign y[351] = (x[175]);
  assign y[352] = (x[176]);
  assign y[353] = (x[176]);
  assign y[354] = (x[177]);
  assign y[355] = (x[177]);
  assign y[356] = (x[178]);
  assign y[357] = (x[178]);
  assign y[358] = (x[179]);
  assign y[359] = (x[179]);
  assign y[360] = (x[180]);
  assign y[361] = (x[180]);
  assign y[362] = (x[181]);
  assign y[363] = (x[181]);
  assign y[364] = (x[182]);
  assign y[365] = (x[182]);
  assign y[366] = (x[183]);
  assign y[367] = (x[183]);
  assign y[368] = (x[184]);
  assign y[369] = (x[184]);
  assign y[370] = (x[185]);
  assign y[371] = (x[185]);
  assign y[372] = (x[186]);
  assign y[373] = (x[186]);
  assign y[374] = (x[187]);
  assign y[375] = (x[187]);
  assign y[376] = (x[188]);
  assign y[377] = (x[188]);
  assign y[378] = (x[189]);
  assign y[379] = (x[189]);
  assign y[380] = (x[190]);
  assign y[381] = (x[190]);
  assign y[382] = (x[191]);
  assign y[383] = (x[191]);
  assign y[384] = (x[192]);
  assign y[385] = (x[192]);
endmodule

module Fx0(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx1(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx2(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx3(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx4(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx5(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx6(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx7(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx8(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx9(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx10(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx11(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx12(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx13(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx14(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx15(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx16(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx17(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx18(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx19(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx20(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx21(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx22(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx23(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx24(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx25(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx26(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx27(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx28(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx29(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx30(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx31(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx32(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx33(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx34(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx35(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx36(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx37(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx38(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx39(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx40(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx41(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx42(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx43(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx44(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx45(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx46(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx47(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx48(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx49(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx50(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx51(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx52(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx53(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx54(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx55(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx56(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx57(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx58(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx59(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx60(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx61(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx62(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx63(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx64(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx65(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx66(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx67(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx68(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx69(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx70(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx71(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx72(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx73(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx74(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx75(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx76(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx77(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx78(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx79(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx80(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx81(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx82(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx83(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx84(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx85(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx86(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx87(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx88(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx89(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx90(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx91(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx92(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx93(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx94(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx95(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx96(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx97(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx98(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx99(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx100(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx101(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx102(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx103(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx104(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx105(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx106(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx107(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx108(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx109(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx110(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx111(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx112(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx113(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx114(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx115(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx116(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx117(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx118(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx119(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx120(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx121(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx122(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx123(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx124(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx125(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx126(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx127(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx128(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx129(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx130(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx131(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx132(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx133(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx134(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx135(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx136(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx137(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx138(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx139(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx140(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx141(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx142(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx143(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx144(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx145(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx146(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx147(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx148(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx149(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module FX(x, y);
 input [224:0] x;
 output [149:0] y;

  Fx0 Fx0_inst(.x({x[1], x[0]}), .y(y[0]));
  Fx1 Fx1_inst(.x({x[2], x[0]}), .y(y[1]));
  Fx2 Fx2_inst(.x({x[4], x[3]}), .y(y[2]));
  Fx3 Fx3_inst(.x({x[5], x[3]}), .y(y[3]));
  Fx4 Fx4_inst(.x({x[7], x[6]}), .y(y[4]));
  Fx5 Fx5_inst(.x({x[8], x[6]}), .y(y[5]));
  Fx6 Fx6_inst(.x({x[10], x[9]}), .y(y[6]));
  Fx7 Fx7_inst(.x({x[11], x[9]}), .y(y[7]));
  Fx8 Fx8_inst(.x({x[13], x[12]}), .y(y[8]));
  Fx9 Fx9_inst(.x({x[14], x[12]}), .y(y[9]));
  Fx10 Fx10_inst(.x({x[16], x[15]}), .y(y[10]));
  Fx11 Fx11_inst(.x({x[17], x[15]}), .y(y[11]));
  Fx12 Fx12_inst(.x({x[19], x[18]}), .y(y[12]));
  Fx13 Fx13_inst(.x({x[20], x[18]}), .y(y[13]));
  Fx14 Fx14_inst(.x({x[22], x[21]}), .y(y[14]));
  Fx15 Fx15_inst(.x({x[23], x[21]}), .y(y[15]));
  Fx16 Fx16_inst(.x({x[25], x[24]}), .y(y[16]));
  Fx17 Fx17_inst(.x({x[26], x[24]}), .y(y[17]));
  Fx18 Fx18_inst(.x({x[28], x[27]}), .y(y[18]));
  Fx19 Fx19_inst(.x({x[29], x[27]}), .y(y[19]));
  Fx20 Fx20_inst(.x({x[31], x[30]}), .y(y[20]));
  Fx21 Fx21_inst(.x({x[32], x[30]}), .y(y[21]));
  Fx22 Fx22_inst(.x({x[34], x[33]}), .y(y[22]));
  Fx23 Fx23_inst(.x({x[35], x[33]}), .y(y[23]));
  Fx24 Fx24_inst(.x({x[37], x[36]}), .y(y[24]));
  Fx25 Fx25_inst(.x({x[38], x[36]}), .y(y[25]));
  Fx26 Fx26_inst(.x({x[40], x[39]}), .y(y[26]));
  Fx27 Fx27_inst(.x({x[41], x[39]}), .y(y[27]));
  Fx28 Fx28_inst(.x({x[43], x[42]}), .y(y[28]));
  Fx29 Fx29_inst(.x({x[44], x[42]}), .y(y[29]));
  Fx30 Fx30_inst(.x({x[46], x[45]}), .y(y[30]));
  Fx31 Fx31_inst(.x({x[47], x[45]}), .y(y[31]));
  Fx32 Fx32_inst(.x({x[49], x[48]}), .y(y[32]));
  Fx33 Fx33_inst(.x({x[50], x[48]}), .y(y[33]));
  Fx34 Fx34_inst(.x({x[52], x[51]}), .y(y[34]));
  Fx35 Fx35_inst(.x({x[53], x[51]}), .y(y[35]));
  Fx36 Fx36_inst(.x({x[55], x[54]}), .y(y[36]));
  Fx37 Fx37_inst(.x({x[56], x[54]}), .y(y[37]));
  Fx38 Fx38_inst(.x({x[58], x[57]}), .y(y[38]));
  Fx39 Fx39_inst(.x({x[59], x[57]}), .y(y[39]));
  Fx40 Fx40_inst(.x({x[61], x[60]}), .y(y[40]));
  Fx41 Fx41_inst(.x({x[62], x[60]}), .y(y[41]));
  Fx42 Fx42_inst(.x({x[64], x[63]}), .y(y[42]));
  Fx43 Fx43_inst(.x({x[65], x[63]}), .y(y[43]));
  Fx44 Fx44_inst(.x({x[67], x[66]}), .y(y[44]));
  Fx45 Fx45_inst(.x({x[68], x[66]}), .y(y[45]));
  Fx46 Fx46_inst(.x({x[70], x[69]}), .y(y[46]));
  Fx47 Fx47_inst(.x({x[71], x[69]}), .y(y[47]));
  Fx48 Fx48_inst(.x({x[73], x[72]}), .y(y[48]));
  Fx49 Fx49_inst(.x({x[74], x[72]}), .y(y[49]));
  Fx50 Fx50_inst(.x({x[76], x[75]}), .y(y[50]));
  Fx51 Fx51_inst(.x({x[77], x[75]}), .y(y[51]));
  Fx52 Fx52_inst(.x({x[79], x[78]}), .y(y[52]));
  Fx53 Fx53_inst(.x({x[80], x[78]}), .y(y[53]));
  Fx54 Fx54_inst(.x({x[82], x[81]}), .y(y[54]));
  Fx55 Fx55_inst(.x({x[83], x[81]}), .y(y[55]));
  Fx56 Fx56_inst(.x({x[85], x[84]}), .y(y[56]));
  Fx57 Fx57_inst(.x({x[86], x[84]}), .y(y[57]));
  Fx58 Fx58_inst(.x({x[88], x[87]}), .y(y[58]));
  Fx59 Fx59_inst(.x({x[89], x[87]}), .y(y[59]));
  Fx60 Fx60_inst(.x({x[91], x[90]}), .y(y[60]));
  Fx61 Fx61_inst(.x({x[92], x[90]}), .y(y[61]));
  Fx62 Fx62_inst(.x({x[94], x[93]}), .y(y[62]));
  Fx63 Fx63_inst(.x({x[95], x[93]}), .y(y[63]));
  Fx64 Fx64_inst(.x({x[97], x[96]}), .y(y[64]));
  Fx65 Fx65_inst(.x({x[98], x[96]}), .y(y[65]));
  Fx66 Fx66_inst(.x({x[100], x[99]}), .y(y[66]));
  Fx67 Fx67_inst(.x({x[101], x[99]}), .y(y[67]));
  Fx68 Fx68_inst(.x({x[103], x[102]}), .y(y[68]));
  Fx69 Fx69_inst(.x({x[104], x[102]}), .y(y[69]));
  Fx70 Fx70_inst(.x({x[106], x[105]}), .y(y[70]));
  Fx71 Fx71_inst(.x({x[107], x[105]}), .y(y[71]));
  Fx72 Fx72_inst(.x({x[109], x[108]}), .y(y[72]));
  Fx73 Fx73_inst(.x({x[110], x[108]}), .y(y[73]));
  Fx74 Fx74_inst(.x({x[112], x[111]}), .y(y[74]));
  Fx75 Fx75_inst(.x({x[113], x[111]}), .y(y[75]));
  Fx76 Fx76_inst(.x({x[115], x[114]}), .y(y[76]));
  Fx77 Fx77_inst(.x({x[116], x[114]}), .y(y[77]));
  Fx78 Fx78_inst(.x({x[118], x[117]}), .y(y[78]));
  Fx79 Fx79_inst(.x({x[119], x[117]}), .y(y[79]));
  Fx80 Fx80_inst(.x({x[121], x[120]}), .y(y[80]));
  Fx81 Fx81_inst(.x({x[122], x[120]}), .y(y[81]));
  Fx82 Fx82_inst(.x({x[124], x[123]}), .y(y[82]));
  Fx83 Fx83_inst(.x({x[125], x[123]}), .y(y[83]));
  Fx84 Fx84_inst(.x({x[127], x[126]}), .y(y[84]));
  Fx85 Fx85_inst(.x({x[128], x[126]}), .y(y[85]));
  Fx86 Fx86_inst(.x({x[130], x[129]}), .y(y[86]));
  Fx87 Fx87_inst(.x({x[131], x[129]}), .y(y[87]));
  Fx88 Fx88_inst(.x({x[133], x[132]}), .y(y[88]));
  Fx89 Fx89_inst(.x({x[134], x[132]}), .y(y[89]));
  Fx90 Fx90_inst(.x({x[136], x[135]}), .y(y[90]));
  Fx91 Fx91_inst(.x({x[137], x[135]}), .y(y[91]));
  Fx92 Fx92_inst(.x({x[139], x[138]}), .y(y[92]));
  Fx93 Fx93_inst(.x({x[140], x[138]}), .y(y[93]));
  Fx94 Fx94_inst(.x({x[142], x[141]}), .y(y[94]));
  Fx95 Fx95_inst(.x({x[143], x[141]}), .y(y[95]));
  Fx96 Fx96_inst(.x({x[145], x[144]}), .y(y[96]));
  Fx97 Fx97_inst(.x({x[146], x[144]}), .y(y[97]));
  Fx98 Fx98_inst(.x({x[148], x[147]}), .y(y[98]));
  Fx99 Fx99_inst(.x({x[149], x[147]}), .y(y[99]));
  Fx100 Fx100_inst(.x({x[151], x[150]}), .y(y[100]));
  Fx101 Fx101_inst(.x({x[152], x[150]}), .y(y[101]));
  Fx102 Fx102_inst(.x({x[154], x[153]}), .y(y[102]));
  Fx103 Fx103_inst(.x({x[155], x[153]}), .y(y[103]));
  Fx104 Fx104_inst(.x({x[157], x[156]}), .y(y[104]));
  Fx105 Fx105_inst(.x({x[158], x[156]}), .y(y[105]));
  Fx106 Fx106_inst(.x({x[160], x[159]}), .y(y[106]));
  Fx107 Fx107_inst(.x({x[161], x[159]}), .y(y[107]));
  Fx108 Fx108_inst(.x({x[163], x[162]}), .y(y[108]));
  Fx109 Fx109_inst(.x({x[164], x[162]}), .y(y[109]));
  Fx110 Fx110_inst(.x({x[166], x[165]}), .y(y[110]));
  Fx111 Fx111_inst(.x({x[167], x[165]}), .y(y[111]));
  Fx112 Fx112_inst(.x({x[169], x[168]}), .y(y[112]));
  Fx113 Fx113_inst(.x({x[170], x[168]}), .y(y[113]));
  Fx114 Fx114_inst(.x({x[172], x[171]}), .y(y[114]));
  Fx115 Fx115_inst(.x({x[173], x[171]}), .y(y[115]));
  Fx116 Fx116_inst(.x({x[175], x[174]}), .y(y[116]));
  Fx117 Fx117_inst(.x({x[176], x[174]}), .y(y[117]));
  Fx118 Fx118_inst(.x({x[178], x[177]}), .y(y[118]));
  Fx119 Fx119_inst(.x({x[179], x[177]}), .y(y[119]));
  Fx120 Fx120_inst(.x({x[181], x[180]}), .y(y[120]));
  Fx121 Fx121_inst(.x({x[182], x[180]}), .y(y[121]));
  Fx122 Fx122_inst(.x({x[184], x[183]}), .y(y[122]));
  Fx123 Fx123_inst(.x({x[185], x[183]}), .y(y[123]));
  Fx124 Fx124_inst(.x({x[187], x[186]}), .y(y[124]));
  Fx125 Fx125_inst(.x({x[188], x[186]}), .y(y[125]));
  Fx126 Fx126_inst(.x({x[190], x[189]}), .y(y[126]));
  Fx127 Fx127_inst(.x({x[191], x[189]}), .y(y[127]));
  Fx128 Fx128_inst(.x({x[193], x[192]}), .y(y[128]));
  Fx129 Fx129_inst(.x({x[194], x[192]}), .y(y[129]));
  Fx130 Fx130_inst(.x({x[196], x[195]}), .y(y[130]));
  Fx131 Fx131_inst(.x({x[197], x[195]}), .y(y[131]));
  Fx132 Fx132_inst(.x({x[199], x[198]}), .y(y[132]));
  Fx133 Fx133_inst(.x({x[200], x[198]}), .y(y[133]));
  Fx134 Fx134_inst(.x({x[202], x[201]}), .y(y[134]));
  Fx135 Fx135_inst(.x({x[203], x[201]}), .y(y[135]));
  Fx136 Fx136_inst(.x({x[205], x[204]}), .y(y[136]));
  Fx137 Fx137_inst(.x({x[206], x[204]}), .y(y[137]));
  Fx138 Fx138_inst(.x({x[208], x[207]}), .y(y[138]));
  Fx139 Fx139_inst(.x({x[209], x[207]}), .y(y[139]));
  Fx140 Fx140_inst(.x({x[211], x[210]}), .y(y[140]));
  Fx141 Fx141_inst(.x({x[212], x[210]}), .y(y[141]));
  Fx142 Fx142_inst(.x({x[214], x[213]}), .y(y[142]));
  Fx143 Fx143_inst(.x({x[215], x[213]}), .y(y[143]));
  Fx144 Fx144_inst(.x({x[217], x[216]}), .y(y[144]));
  Fx145 Fx145_inst(.x({x[218], x[216]}), .y(y[145]));
  Fx146 Fx146_inst(.x({x[220], x[219]}), .y(y[146]));
  Fx147 Fx147_inst(.x({x[221], x[219]}), .y(y[147]));
  Fx148 Fx148_inst(.x({x[223], x[222]}), .y(y[148]));
  Fx149 Fx149_inst(.x({x[224], x[222]}), .y(y[149]));
endmodule

module R1ind0(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind1(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind2(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind3(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind4(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind5(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind6(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind7(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind8(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind9(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind10(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind11(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind12(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind13(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind14(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind15(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind16(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind17(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind18(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind19(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind20(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind21(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind22(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind23(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind24(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind25(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind26(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind27(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind28(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind29(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind30(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind31(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind32(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind33(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind34(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind35(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind36(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind37(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind38(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind39(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind40(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind41(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind42(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind43(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind44(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind45(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind46(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind47(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind48(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind49(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind50(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind51(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind52(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind53(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind54(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind55(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind56(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind57(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind58(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind59(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind60(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind61(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind62(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind63(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind64(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind65(x, y);
 input [21:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = ~x[0] & t[12];
  assign t[10] = ~x[0] & t[17];
  assign t[11] = ~x[0] & t[18];
  assign t[12] = t[19] ^ x[3];
  assign t[13] = t[20] ^ x[6];
  assign t[14] = t[21] ^ x[9];
  assign t[15] = t[22] ^ x[12];
  assign t[16] = t[23] ^ x[15];
  assign t[17] = t[24] ^ x[18];
  assign t[18] = t[25] ^ x[21];
  assign t[19] = (x[1] & x[2]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[20] = (x[4] & x[5]);
  assign t[21] = (x[7] & x[8]);
  assign t[22] = (x[10] & x[11]);
  assign t[23] = (x[13] & x[14]);
  assign t[24] = (x[16] & x[17]);
  assign t[25] = (x[19] & x[20]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[7]);
  assign t[4] = ~(~x[0] & ~t[13]);
  assign t[5] = ~x[0] & t[14];
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~x[0] & t[15];
  assign t[9] = ~(~x[0] & ~t[16]);
  assign y = t[0] & t[1];
endmodule

module R1ind66(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = ~(t[0]);
endmodule

module R1ind67(x, y);
 input [6:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = ~t[2];
  assign t[1] = ~x[3] & t[3];
  assign t[2] = t[4] ^ x[2];
  assign t[3] = t[5] ^ x[6];
  assign t[4] = (x[0] & x[1]);
  assign t[5] = (x[4] & x[5]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind68(x, y);
 input [3:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = ~x[0] & t[2];
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (x[1] & x[2]);
  assign y = ~(t[0]);
endmodule

module R1ind69(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = ~x[0] & t[0];
endmodule

module R1ind70(x, y);
 input [6:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = ~x[0] & t[2];
  assign t[1] = ~(~x[0] & ~t[3]);
  assign t[2] = t[4] ^ x[3];
  assign t[3] = t[5] ^ x[6];
  assign t[4] = (x[1] & x[2]);
  assign t[5] = (x[4] & x[5]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind71(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = ~x[0] & t[0];
endmodule

module R1ind72(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = ~x[0] & t[0];
endmodule

module R1ind73(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = ~x[0] & t[0];
endmodule

module R1ind74(x, y);
 input [6:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = ~(~x[0] & ~t[2]);
  assign t[1] = ~x[0] & t[3];
  assign t[2] = t[4] ^ x[3];
  assign t[3] = t[5] ^ x[6];
  assign t[4] = (x[1] & x[2]);
  assign t[5] = (x[4] & x[5]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind75(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[1] ? x[3] : x[2];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind76(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[1] ? x[3] : x[2];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind77(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[1] ? x[3] : x[2];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind78(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[1] ? x[3] : x[2];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind79(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[1] ? x[3] : x[2];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind80(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[1] ? x[3] : x[2];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind81(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[1] ? x[3] : x[2];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind82(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[1] ? x[3] : x[2];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind83(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[1] ? x[3] : x[2];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind84(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[1] ? x[3] : x[2];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind85(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[1] ? x[3] : x[2];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind86(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[1] ? x[3] : x[2];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind87(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[1] ? x[3] : x[2];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind88(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[1] ? x[3] : x[2];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind89(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[1] ? x[3] : x[2];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind90(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[1] ? x[3] : x[2];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind91(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[1] ? x[3] : x[2];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind92(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[1] ? x[3] : x[2];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind93(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[1] ? x[3] : x[2];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind94(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[1] ? x[3] : x[2];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind95(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[1] ? x[3] : x[2];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind96(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[1] ? x[3] : x[2];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind97(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[1] ? x[3] : x[2];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind98(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[1] ? x[3] : x[2];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind99(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[1] ? x[3] : x[2];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind100(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[1] ? x[3] : x[2];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind101(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[1] ? x[3] : x[2];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind102(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[1] ? x[3] : x[2];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind103(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[1] ? x[3] : x[2];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind104(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[1] ? x[3] : x[2];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind105(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[1] ? x[3] : x[2];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind106(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[1] ? x[3] : x[2];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind107(x, y);
 input [5:0] x;
 output y;

 wire [4:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[1] ? x[3] : x[2];
  assign t[4] = x[1] ? x[5] : x[4];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind108(x, y);
 input [5:0] x;
 output y;

 wire [4:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[1] ? x[3] : x[2];
  assign t[4] = x[1] ? x[5] : x[4];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind109(x, y);
 input [5:0] x;
 output y;

 wire [4:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[1] ? x[3] : x[2];
  assign t[4] = x[1] ? x[5] : x[4];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind110(x, y);
 input [5:0] x;
 output y;

 wire [4:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[1] ? x[3] : x[2];
  assign t[4] = x[1] ? x[5] : x[4];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind111(x, y);
 input [5:0] x;
 output y;

 wire [4:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[1] ? x[3] : x[2];
  assign t[4] = x[1] ? x[5] : x[4];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind112(x, y);
 input [5:0] x;
 output y;

 wire [4:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[1] ? x[3] : x[2];
  assign t[4] = x[1] ? x[5] : x[4];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind113(x, y);
 input [5:0] x;
 output y;

 wire [4:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[1] ? x[3] : x[2];
  assign t[4] = x[1] ? x[5] : x[4];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind114(x, y);
 input [5:0] x;
 output y;

 wire [4:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[1] ? x[3] : x[2];
  assign t[4] = x[1] ? x[5] : x[4];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind115(x, y);
 input [5:0] x;
 output y;

 wire [4:0] t;
  assign t[0] = t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[1] ? x[3] : x[2];
  assign t[4] = x[1] ? x[5] : x[4];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind116(x, y);
 input [5:0] x;
 output y;

 wire [4:0] t;
  assign t[0] = t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[1] ? x[3] : x[2];
  assign t[4] = x[1] ? x[5] : x[4];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind117(x, y);
 input [5:0] x;
 output y;

 wire [4:0] t;
  assign t[0] = t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[1] ? x[3] : x[2];
  assign t[4] = x[1] ? x[5] : x[4];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind118(x, y);
 input [5:0] x;
 output y;

 wire [4:0] t;
  assign t[0] = t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[1] ? x[3] : x[2];
  assign t[4] = x[1] ? x[5] : x[4];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind119(x, y);
 input [5:0] x;
 output y;

 wire [4:0] t;
  assign t[0] = t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[1] ? x[3] : x[2];
  assign t[4] = x[1] ? x[5] : x[4];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind120(x, y);
 input [5:0] x;
 output y;

 wire [4:0] t;
  assign t[0] = t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[1] ? x[3] : x[2];
  assign t[4] = x[1] ? x[5] : x[4];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind121(x, y);
 input [5:0] x;
 output y;

 wire [4:0] t;
  assign t[0] = t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[1] ? x[3] : x[2];
  assign t[4] = x[1] ? x[5] : x[4];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind122(x, y);
 input [5:0] x;
 output y;

 wire [4:0] t;
  assign t[0] = t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[1] ? x[3] : x[2];
  assign t[4] = x[1] ? x[5] : x[4];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind123(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[1] ? x[3] : x[2];
  assign t[5] = x[1] ? x[5] : x[4];
  assign t[6] = x[1] ? x[7] : x[6];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind124(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[1] ? x[3] : x[2];
  assign t[5] = x[1] ? x[5] : x[4];
  assign t[6] = x[1] ? x[7] : x[6];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind125(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[1] ? x[3] : x[2];
  assign t[5] = x[1] ? x[5] : x[4];
  assign t[6] = x[1] ? x[7] : x[6];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind126(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[1] ? x[3] : x[2];
  assign t[5] = x[1] ? x[5] : x[4];
  assign t[6] = x[1] ? x[7] : x[6];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind127(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[1] ? x[3] : x[2];
  assign t[5] = x[1] ? x[5] : x[4];
  assign t[6] = x[1] ? x[7] : x[6];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind128(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[1] ? x[3] : x[2];
  assign t[5] = x[1] ? x[5] : x[4];
  assign t[6] = x[1] ? x[7] : x[6];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind129(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[1] ? x[3] : x[2];
  assign t[5] = x[1] ? x[5] : x[4];
  assign t[6] = x[1] ? x[7] : x[6];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind130(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[1] ? x[3] : x[2];
  assign t[5] = x[1] ? x[5] : x[4];
  assign t[6] = x[1] ? x[7] : x[6];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind131(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[1] ? x[3] : x[2];
  assign t[5] = x[1] ? x[5] : x[4];
  assign t[6] = x[1] ? x[7] : x[6];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind132(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[1] ? x[3] : x[2];
  assign t[5] = x[1] ? x[5] : x[4];
  assign t[6] = x[1] ? x[7] : x[6];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind133(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[1] ? x[3] : x[2];
  assign t[5] = x[1] ? x[5] : x[4];
  assign t[6] = x[1] ? x[7] : x[6];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind134(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[1] ? x[3] : x[2];
  assign t[5] = x[1] ? x[5] : x[4];
  assign t[6] = x[1] ? x[7] : x[6];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind135(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[1] ? x[3] : x[2];
  assign t[5] = x[1] ? x[5] : x[4];
  assign t[6] = x[1] ? x[7] : x[6];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind136(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[1] ? x[3] : x[2];
  assign t[5] = x[1] ? x[5] : x[4];
  assign t[6] = x[1] ? x[7] : x[6];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind137(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[1] ? x[3] : x[2];
  assign t[5] = x[1] ? x[5] : x[4];
  assign t[6] = x[1] ? x[7] : x[6];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind138(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[1] ? x[3] : x[2];
  assign t[5] = x[1] ? x[5] : x[4];
  assign t[6] = x[1] ? x[7] : x[6];
  assign y = ~(t[0] ^ x[0]);
endmodule

module R1ind139(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = ~x[0] & t[0];
endmodule

module R1ind140(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind141(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[12] ^ t[3];
  assign t[11] = t[13] & t[14];
  assign t[12] = t[15] & t[16];
  assign t[13] = ~(t[12] ^ t[17]);
  assign t[14] = t[2] ^ t[18];
  assign t[15] = ~(t[18]);
  assign t[16] = ~(t[6]);
  assign t[17] = t[4] ^ t[6];
  assign t[18] = t[9] ^ t[19];
  assign t[19] = t[23] ^ x[2];
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[24] ^ x[5];
  assign t[21] = t[25] ^ x[8];
  assign t[22] = t[26] ^ x[11];
  assign t[23] = (x[0] & x[1]);
  assign t[24] = (x[3] & x[4]);
  assign t[25] = (x[6] & x[7]);
  assign t[26] = (x[9] & x[10]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] & t[9];
  assign t[4] = t[19] ^ t[7];
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[20] ^ t[19];
  assign t[7] = ~(t[21]);
  assign t[8] = ~(t[19]);
  assign t[9] = t[6] ^ t[22];
  assign y = t[0] ^ t[1];
endmodule

module R1ind142(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind143(x, y);
 input [11:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[23] ^ t[21];
  assign t[11] = ~(t[21]);
  assign t[12] = t[10] ^ t[24];
  assign t[13] = ~(t[6] ^ t[15]);
  assign t[14] = t[16] ^ t[12];
  assign t[15] = t[17] ^ t[5];
  assign t[16] = t[21] ^ t[8];
  assign t[17] = t[18] & t[19];
  assign t[18] = ~(t[20]);
  assign t[19] = ~(t[10]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[12] ^ t[21];
  assign t[21] = t[25] ^ x[2];
  assign t[22] = t[26] ^ x[5];
  assign t[23] = t[27] ^ x[8];
  assign t[24] = t[28] ^ x[11];
  assign t[25] = (x[0] & x[1]);
  assign t[26] = (x[3] & x[4]);
  assign t[27] = (x[6] & x[7]);
  assign t[28] = (x[9] & x[10]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[10] ^ t[8];
  assign t[5] = t[11] & t[12];
  assign t[6] = t[10] ^ t[21];
  assign t[7] = t[13] & t[14];
  assign t[8] = ~(t[22]);
  assign t[9] = t[15] ^ t[7];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind144(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind145(x, y);
 input [11:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[14] ^ t[28];
  assign t[11] = t[19] & t[20];
  assign t[12] = ~(t[29]);
  assign t[13] = t[17] ^ t[11];
  assign t[14] = t[30] ^ t[28];
  assign t[15] = ~(t[28]);
  assign t[16] = t[14] ^ t[31];
  assign t[17] = t[21] ^ t[7];
  assign t[18] = t[22] & t[23];
  assign t[19] = ~(t[10] ^ t[17]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[8] ^ t[16];
  assign t[21] = t[24] & t[25];
  assign t[22] = ~(t[21] ^ t[26]);
  assign t[23] = t[6] ^ t[27];
  assign t[24] = ~(t[27]);
  assign t[25] = ~(t[14]);
  assign t[26] = t[8] ^ t[14];
  assign t[27] = t[16] ^ t[28];
  assign t[28] = t[32] ^ x[2];
  assign t[29] = t[33] ^ x[5];
  assign t[2] = t[6] ^ t[7];
  assign t[30] = t[34] ^ x[8];
  assign t[31] = t[35] ^ x[11];
  assign t[32] = (x[0] & x[1]);
  assign t[33] = (x[3] & x[4]);
  assign t[34] = (x[6] & x[7]);
  assign t[35] = (x[9] & x[10]);
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[10] ^ t[11];
  assign t[5] = t[12] ^ t[13];
  assign t[6] = t[14] ^ t[12];
  assign t[7] = t[15] & t[16];
  assign t[8] = t[28] ^ t[12];
  assign t[9] = t[17] ^ t[18];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind146(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind147(x, y);
 input [11:0] x;
 output y;

 wire [33:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[16] ^ t[7];
  assign t[11] = t[17] & t[18];
  assign t[12] = t[28] ^ t[27];
  assign t[13] = ~(t[27]);
  assign t[14] = t[12] ^ t[29];
  assign t[15] = t[19] & t[20];
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[23] ^ t[10]);
  assign t[18] = t[8] ^ t[14];
  assign t[19] = ~(t[16] ^ t[24]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[6] ^ t[25];
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[12]);
  assign t[23] = t[12] ^ t[27];
  assign t[24] = t[8] ^ t[12];
  assign t[25] = t[14] ^ t[27];
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[6] ^ t[7];
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[3] & x[4]);
  assign t[32] = (x[6] & x[7]);
  assign t[33] = (x[9] & x[10]);
  assign t[3] = t[8] ^ t[9];
  assign t[4] = ~(t[26]);
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[12] ^ t[4];
  assign t[7] = t[13] & t[14];
  assign t[8] = t[27] ^ t[4];
  assign t[9] = t[10] ^ t[15];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind148(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind149(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[12] ^ t[3];
  assign t[11] = t[13] & t[14];
  assign t[12] = t[15] & t[16];
  assign t[13] = ~(t[12] ^ t[17]);
  assign t[14] = t[2] ^ t[18];
  assign t[15] = ~(t[18]);
  assign t[16] = ~(t[6]);
  assign t[17] = t[4] ^ t[6];
  assign t[18] = t[9] ^ t[19];
  assign t[19] = t[23] ^ x[2];
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[24] ^ x[5];
  assign t[21] = t[25] ^ x[8];
  assign t[22] = t[26] ^ x[11];
  assign t[23] = (x[0] & x[1]);
  assign t[24] = (x[3] & x[4]);
  assign t[25] = (x[6] & x[7]);
  assign t[26] = (x[9] & x[10]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] & t[9];
  assign t[4] = t[19] ^ t[7];
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[20] ^ t[19];
  assign t[7] = ~(t[21]);
  assign t[8] = ~(t[19]);
  assign t[9] = t[6] ^ t[22];
  assign y = t[0] ^ t[1];
endmodule

module R1ind150(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind151(x, y);
 input [11:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[23] ^ t[21];
  assign t[11] = ~(t[21]);
  assign t[12] = t[10] ^ t[24];
  assign t[13] = ~(t[6] ^ t[15]);
  assign t[14] = t[16] ^ t[12];
  assign t[15] = t[17] ^ t[5];
  assign t[16] = t[21] ^ t[8];
  assign t[17] = t[18] & t[19];
  assign t[18] = ~(t[20]);
  assign t[19] = ~(t[10]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[12] ^ t[21];
  assign t[21] = t[25] ^ x[2];
  assign t[22] = t[26] ^ x[5];
  assign t[23] = t[27] ^ x[8];
  assign t[24] = t[28] ^ x[11];
  assign t[25] = (x[0] & x[1]);
  assign t[26] = (x[3] & x[4]);
  assign t[27] = (x[6] & x[7]);
  assign t[28] = (x[9] & x[10]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[10] ^ t[8];
  assign t[5] = t[11] & t[12];
  assign t[6] = t[10] ^ t[21];
  assign t[7] = t[13] & t[14];
  assign t[8] = ~(t[22]);
  assign t[9] = t[15] ^ t[7];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind152(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind153(x, y);
 input [11:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[14] ^ t[28];
  assign t[11] = t[19] & t[20];
  assign t[12] = ~(t[29]);
  assign t[13] = t[17] ^ t[11];
  assign t[14] = t[30] ^ t[28];
  assign t[15] = ~(t[28]);
  assign t[16] = t[14] ^ t[31];
  assign t[17] = t[21] ^ t[7];
  assign t[18] = t[22] & t[23];
  assign t[19] = ~(t[10] ^ t[17]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[8] ^ t[16];
  assign t[21] = t[24] & t[25];
  assign t[22] = ~(t[21] ^ t[26]);
  assign t[23] = t[6] ^ t[27];
  assign t[24] = ~(t[27]);
  assign t[25] = ~(t[14]);
  assign t[26] = t[8] ^ t[14];
  assign t[27] = t[16] ^ t[28];
  assign t[28] = t[32] ^ x[2];
  assign t[29] = t[33] ^ x[5];
  assign t[2] = t[6] ^ t[7];
  assign t[30] = t[34] ^ x[8];
  assign t[31] = t[35] ^ x[11];
  assign t[32] = (x[0] & x[1]);
  assign t[33] = (x[3] & x[4]);
  assign t[34] = (x[6] & x[7]);
  assign t[35] = (x[9] & x[10]);
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[10] ^ t[11];
  assign t[5] = t[12] ^ t[13];
  assign t[6] = t[14] ^ t[12];
  assign t[7] = t[15] & t[16];
  assign t[8] = t[28] ^ t[12];
  assign t[9] = t[17] ^ t[18];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind154(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind155(x, y);
 input [11:0] x;
 output y;

 wire [33:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[16] ^ t[7];
  assign t[11] = t[17] & t[18];
  assign t[12] = t[28] ^ t[27];
  assign t[13] = ~(t[27]);
  assign t[14] = t[12] ^ t[29];
  assign t[15] = t[19] & t[20];
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[23] ^ t[10]);
  assign t[18] = t[8] ^ t[14];
  assign t[19] = ~(t[16] ^ t[24]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[6] ^ t[25];
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[12]);
  assign t[23] = t[12] ^ t[27];
  assign t[24] = t[8] ^ t[12];
  assign t[25] = t[14] ^ t[27];
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[6] ^ t[7];
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[3] & x[4]);
  assign t[32] = (x[6] & x[7]);
  assign t[33] = (x[9] & x[10]);
  assign t[3] = t[8] ^ t[9];
  assign t[4] = ~(t[26]);
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[12] ^ t[4];
  assign t[7] = t[13] & t[14];
  assign t[8] = t[27] ^ t[4];
  assign t[9] = t[10] ^ t[15];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind156(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind157(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[12] ^ t[3];
  assign t[11] = t[13] & t[14];
  assign t[12] = t[15] & t[16];
  assign t[13] = ~(t[12] ^ t[17]);
  assign t[14] = t[2] ^ t[18];
  assign t[15] = ~(t[18]);
  assign t[16] = ~(t[6]);
  assign t[17] = t[4] ^ t[6];
  assign t[18] = t[9] ^ t[19];
  assign t[19] = t[23] ^ x[2];
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[24] ^ x[5];
  assign t[21] = t[25] ^ x[8];
  assign t[22] = t[26] ^ x[11];
  assign t[23] = (x[0] & x[1]);
  assign t[24] = (x[3] & x[4]);
  assign t[25] = (x[6] & x[7]);
  assign t[26] = (x[9] & x[10]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] & t[9];
  assign t[4] = t[19] ^ t[7];
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[20] ^ t[19];
  assign t[7] = ~(t[21]);
  assign t[8] = ~(t[19]);
  assign t[9] = t[6] ^ t[22];
  assign y = t[0] ^ t[1];
endmodule

module R1ind158(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind159(x, y);
 input [11:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[23] ^ t[21];
  assign t[11] = ~(t[21]);
  assign t[12] = t[10] ^ t[24];
  assign t[13] = ~(t[6] ^ t[15]);
  assign t[14] = t[16] ^ t[12];
  assign t[15] = t[17] ^ t[5];
  assign t[16] = t[21] ^ t[8];
  assign t[17] = t[18] & t[19];
  assign t[18] = ~(t[20]);
  assign t[19] = ~(t[10]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[12] ^ t[21];
  assign t[21] = t[25] ^ x[2];
  assign t[22] = t[26] ^ x[5];
  assign t[23] = t[27] ^ x[8];
  assign t[24] = t[28] ^ x[11];
  assign t[25] = (x[0] & x[1]);
  assign t[26] = (x[3] & x[4]);
  assign t[27] = (x[6] & x[7]);
  assign t[28] = (x[9] & x[10]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[10] ^ t[8];
  assign t[5] = t[11] & t[12];
  assign t[6] = t[10] ^ t[21];
  assign t[7] = t[13] & t[14];
  assign t[8] = ~(t[22]);
  assign t[9] = t[15] ^ t[7];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind160(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind161(x, y);
 input [11:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[14] ^ t[28];
  assign t[11] = t[19] & t[20];
  assign t[12] = ~(t[29]);
  assign t[13] = t[17] ^ t[11];
  assign t[14] = t[30] ^ t[28];
  assign t[15] = ~(t[28]);
  assign t[16] = t[14] ^ t[31];
  assign t[17] = t[21] ^ t[7];
  assign t[18] = t[22] & t[23];
  assign t[19] = ~(t[10] ^ t[17]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[8] ^ t[16];
  assign t[21] = t[24] & t[25];
  assign t[22] = ~(t[21] ^ t[26]);
  assign t[23] = t[6] ^ t[27];
  assign t[24] = ~(t[27]);
  assign t[25] = ~(t[14]);
  assign t[26] = t[8] ^ t[14];
  assign t[27] = t[16] ^ t[28];
  assign t[28] = t[32] ^ x[2];
  assign t[29] = t[33] ^ x[5];
  assign t[2] = t[6] ^ t[7];
  assign t[30] = t[34] ^ x[8];
  assign t[31] = t[35] ^ x[11];
  assign t[32] = (x[0] & x[1]);
  assign t[33] = (x[3] & x[4]);
  assign t[34] = (x[6] & x[7]);
  assign t[35] = (x[9] & x[10]);
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[10] ^ t[11];
  assign t[5] = t[12] ^ t[13];
  assign t[6] = t[14] ^ t[12];
  assign t[7] = t[15] & t[16];
  assign t[8] = t[28] ^ t[12];
  assign t[9] = t[17] ^ t[18];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind162(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind163(x, y);
 input [11:0] x;
 output y;

 wire [33:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[16] ^ t[7];
  assign t[11] = t[17] & t[18];
  assign t[12] = t[28] ^ t[27];
  assign t[13] = ~(t[27]);
  assign t[14] = t[12] ^ t[29];
  assign t[15] = t[19] & t[20];
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[23] ^ t[10]);
  assign t[18] = t[8] ^ t[14];
  assign t[19] = ~(t[16] ^ t[24]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[6] ^ t[25];
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[12]);
  assign t[23] = t[12] ^ t[27];
  assign t[24] = t[8] ^ t[12];
  assign t[25] = t[14] ^ t[27];
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[6] ^ t[7];
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[3] & x[4]);
  assign t[32] = (x[6] & x[7]);
  assign t[33] = (x[9] & x[10]);
  assign t[3] = t[8] ^ t[9];
  assign t[4] = ~(t[26]);
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[12] ^ t[4];
  assign t[7] = t[13] & t[14];
  assign t[8] = t[27] ^ t[4];
  assign t[9] = t[10] ^ t[15];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind164(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind165(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[12] ^ t[3];
  assign t[11] = t[13] & t[14];
  assign t[12] = t[15] & t[16];
  assign t[13] = ~(t[12] ^ t[17]);
  assign t[14] = t[2] ^ t[18];
  assign t[15] = ~(t[18]);
  assign t[16] = ~(t[6]);
  assign t[17] = t[4] ^ t[6];
  assign t[18] = t[9] ^ t[19];
  assign t[19] = t[23] ^ x[2];
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[24] ^ x[5];
  assign t[21] = t[25] ^ x[8];
  assign t[22] = t[26] ^ x[11];
  assign t[23] = (x[0] & x[1]);
  assign t[24] = (x[3] & x[4]);
  assign t[25] = (x[6] & x[7]);
  assign t[26] = (x[9] & x[10]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] & t[9];
  assign t[4] = t[19] ^ t[7];
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[20] ^ t[19];
  assign t[7] = ~(t[21]);
  assign t[8] = ~(t[19]);
  assign t[9] = t[6] ^ t[22];
  assign y = t[0] ^ t[1];
endmodule

module R1ind166(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind167(x, y);
 input [11:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[23] ^ t[21];
  assign t[11] = ~(t[21]);
  assign t[12] = t[10] ^ t[24];
  assign t[13] = ~(t[6] ^ t[15]);
  assign t[14] = t[16] ^ t[12];
  assign t[15] = t[17] ^ t[5];
  assign t[16] = t[21] ^ t[8];
  assign t[17] = t[18] & t[19];
  assign t[18] = ~(t[20]);
  assign t[19] = ~(t[10]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[12] ^ t[21];
  assign t[21] = t[25] ^ x[2];
  assign t[22] = t[26] ^ x[5];
  assign t[23] = t[27] ^ x[8];
  assign t[24] = t[28] ^ x[11];
  assign t[25] = (x[0] & x[1]);
  assign t[26] = (x[3] & x[4]);
  assign t[27] = (x[6] & x[7]);
  assign t[28] = (x[9] & x[10]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[10] ^ t[8];
  assign t[5] = t[11] & t[12];
  assign t[6] = t[10] ^ t[21];
  assign t[7] = t[13] & t[14];
  assign t[8] = ~(t[22]);
  assign t[9] = t[15] ^ t[7];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind168(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind169(x, y);
 input [11:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[14] ^ t[28];
  assign t[11] = t[19] & t[20];
  assign t[12] = ~(t[29]);
  assign t[13] = t[17] ^ t[11];
  assign t[14] = t[30] ^ t[28];
  assign t[15] = ~(t[28]);
  assign t[16] = t[14] ^ t[31];
  assign t[17] = t[21] ^ t[7];
  assign t[18] = t[22] & t[23];
  assign t[19] = ~(t[10] ^ t[17]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[8] ^ t[16];
  assign t[21] = t[24] & t[25];
  assign t[22] = ~(t[21] ^ t[26]);
  assign t[23] = t[6] ^ t[27];
  assign t[24] = ~(t[27]);
  assign t[25] = ~(t[14]);
  assign t[26] = t[8] ^ t[14];
  assign t[27] = t[16] ^ t[28];
  assign t[28] = t[32] ^ x[2];
  assign t[29] = t[33] ^ x[5];
  assign t[2] = t[6] ^ t[7];
  assign t[30] = t[34] ^ x[8];
  assign t[31] = t[35] ^ x[11];
  assign t[32] = (x[0] & x[1]);
  assign t[33] = (x[3] & x[4]);
  assign t[34] = (x[6] & x[7]);
  assign t[35] = (x[9] & x[10]);
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[10] ^ t[11];
  assign t[5] = t[12] ^ t[13];
  assign t[6] = t[14] ^ t[12];
  assign t[7] = t[15] & t[16];
  assign t[8] = t[28] ^ t[12];
  assign t[9] = t[17] ^ t[18];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind170(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind171(x, y);
 input [11:0] x;
 output y;

 wire [33:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[16] ^ t[7];
  assign t[11] = t[17] & t[18];
  assign t[12] = t[28] ^ t[27];
  assign t[13] = ~(t[27]);
  assign t[14] = t[12] ^ t[29];
  assign t[15] = t[19] & t[20];
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[23] ^ t[10]);
  assign t[18] = t[8] ^ t[14];
  assign t[19] = ~(t[16] ^ t[24]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[6] ^ t[25];
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[12]);
  assign t[23] = t[12] ^ t[27];
  assign t[24] = t[8] ^ t[12];
  assign t[25] = t[14] ^ t[27];
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[6] ^ t[7];
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[3] & x[4]);
  assign t[32] = (x[6] & x[7]);
  assign t[33] = (x[9] & x[10]);
  assign t[3] = t[8] ^ t[9];
  assign t[4] = ~(t[26]);
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[12] ^ t[4];
  assign t[7] = t[13] & t[14];
  assign t[8] = t[27] ^ t[4];
  assign t[9] = t[10] ^ t[15];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind172(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind173(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[12] ^ t[3];
  assign t[11] = t[13] & t[14];
  assign t[12] = t[15] & t[16];
  assign t[13] = ~(t[12] ^ t[17]);
  assign t[14] = t[2] ^ t[18];
  assign t[15] = ~(t[18]);
  assign t[16] = ~(t[6]);
  assign t[17] = t[4] ^ t[6];
  assign t[18] = t[9] ^ t[19];
  assign t[19] = t[23] ^ x[2];
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[24] ^ x[5];
  assign t[21] = t[25] ^ x[8];
  assign t[22] = t[26] ^ x[11];
  assign t[23] = (x[0] & x[1]);
  assign t[24] = (x[3] & x[4]);
  assign t[25] = (x[6] & x[7]);
  assign t[26] = (x[9] & x[10]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] & t[9];
  assign t[4] = t[19] ^ t[7];
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[20] ^ t[19];
  assign t[7] = ~(t[21]);
  assign t[8] = ~(t[19]);
  assign t[9] = t[6] ^ t[22];
  assign y = t[0] ^ t[1];
endmodule

module R1ind174(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind175(x, y);
 input [11:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[23] ^ t[21];
  assign t[11] = ~(t[21]);
  assign t[12] = t[10] ^ t[24];
  assign t[13] = ~(t[6] ^ t[15]);
  assign t[14] = t[16] ^ t[12];
  assign t[15] = t[17] ^ t[5];
  assign t[16] = t[21] ^ t[8];
  assign t[17] = t[18] & t[19];
  assign t[18] = ~(t[20]);
  assign t[19] = ~(t[10]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[12] ^ t[21];
  assign t[21] = t[25] ^ x[2];
  assign t[22] = t[26] ^ x[5];
  assign t[23] = t[27] ^ x[8];
  assign t[24] = t[28] ^ x[11];
  assign t[25] = (x[0] & x[1]);
  assign t[26] = (x[3] & x[4]);
  assign t[27] = (x[6] & x[7]);
  assign t[28] = (x[9] & x[10]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[10] ^ t[8];
  assign t[5] = t[11] & t[12];
  assign t[6] = t[10] ^ t[21];
  assign t[7] = t[13] & t[14];
  assign t[8] = ~(t[22]);
  assign t[9] = t[15] ^ t[7];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind176(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind177(x, y);
 input [11:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[14] ^ t[28];
  assign t[11] = t[19] & t[20];
  assign t[12] = ~(t[29]);
  assign t[13] = t[17] ^ t[11];
  assign t[14] = t[30] ^ t[28];
  assign t[15] = ~(t[28]);
  assign t[16] = t[14] ^ t[31];
  assign t[17] = t[21] ^ t[7];
  assign t[18] = t[22] & t[23];
  assign t[19] = ~(t[10] ^ t[17]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[8] ^ t[16];
  assign t[21] = t[24] & t[25];
  assign t[22] = ~(t[21] ^ t[26]);
  assign t[23] = t[6] ^ t[27];
  assign t[24] = ~(t[27]);
  assign t[25] = ~(t[14]);
  assign t[26] = t[8] ^ t[14];
  assign t[27] = t[16] ^ t[28];
  assign t[28] = t[32] ^ x[2];
  assign t[29] = t[33] ^ x[5];
  assign t[2] = t[6] ^ t[7];
  assign t[30] = t[34] ^ x[8];
  assign t[31] = t[35] ^ x[11];
  assign t[32] = (x[0] & x[1]);
  assign t[33] = (x[3] & x[4]);
  assign t[34] = (x[6] & x[7]);
  assign t[35] = (x[9] & x[10]);
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[10] ^ t[11];
  assign t[5] = t[12] ^ t[13];
  assign t[6] = t[14] ^ t[12];
  assign t[7] = t[15] & t[16];
  assign t[8] = t[28] ^ t[12];
  assign t[9] = t[17] ^ t[18];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind178(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind179(x, y);
 input [11:0] x;
 output y;

 wire [33:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[16] ^ t[7];
  assign t[11] = t[17] & t[18];
  assign t[12] = t[28] ^ t[27];
  assign t[13] = ~(t[27]);
  assign t[14] = t[12] ^ t[29];
  assign t[15] = t[19] & t[20];
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[23] ^ t[10]);
  assign t[18] = t[8] ^ t[14];
  assign t[19] = ~(t[16] ^ t[24]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[6] ^ t[25];
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[12]);
  assign t[23] = t[12] ^ t[27];
  assign t[24] = t[8] ^ t[12];
  assign t[25] = t[14] ^ t[27];
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[6] ^ t[7];
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[3] & x[4]);
  assign t[32] = (x[6] & x[7]);
  assign t[33] = (x[9] & x[10]);
  assign t[3] = t[8] ^ t[9];
  assign t[4] = ~(t[26]);
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[12] ^ t[4];
  assign t[7] = t[13] & t[14];
  assign t[8] = t[27] ^ t[4];
  assign t[9] = t[10] ^ t[15];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind180(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind181(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[12] ^ t[3];
  assign t[11] = t[13] & t[14];
  assign t[12] = t[15] & t[16];
  assign t[13] = ~(t[12] ^ t[17]);
  assign t[14] = t[2] ^ t[18];
  assign t[15] = ~(t[18]);
  assign t[16] = ~(t[6]);
  assign t[17] = t[4] ^ t[6];
  assign t[18] = t[9] ^ t[19];
  assign t[19] = t[23] ^ x[2];
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[24] ^ x[5];
  assign t[21] = t[25] ^ x[8];
  assign t[22] = t[26] ^ x[11];
  assign t[23] = (x[0] & x[1]);
  assign t[24] = (x[3] & x[4]);
  assign t[25] = (x[6] & x[7]);
  assign t[26] = (x[9] & x[10]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] & t[9];
  assign t[4] = t[19] ^ t[7];
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[20] ^ t[19];
  assign t[7] = ~(t[21]);
  assign t[8] = ~(t[19]);
  assign t[9] = t[6] ^ t[22];
  assign y = t[0] ^ t[1];
endmodule

module R1ind182(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind183(x, y);
 input [11:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[23] ^ t[21];
  assign t[11] = ~(t[21]);
  assign t[12] = t[10] ^ t[24];
  assign t[13] = ~(t[6] ^ t[15]);
  assign t[14] = t[16] ^ t[12];
  assign t[15] = t[17] ^ t[5];
  assign t[16] = t[21] ^ t[8];
  assign t[17] = t[18] & t[19];
  assign t[18] = ~(t[20]);
  assign t[19] = ~(t[10]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[12] ^ t[21];
  assign t[21] = t[25] ^ x[2];
  assign t[22] = t[26] ^ x[5];
  assign t[23] = t[27] ^ x[8];
  assign t[24] = t[28] ^ x[11];
  assign t[25] = (x[0] & x[1]);
  assign t[26] = (x[3] & x[4]);
  assign t[27] = (x[6] & x[7]);
  assign t[28] = (x[9] & x[10]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[10] ^ t[8];
  assign t[5] = t[11] & t[12];
  assign t[6] = t[10] ^ t[21];
  assign t[7] = t[13] & t[14];
  assign t[8] = ~(t[22]);
  assign t[9] = t[15] ^ t[7];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind184(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind185(x, y);
 input [11:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[14] ^ t[28];
  assign t[11] = t[19] & t[20];
  assign t[12] = ~(t[29]);
  assign t[13] = t[17] ^ t[11];
  assign t[14] = t[30] ^ t[28];
  assign t[15] = ~(t[28]);
  assign t[16] = t[14] ^ t[31];
  assign t[17] = t[21] ^ t[7];
  assign t[18] = t[22] & t[23];
  assign t[19] = ~(t[10] ^ t[17]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[8] ^ t[16];
  assign t[21] = t[24] & t[25];
  assign t[22] = ~(t[21] ^ t[26]);
  assign t[23] = t[6] ^ t[27];
  assign t[24] = ~(t[27]);
  assign t[25] = ~(t[14]);
  assign t[26] = t[8] ^ t[14];
  assign t[27] = t[16] ^ t[28];
  assign t[28] = t[32] ^ x[2];
  assign t[29] = t[33] ^ x[5];
  assign t[2] = t[6] ^ t[7];
  assign t[30] = t[34] ^ x[8];
  assign t[31] = t[35] ^ x[11];
  assign t[32] = (x[0] & x[1]);
  assign t[33] = (x[3] & x[4]);
  assign t[34] = (x[6] & x[7]);
  assign t[35] = (x[9] & x[10]);
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[10] ^ t[11];
  assign t[5] = t[12] ^ t[13];
  assign t[6] = t[14] ^ t[12];
  assign t[7] = t[15] & t[16];
  assign t[8] = t[28] ^ t[12];
  assign t[9] = t[17] ^ t[18];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind186(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind187(x, y);
 input [11:0] x;
 output y;

 wire [33:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[16] ^ t[7];
  assign t[11] = t[17] & t[18];
  assign t[12] = t[28] ^ t[27];
  assign t[13] = ~(t[27]);
  assign t[14] = t[12] ^ t[29];
  assign t[15] = t[19] & t[20];
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[23] ^ t[10]);
  assign t[18] = t[8] ^ t[14];
  assign t[19] = ~(t[16] ^ t[24]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[6] ^ t[25];
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[12]);
  assign t[23] = t[12] ^ t[27];
  assign t[24] = t[8] ^ t[12];
  assign t[25] = t[14] ^ t[27];
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[6] ^ t[7];
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[3] & x[4]);
  assign t[32] = (x[6] & x[7]);
  assign t[33] = (x[9] & x[10]);
  assign t[3] = t[8] ^ t[9];
  assign t[4] = ~(t[26]);
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[12] ^ t[4];
  assign t[7] = t[13] & t[14];
  assign t[8] = t[27] ^ t[4];
  assign t[9] = t[10] ^ t[15];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind188(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind189(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[12] ^ t[3];
  assign t[11] = t[13] & t[14];
  assign t[12] = t[15] & t[16];
  assign t[13] = ~(t[12] ^ t[17]);
  assign t[14] = t[2] ^ t[18];
  assign t[15] = ~(t[18]);
  assign t[16] = ~(t[6]);
  assign t[17] = t[4] ^ t[6];
  assign t[18] = t[9] ^ t[19];
  assign t[19] = t[23] ^ x[2];
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[24] ^ x[5];
  assign t[21] = t[25] ^ x[8];
  assign t[22] = t[26] ^ x[11];
  assign t[23] = (x[0] & x[1]);
  assign t[24] = (x[3] & x[4]);
  assign t[25] = (x[6] & x[7]);
  assign t[26] = (x[9] & x[10]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] & t[9];
  assign t[4] = t[19] ^ t[7];
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[20] ^ t[19];
  assign t[7] = ~(t[21]);
  assign t[8] = ~(t[19]);
  assign t[9] = t[6] ^ t[22];
  assign y = t[0] ^ t[1];
endmodule

module R1ind190(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind191(x, y);
 input [11:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[23] ^ t[21];
  assign t[11] = ~(t[21]);
  assign t[12] = t[10] ^ t[24];
  assign t[13] = ~(t[6] ^ t[15]);
  assign t[14] = t[16] ^ t[12];
  assign t[15] = t[17] ^ t[5];
  assign t[16] = t[21] ^ t[8];
  assign t[17] = t[18] & t[19];
  assign t[18] = ~(t[20]);
  assign t[19] = ~(t[10]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[12] ^ t[21];
  assign t[21] = t[25] ^ x[2];
  assign t[22] = t[26] ^ x[5];
  assign t[23] = t[27] ^ x[8];
  assign t[24] = t[28] ^ x[11];
  assign t[25] = (x[0] & x[1]);
  assign t[26] = (x[3] & x[4]);
  assign t[27] = (x[6] & x[7]);
  assign t[28] = (x[9] & x[10]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[10] ^ t[8];
  assign t[5] = t[11] & t[12];
  assign t[6] = t[10] ^ t[21];
  assign t[7] = t[13] & t[14];
  assign t[8] = ~(t[22]);
  assign t[9] = t[15] ^ t[7];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind192(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind193(x, y);
 input [11:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[14] ^ t[28];
  assign t[11] = t[19] & t[20];
  assign t[12] = ~(t[29]);
  assign t[13] = t[17] ^ t[11];
  assign t[14] = t[30] ^ t[28];
  assign t[15] = ~(t[28]);
  assign t[16] = t[14] ^ t[31];
  assign t[17] = t[21] ^ t[7];
  assign t[18] = t[22] & t[23];
  assign t[19] = ~(t[10] ^ t[17]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[8] ^ t[16];
  assign t[21] = t[24] & t[25];
  assign t[22] = ~(t[21] ^ t[26]);
  assign t[23] = t[6] ^ t[27];
  assign t[24] = ~(t[27]);
  assign t[25] = ~(t[14]);
  assign t[26] = t[8] ^ t[14];
  assign t[27] = t[16] ^ t[28];
  assign t[28] = t[32] ^ x[2];
  assign t[29] = t[33] ^ x[5];
  assign t[2] = t[6] ^ t[7];
  assign t[30] = t[34] ^ x[8];
  assign t[31] = t[35] ^ x[11];
  assign t[32] = (x[0] & x[1]);
  assign t[33] = (x[3] & x[4]);
  assign t[34] = (x[6] & x[7]);
  assign t[35] = (x[9] & x[10]);
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[10] ^ t[11];
  assign t[5] = t[12] ^ t[13];
  assign t[6] = t[14] ^ t[12];
  assign t[7] = t[15] & t[16];
  assign t[8] = t[28] ^ t[12];
  assign t[9] = t[17] ^ t[18];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind194(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind195(x, y);
 input [11:0] x;
 output y;

 wire [33:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[16] ^ t[7];
  assign t[11] = t[17] & t[18];
  assign t[12] = t[28] ^ t[27];
  assign t[13] = ~(t[27]);
  assign t[14] = t[12] ^ t[29];
  assign t[15] = t[19] & t[20];
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[23] ^ t[10]);
  assign t[18] = t[8] ^ t[14];
  assign t[19] = ~(t[16] ^ t[24]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[6] ^ t[25];
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[12]);
  assign t[23] = t[12] ^ t[27];
  assign t[24] = t[8] ^ t[12];
  assign t[25] = t[14] ^ t[27];
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[6] ^ t[7];
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[3] & x[4]);
  assign t[32] = (x[6] & x[7]);
  assign t[33] = (x[9] & x[10]);
  assign t[3] = t[8] ^ t[9];
  assign t[4] = ~(t[26]);
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[12] ^ t[4];
  assign t[7] = t[13] & t[14];
  assign t[8] = t[27] ^ t[4];
  assign t[9] = t[10] ^ t[15];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind196(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind197(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[12] ^ t[3];
  assign t[11] = t[13] & t[14];
  assign t[12] = t[15] & t[16];
  assign t[13] = ~(t[12] ^ t[17]);
  assign t[14] = t[2] ^ t[18];
  assign t[15] = ~(t[18]);
  assign t[16] = ~(t[6]);
  assign t[17] = t[4] ^ t[6];
  assign t[18] = t[9] ^ t[19];
  assign t[19] = t[23] ^ x[2];
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[24] ^ x[5];
  assign t[21] = t[25] ^ x[8];
  assign t[22] = t[26] ^ x[11];
  assign t[23] = (x[0] & x[1]);
  assign t[24] = (x[3] & x[4]);
  assign t[25] = (x[6] & x[7]);
  assign t[26] = (x[9] & x[10]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] & t[9];
  assign t[4] = t[19] ^ t[7];
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[20] ^ t[19];
  assign t[7] = ~(t[21]);
  assign t[8] = ~(t[19]);
  assign t[9] = t[6] ^ t[22];
  assign y = t[0] ^ t[1];
endmodule

module R1ind198(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind199(x, y);
 input [11:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[23] ^ t[21];
  assign t[11] = ~(t[21]);
  assign t[12] = t[10] ^ t[24];
  assign t[13] = ~(t[6] ^ t[15]);
  assign t[14] = t[16] ^ t[12];
  assign t[15] = t[17] ^ t[5];
  assign t[16] = t[21] ^ t[8];
  assign t[17] = t[18] & t[19];
  assign t[18] = ~(t[20]);
  assign t[19] = ~(t[10]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[12] ^ t[21];
  assign t[21] = t[25] ^ x[2];
  assign t[22] = t[26] ^ x[5];
  assign t[23] = t[27] ^ x[8];
  assign t[24] = t[28] ^ x[11];
  assign t[25] = (x[0] & x[1]);
  assign t[26] = (x[3] & x[4]);
  assign t[27] = (x[6] & x[7]);
  assign t[28] = (x[9] & x[10]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[10] ^ t[8];
  assign t[5] = t[11] & t[12];
  assign t[6] = t[10] ^ t[21];
  assign t[7] = t[13] & t[14];
  assign t[8] = ~(t[22]);
  assign t[9] = t[15] ^ t[7];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind200(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind201(x, y);
 input [11:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[14] ^ t[28];
  assign t[11] = t[19] & t[20];
  assign t[12] = ~(t[29]);
  assign t[13] = t[17] ^ t[11];
  assign t[14] = t[30] ^ t[28];
  assign t[15] = ~(t[28]);
  assign t[16] = t[14] ^ t[31];
  assign t[17] = t[21] ^ t[7];
  assign t[18] = t[22] & t[23];
  assign t[19] = ~(t[10] ^ t[17]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[8] ^ t[16];
  assign t[21] = t[24] & t[25];
  assign t[22] = ~(t[21] ^ t[26]);
  assign t[23] = t[6] ^ t[27];
  assign t[24] = ~(t[27]);
  assign t[25] = ~(t[14]);
  assign t[26] = t[8] ^ t[14];
  assign t[27] = t[16] ^ t[28];
  assign t[28] = t[32] ^ x[2];
  assign t[29] = t[33] ^ x[5];
  assign t[2] = t[6] ^ t[7];
  assign t[30] = t[34] ^ x[8];
  assign t[31] = t[35] ^ x[11];
  assign t[32] = (x[0] & x[1]);
  assign t[33] = (x[3] & x[4]);
  assign t[34] = (x[6] & x[7]);
  assign t[35] = (x[9] & x[10]);
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[10] ^ t[11];
  assign t[5] = t[12] ^ t[13];
  assign t[6] = t[14] ^ t[12];
  assign t[7] = t[15] & t[16];
  assign t[8] = t[28] ^ t[12];
  assign t[9] = t[17] ^ t[18];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind202(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind203(x, y);
 input [11:0] x;
 output y;

 wire [33:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[16] ^ t[7];
  assign t[11] = t[17] & t[18];
  assign t[12] = t[28] ^ t[27];
  assign t[13] = ~(t[27]);
  assign t[14] = t[12] ^ t[29];
  assign t[15] = t[19] & t[20];
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[23] ^ t[10]);
  assign t[18] = t[8] ^ t[14];
  assign t[19] = ~(t[16] ^ t[24]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[6] ^ t[25];
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[12]);
  assign t[23] = t[12] ^ t[27];
  assign t[24] = t[8] ^ t[12];
  assign t[25] = t[14] ^ t[27];
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[6] ^ t[7];
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[3] & x[4]);
  assign t[32] = (x[6] & x[7]);
  assign t[33] = (x[9] & x[10]);
  assign t[3] = t[8] ^ t[9];
  assign t[4] = ~(t[26]);
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[12] ^ t[4];
  assign t[7] = t[13] & t[14];
  assign t[8] = t[27] ^ t[4];
  assign t[9] = t[10] ^ t[15];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind204(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind205(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[12] ^ t[3];
  assign t[11] = t[13] & t[14];
  assign t[12] = t[15] & t[16];
  assign t[13] = ~(t[12] ^ t[17]);
  assign t[14] = t[2] ^ t[18];
  assign t[15] = ~(t[18]);
  assign t[16] = ~(t[6]);
  assign t[17] = t[4] ^ t[6];
  assign t[18] = t[9] ^ t[19];
  assign t[19] = t[23] ^ x[2];
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[24] ^ x[5];
  assign t[21] = t[25] ^ x[8];
  assign t[22] = t[26] ^ x[11];
  assign t[23] = (x[0] & x[1]);
  assign t[24] = (x[3] & x[4]);
  assign t[25] = (x[6] & x[7]);
  assign t[26] = (x[9] & x[10]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] & t[9];
  assign t[4] = t[19] ^ t[7];
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[20] ^ t[19];
  assign t[7] = ~(t[21]);
  assign t[8] = ~(t[19]);
  assign t[9] = t[6] ^ t[22];
  assign y = t[0] ^ t[1];
endmodule

module R1ind206(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind207(x, y);
 input [11:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[23] ^ t[21];
  assign t[11] = ~(t[21]);
  assign t[12] = t[10] ^ t[24];
  assign t[13] = ~(t[6] ^ t[15]);
  assign t[14] = t[16] ^ t[12];
  assign t[15] = t[17] ^ t[5];
  assign t[16] = t[21] ^ t[8];
  assign t[17] = t[18] & t[19];
  assign t[18] = ~(t[20]);
  assign t[19] = ~(t[10]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[12] ^ t[21];
  assign t[21] = t[25] ^ x[2];
  assign t[22] = t[26] ^ x[5];
  assign t[23] = t[27] ^ x[8];
  assign t[24] = t[28] ^ x[11];
  assign t[25] = (x[0] & x[1]);
  assign t[26] = (x[3] & x[4]);
  assign t[27] = (x[6] & x[7]);
  assign t[28] = (x[9] & x[10]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[10] ^ t[8];
  assign t[5] = t[11] & t[12];
  assign t[6] = t[10] ^ t[21];
  assign t[7] = t[13] & t[14];
  assign t[8] = ~(t[22]);
  assign t[9] = t[15] ^ t[7];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind208(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind209(x, y);
 input [11:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[14] ^ t[28];
  assign t[11] = t[19] & t[20];
  assign t[12] = ~(t[29]);
  assign t[13] = t[17] ^ t[11];
  assign t[14] = t[30] ^ t[28];
  assign t[15] = ~(t[28]);
  assign t[16] = t[14] ^ t[31];
  assign t[17] = t[21] ^ t[7];
  assign t[18] = t[22] & t[23];
  assign t[19] = ~(t[10] ^ t[17]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[8] ^ t[16];
  assign t[21] = t[24] & t[25];
  assign t[22] = ~(t[21] ^ t[26]);
  assign t[23] = t[6] ^ t[27];
  assign t[24] = ~(t[27]);
  assign t[25] = ~(t[14]);
  assign t[26] = t[8] ^ t[14];
  assign t[27] = t[16] ^ t[28];
  assign t[28] = t[32] ^ x[2];
  assign t[29] = t[33] ^ x[5];
  assign t[2] = t[6] ^ t[7];
  assign t[30] = t[34] ^ x[8];
  assign t[31] = t[35] ^ x[11];
  assign t[32] = (x[0] & x[1]);
  assign t[33] = (x[3] & x[4]);
  assign t[34] = (x[6] & x[7]);
  assign t[35] = (x[9] & x[10]);
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[10] ^ t[11];
  assign t[5] = t[12] ^ t[13];
  assign t[6] = t[14] ^ t[12];
  assign t[7] = t[15] & t[16];
  assign t[8] = t[28] ^ t[12];
  assign t[9] = t[17] ^ t[18];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind210(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind211(x, y);
 input [11:0] x;
 output y;

 wire [33:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[16] ^ t[7];
  assign t[11] = t[17] & t[18];
  assign t[12] = t[28] ^ t[27];
  assign t[13] = ~(t[27]);
  assign t[14] = t[12] ^ t[29];
  assign t[15] = t[19] & t[20];
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[23] ^ t[10]);
  assign t[18] = t[8] ^ t[14];
  assign t[19] = ~(t[16] ^ t[24]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[6] ^ t[25];
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[12]);
  assign t[23] = t[12] ^ t[27];
  assign t[24] = t[8] ^ t[12];
  assign t[25] = t[14] ^ t[27];
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[6] ^ t[7];
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[3] & x[4]);
  assign t[32] = (x[6] & x[7]);
  assign t[33] = (x[9] & x[10]);
  assign t[3] = t[8] ^ t[9];
  assign t[4] = ~(t[26]);
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[12] ^ t[4];
  assign t[7] = t[13] & t[14];
  assign t[8] = t[27] ^ t[4];
  assign t[9] = t[10] ^ t[15];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind212(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind213(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[12] ^ t[3];
  assign t[11] = t[13] & t[14];
  assign t[12] = t[15] & t[16];
  assign t[13] = ~(t[12] ^ t[17]);
  assign t[14] = t[2] ^ t[18];
  assign t[15] = ~(t[18]);
  assign t[16] = ~(t[6]);
  assign t[17] = t[4] ^ t[6];
  assign t[18] = t[9] ^ t[19];
  assign t[19] = t[23] ^ x[2];
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[24] ^ x[5];
  assign t[21] = t[25] ^ x[8];
  assign t[22] = t[26] ^ x[11];
  assign t[23] = (x[0] & x[1]);
  assign t[24] = (x[3] & x[4]);
  assign t[25] = (x[6] & x[7]);
  assign t[26] = (x[9] & x[10]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] & t[9];
  assign t[4] = t[19] ^ t[7];
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[20] ^ t[19];
  assign t[7] = ~(t[21]);
  assign t[8] = ~(t[19]);
  assign t[9] = t[6] ^ t[22];
  assign y = t[0] ^ t[1];
endmodule

module R1ind214(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind215(x, y);
 input [11:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[23] ^ t[21];
  assign t[11] = ~(t[21]);
  assign t[12] = t[10] ^ t[24];
  assign t[13] = ~(t[6] ^ t[15]);
  assign t[14] = t[16] ^ t[12];
  assign t[15] = t[17] ^ t[5];
  assign t[16] = t[21] ^ t[8];
  assign t[17] = t[18] & t[19];
  assign t[18] = ~(t[20]);
  assign t[19] = ~(t[10]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[12] ^ t[21];
  assign t[21] = t[25] ^ x[2];
  assign t[22] = t[26] ^ x[5];
  assign t[23] = t[27] ^ x[8];
  assign t[24] = t[28] ^ x[11];
  assign t[25] = (x[0] & x[1]);
  assign t[26] = (x[3] & x[4]);
  assign t[27] = (x[6] & x[7]);
  assign t[28] = (x[9] & x[10]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[10] ^ t[8];
  assign t[5] = t[11] & t[12];
  assign t[6] = t[10] ^ t[21];
  assign t[7] = t[13] & t[14];
  assign t[8] = ~(t[22]);
  assign t[9] = t[15] ^ t[7];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind216(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind217(x, y);
 input [11:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[14] ^ t[28];
  assign t[11] = t[19] & t[20];
  assign t[12] = ~(t[29]);
  assign t[13] = t[17] ^ t[11];
  assign t[14] = t[30] ^ t[28];
  assign t[15] = ~(t[28]);
  assign t[16] = t[14] ^ t[31];
  assign t[17] = t[21] ^ t[7];
  assign t[18] = t[22] & t[23];
  assign t[19] = ~(t[10] ^ t[17]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[8] ^ t[16];
  assign t[21] = t[24] & t[25];
  assign t[22] = ~(t[21] ^ t[26]);
  assign t[23] = t[6] ^ t[27];
  assign t[24] = ~(t[27]);
  assign t[25] = ~(t[14]);
  assign t[26] = t[8] ^ t[14];
  assign t[27] = t[16] ^ t[28];
  assign t[28] = t[32] ^ x[2];
  assign t[29] = t[33] ^ x[5];
  assign t[2] = t[6] ^ t[7];
  assign t[30] = t[34] ^ x[8];
  assign t[31] = t[35] ^ x[11];
  assign t[32] = (x[0] & x[1]);
  assign t[33] = (x[3] & x[4]);
  assign t[34] = (x[6] & x[7]);
  assign t[35] = (x[9] & x[10]);
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[10] ^ t[11];
  assign t[5] = t[12] ^ t[13];
  assign t[6] = t[14] ^ t[12];
  assign t[7] = t[15] & t[16];
  assign t[8] = t[28] ^ t[12];
  assign t[9] = t[17] ^ t[18];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind218(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind219(x, y);
 input [11:0] x;
 output y;

 wire [33:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[16] ^ t[7];
  assign t[11] = t[17] & t[18];
  assign t[12] = t[28] ^ t[27];
  assign t[13] = ~(t[27]);
  assign t[14] = t[12] ^ t[29];
  assign t[15] = t[19] & t[20];
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[23] ^ t[10]);
  assign t[18] = t[8] ^ t[14];
  assign t[19] = ~(t[16] ^ t[24]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[6] ^ t[25];
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[12]);
  assign t[23] = t[12] ^ t[27];
  assign t[24] = t[8] ^ t[12];
  assign t[25] = t[14] ^ t[27];
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[6] ^ t[7];
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[3] & x[4]);
  assign t[32] = (x[6] & x[7]);
  assign t[33] = (x[9] & x[10]);
  assign t[3] = t[8] ^ t[9];
  assign t[4] = ~(t[26]);
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[12] ^ t[4];
  assign t[7] = t[13] & t[14];
  assign t[8] = t[27] ^ t[4];
  assign t[9] = t[10] ^ t[15];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind220(x, y);
 input [8:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[2] ? x[4] : x[3];
  assign t[1] = ~(~x[5] & ~t[3]);
  assign t[2] = t[4] ^ x[2];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (x[0] & x[1]);
  assign t[5] = (x[6] & x[7]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind221(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[12] ^ t[3];
  assign t[11] = t[13] & t[14];
  assign t[12] = t[15] & t[16];
  assign t[13] = ~(t[12] ^ t[17]);
  assign t[14] = t[2] ^ t[18];
  assign t[15] = ~(t[18]);
  assign t[16] = ~(t[6]);
  assign t[17] = t[4] ^ t[6];
  assign t[18] = t[9] ^ t[19];
  assign t[19] = t[23] ^ x[2];
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[24] ^ x[5];
  assign t[21] = t[25] ^ x[8];
  assign t[22] = t[26] ^ x[11];
  assign t[23] = (x[0] & x[1]);
  assign t[24] = (x[3] & x[4]);
  assign t[25] = (x[6] & x[7]);
  assign t[26] = (x[9] & x[10]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] & t[9];
  assign t[4] = t[19] ^ t[7];
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[20] ^ t[19];
  assign t[7] = ~(t[21]);
  assign t[8] = ~(t[19]);
  assign t[9] = t[6] ^ t[22];
  assign y = t[0] ^ t[1];
endmodule

module R1ind222(x, y);
 input [8:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[4] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[3]);
  assign t[3] = ~x[5] & t[5];
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[8];
  assign t[6] = (x[0] & x[1]);
  assign t[7] = (x[6] & x[7]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind223(x, y);
 input [11:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[23] ^ t[21];
  assign t[11] = ~(t[21]);
  assign t[12] = t[10] ^ t[24];
  assign t[13] = ~(t[6] ^ t[15]);
  assign t[14] = t[16] ^ t[12];
  assign t[15] = t[17] ^ t[5];
  assign t[16] = t[21] ^ t[8];
  assign t[17] = t[18] & t[19];
  assign t[18] = ~(t[20]);
  assign t[19] = ~(t[10]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[12] ^ t[21];
  assign t[21] = t[25] ^ x[2];
  assign t[22] = t[26] ^ x[5];
  assign t[23] = t[27] ^ x[8];
  assign t[24] = t[28] ^ x[11];
  assign t[25] = (x[0] & x[1]);
  assign t[26] = (x[3] & x[4]);
  assign t[27] = (x[6] & x[7]);
  assign t[28] = (x[9] & x[10]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[10] ^ t[8];
  assign t[5] = t[11] & t[12];
  assign t[6] = t[10] ^ t[21];
  assign t[7] = t[13] & t[14];
  assign t[8] = ~(t[22]);
  assign t[9] = t[15] ^ t[7];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind224(x, y);
 input [8:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[2] ? x[4] : x[3];
  assign t[1] = ~x[5] & t[3];
  assign t[2] = t[4] ^ x[2];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (x[0] & x[1]);
  assign t[5] = (x[6] & x[7]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind225(x, y);
 input [11:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[14] ^ t[28];
  assign t[11] = t[19] & t[20];
  assign t[12] = ~(t[29]);
  assign t[13] = t[17] ^ t[11];
  assign t[14] = t[30] ^ t[28];
  assign t[15] = ~(t[28]);
  assign t[16] = t[14] ^ t[31];
  assign t[17] = t[21] ^ t[7];
  assign t[18] = t[22] & t[23];
  assign t[19] = ~(t[10] ^ t[17]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[8] ^ t[16];
  assign t[21] = t[24] & t[25];
  assign t[22] = ~(t[21] ^ t[26]);
  assign t[23] = t[6] ^ t[27];
  assign t[24] = ~(t[27]);
  assign t[25] = ~(t[14]);
  assign t[26] = t[8] ^ t[14];
  assign t[27] = t[16] ^ t[28];
  assign t[28] = t[32] ^ x[2];
  assign t[29] = t[33] ^ x[5];
  assign t[2] = t[6] ^ t[7];
  assign t[30] = t[34] ^ x[8];
  assign t[31] = t[35] ^ x[11];
  assign t[32] = (x[0] & x[1]);
  assign t[33] = (x[3] & x[4]);
  assign t[34] = (x[6] & x[7]);
  assign t[35] = (x[9] & x[10]);
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[10] ^ t[11];
  assign t[5] = t[12] ^ t[13];
  assign t[6] = t[14] ^ t[12];
  assign t[7] = t[15] & t[16];
  assign t[8] = t[28] ^ t[12];
  assign t[9] = t[17] ^ t[18];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind226(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = ~t[0];
endmodule

module R1ind227(x, y);
 input [11:0] x;
 output y;

 wire [33:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[16] ^ t[7];
  assign t[11] = t[17] & t[18];
  assign t[12] = t[28] ^ t[27];
  assign t[13] = ~(t[27]);
  assign t[14] = t[12] ^ t[29];
  assign t[15] = t[19] & t[20];
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[23] ^ t[10]);
  assign t[18] = t[8] ^ t[14];
  assign t[19] = ~(t[16] ^ t[24]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[6] ^ t[25];
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[12]);
  assign t[23] = t[12] ^ t[27];
  assign t[24] = t[8] ^ t[12];
  assign t[25] = t[14] ^ t[27];
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[6] ^ t[7];
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[3] & x[4]);
  assign t[32] = (x[6] & x[7]);
  assign t[33] = (x[9] & x[10]);
  assign t[3] = t[8] ^ t[9];
  assign t[4] = ~(t[26]);
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[12] ^ t[4];
  assign t[7] = t[13] & t[14];
  assign t[8] = t[27] ^ t[4];
  assign t[9] = t[10] ^ t[15];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind228(x, y);
 input [8:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[2] ? x[4] : x[3];
  assign t[1] = ~(~x[5] & ~t[3]);
  assign t[2] = t[4] ^ x[2];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (x[0] & x[1]);
  assign t[5] = (x[6] & x[7]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind229(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[12] ^ t[3];
  assign t[11] = t[13] & t[14];
  assign t[12] = t[15] & t[16];
  assign t[13] = ~(t[12] ^ t[17]);
  assign t[14] = t[2] ^ t[18];
  assign t[15] = ~(t[18]);
  assign t[16] = ~(t[6]);
  assign t[17] = t[4] ^ t[6];
  assign t[18] = t[9] ^ t[19];
  assign t[19] = t[23] ^ x[2];
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[24] ^ x[5];
  assign t[21] = t[25] ^ x[8];
  assign t[22] = t[26] ^ x[11];
  assign t[23] = (x[0] & x[1]);
  assign t[24] = (x[3] & x[4]);
  assign t[25] = (x[6] & x[7]);
  assign t[26] = (x[9] & x[10]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] & t[9];
  assign t[4] = t[19] ^ t[7];
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[20] ^ t[19];
  assign t[7] = ~(t[21]);
  assign t[8] = ~(t[19]);
  assign t[9] = t[6] ^ t[22];
  assign y = t[0] ^ t[1];
endmodule

module R1ind230(x, y);
 input [8:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[2] ? x[4] : x[3];
  assign t[1] = ~x[5] & t[3];
  assign t[2] = t[4] ^ x[2];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (x[0] & x[1]);
  assign t[5] = (x[6] & x[7]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind231(x, y);
 input [11:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[23] ^ t[21];
  assign t[11] = ~(t[21]);
  assign t[12] = t[10] ^ t[24];
  assign t[13] = ~(t[6] ^ t[15]);
  assign t[14] = t[16] ^ t[12];
  assign t[15] = t[17] ^ t[5];
  assign t[16] = t[21] ^ t[8];
  assign t[17] = t[18] & t[19];
  assign t[18] = ~(t[20]);
  assign t[19] = ~(t[10]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[12] ^ t[21];
  assign t[21] = t[25] ^ x[2];
  assign t[22] = t[26] ^ x[5];
  assign t[23] = t[27] ^ x[8];
  assign t[24] = t[28] ^ x[11];
  assign t[25] = (x[0] & x[1]);
  assign t[26] = (x[3] & x[4]);
  assign t[27] = (x[6] & x[7]);
  assign t[28] = (x[9] & x[10]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[10] ^ t[8];
  assign t[5] = t[11] & t[12];
  assign t[6] = t[10] ^ t[21];
  assign t[7] = t[13] & t[14];
  assign t[8] = ~(t[22]);
  assign t[9] = t[15] ^ t[7];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind232(x, y);
 input [8:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[2] ? x[4] : x[3];
  assign t[1] = ~x[5] & t[3];
  assign t[2] = t[4] ^ x[2];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (x[0] & x[1]);
  assign t[5] = (x[6] & x[7]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind233(x, y);
 input [11:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[14] ^ t[28];
  assign t[11] = t[19] & t[20];
  assign t[12] = ~(t[29]);
  assign t[13] = t[17] ^ t[11];
  assign t[14] = t[30] ^ t[28];
  assign t[15] = ~(t[28]);
  assign t[16] = t[14] ^ t[31];
  assign t[17] = t[21] ^ t[7];
  assign t[18] = t[22] & t[23];
  assign t[19] = ~(t[10] ^ t[17]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[8] ^ t[16];
  assign t[21] = t[24] & t[25];
  assign t[22] = ~(t[21] ^ t[26]);
  assign t[23] = t[6] ^ t[27];
  assign t[24] = ~(t[27]);
  assign t[25] = ~(t[14]);
  assign t[26] = t[8] ^ t[14];
  assign t[27] = t[16] ^ t[28];
  assign t[28] = t[32] ^ x[2];
  assign t[29] = t[33] ^ x[5];
  assign t[2] = t[6] ^ t[7];
  assign t[30] = t[34] ^ x[8];
  assign t[31] = t[35] ^ x[11];
  assign t[32] = (x[0] & x[1]);
  assign t[33] = (x[3] & x[4]);
  assign t[34] = (x[6] & x[7]);
  assign t[35] = (x[9] & x[10]);
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[10] ^ t[11];
  assign t[5] = t[12] ^ t[13];
  assign t[6] = t[14] ^ t[12];
  assign t[7] = t[15] & t[16];
  assign t[8] = t[28] ^ t[12];
  assign t[9] = t[17] ^ t[18];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind234(x, y);
 input [8:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[2] ? x[4] : x[3];
  assign t[1] = ~x[5] & t[3];
  assign t[2] = t[4] ^ x[2];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (x[0] & x[1]);
  assign t[5] = (x[6] & x[7]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind235(x, y);
 input [11:0] x;
 output y;

 wire [33:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[16] ^ t[7];
  assign t[11] = t[17] & t[18];
  assign t[12] = t[28] ^ t[27];
  assign t[13] = ~(t[27]);
  assign t[14] = t[12] ^ t[29];
  assign t[15] = t[19] & t[20];
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[23] ^ t[10]);
  assign t[18] = t[8] ^ t[14];
  assign t[19] = ~(t[16] ^ t[24]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[6] ^ t[25];
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[12]);
  assign t[23] = t[12] ^ t[27];
  assign t[24] = t[8] ^ t[12];
  assign t[25] = t[14] ^ t[27];
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[6] ^ t[7];
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[3] & x[4]);
  assign t[32] = (x[6] & x[7]);
  assign t[33] = (x[9] & x[10]);
  assign t[3] = t[8] ^ t[9];
  assign t[4] = ~(t[26]);
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[12] ^ t[4];
  assign t[7] = t[13] & t[14];
  assign t[8] = t[27] ^ t[4];
  assign t[9] = t[10] ^ t[15];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind236(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind237(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[12] ^ t[3];
  assign t[11] = t[13] & t[14];
  assign t[12] = t[15] & t[16];
  assign t[13] = ~(t[12] ^ t[17]);
  assign t[14] = t[2] ^ t[18];
  assign t[15] = ~(t[18]);
  assign t[16] = ~(t[6]);
  assign t[17] = t[4] ^ t[6];
  assign t[18] = t[9] ^ t[19];
  assign t[19] = t[23] ^ x[2];
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[24] ^ x[5];
  assign t[21] = t[25] ^ x[8];
  assign t[22] = t[26] ^ x[11];
  assign t[23] = (x[0] & x[1]);
  assign t[24] = (x[3] & x[4]);
  assign t[25] = (x[6] & x[7]);
  assign t[26] = (x[9] & x[10]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] & t[9];
  assign t[4] = t[19] ^ t[7];
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[20] ^ t[19];
  assign t[7] = ~(t[21]);
  assign t[8] = ~(t[19]);
  assign t[9] = t[6] ^ t[22];
  assign y = t[0] ^ t[1];
endmodule

module R1ind238(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind239(x, y);
 input [11:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[23] ^ t[21];
  assign t[11] = ~(t[21]);
  assign t[12] = t[10] ^ t[24];
  assign t[13] = ~(t[6] ^ t[15]);
  assign t[14] = t[16] ^ t[12];
  assign t[15] = t[17] ^ t[5];
  assign t[16] = t[21] ^ t[8];
  assign t[17] = t[18] & t[19];
  assign t[18] = ~(t[20]);
  assign t[19] = ~(t[10]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[12] ^ t[21];
  assign t[21] = t[25] ^ x[2];
  assign t[22] = t[26] ^ x[5];
  assign t[23] = t[27] ^ x[8];
  assign t[24] = t[28] ^ x[11];
  assign t[25] = (x[0] & x[1]);
  assign t[26] = (x[3] & x[4]);
  assign t[27] = (x[6] & x[7]);
  assign t[28] = (x[9] & x[10]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[10] ^ t[8];
  assign t[5] = t[11] & t[12];
  assign t[6] = t[10] ^ t[21];
  assign t[7] = t[13] & t[14];
  assign t[8] = ~(t[22]);
  assign t[9] = t[15] ^ t[7];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind240(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind241(x, y);
 input [11:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[14] ^ t[28];
  assign t[11] = t[19] & t[20];
  assign t[12] = ~(t[29]);
  assign t[13] = t[17] ^ t[11];
  assign t[14] = t[30] ^ t[28];
  assign t[15] = ~(t[28]);
  assign t[16] = t[14] ^ t[31];
  assign t[17] = t[21] ^ t[7];
  assign t[18] = t[22] & t[23];
  assign t[19] = ~(t[10] ^ t[17]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[8] ^ t[16];
  assign t[21] = t[24] & t[25];
  assign t[22] = ~(t[21] ^ t[26]);
  assign t[23] = t[6] ^ t[27];
  assign t[24] = ~(t[27]);
  assign t[25] = ~(t[14]);
  assign t[26] = t[8] ^ t[14];
  assign t[27] = t[16] ^ t[28];
  assign t[28] = t[32] ^ x[2];
  assign t[29] = t[33] ^ x[5];
  assign t[2] = t[6] ^ t[7];
  assign t[30] = t[34] ^ x[8];
  assign t[31] = t[35] ^ x[11];
  assign t[32] = (x[0] & x[1]);
  assign t[33] = (x[3] & x[4]);
  assign t[34] = (x[6] & x[7]);
  assign t[35] = (x[9] & x[10]);
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[10] ^ t[11];
  assign t[5] = t[12] ^ t[13];
  assign t[6] = t[14] ^ t[12];
  assign t[7] = t[15] & t[16];
  assign t[8] = t[28] ^ t[12];
  assign t[9] = t[17] ^ t[18];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind242(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind243(x, y);
 input [11:0] x;
 output y;

 wire [33:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[16] ^ t[7];
  assign t[11] = t[17] & t[18];
  assign t[12] = t[28] ^ t[27];
  assign t[13] = ~(t[27]);
  assign t[14] = t[12] ^ t[29];
  assign t[15] = t[19] & t[20];
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[23] ^ t[10]);
  assign t[18] = t[8] ^ t[14];
  assign t[19] = ~(t[16] ^ t[24]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[6] ^ t[25];
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[12]);
  assign t[23] = t[12] ^ t[27];
  assign t[24] = t[8] ^ t[12];
  assign t[25] = t[14] ^ t[27];
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[6] ^ t[7];
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[3] & x[4]);
  assign t[32] = (x[6] & x[7]);
  assign t[33] = (x[9] & x[10]);
  assign t[3] = t[8] ^ t[9];
  assign t[4] = ~(t[26]);
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[12] ^ t[4];
  assign t[7] = t[13] & t[14];
  assign t[8] = t[27] ^ t[4];
  assign t[9] = t[10] ^ t[15];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind244(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind245(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[12] ^ t[3];
  assign t[11] = t[13] & t[14];
  assign t[12] = t[15] & t[16];
  assign t[13] = ~(t[12] ^ t[17]);
  assign t[14] = t[2] ^ t[18];
  assign t[15] = ~(t[18]);
  assign t[16] = ~(t[6]);
  assign t[17] = t[4] ^ t[6];
  assign t[18] = t[9] ^ t[19];
  assign t[19] = t[23] ^ x[2];
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[24] ^ x[5];
  assign t[21] = t[25] ^ x[8];
  assign t[22] = t[26] ^ x[11];
  assign t[23] = (x[0] & x[1]);
  assign t[24] = (x[3] & x[4]);
  assign t[25] = (x[6] & x[7]);
  assign t[26] = (x[9] & x[10]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] & t[9];
  assign t[4] = t[19] ^ t[7];
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[20] ^ t[19];
  assign t[7] = ~(t[21]);
  assign t[8] = ~(t[19]);
  assign t[9] = t[6] ^ t[22];
  assign y = t[0] ^ t[1];
endmodule

module R1ind246(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind247(x, y);
 input [11:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[23] ^ t[21];
  assign t[11] = ~(t[21]);
  assign t[12] = t[10] ^ t[24];
  assign t[13] = ~(t[6] ^ t[15]);
  assign t[14] = t[16] ^ t[12];
  assign t[15] = t[17] ^ t[5];
  assign t[16] = t[21] ^ t[8];
  assign t[17] = t[18] & t[19];
  assign t[18] = ~(t[20]);
  assign t[19] = ~(t[10]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[12] ^ t[21];
  assign t[21] = t[25] ^ x[2];
  assign t[22] = t[26] ^ x[5];
  assign t[23] = t[27] ^ x[8];
  assign t[24] = t[28] ^ x[11];
  assign t[25] = (x[0] & x[1]);
  assign t[26] = (x[3] & x[4]);
  assign t[27] = (x[6] & x[7]);
  assign t[28] = (x[9] & x[10]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[10] ^ t[8];
  assign t[5] = t[11] & t[12];
  assign t[6] = t[10] ^ t[21];
  assign t[7] = t[13] & t[14];
  assign t[8] = ~(t[22]);
  assign t[9] = t[15] ^ t[7];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind248(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind249(x, y);
 input [11:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[14] ^ t[28];
  assign t[11] = t[19] & t[20];
  assign t[12] = ~(t[29]);
  assign t[13] = t[17] ^ t[11];
  assign t[14] = t[30] ^ t[28];
  assign t[15] = ~(t[28]);
  assign t[16] = t[14] ^ t[31];
  assign t[17] = t[21] ^ t[7];
  assign t[18] = t[22] & t[23];
  assign t[19] = ~(t[10] ^ t[17]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[8] ^ t[16];
  assign t[21] = t[24] & t[25];
  assign t[22] = ~(t[21] ^ t[26]);
  assign t[23] = t[6] ^ t[27];
  assign t[24] = ~(t[27]);
  assign t[25] = ~(t[14]);
  assign t[26] = t[8] ^ t[14];
  assign t[27] = t[16] ^ t[28];
  assign t[28] = t[32] ^ x[2];
  assign t[29] = t[33] ^ x[5];
  assign t[2] = t[6] ^ t[7];
  assign t[30] = t[34] ^ x[8];
  assign t[31] = t[35] ^ x[11];
  assign t[32] = (x[0] & x[1]);
  assign t[33] = (x[3] & x[4]);
  assign t[34] = (x[6] & x[7]);
  assign t[35] = (x[9] & x[10]);
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[10] ^ t[11];
  assign t[5] = t[12] ^ t[13];
  assign t[6] = t[14] ^ t[12];
  assign t[7] = t[15] & t[16];
  assign t[8] = t[28] ^ t[12];
  assign t[9] = t[17] ^ t[18];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind250(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind251(x, y);
 input [11:0] x;
 output y;

 wire [33:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[16] ^ t[7];
  assign t[11] = t[17] & t[18];
  assign t[12] = t[28] ^ t[27];
  assign t[13] = ~(t[27]);
  assign t[14] = t[12] ^ t[29];
  assign t[15] = t[19] & t[20];
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[23] ^ t[10]);
  assign t[18] = t[8] ^ t[14];
  assign t[19] = ~(t[16] ^ t[24]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[6] ^ t[25];
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[12]);
  assign t[23] = t[12] ^ t[27];
  assign t[24] = t[8] ^ t[12];
  assign t[25] = t[14] ^ t[27];
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[6] ^ t[7];
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[3] & x[4]);
  assign t[32] = (x[6] & x[7]);
  assign t[33] = (x[9] & x[10]);
  assign t[3] = t[8] ^ t[9];
  assign t[4] = ~(t[26]);
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[12] ^ t[4];
  assign t[7] = t[13] & t[14];
  assign t[8] = t[27] ^ t[4];
  assign t[9] = t[10] ^ t[15];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind252(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind253(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[12] ^ t[3];
  assign t[11] = t[13] & t[14];
  assign t[12] = t[15] & t[16];
  assign t[13] = ~(t[12] ^ t[17]);
  assign t[14] = t[2] ^ t[18];
  assign t[15] = ~(t[18]);
  assign t[16] = ~(t[6]);
  assign t[17] = t[4] ^ t[6];
  assign t[18] = t[9] ^ t[19];
  assign t[19] = t[23] ^ x[2];
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[24] ^ x[5];
  assign t[21] = t[25] ^ x[8];
  assign t[22] = t[26] ^ x[11];
  assign t[23] = (x[0] & x[1]);
  assign t[24] = (x[3] & x[4]);
  assign t[25] = (x[6] & x[7]);
  assign t[26] = (x[9] & x[10]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] & t[9];
  assign t[4] = t[19] ^ t[7];
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[20] ^ t[19];
  assign t[7] = ~(t[21]);
  assign t[8] = ~(t[19]);
  assign t[9] = t[6] ^ t[22];
  assign y = t[0] ^ t[1];
endmodule

module R1ind254(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind255(x, y);
 input [11:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[23] ^ t[21];
  assign t[11] = ~(t[21]);
  assign t[12] = t[10] ^ t[24];
  assign t[13] = ~(t[6] ^ t[15]);
  assign t[14] = t[16] ^ t[12];
  assign t[15] = t[17] ^ t[5];
  assign t[16] = t[21] ^ t[8];
  assign t[17] = t[18] & t[19];
  assign t[18] = ~(t[20]);
  assign t[19] = ~(t[10]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[12] ^ t[21];
  assign t[21] = t[25] ^ x[2];
  assign t[22] = t[26] ^ x[5];
  assign t[23] = t[27] ^ x[8];
  assign t[24] = t[28] ^ x[11];
  assign t[25] = (x[0] & x[1]);
  assign t[26] = (x[3] & x[4]);
  assign t[27] = (x[6] & x[7]);
  assign t[28] = (x[9] & x[10]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[10] ^ t[8];
  assign t[5] = t[11] & t[12];
  assign t[6] = t[10] ^ t[21];
  assign t[7] = t[13] & t[14];
  assign t[8] = ~(t[22]);
  assign t[9] = t[15] ^ t[7];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind256(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind257(x, y);
 input [11:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[14] ^ t[28];
  assign t[11] = t[19] & t[20];
  assign t[12] = ~(t[29]);
  assign t[13] = t[17] ^ t[11];
  assign t[14] = t[30] ^ t[28];
  assign t[15] = ~(t[28]);
  assign t[16] = t[14] ^ t[31];
  assign t[17] = t[21] ^ t[7];
  assign t[18] = t[22] & t[23];
  assign t[19] = ~(t[10] ^ t[17]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[8] ^ t[16];
  assign t[21] = t[24] & t[25];
  assign t[22] = ~(t[21] ^ t[26]);
  assign t[23] = t[6] ^ t[27];
  assign t[24] = ~(t[27]);
  assign t[25] = ~(t[14]);
  assign t[26] = t[8] ^ t[14];
  assign t[27] = t[16] ^ t[28];
  assign t[28] = t[32] ^ x[2];
  assign t[29] = t[33] ^ x[5];
  assign t[2] = t[6] ^ t[7];
  assign t[30] = t[34] ^ x[8];
  assign t[31] = t[35] ^ x[11];
  assign t[32] = (x[0] & x[1]);
  assign t[33] = (x[3] & x[4]);
  assign t[34] = (x[6] & x[7]);
  assign t[35] = (x[9] & x[10]);
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[10] ^ t[11];
  assign t[5] = t[12] ^ t[13];
  assign t[6] = t[14] ^ t[12];
  assign t[7] = t[15] & t[16];
  assign t[8] = t[28] ^ t[12];
  assign t[9] = t[17] ^ t[18];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind258(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind259(x, y);
 input [11:0] x;
 output y;

 wire [33:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[16] ^ t[7];
  assign t[11] = t[17] & t[18];
  assign t[12] = t[28] ^ t[27];
  assign t[13] = ~(t[27]);
  assign t[14] = t[12] ^ t[29];
  assign t[15] = t[19] & t[20];
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[23] ^ t[10]);
  assign t[18] = t[8] ^ t[14];
  assign t[19] = ~(t[16] ^ t[24]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[6] ^ t[25];
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[12]);
  assign t[23] = t[12] ^ t[27];
  assign t[24] = t[8] ^ t[12];
  assign t[25] = t[14] ^ t[27];
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[6] ^ t[7];
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[3] & x[4]);
  assign t[32] = (x[6] & x[7]);
  assign t[33] = (x[9] & x[10]);
  assign t[3] = t[8] ^ t[9];
  assign t[4] = ~(t[26]);
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[12] ^ t[4];
  assign t[7] = t[13] & t[14];
  assign t[8] = t[27] ^ t[4];
  assign t[9] = t[10] ^ t[15];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind260(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind261(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[12] ^ t[3];
  assign t[11] = t[13] & t[14];
  assign t[12] = t[15] & t[16];
  assign t[13] = ~(t[12] ^ t[17]);
  assign t[14] = t[2] ^ t[18];
  assign t[15] = ~(t[18]);
  assign t[16] = ~(t[6]);
  assign t[17] = t[4] ^ t[6];
  assign t[18] = t[9] ^ t[19];
  assign t[19] = t[23] ^ x[2];
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[24] ^ x[5];
  assign t[21] = t[25] ^ x[8];
  assign t[22] = t[26] ^ x[11];
  assign t[23] = (x[0] & x[1]);
  assign t[24] = (x[3] & x[4]);
  assign t[25] = (x[6] & x[7]);
  assign t[26] = (x[9] & x[10]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] & t[9];
  assign t[4] = t[19] ^ t[7];
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[20] ^ t[19];
  assign t[7] = ~(t[21]);
  assign t[8] = ~(t[19]);
  assign t[9] = t[6] ^ t[22];
  assign y = t[0] ^ t[1];
endmodule

module R1ind262(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind263(x, y);
 input [11:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[23] ^ t[21];
  assign t[11] = ~(t[21]);
  assign t[12] = t[10] ^ t[24];
  assign t[13] = ~(t[6] ^ t[15]);
  assign t[14] = t[16] ^ t[12];
  assign t[15] = t[17] ^ t[5];
  assign t[16] = t[21] ^ t[8];
  assign t[17] = t[18] & t[19];
  assign t[18] = ~(t[20]);
  assign t[19] = ~(t[10]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[12] ^ t[21];
  assign t[21] = t[25] ^ x[2];
  assign t[22] = t[26] ^ x[5];
  assign t[23] = t[27] ^ x[8];
  assign t[24] = t[28] ^ x[11];
  assign t[25] = (x[0] & x[1]);
  assign t[26] = (x[3] & x[4]);
  assign t[27] = (x[6] & x[7]);
  assign t[28] = (x[9] & x[10]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[10] ^ t[8];
  assign t[5] = t[11] & t[12];
  assign t[6] = t[10] ^ t[21];
  assign t[7] = t[13] & t[14];
  assign t[8] = ~(t[22]);
  assign t[9] = t[15] ^ t[7];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind264(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind265(x, y);
 input [11:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[14] ^ t[28];
  assign t[11] = t[19] & t[20];
  assign t[12] = ~(t[29]);
  assign t[13] = t[17] ^ t[11];
  assign t[14] = t[30] ^ t[28];
  assign t[15] = ~(t[28]);
  assign t[16] = t[14] ^ t[31];
  assign t[17] = t[21] ^ t[7];
  assign t[18] = t[22] & t[23];
  assign t[19] = ~(t[10] ^ t[17]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[8] ^ t[16];
  assign t[21] = t[24] & t[25];
  assign t[22] = ~(t[21] ^ t[26]);
  assign t[23] = t[6] ^ t[27];
  assign t[24] = ~(t[27]);
  assign t[25] = ~(t[14]);
  assign t[26] = t[8] ^ t[14];
  assign t[27] = t[16] ^ t[28];
  assign t[28] = t[32] ^ x[2];
  assign t[29] = t[33] ^ x[5];
  assign t[2] = t[6] ^ t[7];
  assign t[30] = t[34] ^ x[8];
  assign t[31] = t[35] ^ x[11];
  assign t[32] = (x[0] & x[1]);
  assign t[33] = (x[3] & x[4]);
  assign t[34] = (x[6] & x[7]);
  assign t[35] = (x[9] & x[10]);
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[10] ^ t[11];
  assign t[5] = t[12] ^ t[13];
  assign t[6] = t[14] ^ t[12];
  assign t[7] = t[15] & t[16];
  assign t[8] = t[28] ^ t[12];
  assign t[9] = t[17] ^ t[18];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind266(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0] ? x[4] : x[3];
endmodule

module R1ind267(x, y);
 input [11:0] x;
 output y;

 wire [33:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[16] ^ t[7];
  assign t[11] = t[17] & t[18];
  assign t[12] = t[28] ^ t[27];
  assign t[13] = ~(t[27]);
  assign t[14] = t[12] ^ t[29];
  assign t[15] = t[19] & t[20];
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[23] ^ t[10]);
  assign t[18] = t[8] ^ t[14];
  assign t[19] = ~(t[16] ^ t[24]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = t[6] ^ t[25];
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[12]);
  assign t[23] = t[12] ^ t[27];
  assign t[24] = t[8] ^ t[12];
  assign t[25] = t[14] ^ t[27];
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[6] ^ t[7];
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[3] & x[4]);
  assign t[32] = (x[6] & x[7]);
  assign t[33] = (x[9] & x[10]);
  assign t[3] = t[8] ^ t[9];
  assign t[4] = ~(t[26]);
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[12] ^ t[4];
  assign t[7] = t[13] & t[14];
  assign t[8] = t[27] ^ t[4];
  assign t[9] = t[10] ^ t[15];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1_ind(x, y);
 input [545:0] x;
 output [267:0] y;

  R1ind0 R1ind0_inst(.x({x[2], x[1], x[0]}), .y(y[0]));
  R1ind1 R1ind1_inst(.x({x[5], x[4], x[3]}), .y(y[1]));
  R1ind2 R1ind2_inst(.x({x[8], x[7], x[6]}), .y(y[2]));
  R1ind3 R1ind3_inst(.x({x[11], x[10], x[9]}), .y(y[3]));
  R1ind4 R1ind4_inst(.x({x[14], x[13], x[12]}), .y(y[4]));
  R1ind5 R1ind5_inst(.x({x[17], x[16], x[15]}), .y(y[5]));
  R1ind6 R1ind6_inst(.x({x[20], x[19], x[18]}), .y(y[6]));
  R1ind7 R1ind7_inst(.x({x[23], x[22], x[21]}), .y(y[7]));
  R1ind8 R1ind8_inst(.x({x[26], x[25], x[24]}), .y(y[8]));
  R1ind9 R1ind9_inst(.x({x[29], x[28], x[27]}), .y(y[9]));
  R1ind10 R1ind10_inst(.x({x[32], x[31], x[30]}), .y(y[10]));
  R1ind11 R1ind11_inst(.x({x[35], x[34], x[33]}), .y(y[11]));
  R1ind12 R1ind12_inst(.x({x[38], x[37], x[36]}), .y(y[12]));
  R1ind13 R1ind13_inst(.x({x[41], x[40], x[39]}), .y(y[13]));
  R1ind14 R1ind14_inst(.x({x[44], x[43], x[42]}), .y(y[14]));
  R1ind15 R1ind15_inst(.x({x[47], x[46], x[45]}), .y(y[15]));
  R1ind16 R1ind16_inst(.x({x[50], x[49], x[48]}), .y(y[16]));
  R1ind17 R1ind17_inst(.x({x[53], x[52], x[51]}), .y(y[17]));
  R1ind18 R1ind18_inst(.x({x[56], x[55], x[54]}), .y(y[18]));
  R1ind19 R1ind19_inst(.x({x[59], x[58], x[57]}), .y(y[19]));
  R1ind20 R1ind20_inst(.x({x[62], x[61], x[60]}), .y(y[20]));
  R1ind21 R1ind21_inst(.x({x[65], x[64], x[63]}), .y(y[21]));
  R1ind22 R1ind22_inst(.x({x[68], x[67], x[66]}), .y(y[22]));
  R1ind23 R1ind23_inst(.x({x[71], x[70], x[69]}), .y(y[23]));
  R1ind24 R1ind24_inst(.x({x[74], x[73], x[72]}), .y(y[24]));
  R1ind25 R1ind25_inst(.x({x[77], x[76], x[75]}), .y(y[25]));
  R1ind26 R1ind26_inst(.x({x[80], x[79], x[78]}), .y(y[26]));
  R1ind27 R1ind27_inst(.x({x[83], x[82], x[81]}), .y(y[27]));
  R1ind28 R1ind28_inst(.x({x[86], x[85], x[84]}), .y(y[28]));
  R1ind29 R1ind29_inst(.x({x[89], x[88], x[87]}), .y(y[29]));
  R1ind30 R1ind30_inst(.x({x[92], x[91], x[90]}), .y(y[30]));
  R1ind31 R1ind31_inst(.x({x[95], x[94], x[93]}), .y(y[31]));
  R1ind32 R1ind32_inst(.x({x[98], x[97], x[96]}), .y(y[32]));
  R1ind33 R1ind33_inst(.x({x[101], x[100], x[99]}), .y(y[33]));
  R1ind34 R1ind34_inst(.x({x[104], x[103], x[102]}), .y(y[34]));
  R1ind35 R1ind35_inst(.x({x[107], x[106], x[105]}), .y(y[35]));
  R1ind36 R1ind36_inst(.x({x[110], x[109], x[108]}), .y(y[36]));
  R1ind37 R1ind37_inst(.x({x[113], x[112], x[111]}), .y(y[37]));
  R1ind38 R1ind38_inst(.x({x[116], x[115], x[114]}), .y(y[38]));
  R1ind39 R1ind39_inst(.x({x[119], x[118], x[117]}), .y(y[39]));
  R1ind40 R1ind40_inst(.x({x[122], x[121], x[120]}), .y(y[40]));
  R1ind41 R1ind41_inst(.x({x[125], x[124], x[123]}), .y(y[41]));
  R1ind42 R1ind42_inst(.x({x[128], x[127], x[126]}), .y(y[42]));
  R1ind43 R1ind43_inst(.x({x[131], x[130], x[129]}), .y(y[43]));
  R1ind44 R1ind44_inst(.x({x[134], x[133], x[132]}), .y(y[44]));
  R1ind45 R1ind45_inst(.x({x[137], x[136], x[135]}), .y(y[45]));
  R1ind46 R1ind46_inst(.x({x[140], x[139], x[138]}), .y(y[46]));
  R1ind47 R1ind47_inst(.x({x[143], x[142], x[141]}), .y(y[47]));
  R1ind48 R1ind48_inst(.x({x[146], x[145], x[144]}), .y(y[48]));
  R1ind49 R1ind49_inst(.x({x[149], x[148], x[147]}), .y(y[49]));
  R1ind50 R1ind50_inst(.x({x[152], x[151], x[150]}), .y(y[50]));
  R1ind51 R1ind51_inst(.x({x[155], x[154], x[153]}), .y(y[51]));
  R1ind52 R1ind52_inst(.x({x[158], x[157], x[156]}), .y(y[52]));
  R1ind53 R1ind53_inst(.x({x[161], x[160], x[159]}), .y(y[53]));
  R1ind54 R1ind54_inst(.x({x[164], x[163], x[162]}), .y(y[54]));
  R1ind55 R1ind55_inst(.x({x[167], x[166], x[165]}), .y(y[55]));
  R1ind56 R1ind56_inst(.x({x[170], x[169], x[168]}), .y(y[56]));
  R1ind57 R1ind57_inst(.x({x[173], x[172], x[171]}), .y(y[57]));
  R1ind58 R1ind58_inst(.x({x[176], x[175], x[174]}), .y(y[58]));
  R1ind59 R1ind59_inst(.x({x[179], x[178], x[177]}), .y(y[59]));
  R1ind60 R1ind60_inst(.x({x[182], x[181], x[180]}), .y(y[60]));
  R1ind61 R1ind61_inst(.x({x[185], x[184], x[183]}), .y(y[61]));
  R1ind62 R1ind62_inst(.x({x[188], x[187], x[186]}), .y(y[62]));
  R1ind63 R1ind63_inst(.x({x[191], x[190], x[189]}), .y(y[63]));
  R1ind64 R1ind64_inst(.x({x[194], x[193], x[192]}), .y(y[64]));
  R1ind65 R1ind65_inst(.x({x[216], x[215], x[214], x[213], x[212], x[211], x[210], x[209], x[208], x[207], x[206], x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[197], x[196], x[195]}), .y(y[65]));
  R1ind66 R1ind66_inst(.x({x[219], x[218], x[217]}), .y(y[66]));
  R1ind67 R1ind67_inst(.x({x[222], x[221], x[220], x[195], x[219], x[218], x[217]}), .y(y[67]));
  R1ind68 R1ind68_inst(.x({x[207], x[206], x[205], x[195]}), .y(y[68]));
  R1ind69 R1ind69_inst(.x({x[204], x[203], x[202], x[195]}), .y(y[69]));
  R1ind70 R1ind70_inst(.x({x[201], x[200], x[199], x[207], x[206], x[205], x[195]}), .y(y[70]));
  R1ind71 R1ind71_inst(.x({x[213], x[212], x[211], x[195]}), .y(y[71]));
  R1ind72 R1ind72_inst(.x({x[216], x[215], x[214], x[195]}), .y(y[72]));
  R1ind73 R1ind73_inst(.x({x[198], x[197], x[196], x[195]}), .y(y[73]));
  R1ind74 R1ind74_inst(.x({x[213], x[212], x[211], x[210], x[209], x[208], x[195]}), .y(y[74]));
  R1ind75 R1ind75_inst(.x({x[225], x[224], x[195], x[223]}), .y(y[75]));
  R1ind76 R1ind76_inst(.x({x[228], x[227], x[195], x[226]}), .y(y[76]));
  R1ind77 R1ind77_inst(.x({x[231], x[230], x[195], x[229]}), .y(y[77]));
  R1ind78 R1ind78_inst(.x({x[234], x[233], x[195], x[232]}), .y(y[78]));
  R1ind79 R1ind79_inst(.x({x[237], x[236], x[195], x[235]}), .y(y[79]));
  R1ind80 R1ind80_inst(.x({x[240], x[239], x[195], x[238]}), .y(y[80]));
  R1ind81 R1ind81_inst(.x({x[243], x[242], x[195], x[241]}), .y(y[81]));
  R1ind82 R1ind82_inst(.x({x[246], x[245], x[195], x[244]}), .y(y[82]));
  R1ind83 R1ind83_inst(.x({x[249], x[248], x[195], x[247]}), .y(y[83]));
  R1ind84 R1ind84_inst(.x({x[252], x[251], x[195], x[250]}), .y(y[84]));
  R1ind85 R1ind85_inst(.x({x[255], x[254], x[195], x[253]}), .y(y[85]));
  R1ind86 R1ind86_inst(.x({x[258], x[257], x[195], x[256]}), .y(y[86]));
  R1ind87 R1ind87_inst(.x({x[261], x[260], x[195], x[259]}), .y(y[87]));
  R1ind88 R1ind88_inst(.x({x[264], x[263], x[195], x[262]}), .y(y[88]));
  R1ind89 R1ind89_inst(.x({x[267], x[266], x[195], x[265]}), .y(y[89]));
  R1ind90 R1ind90_inst(.x({x[270], x[269], x[195], x[268]}), .y(y[90]));
  R1ind91 R1ind91_inst(.x({x[273], x[272], x[195], x[271]}), .y(y[91]));
  R1ind92 R1ind92_inst(.x({x[276], x[275], x[195], x[274]}), .y(y[92]));
  R1ind93 R1ind93_inst(.x({x[279], x[278], x[195], x[277]}), .y(y[93]));
  R1ind94 R1ind94_inst(.x({x[282], x[281], x[195], x[280]}), .y(y[94]));
  R1ind95 R1ind95_inst(.x({x[285], x[284], x[195], x[283]}), .y(y[95]));
  R1ind96 R1ind96_inst(.x({x[288], x[287], x[195], x[286]}), .y(y[96]));
  R1ind97 R1ind97_inst(.x({x[291], x[290], x[195], x[289]}), .y(y[97]));
  R1ind98 R1ind98_inst(.x({x[294], x[293], x[195], x[292]}), .y(y[98]));
  R1ind99 R1ind99_inst(.x({x[297], x[296], x[195], x[295]}), .y(y[99]));
  R1ind100 R1ind100_inst(.x({x[300], x[299], x[195], x[298]}), .y(y[100]));
  R1ind101 R1ind101_inst(.x({x[303], x[302], x[195], x[301]}), .y(y[101]));
  R1ind102 R1ind102_inst(.x({x[306], x[305], x[195], x[304]}), .y(y[102]));
  R1ind103 R1ind103_inst(.x({x[309], x[308], x[195], x[307]}), .y(y[103]));
  R1ind104 R1ind104_inst(.x({x[312], x[311], x[195], x[310]}), .y(y[104]));
  R1ind105 R1ind105_inst(.x({x[315], x[314], x[195], x[313]}), .y(y[105]));
  R1ind106 R1ind106_inst(.x({x[318], x[317], x[195], x[316]}), .y(y[106]));
  R1ind107 R1ind107_inst(.x({x[321], x[320], x[225], x[224], x[195], x[319]}), .y(y[107]));
  R1ind108 R1ind108_inst(.x({x[324], x[323], x[228], x[227], x[195], x[322]}), .y(y[108]));
  R1ind109 R1ind109_inst(.x({x[327], x[326], x[231], x[230], x[195], x[325]}), .y(y[109]));
  R1ind110 R1ind110_inst(.x({x[330], x[329], x[234], x[233], x[195], x[328]}), .y(y[110]));
  R1ind111 R1ind111_inst(.x({x[333], x[332], x[237], x[236], x[195], x[331]}), .y(y[111]));
  R1ind112 R1ind112_inst(.x({x[336], x[335], x[240], x[239], x[195], x[334]}), .y(y[112]));
  R1ind113 R1ind113_inst(.x({x[339], x[338], x[243], x[242], x[195], x[337]}), .y(y[113]));
  R1ind114 R1ind114_inst(.x({x[342], x[341], x[246], x[245], x[195], x[340]}), .y(y[114]));
  R1ind115 R1ind115_inst(.x({x[345], x[344], x[249], x[248], x[195], x[343]}), .y(y[115]));
  R1ind116 R1ind116_inst(.x({x[348], x[347], x[252], x[251], x[195], x[346]}), .y(y[116]));
  R1ind117 R1ind117_inst(.x({x[351], x[350], x[255], x[254], x[195], x[349]}), .y(y[117]));
  R1ind118 R1ind118_inst(.x({x[354], x[353], x[258], x[257], x[195], x[352]}), .y(y[118]));
  R1ind119 R1ind119_inst(.x({x[357], x[356], x[261], x[260], x[195], x[355]}), .y(y[119]));
  R1ind120 R1ind120_inst(.x({x[360], x[359], x[264], x[263], x[195], x[358]}), .y(y[120]));
  R1ind121 R1ind121_inst(.x({x[363], x[362], x[267], x[266], x[195], x[361]}), .y(y[121]));
  R1ind122 R1ind122_inst(.x({x[366], x[365], x[270], x[269], x[195], x[364]}), .y(y[122]));
  R1ind123 R1ind123_inst(.x({x[225], x[224], x[273], x[272], x[369], x[368], x[195], x[367]}), .y(y[123]));
  R1ind124 R1ind124_inst(.x({x[228], x[227], x[276], x[275], x[372], x[371], x[195], x[370]}), .y(y[124]));
  R1ind125 R1ind125_inst(.x({x[231], x[230], x[279], x[278], x[375], x[374], x[195], x[373]}), .y(y[125]));
  R1ind126 R1ind126_inst(.x({x[234], x[233], x[282], x[281], x[378], x[377], x[195], x[376]}), .y(y[126]));
  R1ind127 R1ind127_inst(.x({x[237], x[236], x[285], x[284], x[381], x[380], x[195], x[379]}), .y(y[127]));
  R1ind128 R1ind128_inst(.x({x[240], x[239], x[288], x[287], x[384], x[383], x[195], x[382]}), .y(y[128]));
  R1ind129 R1ind129_inst(.x({x[243], x[242], x[291], x[290], x[387], x[386], x[195], x[385]}), .y(y[129]));
  R1ind130 R1ind130_inst(.x({x[246], x[245], x[294], x[293], x[390], x[389], x[195], x[388]}), .y(y[130]));
  R1ind131 R1ind131_inst(.x({x[249], x[248], x[297], x[296], x[393], x[392], x[195], x[391]}), .y(y[131]));
  R1ind132 R1ind132_inst(.x({x[252], x[251], x[300], x[299], x[396], x[395], x[195], x[394]}), .y(y[132]));
  R1ind133 R1ind133_inst(.x({x[255], x[254], x[303], x[302], x[399], x[398], x[195], x[397]}), .y(y[133]));
  R1ind134 R1ind134_inst(.x({x[258], x[257], x[306], x[305], x[402], x[401], x[195], x[400]}), .y(y[134]));
  R1ind135 R1ind135_inst(.x({x[261], x[260], x[309], x[308], x[405], x[404], x[195], x[403]}), .y(y[135]));
  R1ind136 R1ind136_inst(.x({x[264], x[263], x[312], x[311], x[408], x[407], x[195], x[406]}), .y(y[136]));
  R1ind137 R1ind137_inst(.x({x[267], x[266], x[315], x[314], x[411], x[410], x[195], x[409]}), .y(y[137]));
  R1ind138 R1ind138_inst(.x({x[270], x[269], x[318], x[317], x[414], x[413], x[195], x[412]}), .y(y[138]));
  R1ind139 R1ind139_inst(.x({x[417], x[416], x[415], x[195]}), .y(y[139]));
  R1ind140 R1ind140_inst(.x({x[419], x[418], x[219], x[218], x[217]}), .y(y[140]));
  R1ind141 R1ind141_inst(.x({x[191], x[190], x[189], x[188], x[187], x[186], x[185], x[184], x[183], x[194], x[193], x[192]}), .y(y[141]));
  R1ind142 R1ind142_inst(.x({x[421], x[420], x[219], x[218], x[217]}), .y(y[142]));
  R1ind143 R1ind143_inst(.x({x[191], x[190], x[189], x[185], x[184], x[183], x[188], x[187], x[186], x[194], x[193], x[192]}), .y(y[143]));
  R1ind144 R1ind144_inst(.x({x[423], x[422], x[219], x[218], x[217]}), .y(y[144]));
  R1ind145 R1ind145_inst(.x({x[191], x[190], x[189], x[185], x[184], x[183], x[188], x[187], x[186], x[194], x[193], x[192]}), .y(y[145]));
  R1ind146 R1ind146_inst(.x({x[425], x[424], x[219], x[218], x[217]}), .y(y[146]));
  R1ind147 R1ind147_inst(.x({x[191], x[190], x[189], x[185], x[184], x[183], x[194], x[193], x[192], x[188], x[187], x[186]}), .y(y[147]));
  R1ind148 R1ind148_inst(.x({x[427], x[426], x[219], x[218], x[217]}), .y(y[148]));
  R1ind149 R1ind149_inst(.x({x[155], x[154], x[153], x[152], x[151], x[150], x[149], x[148], x[147], x[158], x[157], x[156]}), .y(y[149]));
  R1ind150 R1ind150_inst(.x({x[429], x[428], x[219], x[218], x[217]}), .y(y[150]));
  R1ind151 R1ind151_inst(.x({x[155], x[154], x[153], x[149], x[148], x[147], x[152], x[151], x[150], x[158], x[157], x[156]}), .y(y[151]));
  R1ind152 R1ind152_inst(.x({x[431], x[430], x[219], x[218], x[217]}), .y(y[152]));
  R1ind153 R1ind153_inst(.x({x[155], x[154], x[153], x[149], x[148], x[147], x[152], x[151], x[150], x[158], x[157], x[156]}), .y(y[153]));
  R1ind154 R1ind154_inst(.x({x[433], x[432], x[219], x[218], x[217]}), .y(y[154]));
  R1ind155 R1ind155_inst(.x({x[155], x[154], x[153], x[149], x[148], x[147], x[158], x[157], x[156], x[152], x[151], x[150]}), .y(y[155]));
  R1ind156 R1ind156_inst(.x({x[435], x[434], x[219], x[218], x[217]}), .y(y[156]));
  R1ind157 R1ind157_inst(.x({x[167], x[166], x[165], x[164], x[163], x[162], x[161], x[160], x[159], x[170], x[169], x[168]}), .y(y[157]));
  R1ind158 R1ind158_inst(.x({x[437], x[436], x[219], x[218], x[217]}), .y(y[158]));
  R1ind159 R1ind159_inst(.x({x[167], x[166], x[165], x[161], x[160], x[159], x[164], x[163], x[162], x[170], x[169], x[168]}), .y(y[159]));
  R1ind160 R1ind160_inst(.x({x[439], x[438], x[219], x[218], x[217]}), .y(y[160]));
  R1ind161 R1ind161_inst(.x({x[167], x[166], x[165], x[161], x[160], x[159], x[164], x[163], x[162], x[170], x[169], x[168]}), .y(y[161]));
  R1ind162 R1ind162_inst(.x({x[441], x[440], x[219], x[218], x[217]}), .y(y[162]));
  R1ind163 R1ind163_inst(.x({x[167], x[166], x[165], x[161], x[160], x[159], x[170], x[169], x[168], x[164], x[163], x[162]}), .y(y[163]));
  R1ind164 R1ind164_inst(.x({x[443], x[442], x[219], x[218], x[217]}), .y(y[164]));
  R1ind165 R1ind165_inst(.x({x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[172], x[171], x[182], x[181], x[180]}), .y(y[165]));
  R1ind166 R1ind166_inst(.x({x[445], x[444], x[219], x[218], x[217]}), .y(y[166]));
  R1ind167 R1ind167_inst(.x({x[179], x[178], x[177], x[173], x[172], x[171], x[176], x[175], x[174], x[182], x[181], x[180]}), .y(y[167]));
  R1ind168 R1ind168_inst(.x({x[447], x[446], x[219], x[218], x[217]}), .y(y[168]));
  R1ind169 R1ind169_inst(.x({x[179], x[178], x[177], x[173], x[172], x[171], x[176], x[175], x[174], x[182], x[181], x[180]}), .y(y[169]));
  R1ind170 R1ind170_inst(.x({x[449], x[448], x[219], x[218], x[217]}), .y(y[170]));
  R1ind171 R1ind171_inst(.x({x[179], x[178], x[177], x[173], x[172], x[171], x[182], x[181], x[180], x[176], x[175], x[174]}), .y(y[171]));
  R1ind172 R1ind172_inst(.x({x[451], x[450], x[219], x[218], x[217]}), .y(y[172]));
  R1ind173 R1ind173_inst(.x({x[107], x[106], x[105], x[104], x[103], x[102], x[101], x[100], x[99], x[110], x[109], x[108]}), .y(y[173]));
  R1ind174 R1ind174_inst(.x({x[453], x[452], x[219], x[218], x[217]}), .y(y[174]));
  R1ind175 R1ind175_inst(.x({x[107], x[106], x[105], x[101], x[100], x[99], x[104], x[103], x[102], x[110], x[109], x[108]}), .y(y[175]));
  R1ind176 R1ind176_inst(.x({x[455], x[454], x[219], x[218], x[217]}), .y(y[176]));
  R1ind177 R1ind177_inst(.x({x[107], x[106], x[105], x[101], x[100], x[99], x[104], x[103], x[102], x[110], x[109], x[108]}), .y(y[177]));
  R1ind178 R1ind178_inst(.x({x[457], x[456], x[219], x[218], x[217]}), .y(y[178]));
  R1ind179 R1ind179_inst(.x({x[107], x[106], x[105], x[101], x[100], x[99], x[110], x[109], x[108], x[104], x[103], x[102]}), .y(y[179]));
  R1ind180 R1ind180_inst(.x({x[459], x[458], x[219], x[218], x[217]}), .y(y[180]));
  R1ind181 R1ind181_inst(.x({x[143], x[142], x[141], x[140], x[139], x[138], x[137], x[136], x[135], x[146], x[145], x[144]}), .y(y[181]));
  R1ind182 R1ind182_inst(.x({x[461], x[460], x[219], x[218], x[217]}), .y(y[182]));
  R1ind183 R1ind183_inst(.x({x[143], x[142], x[141], x[137], x[136], x[135], x[140], x[139], x[138], x[146], x[145], x[144]}), .y(y[183]));
  R1ind184 R1ind184_inst(.x({x[463], x[462], x[219], x[218], x[217]}), .y(y[184]));
  R1ind185 R1ind185_inst(.x({x[143], x[142], x[141], x[137], x[136], x[135], x[140], x[139], x[138], x[146], x[145], x[144]}), .y(y[185]));
  R1ind186 R1ind186_inst(.x({x[465], x[464], x[219], x[218], x[217]}), .y(y[186]));
  R1ind187 R1ind187_inst(.x({x[143], x[142], x[141], x[137], x[136], x[135], x[146], x[145], x[144], x[140], x[139], x[138]}), .y(y[187]));
  R1ind188 R1ind188_inst(.x({x[467], x[466], x[219], x[218], x[217]}), .y(y[188]));
  R1ind189 R1ind189_inst(.x({x[131], x[130], x[129], x[128], x[127], x[126], x[125], x[124], x[123], x[134], x[133], x[132]}), .y(y[189]));
  R1ind190 R1ind190_inst(.x({x[469], x[468], x[219], x[218], x[217]}), .y(y[190]));
  R1ind191 R1ind191_inst(.x({x[131], x[130], x[129], x[125], x[124], x[123], x[128], x[127], x[126], x[134], x[133], x[132]}), .y(y[191]));
  R1ind192 R1ind192_inst(.x({x[471], x[470], x[219], x[218], x[217]}), .y(y[192]));
  R1ind193 R1ind193_inst(.x({x[131], x[130], x[129], x[125], x[124], x[123], x[128], x[127], x[126], x[134], x[133], x[132]}), .y(y[193]));
  R1ind194 R1ind194_inst(.x({x[473], x[472], x[219], x[218], x[217]}), .y(y[194]));
  R1ind195 R1ind195_inst(.x({x[131], x[130], x[129], x[125], x[124], x[123], x[134], x[133], x[132], x[128], x[127], x[126]}), .y(y[195]));
  R1ind196 R1ind196_inst(.x({x[475], x[474], x[219], x[218], x[217]}), .y(y[196]));
  R1ind197 R1ind197_inst(.x({x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[112], x[111], x[122], x[121], x[120]}), .y(y[197]));
  R1ind198 R1ind198_inst(.x({x[477], x[476], x[219], x[218], x[217]}), .y(y[198]));
  R1ind199 R1ind199_inst(.x({x[119], x[118], x[117], x[113], x[112], x[111], x[116], x[115], x[114], x[122], x[121], x[120]}), .y(y[199]));
  R1ind200 R1ind200_inst(.x({x[479], x[478], x[219], x[218], x[217]}), .y(y[200]));
  R1ind201 R1ind201_inst(.x({x[119], x[118], x[117], x[113], x[112], x[111], x[116], x[115], x[114], x[122], x[121], x[120]}), .y(y[201]));
  R1ind202 R1ind202_inst(.x({x[481], x[480], x[219], x[218], x[217]}), .y(y[202]));
  R1ind203 R1ind203_inst(.x({x[119], x[118], x[117], x[113], x[112], x[111], x[122], x[121], x[120], x[116], x[115], x[114]}), .y(y[203]));
  R1ind204 R1ind204_inst(.x({x[483], x[482], x[219], x[218], x[217]}), .y(y[204]));
  R1ind205 R1ind205_inst(.x({x[59], x[58], x[57], x[56], x[55], x[54], x[53], x[52], x[51], x[62], x[61], x[60]}), .y(y[205]));
  R1ind206 R1ind206_inst(.x({x[485], x[484], x[219], x[218], x[217]}), .y(y[206]));
  R1ind207 R1ind207_inst(.x({x[59], x[58], x[57], x[53], x[52], x[51], x[56], x[55], x[54], x[62], x[61], x[60]}), .y(y[207]));
  R1ind208 R1ind208_inst(.x({x[487], x[486], x[219], x[218], x[217]}), .y(y[208]));
  R1ind209 R1ind209_inst(.x({x[59], x[58], x[57], x[53], x[52], x[51], x[56], x[55], x[54], x[62], x[61], x[60]}), .y(y[209]));
  R1ind210 R1ind210_inst(.x({x[489], x[488], x[219], x[218], x[217]}), .y(y[210]));
  R1ind211 R1ind211_inst(.x({x[59], x[58], x[57], x[53], x[52], x[51], x[62], x[61], x[60], x[56], x[55], x[54]}), .y(y[211]));
  R1ind212 R1ind212_inst(.x({x[491], x[490], x[219], x[218], x[217]}), .y(y[212]));
  R1ind213 R1ind213_inst(.x({x[95], x[94], x[93], x[92], x[91], x[90], x[89], x[88], x[87], x[98], x[97], x[96]}), .y(y[213]));
  R1ind214 R1ind214_inst(.x({x[493], x[492], x[219], x[218], x[217]}), .y(y[214]));
  R1ind215 R1ind215_inst(.x({x[95], x[94], x[93], x[89], x[88], x[87], x[92], x[91], x[90], x[98], x[97], x[96]}), .y(y[215]));
  R1ind216 R1ind216_inst(.x({x[495], x[494], x[219], x[218], x[217]}), .y(y[216]));
  R1ind217 R1ind217_inst(.x({x[95], x[94], x[93], x[89], x[88], x[87], x[92], x[91], x[90], x[98], x[97], x[96]}), .y(y[217]));
  R1ind218 R1ind218_inst(.x({x[497], x[496], x[219], x[218], x[217]}), .y(y[218]));
  R1ind219 R1ind219_inst(.x({x[95], x[94], x[93], x[89], x[88], x[87], x[98], x[97], x[96], x[92], x[91], x[90]}), .y(y[219]));
  R1ind220 R1ind220_inst(.x({x[201], x[200], x[199], x[195], x[499], x[498], x[219], x[218], x[217]}), .y(y[220]));
  R1ind221 R1ind221_inst(.x({x[83], x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[86], x[85], x[84]}), .y(y[221]));
  R1ind222 R1ind222_inst(.x({x[207], x[206], x[205], x[195], x[501], x[500], x[219], x[218], x[217]}), .y(y[222]));
  R1ind223 R1ind223_inst(.x({x[83], x[82], x[81], x[77], x[76], x[75], x[80], x[79], x[78], x[86], x[85], x[84]}), .y(y[223]));
  R1ind224 R1ind224_inst(.x({x[204], x[203], x[202], x[195], x[503], x[502], x[219], x[218], x[217]}), .y(y[224]));
  R1ind225 R1ind225_inst(.x({x[83], x[82], x[81], x[77], x[76], x[75], x[80], x[79], x[78], x[86], x[85], x[84]}), .y(y[225]));
  R1ind226 R1ind226_inst(.x({x[505], x[504], x[219], x[218], x[217]}), .y(y[226]));
  R1ind227 R1ind227_inst(.x({x[83], x[82], x[81], x[77], x[76], x[75], x[86], x[85], x[84], x[80], x[79], x[78]}), .y(y[227]));
  R1ind228 R1ind228_inst(.x({x[210], x[209], x[208], x[195], x[507], x[506], x[219], x[218], x[217]}), .y(y[228]));
  R1ind229 R1ind229_inst(.x({x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[74], x[73], x[72]}), .y(y[229]));
  R1ind230 R1ind230_inst(.x({x[213], x[212], x[211], x[195], x[509], x[508], x[219], x[218], x[217]}), .y(y[230]));
  R1ind231 R1ind231_inst(.x({x[71], x[70], x[69], x[65], x[64], x[63], x[68], x[67], x[66], x[74], x[73], x[72]}), .y(y[231]));
  R1ind232 R1ind232_inst(.x({x[216], x[215], x[214], x[195], x[511], x[510], x[219], x[218], x[217]}), .y(y[232]));
  R1ind233 R1ind233_inst(.x({x[71], x[70], x[69], x[65], x[64], x[63], x[68], x[67], x[66], x[74], x[73], x[72]}), .y(y[233]));
  R1ind234 R1ind234_inst(.x({x[198], x[197], x[196], x[195], x[513], x[512], x[219], x[218], x[217]}), .y(y[234]));
  R1ind235 R1ind235_inst(.x({x[71], x[70], x[69], x[65], x[64], x[63], x[74], x[73], x[72], x[68], x[67], x[66]}), .y(y[235]));
  R1ind236 R1ind236_inst(.x({x[515], x[514], x[219], x[218], x[217]}), .y(y[236]));
  R1ind237 R1ind237_inst(.x({x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[26], x[25], x[24]}), .y(y[237]));
  R1ind238 R1ind238_inst(.x({x[517], x[516], x[219], x[218], x[217]}), .y(y[238]));
  R1ind239 R1ind239_inst(.x({x[23], x[22], x[21], x[17], x[16], x[15], x[20], x[19], x[18], x[26], x[25], x[24]}), .y(y[239]));
  R1ind240 R1ind240_inst(.x({x[519], x[518], x[219], x[218], x[217]}), .y(y[240]));
  R1ind241 R1ind241_inst(.x({x[23], x[22], x[21], x[17], x[16], x[15], x[20], x[19], x[18], x[26], x[25], x[24]}), .y(y[241]));
  R1ind242 R1ind242_inst(.x({x[521], x[520], x[219], x[218], x[217]}), .y(y[242]));
  R1ind243 R1ind243_inst(.x({x[23], x[22], x[21], x[17], x[16], x[15], x[26], x[25], x[24], x[20], x[19], x[18]}), .y(y[243]));
  R1ind244 R1ind244_inst(.x({x[523], x[522], x[219], x[218], x[217]}), .y(y[244]));
  R1ind245 R1ind245_inst(.x({x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[38], x[37], x[36]}), .y(y[245]));
  R1ind246 R1ind246_inst(.x({x[525], x[524], x[219], x[218], x[217]}), .y(y[246]));
  R1ind247 R1ind247_inst(.x({x[35], x[34], x[33], x[29], x[28], x[27], x[32], x[31], x[30], x[38], x[37], x[36]}), .y(y[247]));
  R1ind248 R1ind248_inst(.x({x[527], x[526], x[219], x[218], x[217]}), .y(y[248]));
  R1ind249 R1ind249_inst(.x({x[35], x[34], x[33], x[29], x[28], x[27], x[32], x[31], x[30], x[38], x[37], x[36]}), .y(y[249]));
  R1ind250 R1ind250_inst(.x({x[529], x[528], x[219], x[218], x[217]}), .y(y[250]));
  R1ind251 R1ind251_inst(.x({x[35], x[34], x[33], x[29], x[28], x[27], x[38], x[37], x[36], x[32], x[31], x[30]}), .y(y[251]));
  R1ind252 R1ind252_inst(.x({x[531], x[530], x[219], x[218], x[217]}), .y(y[252]));
  R1ind253 R1ind253_inst(.x({x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[50], x[49], x[48]}), .y(y[253]));
  R1ind254 R1ind254_inst(.x({x[533], x[532], x[219], x[218], x[217]}), .y(y[254]));
  R1ind255 R1ind255_inst(.x({x[47], x[46], x[45], x[41], x[40], x[39], x[44], x[43], x[42], x[50], x[49], x[48]}), .y(y[255]));
  R1ind256 R1ind256_inst(.x({x[535], x[534], x[219], x[218], x[217]}), .y(y[256]));
  R1ind257 R1ind257_inst(.x({x[47], x[46], x[45], x[41], x[40], x[39], x[44], x[43], x[42], x[50], x[49], x[48]}), .y(y[257]));
  R1ind258 R1ind258_inst(.x({x[537], x[536], x[219], x[218], x[217]}), .y(y[258]));
  R1ind259 R1ind259_inst(.x({x[47], x[46], x[45], x[41], x[40], x[39], x[50], x[49], x[48], x[44], x[43], x[42]}), .y(y[259]));
  R1ind260 R1ind260_inst(.x({x[539], x[538], x[219], x[218], x[217]}), .y(y[260]));
  R1ind261 R1ind261_inst(.x({x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[14], x[13], x[12]}), .y(y[261]));
  R1ind262 R1ind262_inst(.x({x[541], x[540], x[219], x[218], x[217]}), .y(y[262]));
  R1ind263 R1ind263_inst(.x({x[11], x[10], x[9], x[5], x[4], x[3], x[8], x[7], x[6], x[14], x[13], x[12]}), .y(y[263]));
  R1ind264 R1ind264_inst(.x({x[543], x[542], x[219], x[218], x[217]}), .y(y[264]));
  R1ind265 R1ind265_inst(.x({x[11], x[10], x[9], x[5], x[4], x[3], x[8], x[7], x[6], x[14], x[13], x[12]}), .y(y[265]));
  R1ind266 R1ind266_inst(.x({x[545], x[544], x[219], x[218], x[217]}), .y(y[266]));
  R1ind267 R1ind267_inst(.x({x[11], x[10], x[9], x[5], x[4], x[3], x[14], x[13], x[12], x[8], x[7], x[6]}), .y(y[267]));
endmodule

module R2ind0(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (t[2] & ~t[3]);
  assign t[2] = t[4] ^ x[2];
  assign t[3] = t[5] ^ x[1];
  assign t[4] = (x[0]);
  assign t[5] = (x[0]);
  assign y = t[0];
endmodule

module R2ind1(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0]);
  assign t[5] = (x[0]);
  assign y = t[0];
endmodule

module R2ind2(x, y);
 input [21:0] x;
 output y;

 wire [61:0] t;
  assign t[0] = t[1] & t[2];
  assign t[10] = ~(~x[0] & ~t[17]);
  assign t[11] = ~x[0] & t[18];
  assign t[12] = ~x[0] & t[19];
  assign t[13] = (t[20]);
  assign t[14] = (t[21]);
  assign t[15] = (t[22]);
  assign t[16] = (t[23]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~x[0] & t[13];
  assign t[20] = t[27] ^ x[3];
  assign t[21] = t[28] ^ x[6];
  assign t[22] = t[29] ^ x[9];
  assign t[23] = t[30] ^ x[12];
  assign t[24] = t[31] ^ x[15];
  assign t[25] = t[32] ^ x[18];
  assign t[26] = t[33] ^ x[21];
  assign t[27] = (t[34] & ~t[35]);
  assign t[28] = (t[36] & ~t[37]);
  assign t[29] = (t[38] & ~t[39]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (t[40] & ~t[41]);
  assign t[31] = (t[42] & ~t[43]);
  assign t[32] = (t[44] & ~t[45]);
  assign t[33] = (t[46] & ~t[47]);
  assign t[34] = t[48] ^ x[3];
  assign t[35] = t[49] ^ x[2];
  assign t[36] = t[50] ^ x[6];
  assign t[37] = t[51] ^ x[5];
  assign t[38] = t[52] ^ x[9];
  assign t[39] = t[53] ^ x[8];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[54] ^ x[12];
  assign t[41] = t[55] ^ x[11];
  assign t[42] = t[56] ^ x[15];
  assign t[43] = t[57] ^ x[14];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[17];
  assign t[46] = t[60] ^ x[21];
  assign t[47] = t[61] ^ x[20];
  assign t[48] = (x[1]);
  assign t[49] = (x[1]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[50] = (x[4]);
  assign t[51] = (x[4]);
  assign t[52] = (x[7]);
  assign t[53] = (x[7]);
  assign t[54] = (x[10]);
  assign t[55] = (x[10]);
  assign t[56] = (x[13]);
  assign t[57] = (x[13]);
  assign t[58] = (x[16]);
  assign t[59] = (x[16]);
  assign t[5] = ~(~x[0] & ~t[14]);
  assign t[60] = (x[19]);
  assign t[61] = (x[19]);
  assign t[6] = ~x[0] & t[15];
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = ~(t[11] | t[12]);
  assign t[9] = ~x[0] & t[16];
  assign y = (t[0]);
endmodule

module R2ind3(x, y);
 input [21:0] x;
 output y;

 wire [61:0] t;
  assign t[0] = t[1] & t[2];
  assign t[10] = ~(~x[0] & ~t[17]);
  assign t[11] = ~x[0] & t[18];
  assign t[12] = ~x[0] & t[19];
  assign t[13] = (t[20]);
  assign t[14] = (t[21]);
  assign t[15] = (t[22]);
  assign t[16] = (t[23]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~x[0] & t[13];
  assign t[20] = t[27] ^ x[3];
  assign t[21] = t[28] ^ x[6];
  assign t[22] = t[29] ^ x[9];
  assign t[23] = t[30] ^ x[12];
  assign t[24] = t[31] ^ x[15];
  assign t[25] = t[32] ^ x[18];
  assign t[26] = t[33] ^ x[21];
  assign t[27] = (t[34] & ~t[35]);
  assign t[28] = (t[36] & ~t[37]);
  assign t[29] = (t[38] & ~t[39]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (t[40] & ~t[41]);
  assign t[31] = (t[42] & ~t[43]);
  assign t[32] = (t[44] & ~t[45]);
  assign t[33] = (t[46] & ~t[47]);
  assign t[34] = t[48] ^ x[3];
  assign t[35] = t[49] ^ x[2];
  assign t[36] = t[50] ^ x[6];
  assign t[37] = t[51] ^ x[5];
  assign t[38] = t[52] ^ x[9];
  assign t[39] = t[53] ^ x[8];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[54] ^ x[12];
  assign t[41] = t[55] ^ x[11];
  assign t[42] = t[56] ^ x[15];
  assign t[43] = t[57] ^ x[14];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[17];
  assign t[46] = t[60] ^ x[21];
  assign t[47] = t[61] ^ x[20];
  assign t[48] = (x[1]);
  assign t[49] = (x[1]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[50] = (x[4]);
  assign t[51] = (x[4]);
  assign t[52] = (x[7]);
  assign t[53] = (x[7]);
  assign t[54] = (x[10]);
  assign t[55] = (x[10]);
  assign t[56] = (x[13]);
  assign t[57] = (x[13]);
  assign t[58] = (x[16]);
  assign t[59] = (x[16]);
  assign t[5] = ~(~x[0] & ~t[14]);
  assign t[60] = (x[19]);
  assign t[61] = (x[19]);
  assign t[6] = ~x[0] & t[15];
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = ~(t[11] | t[12]);
  assign t[9] = ~x[0] & t[16];
  assign y = (t[0]);
endmodule

module R2ind4(x, y);
 input [3:0] x;
 output y;

 wire [9:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = ~(t[2]);
  assign t[2] = ~x[0] & t[3];
  assign t[3] = (t[4]);
  assign t[4] = t[5] ^ x[3];
  assign t[5] = (t[6] & ~t[7]);
  assign t[6] = t[8] ^ x[3];
  assign t[7] = t[9] ^ x[2];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind5(x, y);
 input [3:0] x;
 output y;

 wire [9:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = ~(t[2]);
  assign t[2] = ~x[0] & t[3];
  assign t[3] = (t[4]);
  assign t[4] = t[5] ^ x[3];
  assign t[5] = (t[6] & ~t[7]);
  assign t[6] = t[8] ^ x[3];
  assign t[7] = t[9] ^ x[2];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind6(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[3];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[1]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind7(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[3];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[1]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind8(x, y);
 input [6:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[14] ^ x[2];
  assign t[11] = t[15] ^ x[6];
  assign t[12] = t[16] ^ x[5];
  assign t[13] = (x[1]);
  assign t[14] = (x[1]);
  assign t[15] = (x[4]);
  assign t[16] = (x[4]);
  assign t[1] = ~x[0] & t[3];
  assign t[2] = ~(~x[0] & ~t[4]);
  assign t[3] = (t[5]);
  assign t[4] = (t[6]);
  assign t[5] = t[7] ^ x[3];
  assign t[6] = t[8] ^ x[6];
  assign t[7] = (t[9] & ~t[10]);
  assign t[8] = (t[11] & ~t[12]);
  assign t[9] = t[13] ^ x[3];
  assign y = (t[0]);
endmodule

module R2ind9(x, y);
 input [6:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[14] ^ x[2];
  assign t[11] = t[15] ^ x[6];
  assign t[12] = t[16] ^ x[5];
  assign t[13] = (x[1]);
  assign t[14] = (x[1]);
  assign t[15] = (x[4]);
  assign t[16] = (x[4]);
  assign t[1] = ~x[0] & t[3];
  assign t[2] = ~(~x[0] & ~t[4]);
  assign t[3] = (t[5]);
  assign t[4] = (t[6]);
  assign t[5] = t[7] ^ x[3];
  assign t[6] = t[8] ^ x[6];
  assign t[7] = (t[9] & ~t[10]);
  assign t[8] = (t[11] & ~t[12]);
  assign t[9] = t[13] ^ x[3];
  assign y = (t[0]);
endmodule

module R2ind10(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[3];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[1]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind11(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[3];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[1]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind12(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[3];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[1]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind13(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[3];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[1]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind14(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[3];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[1]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind15(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[3];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[1]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind16(x, y);
 input [6:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[14] ^ x[2];
  assign t[11] = t[15] ^ x[6];
  assign t[12] = t[16] ^ x[5];
  assign t[13] = (x[1]);
  assign t[14] = (x[1]);
  assign t[15] = (x[4]);
  assign t[16] = (x[4]);
  assign t[1] = ~(~x[0] & ~t[3]);
  assign t[2] = ~x[0] & t[4];
  assign t[3] = (t[5]);
  assign t[4] = (t[6]);
  assign t[5] = t[7] ^ x[3];
  assign t[6] = t[8] ^ x[6];
  assign t[7] = (t[9] & ~t[10]);
  assign t[8] = (t[11] & ~t[12]);
  assign t[9] = t[13] ^ x[3];
  assign y = (t[0]);
endmodule

module R2ind17(x, y);
 input [6:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[14] ^ x[2];
  assign t[11] = t[15] ^ x[6];
  assign t[12] = t[16] ^ x[5];
  assign t[13] = (x[1]);
  assign t[14] = (x[1]);
  assign t[15] = (x[4]);
  assign t[16] = (x[4]);
  assign t[1] = ~(~x[0] & ~t[3]);
  assign t[2] = ~x[0] & t[4];
  assign t[3] = (t[5]);
  assign t[4] = (t[6]);
  assign t[5] = t[7] ^ x[3];
  assign t[6] = t[8] ^ x[6];
  assign t[7] = (t[9] & ~t[10]);
  assign t[8] = (t[11] & ~t[12]);
  assign t[9] = t[13] ^ x[3];
  assign y = (t[0]);
endmodule

module R2ind18(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind19(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind20(x, y);
 input [6:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[14] ^ x[1];
  assign t[11] = t[15] ^ x[6];
  assign t[12] = t[16] ^ x[5];
  assign t[13] = (x[0]);
  assign t[14] = (x[0]);
  assign t[15] = (x[4]);
  assign t[16] = (x[4]);
  assign t[1] = ~t[3];
  assign t[2] = ~x[3] & t[4];
  assign t[3] = (t[5]);
  assign t[4] = (t[6]);
  assign t[5] = t[7] ^ x[2];
  assign t[6] = t[8] ^ x[6];
  assign t[7] = (t[9] & ~t[10]);
  assign t[8] = (t[11] & ~t[12]);
  assign t[9] = t[13] ^ x[2];
  assign y = (t[0]);
endmodule

module R2ind21(x, y);
 input [6:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[14] ^ x[1];
  assign t[11] = t[15] ^ x[6];
  assign t[12] = t[16] ^ x[5];
  assign t[13] = (x[0]);
  assign t[14] = (x[0]);
  assign t[15] = (x[4]);
  assign t[16] = (x[4]);
  assign t[1] = ~t[3];
  assign t[2] = ~x[3] & t[4];
  assign t[3] = (t[5]);
  assign t[4] = (t[6]);
  assign t[5] = t[7] ^ x[2];
  assign t[6] = t[8] ^ x[6];
  assign t[7] = (t[9] & ~t[10]);
  assign t[8] = (t[11] & ~t[12]);
  assign t[9] = t[13] ^ x[2];
  assign y = (t[0]);
endmodule

module R2ind22(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[3];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[1]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind23(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[3];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[1]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind24(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind25(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind26(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind27(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind28(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind29(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind30(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind31(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind32(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind33(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind34(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind35(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind36(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind37(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind38(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind39(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind40(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind41(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind42(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind43(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind44(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind45(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind46(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind47(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind48(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind49(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind50(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind51(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind52(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind53(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind54(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind55(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind56(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind57(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind58(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind59(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind60(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind61(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind62(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind63(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind64(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind65(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind66(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind67(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind68(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind69(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind70(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind71(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind72(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind73(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind74(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind75(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind76(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind77(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind78(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind79(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind80(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind81(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind82(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind83(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind84(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind85(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind86(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind87(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~t[1];
  assign t[1] = x[3] ? x[2] : x[0];
  assign t[2] = ~(t[0] ^ x[1]);
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind88(x, y);
 input [5:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[5] ? x[3] : x[0];
  assign t[4] = x[5] ? x[4] : x[1];
  assign t[5] = ~(t[0] ^ x[2]);
  assign y = t[5] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind89(x, y);
 input [5:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[5] ? x[3] : x[0];
  assign t[4] = x[5] ? x[4] : x[1];
  assign t[5] = ~(t[0] ^ x[2]);
  assign y = t[5] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind90(x, y);
 input [5:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[5] ? x[3] : x[0];
  assign t[4] = x[5] ? x[4] : x[1];
  assign t[5] = ~(t[0] ^ x[2]);
  assign y = t[5] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind91(x, y);
 input [5:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[5] ? x[3] : x[0];
  assign t[4] = x[5] ? x[4] : x[1];
  assign t[5] = ~(t[0] ^ x[2]);
  assign y = t[5] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind92(x, y);
 input [5:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[5] ? x[3] : x[0];
  assign t[4] = x[5] ? x[4] : x[1];
  assign t[5] = ~(t[0] ^ x[2]);
  assign y = t[5] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind93(x, y);
 input [5:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[5] ? x[3] : x[0];
  assign t[4] = x[5] ? x[4] : x[1];
  assign t[5] = ~(t[0] ^ x[2]);
  assign y = t[5] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind94(x, y);
 input [5:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[5] ? x[4] : x[1];
  assign t[4] = x[5] ? x[3] : x[0];
  assign t[5] = ~(t[0] ^ x[2]);
  assign y = t[5] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind95(x, y);
 input [5:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[5] ? x[4] : x[1];
  assign t[4] = x[5] ? x[3] : x[0];
  assign t[5] = ~(t[0] ^ x[2]);
  assign y = t[5] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind96(x, y);
 input [5:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[5] ? x[4] : x[1];
  assign t[4] = x[5] ? x[3] : x[0];
  assign t[5] = ~(t[0] ^ x[2]);
  assign y = t[5] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind97(x, y);
 input [5:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[5] ? x[4] : x[1];
  assign t[4] = x[5] ? x[3] : x[0];
  assign t[5] = ~(t[0] ^ x[2]);
  assign y = t[5] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind98(x, y);
 input [5:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[5] ? x[4] : x[1];
  assign t[4] = x[5] ? x[3] : x[0];
  assign t[5] = ~(t[0] ^ x[2]);
  assign y = t[5] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind99(x, y);
 input [5:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[5] ? x[4] : x[1];
  assign t[4] = x[5] ? x[3] : x[0];
  assign t[5] = ~(t[0] ^ x[2]);
  assign y = t[5] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind100(x, y);
 input [5:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[5] ? x[4] : x[1];
  assign t[4] = x[5] ? x[3] : x[0];
  assign t[5] = ~(t[0] ^ x[2]);
  assign y = t[5] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind101(x, y);
 input [5:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[5] ? x[4] : x[1];
  assign t[4] = x[5] ? x[3] : x[0];
  assign t[5] = ~(t[0] ^ x[2]);
  assign y = t[5] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind102(x, y);
 input [5:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[5] ? x[4] : x[1];
  assign t[4] = x[5] ? x[3] : x[0];
  assign t[5] = ~(t[0] ^ x[2]);
  assign y = t[5] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind103(x, y);
 input [5:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[5] ? x[4] : x[1];
  assign t[4] = x[5] ? x[3] : x[0];
  assign t[5] = ~(t[0] ^ x[2]);
  assign y = t[5] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind104(x, y);
 input [5:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[5] ? x[4] : x[1];
  assign t[4] = x[5] ? x[3] : x[0];
  assign t[5] = ~(t[0] ^ x[2]);
  assign y = t[5] ^ 1'b1 ^ 1'b1;
endmodule

module R2ind105(x, y);
 input [5:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[5] ? x[4] : x[1];
  assign t[4] = x[5] ? x[3] : x[0];
  assign t[5] = ~(t[0] ^ x[2]);
  assign y = t[5] ^ 1'b1 ^ 1'b1;
endmodule

module R2ind106(x, y);
 input [5:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[5] ? x[4] : x[1];
  assign t[4] = x[5] ? x[3] : x[0];
  assign t[5] = ~(t[0] ^ x[2]);
  assign y = t[5] ^ 1'b1 ^ 1'b1;
endmodule

module R2ind107(x, y);
 input [5:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[5] ? x[4] : x[1];
  assign t[4] = x[5] ? x[3] : x[0];
  assign t[5] = ~(t[0] ^ x[2]);
  assign y = t[5] ^ 1'b1 ^ 1'b1;
endmodule

module R2ind108(x, y);
 input [5:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[5] ? x[3] : x[0];
  assign t[4] = x[5] ? x[4] : x[1];
  assign t[5] = ~(t[0] ^ x[2]);
  assign y = t[5] ^ 1'b1 ^ 1'b1;
endmodule

module R2ind109(x, y);
 input [5:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[5] ? x[3] : x[0];
  assign t[4] = x[5] ? x[4] : x[1];
  assign t[5] = ~(t[0] ^ x[2]);
  assign y = t[5] ^ 1'b1 ^ 1'b1;
endmodule

module R2ind110(x, y);
 input [5:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[5] ? x[3] : x[0];
  assign t[4] = x[5] ? x[4] : x[1];
  assign t[5] = ~(t[0] ^ x[2]);
  assign y = t[5] ^ 1'b1 ^ 1'b1;
endmodule

module R2ind111(x, y);
 input [5:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[5] ? x[3] : x[0];
  assign t[4] = x[5] ? x[4] : x[1];
  assign t[5] = ~(t[0] ^ x[2]);
  assign y = t[5] ^ 1'b1 ^ 1'b1;
endmodule

module R2ind112(x, y);
 input [5:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[5] ? x[3] : x[0];
  assign t[4] = x[5] ? x[4] : x[1];
  assign t[5] = ~(t[0] ^ x[2]);
  assign y = t[5] ^ 1'b1 ^ 1'b1;
endmodule

module R2ind113(x, y);
 input [5:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[5] ? x[3] : x[0];
  assign t[4] = x[5] ? x[4] : x[1];
  assign t[5] = ~(t[0] ^ x[2]);
  assign y = t[5] ^ 1'b1 ^ 1'b1;
endmodule

module R2ind114(x, y);
 input [5:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[5] ? x[3] : x[0];
  assign t[4] = x[5] ? x[4] : x[1];
  assign t[5] = ~(t[0] ^ x[2]);
  assign y = t[5] ^ 1'b1 ^ 1'b1;
endmodule

module R2ind115(x, y);
 input [5:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[5] ? x[3] : x[0];
  assign t[4] = x[5] ? x[4] : x[1];
  assign t[5] = ~(t[0] ^ x[2]);
  assign y = t[5] ^ 1'b1 ^ 1'b1;
endmodule

module R2ind116(x, y);
 input [5:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[5] ? x[3] : x[0];
  assign t[4] = x[5] ? x[4] : x[1];
  assign t[5] = ~(t[0] ^ x[2]);
  assign y = t[5] ^ 1'b1 ^ 1'b1;
endmodule

module R2ind117(x, y);
 input [5:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[5] ? x[3] : x[0];
  assign t[4] = x[5] ? x[4] : x[1];
  assign t[5] = ~(t[0] ^ x[2]);
  assign y = t[5] ^ 1'b1 ^ 1'b1;
endmodule

module R2ind118(x, y);
 input [5:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[5] ? x[3] : x[0];
  assign t[4] = x[5] ? x[4] : x[1];
  assign t[5] = ~(t[0] ^ x[2]);
  assign y = t[5] ^ 1'b1 ^ 1'b1;
endmodule

module R2ind119(x, y);
 input [5:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = ~t[4];
  assign t[3] = x[5] ? x[3] : x[0];
  assign t[4] = x[5] ? x[4] : x[1];
  assign t[5] = ~(t[0] ^ x[2]);
  assign y = t[5] ^ 1'b1 ^ 1'b1;
endmodule

module R2ind120(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[7] ? x[6] : x[2];
  assign t[5] = x[7] ? x[5] : x[1];
  assign t[6] = x[7] ? x[4] : x[0];
  assign t[7] = ~(t[0] ^ x[3]);
  assign y = t[7] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind121(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[7] ? x[6] : x[2];
  assign t[5] = x[7] ? x[5] : x[1];
  assign t[6] = x[7] ? x[4] : x[0];
  assign t[7] = ~(t[0] ^ x[3]);
  assign y = t[7] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind122(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[7] ? x[6] : x[2];
  assign t[5] = x[7] ? x[4] : x[0];
  assign t[6] = x[7] ? x[5] : x[1];
  assign t[7] = ~(t[0] ^ x[3]);
  assign y = t[7] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind123(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[7] ? x[6] : x[2];
  assign t[5] = x[7] ? x[4] : x[0];
  assign t[6] = x[7] ? x[5] : x[1];
  assign t[7] = ~(t[0] ^ x[3]);
  assign y = t[7] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind124(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[7] ? x[6] : x[2];
  assign t[5] = x[7] ? x[4] : x[0];
  assign t[6] = x[7] ? x[5] : x[1];
  assign t[7] = ~(t[0] ^ x[3]);
  assign y = t[7] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind125(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[7] ? x[6] : x[2];
  assign t[5] = x[7] ? x[4] : x[0];
  assign t[6] = x[7] ? x[5] : x[1];
  assign t[7] = ~(t[0] ^ x[3]);
  assign y = t[7] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind126(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[7] ? x[6] : x[2];
  assign t[5] = x[7] ? x[4] : x[0];
  assign t[6] = x[7] ? x[5] : x[1];
  assign t[7] = ~(t[0] ^ x[3]);
  assign y = t[7] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind127(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[7] ? x[6] : x[2];
  assign t[5] = x[7] ? x[4] : x[0];
  assign t[6] = x[7] ? x[5] : x[1];
  assign t[7] = ~(t[0] ^ x[3]);
  assign y = t[7] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind128(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[7] ? x[6] : x[2];
  assign t[5] = x[7] ? x[4] : x[0];
  assign t[6] = x[7] ? x[5] : x[1];
  assign t[7] = ~(t[0] ^ x[3]);
  assign y = t[7] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind129(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[7] ? x[6] : x[2];
  assign t[5] = x[7] ? x[4] : x[0];
  assign t[6] = x[7] ? x[5] : x[1];
  assign t[7] = ~(t[0] ^ x[3]);
  assign y = t[7] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind130(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[7] ? x[5] : x[1];
  assign t[5] = x[7] ? x[4] : x[0];
  assign t[6] = x[7] ? x[6] : x[2];
  assign t[7] = ~(t[0] ^ x[3]);
  assign y = t[7] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind131(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[7] ? x[5] : x[1];
  assign t[5] = x[7] ? x[4] : x[0];
  assign t[6] = x[7] ? x[6] : x[2];
  assign t[7] = ~(t[0] ^ x[3]);
  assign y = t[7] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind132(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[7] ? x[5] : x[1];
  assign t[5] = x[7] ? x[4] : x[0];
  assign t[6] = x[7] ? x[6] : x[2];
  assign t[7] = ~(t[0] ^ x[3]);
  assign y = t[7] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind133(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[7] ? x[5] : x[1];
  assign t[5] = x[7] ? x[4] : x[0];
  assign t[6] = x[7] ? x[6] : x[2];
  assign t[7] = ~(t[0] ^ x[3]);
  assign y = t[7] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind134(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[7] ? x[5] : x[1];
  assign t[5] = x[7] ? x[4] : x[0];
  assign t[6] = x[7] ? x[6] : x[2];
  assign t[7] = ~(t[0] ^ x[3]);
  assign y = t[7] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind135(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[7] ? x[5] : x[1];
  assign t[5] = x[7] ? x[4] : x[0];
  assign t[6] = x[7] ? x[6] : x[2];
  assign t[7] = ~(t[0] ^ x[3]);
  assign y = t[7] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind136(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[7] ? x[5] : x[1];
  assign t[5] = x[7] ? x[4] : x[0];
  assign t[6] = x[7] ? x[6] : x[2];
  assign t[7] = ~(t[0] ^ x[3]);
  assign y = t[7] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind137(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[7] ? x[5] : x[1];
  assign t[5] = x[7] ? x[4] : x[0];
  assign t[6] = x[7] ? x[6] : x[2];
  assign t[7] = ~(t[0] ^ x[3]);
  assign y = t[7] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind138(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[7] ? x[5] : x[1];
  assign t[5] = x[7] ? x[4] : x[0];
  assign t[6] = x[7] ? x[6] : x[2];
  assign t[7] = ~(t[0] ^ x[3]);
  assign y = t[7] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind139(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[7] ? x[5] : x[1];
  assign t[5] = x[7] ? x[4] : x[0];
  assign t[6] = x[7] ? x[6] : x[2];
  assign t[7] = ~(t[0] ^ x[3]);
  assign y = t[7] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind140(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[7] ? x[6] : x[2];
  assign t[5] = x[7] ? x[5] : x[1];
  assign t[6] = x[7] ? x[4] : x[0];
  assign t[7] = ~(t[0] ^ x[3]);
  assign y = t[7] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind141(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[7] ? x[6] : x[2];
  assign t[5] = x[7] ? x[5] : x[1];
  assign t[6] = x[7] ? x[4] : x[0];
  assign t[7] = ~(t[0] ^ x[3]);
  assign y = t[7] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind142(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[7] ? x[6] : x[2];
  assign t[5] = x[7] ? x[5] : x[1];
  assign t[6] = x[7] ? x[4] : x[0];
  assign t[7] = ~(t[0] ^ x[3]);
  assign y = t[7] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind143(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[7] ? x[6] : x[2];
  assign t[5] = x[7] ? x[5] : x[1];
  assign t[6] = x[7] ? x[4] : x[0];
  assign t[7] = ~(t[0] ^ x[3]);
  assign y = t[7] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind144(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[7] ? x[6] : x[2];
  assign t[5] = x[7] ? x[5] : x[1];
  assign t[6] = x[7] ? x[4] : x[0];
  assign t[7] = ~(t[0] ^ x[3]);
  assign y = t[7] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind145(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[7] ? x[6] : x[2];
  assign t[5] = x[7] ? x[5] : x[1];
  assign t[6] = x[7] ? x[4] : x[0];
  assign t[7] = ~(t[0] ^ x[3]);
  assign y = t[7] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind146(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[7] ? x[6] : x[2];
  assign t[5] = x[7] ? x[5] : x[1];
  assign t[6] = x[7] ? x[4] : x[0];
  assign t[7] = ~(t[0] ^ x[3]);
  assign y = t[7] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind147(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[7] ? x[6] : x[2];
  assign t[5] = x[7] ? x[5] : x[1];
  assign t[6] = x[7] ? x[4] : x[0];
  assign t[7] = ~(t[0] ^ x[3]);
  assign y = t[7] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind148(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[7] ? x[6] : x[2];
  assign t[5] = x[7] ? x[5] : x[1];
  assign t[6] = x[7] ? x[4] : x[0];
  assign t[7] = ~(t[0] ^ x[3]);
  assign y = t[7] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind149(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[7] ? x[6] : x[2];
  assign t[5] = x[7] ? x[5] : x[1];
  assign t[6] = x[7] ? x[4] : x[0];
  assign t[7] = ~(t[0] ^ x[3]);
  assign y = t[7] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind150(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[7] ? x[6] : x[2];
  assign t[5] = x[7] ? x[5] : x[1];
  assign t[6] = x[7] ? x[4] : x[0];
  assign t[7] = ~(t[0] ^ x[3]);
  assign y = t[7] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind151(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~t[1];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[2] = t[4];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[4] = x[7] ? x[6] : x[2];
  assign t[5] = x[7] ? x[5] : x[1];
  assign t[6] = x[7] ? x[4] : x[0];
  assign t[7] = ~(t[0] ^ x[3]);
  assign y = t[7] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind152(x, y);
 input [11:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[7] ^ t[23];
  assign t[11] = t[13] ^ t[4];
  assign t[12] = t[14] & t[15];
  assign t[13] = t[16] & t[17];
  assign t[14] = ~(t[13] ^ t[18]);
  assign t[15] = t[3] ^ t[19];
  assign t[16] = ~(t[19]);
  assign t[17] = ~(t[7]);
  assign t[18] = t[5] ^ t[7];
  assign t[19] = t[10] ^ t[20];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = t[28] ^ x[2];
  assign t[25] = t[29] ^ x[5];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = t[31] ^ x[11];
  assign t[28] = (t[32] & ~t[33]);
  assign t[29] = (t[34] & ~t[35]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[36] & ~t[37]);
  assign t[31] = (t[38] & ~t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[1];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[4];
  assign t[36] = t[44] ^ x[8];
  assign t[37] = t[45] ^ x[7];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[10];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[4] = t[9] & t[10];
  assign t[5] = t[20] ^ t[8];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[21] ^ t[20];
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind153(x, y);
 input [11:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[7] ^ t[23];
  assign t[11] = t[13] ^ t[4];
  assign t[12] = t[14] & t[15];
  assign t[13] = t[16] & t[17];
  assign t[14] = ~(t[13] ^ t[18]);
  assign t[15] = t[3] ^ t[19];
  assign t[16] = ~(t[19]);
  assign t[17] = ~(t[7]);
  assign t[18] = t[5] ^ t[7];
  assign t[19] = t[10] ^ t[20];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = t[28] ^ x[2];
  assign t[25] = t[29] ^ x[5];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = t[31] ^ x[11];
  assign t[28] = (t[32] & ~t[33]);
  assign t[29] = (t[34] & ~t[35]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[36] & ~t[37]);
  assign t[31] = (t[38] & ~t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[1];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[4];
  assign t[36] = t[44] ^ x[8];
  assign t[37] = t[45] ^ x[7];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[10];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[4] = t[9] & t[10];
  assign t[5] = t[20] ^ t[8];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[21] ^ t[20];
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind154(x, y);
 input [11:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[24] ^ t[22];
  assign t[12] = ~(t[22]);
  assign t[13] = t[11] ^ t[25];
  assign t[14] = ~(t[7] ^ t[16]);
  assign t[15] = t[17] ^ t[13];
  assign t[16] = t[18] ^ t[6];
  assign t[17] = t[22] ^ t[9];
  assign t[18] = t[19] & t[20];
  assign t[19] = ~(t[21]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11]);
  assign t[21] = t[13] ^ t[22];
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34] & ~t[35]);
  assign t[31] = (t[36] & ~t[37]);
  assign t[32] = (t[38] & ~t[39]);
  assign t[33] = (t[40] & ~t[41]);
  assign t[34] = t[42] ^ x[2];
  assign t[35] = t[43] ^ x[1];
  assign t[36] = t[44] ^ x[5];
  assign t[37] = t[45] ^ x[4];
  assign t[38] = t[46] ^ x[8];
  assign t[39] = t[47] ^ x[7];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[11];
  assign t[41] = t[49] ^ x[10];
  assign t[42] = (x[0]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[3]);
  assign t[46] = (x[6]);
  assign t[47] = (x[6]);
  assign t[48] = (x[9]);
  assign t[49] = (x[9]);
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[11] ^ t[9];
  assign t[6] = t[12] & t[13];
  assign t[7] = t[11] ^ t[22];
  assign t[8] = t[14] & t[15];
  assign t[9] = ~(t[23]);
  assign y = (t[0]);
endmodule

module R2ind155(x, y);
 input [11:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[24] ^ t[22];
  assign t[12] = ~(t[22]);
  assign t[13] = t[11] ^ t[25];
  assign t[14] = ~(t[7] ^ t[16]);
  assign t[15] = t[17] ^ t[13];
  assign t[16] = t[18] ^ t[6];
  assign t[17] = t[22] ^ t[9];
  assign t[18] = t[19] & t[20];
  assign t[19] = ~(t[21]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11]);
  assign t[21] = t[13] ^ t[22];
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34] & ~t[35]);
  assign t[31] = (t[36] & ~t[37]);
  assign t[32] = (t[38] & ~t[39]);
  assign t[33] = (t[40] & ~t[41]);
  assign t[34] = t[42] ^ x[2];
  assign t[35] = t[43] ^ x[1];
  assign t[36] = t[44] ^ x[5];
  assign t[37] = t[45] ^ x[4];
  assign t[38] = t[46] ^ x[8];
  assign t[39] = t[47] ^ x[7];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[11];
  assign t[41] = t[49] ^ x[10];
  assign t[42] = (x[0]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[3]);
  assign t[46] = (x[6]);
  assign t[47] = (x[6]);
  assign t[48] = (x[9]);
  assign t[49] = (x[9]);
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[11] ^ t[9];
  assign t[6] = t[12] & t[13];
  assign t[7] = t[11] ^ t[22];
  assign t[8] = t[14] & t[15];
  assign t[9] = ~(t[23]);
  assign y = (t[0]);
endmodule

module R2ind156(x, y);
 input [11:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[15] ^ t[29];
  assign t[12] = t[20] & t[21];
  assign t[13] = ~(t[30]);
  assign t[14] = t[18] ^ t[12];
  assign t[15] = t[31] ^ t[29];
  assign t[16] = ~(t[29]);
  assign t[17] = t[15] ^ t[32];
  assign t[18] = t[22] ^ t[8];
  assign t[19] = t[23] & t[24];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11] ^ t[18]);
  assign t[21] = t[9] ^ t[17];
  assign t[22] = t[25] & t[26];
  assign t[23] = ~(t[22] ^ t[27]);
  assign t[24] = t[7] ^ t[28];
  assign t[25] = ~(t[28]);
  assign t[26] = ~(t[15]);
  assign t[27] = t[9] ^ t[15];
  assign t[28] = t[17] ^ t[29];
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = (t[35]);
  assign t[32] = (t[36]);
  assign t[33] = t[37] ^ x[2];
  assign t[34] = t[38] ^ x[5];
  assign t[35] = t[39] ^ x[8];
  assign t[36] = t[40] ^ x[11];
  assign t[37] = (t[41] & ~t[42]);
  assign t[38] = (t[43] & ~t[44]);
  assign t[39] = (t[45] & ~t[46]);
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (t[47] & ~t[48]);
  assign t[41] = t[49] ^ x[2];
  assign t[42] = t[50] ^ x[1];
  assign t[43] = t[51] ^ x[5];
  assign t[44] = t[52] ^ x[4];
  assign t[45] = t[53] ^ x[8];
  assign t[46] = t[54] ^ x[7];
  assign t[47] = t[55] ^ x[11];
  assign t[48] = t[56] ^ x[10];
  assign t[49] = (x[0]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[0]);
  assign t[51] = (x[3]);
  assign t[52] = (x[3]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[9]);
  assign t[56] = (x[9]);
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[15] ^ t[13];
  assign t[8] = t[16] & t[17];
  assign t[9] = t[29] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind157(x, y);
 input [11:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[15] ^ t[29];
  assign t[12] = t[20] & t[21];
  assign t[13] = ~(t[30]);
  assign t[14] = t[18] ^ t[12];
  assign t[15] = t[31] ^ t[29];
  assign t[16] = ~(t[29]);
  assign t[17] = t[15] ^ t[32];
  assign t[18] = t[22] ^ t[8];
  assign t[19] = t[23] & t[24];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11] ^ t[18]);
  assign t[21] = t[9] ^ t[17];
  assign t[22] = t[25] & t[26];
  assign t[23] = ~(t[22] ^ t[27]);
  assign t[24] = t[7] ^ t[28];
  assign t[25] = ~(t[28]);
  assign t[26] = ~(t[15]);
  assign t[27] = t[9] ^ t[15];
  assign t[28] = t[17] ^ t[29];
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = (t[35]);
  assign t[32] = (t[36]);
  assign t[33] = t[37] ^ x[2];
  assign t[34] = t[38] ^ x[5];
  assign t[35] = t[39] ^ x[8];
  assign t[36] = t[40] ^ x[11];
  assign t[37] = (t[41] & ~t[42]);
  assign t[38] = (t[43] & ~t[44]);
  assign t[39] = (t[45] & ~t[46]);
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (t[47] & ~t[48]);
  assign t[41] = t[49] ^ x[2];
  assign t[42] = t[50] ^ x[1];
  assign t[43] = t[51] ^ x[5];
  assign t[44] = t[52] ^ x[4];
  assign t[45] = t[53] ^ x[8];
  assign t[46] = t[54] ^ x[7];
  assign t[47] = t[55] ^ x[11];
  assign t[48] = t[56] ^ x[10];
  assign t[49] = (x[0]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[0]);
  assign t[51] = (x[3]);
  assign t[52] = (x[3]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[9]);
  assign t[56] = (x[9]);
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[15] ^ t[13];
  assign t[8] = t[16] & t[17];
  assign t[9] = t[29] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind158(x, y);
 input [11:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] ^ t[16];
  assign t[11] = t[17] ^ t[8];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[29] ^ t[28];
  assign t[14] = ~(t[28]);
  assign t[15] = t[13] ^ t[30];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[22] & t[23];
  assign t[18] = ~(t[24] ^ t[11]);
  assign t[19] = t[9] ^ t[15];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[17] ^ t[25]);
  assign t[21] = t[7] ^ t[26];
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[13]);
  assign t[24] = t[13] ^ t[28];
  assign t[25] = t[9] ^ t[13];
  assign t[26] = t[15] ^ t[28];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[2];
  assign t[32] = t[36] ^ x[5];
  assign t[33] = t[37] ^ x[8];
  assign t[34] = t[38] ^ x[11];
  assign t[35] = (t[39] & ~t[40]);
  assign t[36] = (t[41] & ~t[42]);
  assign t[37] = (t[43] & ~t[44]);
  assign t[38] = (t[45] & ~t[46]);
  assign t[39] = t[47] ^ x[2];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[1];
  assign t[41] = t[49] ^ x[5];
  assign t[42] = t[50] ^ x[4];
  assign t[43] = t[51] ^ x[8];
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[11];
  assign t[46] = t[54] ^ x[10];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[5] = ~(t[27]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[13] ^ t[5];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[28] ^ t[5];
  assign y = (t[0]);
endmodule

module R2ind159(x, y);
 input [11:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] ^ t[16];
  assign t[11] = t[17] ^ t[8];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[29] ^ t[28];
  assign t[14] = ~(t[28]);
  assign t[15] = t[13] ^ t[30];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[22] & t[23];
  assign t[18] = ~(t[24] ^ t[11]);
  assign t[19] = t[9] ^ t[15];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[17] ^ t[25]);
  assign t[21] = t[7] ^ t[26];
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[13]);
  assign t[24] = t[13] ^ t[28];
  assign t[25] = t[9] ^ t[13];
  assign t[26] = t[15] ^ t[28];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[2];
  assign t[32] = t[36] ^ x[5];
  assign t[33] = t[37] ^ x[8];
  assign t[34] = t[38] ^ x[11];
  assign t[35] = (t[39] & ~t[40]);
  assign t[36] = (t[41] & ~t[42]);
  assign t[37] = (t[43] & ~t[44]);
  assign t[38] = (t[45] & ~t[46]);
  assign t[39] = t[47] ^ x[2];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[1];
  assign t[41] = t[49] ^ x[5];
  assign t[42] = t[50] ^ x[4];
  assign t[43] = t[51] ^ x[8];
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[11];
  assign t[46] = t[54] ^ x[10];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[5] = ~(t[27]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[13] ^ t[5];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[28] ^ t[5];
  assign y = (t[0]);
endmodule

module R2ind160(x, y);
 input [11:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[7] ^ t[23];
  assign t[11] = t[13] ^ t[4];
  assign t[12] = t[14] & t[15];
  assign t[13] = t[16] & t[17];
  assign t[14] = ~(t[13] ^ t[18]);
  assign t[15] = t[3] ^ t[19];
  assign t[16] = ~(t[19]);
  assign t[17] = ~(t[7]);
  assign t[18] = t[5] ^ t[7];
  assign t[19] = t[10] ^ t[20];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = t[28] ^ x[2];
  assign t[25] = t[29] ^ x[5];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = t[31] ^ x[11];
  assign t[28] = (t[32] & ~t[33]);
  assign t[29] = (t[34] & ~t[35]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[36] & ~t[37]);
  assign t[31] = (t[38] & ~t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[1];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[4];
  assign t[36] = t[44] ^ x[8];
  assign t[37] = t[45] ^ x[7];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[10];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[4] = t[9] & t[10];
  assign t[5] = t[20] ^ t[8];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[21] ^ t[20];
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind161(x, y);
 input [11:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[7] ^ t[23];
  assign t[11] = t[13] ^ t[4];
  assign t[12] = t[14] & t[15];
  assign t[13] = t[16] & t[17];
  assign t[14] = ~(t[13] ^ t[18]);
  assign t[15] = t[3] ^ t[19];
  assign t[16] = ~(t[19]);
  assign t[17] = ~(t[7]);
  assign t[18] = t[5] ^ t[7];
  assign t[19] = t[10] ^ t[20];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = t[28] ^ x[2];
  assign t[25] = t[29] ^ x[5];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = t[31] ^ x[11];
  assign t[28] = (t[32] & ~t[33]);
  assign t[29] = (t[34] & ~t[35]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[36] & ~t[37]);
  assign t[31] = (t[38] & ~t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[1];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[4];
  assign t[36] = t[44] ^ x[8];
  assign t[37] = t[45] ^ x[7];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[10];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[4] = t[9] & t[10];
  assign t[5] = t[20] ^ t[8];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[21] ^ t[20];
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind162(x, y);
 input [11:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[24] ^ t[22];
  assign t[12] = ~(t[22]);
  assign t[13] = t[11] ^ t[25];
  assign t[14] = ~(t[7] ^ t[16]);
  assign t[15] = t[17] ^ t[13];
  assign t[16] = t[18] ^ t[6];
  assign t[17] = t[22] ^ t[9];
  assign t[18] = t[19] & t[20];
  assign t[19] = ~(t[21]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11]);
  assign t[21] = t[13] ^ t[22];
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34] & ~t[35]);
  assign t[31] = (t[36] & ~t[37]);
  assign t[32] = (t[38] & ~t[39]);
  assign t[33] = (t[40] & ~t[41]);
  assign t[34] = t[42] ^ x[2];
  assign t[35] = t[43] ^ x[1];
  assign t[36] = t[44] ^ x[5];
  assign t[37] = t[45] ^ x[4];
  assign t[38] = t[46] ^ x[8];
  assign t[39] = t[47] ^ x[7];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[11];
  assign t[41] = t[49] ^ x[10];
  assign t[42] = (x[0]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[3]);
  assign t[46] = (x[6]);
  assign t[47] = (x[6]);
  assign t[48] = (x[9]);
  assign t[49] = (x[9]);
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[11] ^ t[9];
  assign t[6] = t[12] & t[13];
  assign t[7] = t[11] ^ t[22];
  assign t[8] = t[14] & t[15];
  assign t[9] = ~(t[23]);
  assign y = (t[0]);
endmodule

module R2ind163(x, y);
 input [11:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[24] ^ t[22];
  assign t[12] = ~(t[22]);
  assign t[13] = t[11] ^ t[25];
  assign t[14] = ~(t[7] ^ t[16]);
  assign t[15] = t[17] ^ t[13];
  assign t[16] = t[18] ^ t[6];
  assign t[17] = t[22] ^ t[9];
  assign t[18] = t[19] & t[20];
  assign t[19] = ~(t[21]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11]);
  assign t[21] = t[13] ^ t[22];
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34] & ~t[35]);
  assign t[31] = (t[36] & ~t[37]);
  assign t[32] = (t[38] & ~t[39]);
  assign t[33] = (t[40] & ~t[41]);
  assign t[34] = t[42] ^ x[2];
  assign t[35] = t[43] ^ x[1];
  assign t[36] = t[44] ^ x[5];
  assign t[37] = t[45] ^ x[4];
  assign t[38] = t[46] ^ x[8];
  assign t[39] = t[47] ^ x[7];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[11];
  assign t[41] = t[49] ^ x[10];
  assign t[42] = (x[0]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[3]);
  assign t[46] = (x[6]);
  assign t[47] = (x[6]);
  assign t[48] = (x[9]);
  assign t[49] = (x[9]);
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[11] ^ t[9];
  assign t[6] = t[12] & t[13];
  assign t[7] = t[11] ^ t[22];
  assign t[8] = t[14] & t[15];
  assign t[9] = ~(t[23]);
  assign y = (t[0]);
endmodule

module R2ind164(x, y);
 input [11:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[15] ^ t[29];
  assign t[12] = t[20] & t[21];
  assign t[13] = ~(t[30]);
  assign t[14] = t[18] ^ t[12];
  assign t[15] = t[31] ^ t[29];
  assign t[16] = ~(t[29]);
  assign t[17] = t[15] ^ t[32];
  assign t[18] = t[22] ^ t[8];
  assign t[19] = t[23] & t[24];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11] ^ t[18]);
  assign t[21] = t[9] ^ t[17];
  assign t[22] = t[25] & t[26];
  assign t[23] = ~(t[22] ^ t[27]);
  assign t[24] = t[7] ^ t[28];
  assign t[25] = ~(t[28]);
  assign t[26] = ~(t[15]);
  assign t[27] = t[9] ^ t[15];
  assign t[28] = t[17] ^ t[29];
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = (t[35]);
  assign t[32] = (t[36]);
  assign t[33] = t[37] ^ x[2];
  assign t[34] = t[38] ^ x[5];
  assign t[35] = t[39] ^ x[8];
  assign t[36] = t[40] ^ x[11];
  assign t[37] = (t[41] & ~t[42]);
  assign t[38] = (t[43] & ~t[44]);
  assign t[39] = (t[45] & ~t[46]);
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (t[47] & ~t[48]);
  assign t[41] = t[49] ^ x[2];
  assign t[42] = t[50] ^ x[1];
  assign t[43] = t[51] ^ x[5];
  assign t[44] = t[52] ^ x[4];
  assign t[45] = t[53] ^ x[8];
  assign t[46] = t[54] ^ x[7];
  assign t[47] = t[55] ^ x[11];
  assign t[48] = t[56] ^ x[10];
  assign t[49] = (x[0]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[0]);
  assign t[51] = (x[3]);
  assign t[52] = (x[3]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[9]);
  assign t[56] = (x[9]);
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[15] ^ t[13];
  assign t[8] = t[16] & t[17];
  assign t[9] = t[29] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind165(x, y);
 input [11:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[15] ^ t[29];
  assign t[12] = t[20] & t[21];
  assign t[13] = ~(t[30]);
  assign t[14] = t[18] ^ t[12];
  assign t[15] = t[31] ^ t[29];
  assign t[16] = ~(t[29]);
  assign t[17] = t[15] ^ t[32];
  assign t[18] = t[22] ^ t[8];
  assign t[19] = t[23] & t[24];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11] ^ t[18]);
  assign t[21] = t[9] ^ t[17];
  assign t[22] = t[25] & t[26];
  assign t[23] = ~(t[22] ^ t[27]);
  assign t[24] = t[7] ^ t[28];
  assign t[25] = ~(t[28]);
  assign t[26] = ~(t[15]);
  assign t[27] = t[9] ^ t[15];
  assign t[28] = t[17] ^ t[29];
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = (t[35]);
  assign t[32] = (t[36]);
  assign t[33] = t[37] ^ x[2];
  assign t[34] = t[38] ^ x[5];
  assign t[35] = t[39] ^ x[8];
  assign t[36] = t[40] ^ x[11];
  assign t[37] = (t[41] & ~t[42]);
  assign t[38] = (t[43] & ~t[44]);
  assign t[39] = (t[45] & ~t[46]);
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (t[47] & ~t[48]);
  assign t[41] = t[49] ^ x[2];
  assign t[42] = t[50] ^ x[1];
  assign t[43] = t[51] ^ x[5];
  assign t[44] = t[52] ^ x[4];
  assign t[45] = t[53] ^ x[8];
  assign t[46] = t[54] ^ x[7];
  assign t[47] = t[55] ^ x[11];
  assign t[48] = t[56] ^ x[10];
  assign t[49] = (x[0]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[0]);
  assign t[51] = (x[3]);
  assign t[52] = (x[3]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[9]);
  assign t[56] = (x[9]);
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[15] ^ t[13];
  assign t[8] = t[16] & t[17];
  assign t[9] = t[29] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind166(x, y);
 input [11:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] ^ t[16];
  assign t[11] = t[17] ^ t[8];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[29] ^ t[28];
  assign t[14] = ~(t[28]);
  assign t[15] = t[13] ^ t[30];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[22] & t[23];
  assign t[18] = ~(t[24] ^ t[11]);
  assign t[19] = t[9] ^ t[15];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[17] ^ t[25]);
  assign t[21] = t[7] ^ t[26];
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[13]);
  assign t[24] = t[13] ^ t[28];
  assign t[25] = t[9] ^ t[13];
  assign t[26] = t[15] ^ t[28];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[2];
  assign t[32] = t[36] ^ x[5];
  assign t[33] = t[37] ^ x[8];
  assign t[34] = t[38] ^ x[11];
  assign t[35] = (t[39] & ~t[40]);
  assign t[36] = (t[41] & ~t[42]);
  assign t[37] = (t[43] & ~t[44]);
  assign t[38] = (t[45] & ~t[46]);
  assign t[39] = t[47] ^ x[2];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[1];
  assign t[41] = t[49] ^ x[5];
  assign t[42] = t[50] ^ x[4];
  assign t[43] = t[51] ^ x[8];
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[11];
  assign t[46] = t[54] ^ x[10];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[5] = ~(t[27]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[13] ^ t[5];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[28] ^ t[5];
  assign y = (t[0]);
endmodule

module R2ind167(x, y);
 input [11:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] ^ t[16];
  assign t[11] = t[17] ^ t[8];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[29] ^ t[28];
  assign t[14] = ~(t[28]);
  assign t[15] = t[13] ^ t[30];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[22] & t[23];
  assign t[18] = ~(t[24] ^ t[11]);
  assign t[19] = t[9] ^ t[15];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[17] ^ t[25]);
  assign t[21] = t[7] ^ t[26];
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[13]);
  assign t[24] = t[13] ^ t[28];
  assign t[25] = t[9] ^ t[13];
  assign t[26] = t[15] ^ t[28];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[2];
  assign t[32] = t[36] ^ x[5];
  assign t[33] = t[37] ^ x[8];
  assign t[34] = t[38] ^ x[11];
  assign t[35] = (t[39] & ~t[40]);
  assign t[36] = (t[41] & ~t[42]);
  assign t[37] = (t[43] & ~t[44]);
  assign t[38] = (t[45] & ~t[46]);
  assign t[39] = t[47] ^ x[2];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[1];
  assign t[41] = t[49] ^ x[5];
  assign t[42] = t[50] ^ x[4];
  assign t[43] = t[51] ^ x[8];
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[11];
  assign t[46] = t[54] ^ x[10];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[5] = ~(t[27]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[13] ^ t[5];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[28] ^ t[5];
  assign y = (t[0]);
endmodule

module R2ind168(x, y);
 input [11:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[7] ^ t[23];
  assign t[11] = t[13] ^ t[4];
  assign t[12] = t[14] & t[15];
  assign t[13] = t[16] & t[17];
  assign t[14] = ~(t[13] ^ t[18]);
  assign t[15] = t[3] ^ t[19];
  assign t[16] = ~(t[19]);
  assign t[17] = ~(t[7]);
  assign t[18] = t[5] ^ t[7];
  assign t[19] = t[10] ^ t[20];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = t[28] ^ x[2];
  assign t[25] = t[29] ^ x[5];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = t[31] ^ x[11];
  assign t[28] = (t[32] & ~t[33]);
  assign t[29] = (t[34] & ~t[35]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[36] & ~t[37]);
  assign t[31] = (t[38] & ~t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[1];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[4];
  assign t[36] = t[44] ^ x[8];
  assign t[37] = t[45] ^ x[7];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[10];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[4] = t[9] & t[10];
  assign t[5] = t[20] ^ t[8];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[21] ^ t[20];
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind169(x, y);
 input [11:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[7] ^ t[23];
  assign t[11] = t[13] ^ t[4];
  assign t[12] = t[14] & t[15];
  assign t[13] = t[16] & t[17];
  assign t[14] = ~(t[13] ^ t[18]);
  assign t[15] = t[3] ^ t[19];
  assign t[16] = ~(t[19]);
  assign t[17] = ~(t[7]);
  assign t[18] = t[5] ^ t[7];
  assign t[19] = t[10] ^ t[20];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = t[28] ^ x[2];
  assign t[25] = t[29] ^ x[5];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = t[31] ^ x[11];
  assign t[28] = (t[32] & ~t[33]);
  assign t[29] = (t[34] & ~t[35]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[36] & ~t[37]);
  assign t[31] = (t[38] & ~t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[1];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[4];
  assign t[36] = t[44] ^ x[8];
  assign t[37] = t[45] ^ x[7];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[10];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[4] = t[9] & t[10];
  assign t[5] = t[20] ^ t[8];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[21] ^ t[20];
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind170(x, y);
 input [11:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[24] ^ t[22];
  assign t[12] = ~(t[22]);
  assign t[13] = t[11] ^ t[25];
  assign t[14] = ~(t[7] ^ t[16]);
  assign t[15] = t[17] ^ t[13];
  assign t[16] = t[18] ^ t[6];
  assign t[17] = t[22] ^ t[9];
  assign t[18] = t[19] & t[20];
  assign t[19] = ~(t[21]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11]);
  assign t[21] = t[13] ^ t[22];
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34] & ~t[35]);
  assign t[31] = (t[36] & ~t[37]);
  assign t[32] = (t[38] & ~t[39]);
  assign t[33] = (t[40] & ~t[41]);
  assign t[34] = t[42] ^ x[2];
  assign t[35] = t[43] ^ x[1];
  assign t[36] = t[44] ^ x[5];
  assign t[37] = t[45] ^ x[4];
  assign t[38] = t[46] ^ x[8];
  assign t[39] = t[47] ^ x[7];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[11];
  assign t[41] = t[49] ^ x[10];
  assign t[42] = (x[0]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[3]);
  assign t[46] = (x[6]);
  assign t[47] = (x[6]);
  assign t[48] = (x[9]);
  assign t[49] = (x[9]);
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[11] ^ t[9];
  assign t[6] = t[12] & t[13];
  assign t[7] = t[11] ^ t[22];
  assign t[8] = t[14] & t[15];
  assign t[9] = ~(t[23]);
  assign y = (t[0]);
endmodule

module R2ind171(x, y);
 input [11:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[24] ^ t[22];
  assign t[12] = ~(t[22]);
  assign t[13] = t[11] ^ t[25];
  assign t[14] = ~(t[7] ^ t[16]);
  assign t[15] = t[17] ^ t[13];
  assign t[16] = t[18] ^ t[6];
  assign t[17] = t[22] ^ t[9];
  assign t[18] = t[19] & t[20];
  assign t[19] = ~(t[21]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11]);
  assign t[21] = t[13] ^ t[22];
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34] & ~t[35]);
  assign t[31] = (t[36] & ~t[37]);
  assign t[32] = (t[38] & ~t[39]);
  assign t[33] = (t[40] & ~t[41]);
  assign t[34] = t[42] ^ x[2];
  assign t[35] = t[43] ^ x[1];
  assign t[36] = t[44] ^ x[5];
  assign t[37] = t[45] ^ x[4];
  assign t[38] = t[46] ^ x[8];
  assign t[39] = t[47] ^ x[7];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[11];
  assign t[41] = t[49] ^ x[10];
  assign t[42] = (x[0]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[3]);
  assign t[46] = (x[6]);
  assign t[47] = (x[6]);
  assign t[48] = (x[9]);
  assign t[49] = (x[9]);
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[11] ^ t[9];
  assign t[6] = t[12] & t[13];
  assign t[7] = t[11] ^ t[22];
  assign t[8] = t[14] & t[15];
  assign t[9] = ~(t[23]);
  assign y = (t[0]);
endmodule

module R2ind172(x, y);
 input [11:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[15] ^ t[29];
  assign t[12] = t[20] & t[21];
  assign t[13] = ~(t[30]);
  assign t[14] = t[18] ^ t[12];
  assign t[15] = t[31] ^ t[29];
  assign t[16] = ~(t[29]);
  assign t[17] = t[15] ^ t[32];
  assign t[18] = t[22] ^ t[8];
  assign t[19] = t[23] & t[24];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11] ^ t[18]);
  assign t[21] = t[9] ^ t[17];
  assign t[22] = t[25] & t[26];
  assign t[23] = ~(t[22] ^ t[27]);
  assign t[24] = t[7] ^ t[28];
  assign t[25] = ~(t[28]);
  assign t[26] = ~(t[15]);
  assign t[27] = t[9] ^ t[15];
  assign t[28] = t[17] ^ t[29];
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = (t[35]);
  assign t[32] = (t[36]);
  assign t[33] = t[37] ^ x[2];
  assign t[34] = t[38] ^ x[5];
  assign t[35] = t[39] ^ x[8];
  assign t[36] = t[40] ^ x[11];
  assign t[37] = (t[41] & ~t[42]);
  assign t[38] = (t[43] & ~t[44]);
  assign t[39] = (t[45] & ~t[46]);
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (t[47] & ~t[48]);
  assign t[41] = t[49] ^ x[2];
  assign t[42] = t[50] ^ x[1];
  assign t[43] = t[51] ^ x[5];
  assign t[44] = t[52] ^ x[4];
  assign t[45] = t[53] ^ x[8];
  assign t[46] = t[54] ^ x[7];
  assign t[47] = t[55] ^ x[11];
  assign t[48] = t[56] ^ x[10];
  assign t[49] = (x[0]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[0]);
  assign t[51] = (x[3]);
  assign t[52] = (x[3]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[9]);
  assign t[56] = (x[9]);
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[15] ^ t[13];
  assign t[8] = t[16] & t[17];
  assign t[9] = t[29] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind173(x, y);
 input [11:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[15] ^ t[29];
  assign t[12] = t[20] & t[21];
  assign t[13] = ~(t[30]);
  assign t[14] = t[18] ^ t[12];
  assign t[15] = t[31] ^ t[29];
  assign t[16] = ~(t[29]);
  assign t[17] = t[15] ^ t[32];
  assign t[18] = t[22] ^ t[8];
  assign t[19] = t[23] & t[24];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11] ^ t[18]);
  assign t[21] = t[9] ^ t[17];
  assign t[22] = t[25] & t[26];
  assign t[23] = ~(t[22] ^ t[27]);
  assign t[24] = t[7] ^ t[28];
  assign t[25] = ~(t[28]);
  assign t[26] = ~(t[15]);
  assign t[27] = t[9] ^ t[15];
  assign t[28] = t[17] ^ t[29];
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = (t[35]);
  assign t[32] = (t[36]);
  assign t[33] = t[37] ^ x[2];
  assign t[34] = t[38] ^ x[5];
  assign t[35] = t[39] ^ x[8];
  assign t[36] = t[40] ^ x[11];
  assign t[37] = (t[41] & ~t[42]);
  assign t[38] = (t[43] & ~t[44]);
  assign t[39] = (t[45] & ~t[46]);
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (t[47] & ~t[48]);
  assign t[41] = t[49] ^ x[2];
  assign t[42] = t[50] ^ x[1];
  assign t[43] = t[51] ^ x[5];
  assign t[44] = t[52] ^ x[4];
  assign t[45] = t[53] ^ x[8];
  assign t[46] = t[54] ^ x[7];
  assign t[47] = t[55] ^ x[11];
  assign t[48] = t[56] ^ x[10];
  assign t[49] = (x[0]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[0]);
  assign t[51] = (x[3]);
  assign t[52] = (x[3]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[9]);
  assign t[56] = (x[9]);
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[15] ^ t[13];
  assign t[8] = t[16] & t[17];
  assign t[9] = t[29] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind174(x, y);
 input [11:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] ^ t[16];
  assign t[11] = t[17] ^ t[8];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[29] ^ t[28];
  assign t[14] = ~(t[28]);
  assign t[15] = t[13] ^ t[30];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[22] & t[23];
  assign t[18] = ~(t[24] ^ t[11]);
  assign t[19] = t[9] ^ t[15];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[17] ^ t[25]);
  assign t[21] = t[7] ^ t[26];
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[13]);
  assign t[24] = t[13] ^ t[28];
  assign t[25] = t[9] ^ t[13];
  assign t[26] = t[15] ^ t[28];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[2];
  assign t[32] = t[36] ^ x[5];
  assign t[33] = t[37] ^ x[8];
  assign t[34] = t[38] ^ x[11];
  assign t[35] = (t[39] & ~t[40]);
  assign t[36] = (t[41] & ~t[42]);
  assign t[37] = (t[43] & ~t[44]);
  assign t[38] = (t[45] & ~t[46]);
  assign t[39] = t[47] ^ x[2];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[1];
  assign t[41] = t[49] ^ x[5];
  assign t[42] = t[50] ^ x[4];
  assign t[43] = t[51] ^ x[8];
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[11];
  assign t[46] = t[54] ^ x[10];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[5] = ~(t[27]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[13] ^ t[5];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[28] ^ t[5];
  assign y = (t[0]);
endmodule

module R2ind175(x, y);
 input [11:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] ^ t[16];
  assign t[11] = t[17] ^ t[8];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[29] ^ t[28];
  assign t[14] = ~(t[28]);
  assign t[15] = t[13] ^ t[30];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[22] & t[23];
  assign t[18] = ~(t[24] ^ t[11]);
  assign t[19] = t[9] ^ t[15];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[17] ^ t[25]);
  assign t[21] = t[7] ^ t[26];
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[13]);
  assign t[24] = t[13] ^ t[28];
  assign t[25] = t[9] ^ t[13];
  assign t[26] = t[15] ^ t[28];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[2];
  assign t[32] = t[36] ^ x[5];
  assign t[33] = t[37] ^ x[8];
  assign t[34] = t[38] ^ x[11];
  assign t[35] = (t[39] & ~t[40]);
  assign t[36] = (t[41] & ~t[42]);
  assign t[37] = (t[43] & ~t[44]);
  assign t[38] = (t[45] & ~t[46]);
  assign t[39] = t[47] ^ x[2];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[1];
  assign t[41] = t[49] ^ x[5];
  assign t[42] = t[50] ^ x[4];
  assign t[43] = t[51] ^ x[8];
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[11];
  assign t[46] = t[54] ^ x[10];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[5] = ~(t[27]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[13] ^ t[5];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[28] ^ t[5];
  assign y = (t[0]);
endmodule

module R2ind176(x, y);
 input [11:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[7] ^ t[23];
  assign t[11] = t[13] ^ t[4];
  assign t[12] = t[14] & t[15];
  assign t[13] = t[16] & t[17];
  assign t[14] = ~(t[13] ^ t[18]);
  assign t[15] = t[3] ^ t[19];
  assign t[16] = ~(t[19]);
  assign t[17] = ~(t[7]);
  assign t[18] = t[5] ^ t[7];
  assign t[19] = t[10] ^ t[20];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = t[28] ^ x[2];
  assign t[25] = t[29] ^ x[5];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = t[31] ^ x[11];
  assign t[28] = (t[32] & ~t[33]);
  assign t[29] = (t[34] & ~t[35]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[36] & ~t[37]);
  assign t[31] = (t[38] & ~t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[1];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[4];
  assign t[36] = t[44] ^ x[8];
  assign t[37] = t[45] ^ x[7];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[10];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[4] = t[9] & t[10];
  assign t[5] = t[20] ^ t[8];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[21] ^ t[20];
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind177(x, y);
 input [11:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[7] ^ t[23];
  assign t[11] = t[13] ^ t[4];
  assign t[12] = t[14] & t[15];
  assign t[13] = t[16] & t[17];
  assign t[14] = ~(t[13] ^ t[18]);
  assign t[15] = t[3] ^ t[19];
  assign t[16] = ~(t[19]);
  assign t[17] = ~(t[7]);
  assign t[18] = t[5] ^ t[7];
  assign t[19] = t[10] ^ t[20];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = t[28] ^ x[2];
  assign t[25] = t[29] ^ x[5];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = t[31] ^ x[11];
  assign t[28] = (t[32] & ~t[33]);
  assign t[29] = (t[34] & ~t[35]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[36] & ~t[37]);
  assign t[31] = (t[38] & ~t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[1];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[4];
  assign t[36] = t[44] ^ x[8];
  assign t[37] = t[45] ^ x[7];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[10];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[4] = t[9] & t[10];
  assign t[5] = t[20] ^ t[8];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[21] ^ t[20];
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind178(x, y);
 input [11:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[24] ^ t[22];
  assign t[12] = ~(t[22]);
  assign t[13] = t[11] ^ t[25];
  assign t[14] = ~(t[7] ^ t[16]);
  assign t[15] = t[17] ^ t[13];
  assign t[16] = t[18] ^ t[6];
  assign t[17] = t[22] ^ t[9];
  assign t[18] = t[19] & t[20];
  assign t[19] = ~(t[21]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11]);
  assign t[21] = t[13] ^ t[22];
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34] & ~t[35]);
  assign t[31] = (t[36] & ~t[37]);
  assign t[32] = (t[38] & ~t[39]);
  assign t[33] = (t[40] & ~t[41]);
  assign t[34] = t[42] ^ x[2];
  assign t[35] = t[43] ^ x[1];
  assign t[36] = t[44] ^ x[5];
  assign t[37] = t[45] ^ x[4];
  assign t[38] = t[46] ^ x[8];
  assign t[39] = t[47] ^ x[7];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[11];
  assign t[41] = t[49] ^ x[10];
  assign t[42] = (x[0]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[3]);
  assign t[46] = (x[6]);
  assign t[47] = (x[6]);
  assign t[48] = (x[9]);
  assign t[49] = (x[9]);
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[11] ^ t[9];
  assign t[6] = t[12] & t[13];
  assign t[7] = t[11] ^ t[22];
  assign t[8] = t[14] & t[15];
  assign t[9] = ~(t[23]);
  assign y = (t[0]);
endmodule

module R2ind179(x, y);
 input [11:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[24] ^ t[22];
  assign t[12] = ~(t[22]);
  assign t[13] = t[11] ^ t[25];
  assign t[14] = ~(t[7] ^ t[16]);
  assign t[15] = t[17] ^ t[13];
  assign t[16] = t[18] ^ t[6];
  assign t[17] = t[22] ^ t[9];
  assign t[18] = t[19] & t[20];
  assign t[19] = ~(t[21]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11]);
  assign t[21] = t[13] ^ t[22];
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34] & ~t[35]);
  assign t[31] = (t[36] & ~t[37]);
  assign t[32] = (t[38] & ~t[39]);
  assign t[33] = (t[40] & ~t[41]);
  assign t[34] = t[42] ^ x[2];
  assign t[35] = t[43] ^ x[1];
  assign t[36] = t[44] ^ x[5];
  assign t[37] = t[45] ^ x[4];
  assign t[38] = t[46] ^ x[8];
  assign t[39] = t[47] ^ x[7];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[11];
  assign t[41] = t[49] ^ x[10];
  assign t[42] = (x[0]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[3]);
  assign t[46] = (x[6]);
  assign t[47] = (x[6]);
  assign t[48] = (x[9]);
  assign t[49] = (x[9]);
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[11] ^ t[9];
  assign t[6] = t[12] & t[13];
  assign t[7] = t[11] ^ t[22];
  assign t[8] = t[14] & t[15];
  assign t[9] = ~(t[23]);
  assign y = (t[0]);
endmodule

module R2ind180(x, y);
 input [11:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[15] ^ t[29];
  assign t[12] = t[20] & t[21];
  assign t[13] = ~(t[30]);
  assign t[14] = t[18] ^ t[12];
  assign t[15] = t[31] ^ t[29];
  assign t[16] = ~(t[29]);
  assign t[17] = t[15] ^ t[32];
  assign t[18] = t[22] ^ t[8];
  assign t[19] = t[23] & t[24];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11] ^ t[18]);
  assign t[21] = t[9] ^ t[17];
  assign t[22] = t[25] & t[26];
  assign t[23] = ~(t[22] ^ t[27]);
  assign t[24] = t[7] ^ t[28];
  assign t[25] = ~(t[28]);
  assign t[26] = ~(t[15]);
  assign t[27] = t[9] ^ t[15];
  assign t[28] = t[17] ^ t[29];
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = (t[35]);
  assign t[32] = (t[36]);
  assign t[33] = t[37] ^ x[2];
  assign t[34] = t[38] ^ x[5];
  assign t[35] = t[39] ^ x[8];
  assign t[36] = t[40] ^ x[11];
  assign t[37] = (t[41] & ~t[42]);
  assign t[38] = (t[43] & ~t[44]);
  assign t[39] = (t[45] & ~t[46]);
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (t[47] & ~t[48]);
  assign t[41] = t[49] ^ x[2];
  assign t[42] = t[50] ^ x[1];
  assign t[43] = t[51] ^ x[5];
  assign t[44] = t[52] ^ x[4];
  assign t[45] = t[53] ^ x[8];
  assign t[46] = t[54] ^ x[7];
  assign t[47] = t[55] ^ x[11];
  assign t[48] = t[56] ^ x[10];
  assign t[49] = (x[0]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[0]);
  assign t[51] = (x[3]);
  assign t[52] = (x[3]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[9]);
  assign t[56] = (x[9]);
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[15] ^ t[13];
  assign t[8] = t[16] & t[17];
  assign t[9] = t[29] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind181(x, y);
 input [11:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[15] ^ t[29];
  assign t[12] = t[20] & t[21];
  assign t[13] = ~(t[30]);
  assign t[14] = t[18] ^ t[12];
  assign t[15] = t[31] ^ t[29];
  assign t[16] = ~(t[29]);
  assign t[17] = t[15] ^ t[32];
  assign t[18] = t[22] ^ t[8];
  assign t[19] = t[23] & t[24];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11] ^ t[18]);
  assign t[21] = t[9] ^ t[17];
  assign t[22] = t[25] & t[26];
  assign t[23] = ~(t[22] ^ t[27]);
  assign t[24] = t[7] ^ t[28];
  assign t[25] = ~(t[28]);
  assign t[26] = ~(t[15]);
  assign t[27] = t[9] ^ t[15];
  assign t[28] = t[17] ^ t[29];
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = (t[35]);
  assign t[32] = (t[36]);
  assign t[33] = t[37] ^ x[2];
  assign t[34] = t[38] ^ x[5];
  assign t[35] = t[39] ^ x[8];
  assign t[36] = t[40] ^ x[11];
  assign t[37] = (t[41] & ~t[42]);
  assign t[38] = (t[43] & ~t[44]);
  assign t[39] = (t[45] & ~t[46]);
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (t[47] & ~t[48]);
  assign t[41] = t[49] ^ x[2];
  assign t[42] = t[50] ^ x[1];
  assign t[43] = t[51] ^ x[5];
  assign t[44] = t[52] ^ x[4];
  assign t[45] = t[53] ^ x[8];
  assign t[46] = t[54] ^ x[7];
  assign t[47] = t[55] ^ x[11];
  assign t[48] = t[56] ^ x[10];
  assign t[49] = (x[0]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[0]);
  assign t[51] = (x[3]);
  assign t[52] = (x[3]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[9]);
  assign t[56] = (x[9]);
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[15] ^ t[13];
  assign t[8] = t[16] & t[17];
  assign t[9] = t[29] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind182(x, y);
 input [11:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] ^ t[16];
  assign t[11] = t[17] ^ t[8];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[29] ^ t[28];
  assign t[14] = ~(t[28]);
  assign t[15] = t[13] ^ t[30];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[22] & t[23];
  assign t[18] = ~(t[24] ^ t[11]);
  assign t[19] = t[9] ^ t[15];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[17] ^ t[25]);
  assign t[21] = t[7] ^ t[26];
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[13]);
  assign t[24] = t[13] ^ t[28];
  assign t[25] = t[9] ^ t[13];
  assign t[26] = t[15] ^ t[28];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[2];
  assign t[32] = t[36] ^ x[5];
  assign t[33] = t[37] ^ x[8];
  assign t[34] = t[38] ^ x[11];
  assign t[35] = (t[39] & ~t[40]);
  assign t[36] = (t[41] & ~t[42]);
  assign t[37] = (t[43] & ~t[44]);
  assign t[38] = (t[45] & ~t[46]);
  assign t[39] = t[47] ^ x[2];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[1];
  assign t[41] = t[49] ^ x[5];
  assign t[42] = t[50] ^ x[4];
  assign t[43] = t[51] ^ x[8];
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[11];
  assign t[46] = t[54] ^ x[10];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[5] = ~(t[27]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[13] ^ t[5];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[28] ^ t[5];
  assign y = (t[0]);
endmodule

module R2ind183(x, y);
 input [11:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] ^ t[16];
  assign t[11] = t[17] ^ t[8];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[29] ^ t[28];
  assign t[14] = ~(t[28]);
  assign t[15] = t[13] ^ t[30];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[22] & t[23];
  assign t[18] = ~(t[24] ^ t[11]);
  assign t[19] = t[9] ^ t[15];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[17] ^ t[25]);
  assign t[21] = t[7] ^ t[26];
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[13]);
  assign t[24] = t[13] ^ t[28];
  assign t[25] = t[9] ^ t[13];
  assign t[26] = t[15] ^ t[28];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[2];
  assign t[32] = t[36] ^ x[5];
  assign t[33] = t[37] ^ x[8];
  assign t[34] = t[38] ^ x[11];
  assign t[35] = (t[39] & ~t[40]);
  assign t[36] = (t[41] & ~t[42]);
  assign t[37] = (t[43] & ~t[44]);
  assign t[38] = (t[45] & ~t[46]);
  assign t[39] = t[47] ^ x[2];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[1];
  assign t[41] = t[49] ^ x[5];
  assign t[42] = t[50] ^ x[4];
  assign t[43] = t[51] ^ x[8];
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[11];
  assign t[46] = t[54] ^ x[10];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[5] = ~(t[27]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[13] ^ t[5];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[28] ^ t[5];
  assign y = (t[0]);
endmodule

module R2ind184(x, y);
 input [11:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[7] ^ t[23];
  assign t[11] = t[13] ^ t[4];
  assign t[12] = t[14] & t[15];
  assign t[13] = t[16] & t[17];
  assign t[14] = ~(t[13] ^ t[18]);
  assign t[15] = t[3] ^ t[19];
  assign t[16] = ~(t[19]);
  assign t[17] = ~(t[7]);
  assign t[18] = t[5] ^ t[7];
  assign t[19] = t[10] ^ t[20];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = t[28] ^ x[2];
  assign t[25] = t[29] ^ x[5];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = t[31] ^ x[11];
  assign t[28] = (t[32] & ~t[33]);
  assign t[29] = (t[34] & ~t[35]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[36] & ~t[37]);
  assign t[31] = (t[38] & ~t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[1];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[4];
  assign t[36] = t[44] ^ x[8];
  assign t[37] = t[45] ^ x[7];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[10];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[4] = t[9] & t[10];
  assign t[5] = t[20] ^ t[8];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[21] ^ t[20];
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind185(x, y);
 input [11:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[7] ^ t[23];
  assign t[11] = t[13] ^ t[4];
  assign t[12] = t[14] & t[15];
  assign t[13] = t[16] & t[17];
  assign t[14] = ~(t[13] ^ t[18]);
  assign t[15] = t[3] ^ t[19];
  assign t[16] = ~(t[19]);
  assign t[17] = ~(t[7]);
  assign t[18] = t[5] ^ t[7];
  assign t[19] = t[10] ^ t[20];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = t[28] ^ x[2];
  assign t[25] = t[29] ^ x[5];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = t[31] ^ x[11];
  assign t[28] = (t[32] & ~t[33]);
  assign t[29] = (t[34] & ~t[35]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[36] & ~t[37]);
  assign t[31] = (t[38] & ~t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[1];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[4];
  assign t[36] = t[44] ^ x[8];
  assign t[37] = t[45] ^ x[7];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[10];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[4] = t[9] & t[10];
  assign t[5] = t[20] ^ t[8];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[21] ^ t[20];
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind186(x, y);
 input [11:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[24] ^ t[22];
  assign t[12] = ~(t[22]);
  assign t[13] = t[11] ^ t[25];
  assign t[14] = ~(t[7] ^ t[16]);
  assign t[15] = t[17] ^ t[13];
  assign t[16] = t[18] ^ t[6];
  assign t[17] = t[22] ^ t[9];
  assign t[18] = t[19] & t[20];
  assign t[19] = ~(t[21]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11]);
  assign t[21] = t[13] ^ t[22];
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34] & ~t[35]);
  assign t[31] = (t[36] & ~t[37]);
  assign t[32] = (t[38] & ~t[39]);
  assign t[33] = (t[40] & ~t[41]);
  assign t[34] = t[42] ^ x[2];
  assign t[35] = t[43] ^ x[1];
  assign t[36] = t[44] ^ x[5];
  assign t[37] = t[45] ^ x[4];
  assign t[38] = t[46] ^ x[8];
  assign t[39] = t[47] ^ x[7];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[11];
  assign t[41] = t[49] ^ x[10];
  assign t[42] = (x[0]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[3]);
  assign t[46] = (x[6]);
  assign t[47] = (x[6]);
  assign t[48] = (x[9]);
  assign t[49] = (x[9]);
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[11] ^ t[9];
  assign t[6] = t[12] & t[13];
  assign t[7] = t[11] ^ t[22];
  assign t[8] = t[14] & t[15];
  assign t[9] = ~(t[23]);
  assign y = (t[0]);
endmodule

module R2ind187(x, y);
 input [11:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[24] ^ t[22];
  assign t[12] = ~(t[22]);
  assign t[13] = t[11] ^ t[25];
  assign t[14] = ~(t[7] ^ t[16]);
  assign t[15] = t[17] ^ t[13];
  assign t[16] = t[18] ^ t[6];
  assign t[17] = t[22] ^ t[9];
  assign t[18] = t[19] & t[20];
  assign t[19] = ~(t[21]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11]);
  assign t[21] = t[13] ^ t[22];
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34] & ~t[35]);
  assign t[31] = (t[36] & ~t[37]);
  assign t[32] = (t[38] & ~t[39]);
  assign t[33] = (t[40] & ~t[41]);
  assign t[34] = t[42] ^ x[2];
  assign t[35] = t[43] ^ x[1];
  assign t[36] = t[44] ^ x[5];
  assign t[37] = t[45] ^ x[4];
  assign t[38] = t[46] ^ x[8];
  assign t[39] = t[47] ^ x[7];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[11];
  assign t[41] = t[49] ^ x[10];
  assign t[42] = (x[0]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[3]);
  assign t[46] = (x[6]);
  assign t[47] = (x[6]);
  assign t[48] = (x[9]);
  assign t[49] = (x[9]);
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[11] ^ t[9];
  assign t[6] = t[12] & t[13];
  assign t[7] = t[11] ^ t[22];
  assign t[8] = t[14] & t[15];
  assign t[9] = ~(t[23]);
  assign y = (t[0]);
endmodule

module R2ind188(x, y);
 input [11:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[15] ^ t[29];
  assign t[12] = t[20] & t[21];
  assign t[13] = ~(t[30]);
  assign t[14] = t[18] ^ t[12];
  assign t[15] = t[31] ^ t[29];
  assign t[16] = ~(t[29]);
  assign t[17] = t[15] ^ t[32];
  assign t[18] = t[22] ^ t[8];
  assign t[19] = t[23] & t[24];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11] ^ t[18]);
  assign t[21] = t[9] ^ t[17];
  assign t[22] = t[25] & t[26];
  assign t[23] = ~(t[22] ^ t[27]);
  assign t[24] = t[7] ^ t[28];
  assign t[25] = ~(t[28]);
  assign t[26] = ~(t[15]);
  assign t[27] = t[9] ^ t[15];
  assign t[28] = t[17] ^ t[29];
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = (t[35]);
  assign t[32] = (t[36]);
  assign t[33] = t[37] ^ x[2];
  assign t[34] = t[38] ^ x[5];
  assign t[35] = t[39] ^ x[8];
  assign t[36] = t[40] ^ x[11];
  assign t[37] = (t[41] & ~t[42]);
  assign t[38] = (t[43] & ~t[44]);
  assign t[39] = (t[45] & ~t[46]);
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (t[47] & ~t[48]);
  assign t[41] = t[49] ^ x[2];
  assign t[42] = t[50] ^ x[1];
  assign t[43] = t[51] ^ x[5];
  assign t[44] = t[52] ^ x[4];
  assign t[45] = t[53] ^ x[8];
  assign t[46] = t[54] ^ x[7];
  assign t[47] = t[55] ^ x[11];
  assign t[48] = t[56] ^ x[10];
  assign t[49] = (x[0]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[0]);
  assign t[51] = (x[3]);
  assign t[52] = (x[3]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[9]);
  assign t[56] = (x[9]);
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[15] ^ t[13];
  assign t[8] = t[16] & t[17];
  assign t[9] = t[29] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind189(x, y);
 input [11:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[15] ^ t[29];
  assign t[12] = t[20] & t[21];
  assign t[13] = ~(t[30]);
  assign t[14] = t[18] ^ t[12];
  assign t[15] = t[31] ^ t[29];
  assign t[16] = ~(t[29]);
  assign t[17] = t[15] ^ t[32];
  assign t[18] = t[22] ^ t[8];
  assign t[19] = t[23] & t[24];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11] ^ t[18]);
  assign t[21] = t[9] ^ t[17];
  assign t[22] = t[25] & t[26];
  assign t[23] = ~(t[22] ^ t[27]);
  assign t[24] = t[7] ^ t[28];
  assign t[25] = ~(t[28]);
  assign t[26] = ~(t[15]);
  assign t[27] = t[9] ^ t[15];
  assign t[28] = t[17] ^ t[29];
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = (t[35]);
  assign t[32] = (t[36]);
  assign t[33] = t[37] ^ x[2];
  assign t[34] = t[38] ^ x[5];
  assign t[35] = t[39] ^ x[8];
  assign t[36] = t[40] ^ x[11];
  assign t[37] = (t[41] & ~t[42]);
  assign t[38] = (t[43] & ~t[44]);
  assign t[39] = (t[45] & ~t[46]);
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (t[47] & ~t[48]);
  assign t[41] = t[49] ^ x[2];
  assign t[42] = t[50] ^ x[1];
  assign t[43] = t[51] ^ x[5];
  assign t[44] = t[52] ^ x[4];
  assign t[45] = t[53] ^ x[8];
  assign t[46] = t[54] ^ x[7];
  assign t[47] = t[55] ^ x[11];
  assign t[48] = t[56] ^ x[10];
  assign t[49] = (x[0]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[0]);
  assign t[51] = (x[3]);
  assign t[52] = (x[3]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[9]);
  assign t[56] = (x[9]);
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[15] ^ t[13];
  assign t[8] = t[16] & t[17];
  assign t[9] = t[29] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind190(x, y);
 input [11:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] ^ t[16];
  assign t[11] = t[17] ^ t[8];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[29] ^ t[28];
  assign t[14] = ~(t[28]);
  assign t[15] = t[13] ^ t[30];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[22] & t[23];
  assign t[18] = ~(t[24] ^ t[11]);
  assign t[19] = t[9] ^ t[15];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[17] ^ t[25]);
  assign t[21] = t[7] ^ t[26];
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[13]);
  assign t[24] = t[13] ^ t[28];
  assign t[25] = t[9] ^ t[13];
  assign t[26] = t[15] ^ t[28];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[2];
  assign t[32] = t[36] ^ x[5];
  assign t[33] = t[37] ^ x[8];
  assign t[34] = t[38] ^ x[11];
  assign t[35] = (t[39] & ~t[40]);
  assign t[36] = (t[41] & ~t[42]);
  assign t[37] = (t[43] & ~t[44]);
  assign t[38] = (t[45] & ~t[46]);
  assign t[39] = t[47] ^ x[2];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[1];
  assign t[41] = t[49] ^ x[5];
  assign t[42] = t[50] ^ x[4];
  assign t[43] = t[51] ^ x[8];
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[11];
  assign t[46] = t[54] ^ x[10];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[5] = ~(t[27]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[13] ^ t[5];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[28] ^ t[5];
  assign y = (t[0]);
endmodule

module R2ind191(x, y);
 input [11:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] ^ t[16];
  assign t[11] = t[17] ^ t[8];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[29] ^ t[28];
  assign t[14] = ~(t[28]);
  assign t[15] = t[13] ^ t[30];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[22] & t[23];
  assign t[18] = ~(t[24] ^ t[11]);
  assign t[19] = t[9] ^ t[15];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[17] ^ t[25]);
  assign t[21] = t[7] ^ t[26];
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[13]);
  assign t[24] = t[13] ^ t[28];
  assign t[25] = t[9] ^ t[13];
  assign t[26] = t[15] ^ t[28];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[2];
  assign t[32] = t[36] ^ x[5];
  assign t[33] = t[37] ^ x[8];
  assign t[34] = t[38] ^ x[11];
  assign t[35] = (t[39] & ~t[40]);
  assign t[36] = (t[41] & ~t[42]);
  assign t[37] = (t[43] & ~t[44]);
  assign t[38] = (t[45] & ~t[46]);
  assign t[39] = t[47] ^ x[2];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[1];
  assign t[41] = t[49] ^ x[5];
  assign t[42] = t[50] ^ x[4];
  assign t[43] = t[51] ^ x[8];
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[11];
  assign t[46] = t[54] ^ x[10];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[5] = ~(t[27]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[13] ^ t[5];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[28] ^ t[5];
  assign y = (t[0]);
endmodule

module R2ind192(x, y);
 input [11:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[7] ^ t[23];
  assign t[11] = t[13] ^ t[4];
  assign t[12] = t[14] & t[15];
  assign t[13] = t[16] & t[17];
  assign t[14] = ~(t[13] ^ t[18]);
  assign t[15] = t[3] ^ t[19];
  assign t[16] = ~(t[19]);
  assign t[17] = ~(t[7]);
  assign t[18] = t[5] ^ t[7];
  assign t[19] = t[10] ^ t[20];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = t[28] ^ x[2];
  assign t[25] = t[29] ^ x[5];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = t[31] ^ x[11];
  assign t[28] = (t[32] & ~t[33]);
  assign t[29] = (t[34] & ~t[35]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[36] & ~t[37]);
  assign t[31] = (t[38] & ~t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[1];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[4];
  assign t[36] = t[44] ^ x[8];
  assign t[37] = t[45] ^ x[7];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[10];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[4] = t[9] & t[10];
  assign t[5] = t[20] ^ t[8];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[21] ^ t[20];
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind193(x, y);
 input [11:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[7] ^ t[23];
  assign t[11] = t[13] ^ t[4];
  assign t[12] = t[14] & t[15];
  assign t[13] = t[16] & t[17];
  assign t[14] = ~(t[13] ^ t[18]);
  assign t[15] = t[3] ^ t[19];
  assign t[16] = ~(t[19]);
  assign t[17] = ~(t[7]);
  assign t[18] = t[5] ^ t[7];
  assign t[19] = t[10] ^ t[20];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = t[28] ^ x[2];
  assign t[25] = t[29] ^ x[5];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = t[31] ^ x[11];
  assign t[28] = (t[32] & ~t[33]);
  assign t[29] = (t[34] & ~t[35]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[36] & ~t[37]);
  assign t[31] = (t[38] & ~t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[1];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[4];
  assign t[36] = t[44] ^ x[8];
  assign t[37] = t[45] ^ x[7];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[10];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[4] = t[9] & t[10];
  assign t[5] = t[20] ^ t[8];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[21] ^ t[20];
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind194(x, y);
 input [11:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[24] ^ t[22];
  assign t[12] = ~(t[22]);
  assign t[13] = t[11] ^ t[25];
  assign t[14] = ~(t[7] ^ t[16]);
  assign t[15] = t[17] ^ t[13];
  assign t[16] = t[18] ^ t[6];
  assign t[17] = t[22] ^ t[9];
  assign t[18] = t[19] & t[20];
  assign t[19] = ~(t[21]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11]);
  assign t[21] = t[13] ^ t[22];
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34] & ~t[35]);
  assign t[31] = (t[36] & ~t[37]);
  assign t[32] = (t[38] & ~t[39]);
  assign t[33] = (t[40] & ~t[41]);
  assign t[34] = t[42] ^ x[2];
  assign t[35] = t[43] ^ x[1];
  assign t[36] = t[44] ^ x[5];
  assign t[37] = t[45] ^ x[4];
  assign t[38] = t[46] ^ x[8];
  assign t[39] = t[47] ^ x[7];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[11];
  assign t[41] = t[49] ^ x[10];
  assign t[42] = (x[0]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[3]);
  assign t[46] = (x[6]);
  assign t[47] = (x[6]);
  assign t[48] = (x[9]);
  assign t[49] = (x[9]);
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[11] ^ t[9];
  assign t[6] = t[12] & t[13];
  assign t[7] = t[11] ^ t[22];
  assign t[8] = t[14] & t[15];
  assign t[9] = ~(t[23]);
  assign y = (t[0]);
endmodule

module R2ind195(x, y);
 input [11:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[24] ^ t[22];
  assign t[12] = ~(t[22]);
  assign t[13] = t[11] ^ t[25];
  assign t[14] = ~(t[7] ^ t[16]);
  assign t[15] = t[17] ^ t[13];
  assign t[16] = t[18] ^ t[6];
  assign t[17] = t[22] ^ t[9];
  assign t[18] = t[19] & t[20];
  assign t[19] = ~(t[21]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11]);
  assign t[21] = t[13] ^ t[22];
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34] & ~t[35]);
  assign t[31] = (t[36] & ~t[37]);
  assign t[32] = (t[38] & ~t[39]);
  assign t[33] = (t[40] & ~t[41]);
  assign t[34] = t[42] ^ x[2];
  assign t[35] = t[43] ^ x[1];
  assign t[36] = t[44] ^ x[5];
  assign t[37] = t[45] ^ x[4];
  assign t[38] = t[46] ^ x[8];
  assign t[39] = t[47] ^ x[7];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[11];
  assign t[41] = t[49] ^ x[10];
  assign t[42] = (x[0]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[3]);
  assign t[46] = (x[6]);
  assign t[47] = (x[6]);
  assign t[48] = (x[9]);
  assign t[49] = (x[9]);
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[11] ^ t[9];
  assign t[6] = t[12] & t[13];
  assign t[7] = t[11] ^ t[22];
  assign t[8] = t[14] & t[15];
  assign t[9] = ~(t[23]);
  assign y = (t[0]);
endmodule

module R2ind196(x, y);
 input [11:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[15] ^ t[29];
  assign t[12] = t[20] & t[21];
  assign t[13] = ~(t[30]);
  assign t[14] = t[18] ^ t[12];
  assign t[15] = t[31] ^ t[29];
  assign t[16] = ~(t[29]);
  assign t[17] = t[15] ^ t[32];
  assign t[18] = t[22] ^ t[8];
  assign t[19] = t[23] & t[24];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11] ^ t[18]);
  assign t[21] = t[9] ^ t[17];
  assign t[22] = t[25] & t[26];
  assign t[23] = ~(t[22] ^ t[27]);
  assign t[24] = t[7] ^ t[28];
  assign t[25] = ~(t[28]);
  assign t[26] = ~(t[15]);
  assign t[27] = t[9] ^ t[15];
  assign t[28] = t[17] ^ t[29];
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = (t[35]);
  assign t[32] = (t[36]);
  assign t[33] = t[37] ^ x[2];
  assign t[34] = t[38] ^ x[5];
  assign t[35] = t[39] ^ x[8];
  assign t[36] = t[40] ^ x[11];
  assign t[37] = (t[41] & ~t[42]);
  assign t[38] = (t[43] & ~t[44]);
  assign t[39] = (t[45] & ~t[46]);
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (t[47] & ~t[48]);
  assign t[41] = t[49] ^ x[2];
  assign t[42] = t[50] ^ x[1];
  assign t[43] = t[51] ^ x[5];
  assign t[44] = t[52] ^ x[4];
  assign t[45] = t[53] ^ x[8];
  assign t[46] = t[54] ^ x[7];
  assign t[47] = t[55] ^ x[11];
  assign t[48] = t[56] ^ x[10];
  assign t[49] = (x[0]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[0]);
  assign t[51] = (x[3]);
  assign t[52] = (x[3]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[9]);
  assign t[56] = (x[9]);
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[15] ^ t[13];
  assign t[8] = t[16] & t[17];
  assign t[9] = t[29] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind197(x, y);
 input [11:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[15] ^ t[29];
  assign t[12] = t[20] & t[21];
  assign t[13] = ~(t[30]);
  assign t[14] = t[18] ^ t[12];
  assign t[15] = t[31] ^ t[29];
  assign t[16] = ~(t[29]);
  assign t[17] = t[15] ^ t[32];
  assign t[18] = t[22] ^ t[8];
  assign t[19] = t[23] & t[24];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11] ^ t[18]);
  assign t[21] = t[9] ^ t[17];
  assign t[22] = t[25] & t[26];
  assign t[23] = ~(t[22] ^ t[27]);
  assign t[24] = t[7] ^ t[28];
  assign t[25] = ~(t[28]);
  assign t[26] = ~(t[15]);
  assign t[27] = t[9] ^ t[15];
  assign t[28] = t[17] ^ t[29];
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = (t[35]);
  assign t[32] = (t[36]);
  assign t[33] = t[37] ^ x[2];
  assign t[34] = t[38] ^ x[5];
  assign t[35] = t[39] ^ x[8];
  assign t[36] = t[40] ^ x[11];
  assign t[37] = (t[41] & ~t[42]);
  assign t[38] = (t[43] & ~t[44]);
  assign t[39] = (t[45] & ~t[46]);
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (t[47] & ~t[48]);
  assign t[41] = t[49] ^ x[2];
  assign t[42] = t[50] ^ x[1];
  assign t[43] = t[51] ^ x[5];
  assign t[44] = t[52] ^ x[4];
  assign t[45] = t[53] ^ x[8];
  assign t[46] = t[54] ^ x[7];
  assign t[47] = t[55] ^ x[11];
  assign t[48] = t[56] ^ x[10];
  assign t[49] = (x[0]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[0]);
  assign t[51] = (x[3]);
  assign t[52] = (x[3]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[9]);
  assign t[56] = (x[9]);
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[15] ^ t[13];
  assign t[8] = t[16] & t[17];
  assign t[9] = t[29] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind198(x, y);
 input [11:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] ^ t[16];
  assign t[11] = t[17] ^ t[8];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[29] ^ t[28];
  assign t[14] = ~(t[28]);
  assign t[15] = t[13] ^ t[30];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[22] & t[23];
  assign t[18] = ~(t[24] ^ t[11]);
  assign t[19] = t[9] ^ t[15];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[17] ^ t[25]);
  assign t[21] = t[7] ^ t[26];
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[13]);
  assign t[24] = t[13] ^ t[28];
  assign t[25] = t[9] ^ t[13];
  assign t[26] = t[15] ^ t[28];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[2];
  assign t[32] = t[36] ^ x[5];
  assign t[33] = t[37] ^ x[8];
  assign t[34] = t[38] ^ x[11];
  assign t[35] = (t[39] & ~t[40]);
  assign t[36] = (t[41] & ~t[42]);
  assign t[37] = (t[43] & ~t[44]);
  assign t[38] = (t[45] & ~t[46]);
  assign t[39] = t[47] ^ x[2];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[1];
  assign t[41] = t[49] ^ x[5];
  assign t[42] = t[50] ^ x[4];
  assign t[43] = t[51] ^ x[8];
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[11];
  assign t[46] = t[54] ^ x[10];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[5] = ~(t[27]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[13] ^ t[5];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[28] ^ t[5];
  assign y = (t[0]);
endmodule

module R2ind199(x, y);
 input [11:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] ^ t[16];
  assign t[11] = t[17] ^ t[8];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[29] ^ t[28];
  assign t[14] = ~(t[28]);
  assign t[15] = t[13] ^ t[30];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[22] & t[23];
  assign t[18] = ~(t[24] ^ t[11]);
  assign t[19] = t[9] ^ t[15];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[17] ^ t[25]);
  assign t[21] = t[7] ^ t[26];
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[13]);
  assign t[24] = t[13] ^ t[28];
  assign t[25] = t[9] ^ t[13];
  assign t[26] = t[15] ^ t[28];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[2];
  assign t[32] = t[36] ^ x[5];
  assign t[33] = t[37] ^ x[8];
  assign t[34] = t[38] ^ x[11];
  assign t[35] = (t[39] & ~t[40]);
  assign t[36] = (t[41] & ~t[42]);
  assign t[37] = (t[43] & ~t[44]);
  assign t[38] = (t[45] & ~t[46]);
  assign t[39] = t[47] ^ x[2];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[1];
  assign t[41] = t[49] ^ x[5];
  assign t[42] = t[50] ^ x[4];
  assign t[43] = t[51] ^ x[8];
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[11];
  assign t[46] = t[54] ^ x[10];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[5] = ~(t[27]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[13] ^ t[5];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[28] ^ t[5];
  assign y = (t[0]);
endmodule

module R2ind200(x, y);
 input [11:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[7] ^ t[23];
  assign t[11] = t[13] ^ t[4];
  assign t[12] = t[14] & t[15];
  assign t[13] = t[16] & t[17];
  assign t[14] = ~(t[13] ^ t[18]);
  assign t[15] = t[3] ^ t[19];
  assign t[16] = ~(t[19]);
  assign t[17] = ~(t[7]);
  assign t[18] = t[5] ^ t[7];
  assign t[19] = t[10] ^ t[20];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = t[28] ^ x[2];
  assign t[25] = t[29] ^ x[5];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = t[31] ^ x[11];
  assign t[28] = (t[32] & ~t[33]);
  assign t[29] = (t[34] & ~t[35]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[36] & ~t[37]);
  assign t[31] = (t[38] & ~t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[1];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[4];
  assign t[36] = t[44] ^ x[8];
  assign t[37] = t[45] ^ x[7];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[10];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[4] = t[9] & t[10];
  assign t[5] = t[20] ^ t[8];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[21] ^ t[20];
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind201(x, y);
 input [11:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[7] ^ t[23];
  assign t[11] = t[13] ^ t[4];
  assign t[12] = t[14] & t[15];
  assign t[13] = t[16] & t[17];
  assign t[14] = ~(t[13] ^ t[18]);
  assign t[15] = t[3] ^ t[19];
  assign t[16] = ~(t[19]);
  assign t[17] = ~(t[7]);
  assign t[18] = t[5] ^ t[7];
  assign t[19] = t[10] ^ t[20];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = t[28] ^ x[2];
  assign t[25] = t[29] ^ x[5];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = t[31] ^ x[11];
  assign t[28] = (t[32] & ~t[33]);
  assign t[29] = (t[34] & ~t[35]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[36] & ~t[37]);
  assign t[31] = (t[38] & ~t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[1];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[4];
  assign t[36] = t[44] ^ x[8];
  assign t[37] = t[45] ^ x[7];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[10];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[4] = t[9] & t[10];
  assign t[5] = t[20] ^ t[8];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[21] ^ t[20];
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind202(x, y);
 input [11:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[24] ^ t[22];
  assign t[12] = ~(t[22]);
  assign t[13] = t[11] ^ t[25];
  assign t[14] = ~(t[7] ^ t[16]);
  assign t[15] = t[17] ^ t[13];
  assign t[16] = t[18] ^ t[6];
  assign t[17] = t[22] ^ t[9];
  assign t[18] = t[19] & t[20];
  assign t[19] = ~(t[21]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11]);
  assign t[21] = t[13] ^ t[22];
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34] & ~t[35]);
  assign t[31] = (t[36] & ~t[37]);
  assign t[32] = (t[38] & ~t[39]);
  assign t[33] = (t[40] & ~t[41]);
  assign t[34] = t[42] ^ x[2];
  assign t[35] = t[43] ^ x[1];
  assign t[36] = t[44] ^ x[5];
  assign t[37] = t[45] ^ x[4];
  assign t[38] = t[46] ^ x[8];
  assign t[39] = t[47] ^ x[7];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[11];
  assign t[41] = t[49] ^ x[10];
  assign t[42] = (x[0]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[3]);
  assign t[46] = (x[6]);
  assign t[47] = (x[6]);
  assign t[48] = (x[9]);
  assign t[49] = (x[9]);
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[11] ^ t[9];
  assign t[6] = t[12] & t[13];
  assign t[7] = t[11] ^ t[22];
  assign t[8] = t[14] & t[15];
  assign t[9] = ~(t[23]);
  assign y = (t[0]);
endmodule

module R2ind203(x, y);
 input [11:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[24] ^ t[22];
  assign t[12] = ~(t[22]);
  assign t[13] = t[11] ^ t[25];
  assign t[14] = ~(t[7] ^ t[16]);
  assign t[15] = t[17] ^ t[13];
  assign t[16] = t[18] ^ t[6];
  assign t[17] = t[22] ^ t[9];
  assign t[18] = t[19] & t[20];
  assign t[19] = ~(t[21]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11]);
  assign t[21] = t[13] ^ t[22];
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34] & ~t[35]);
  assign t[31] = (t[36] & ~t[37]);
  assign t[32] = (t[38] & ~t[39]);
  assign t[33] = (t[40] & ~t[41]);
  assign t[34] = t[42] ^ x[2];
  assign t[35] = t[43] ^ x[1];
  assign t[36] = t[44] ^ x[5];
  assign t[37] = t[45] ^ x[4];
  assign t[38] = t[46] ^ x[8];
  assign t[39] = t[47] ^ x[7];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[11];
  assign t[41] = t[49] ^ x[10];
  assign t[42] = (x[0]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[3]);
  assign t[46] = (x[6]);
  assign t[47] = (x[6]);
  assign t[48] = (x[9]);
  assign t[49] = (x[9]);
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[11] ^ t[9];
  assign t[6] = t[12] & t[13];
  assign t[7] = t[11] ^ t[22];
  assign t[8] = t[14] & t[15];
  assign t[9] = ~(t[23]);
  assign y = (t[0]);
endmodule

module R2ind204(x, y);
 input [11:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[15] ^ t[29];
  assign t[12] = t[20] & t[21];
  assign t[13] = ~(t[30]);
  assign t[14] = t[18] ^ t[12];
  assign t[15] = t[31] ^ t[29];
  assign t[16] = ~(t[29]);
  assign t[17] = t[15] ^ t[32];
  assign t[18] = t[22] ^ t[8];
  assign t[19] = t[23] & t[24];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11] ^ t[18]);
  assign t[21] = t[9] ^ t[17];
  assign t[22] = t[25] & t[26];
  assign t[23] = ~(t[22] ^ t[27]);
  assign t[24] = t[7] ^ t[28];
  assign t[25] = ~(t[28]);
  assign t[26] = ~(t[15]);
  assign t[27] = t[9] ^ t[15];
  assign t[28] = t[17] ^ t[29];
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = (t[35]);
  assign t[32] = (t[36]);
  assign t[33] = t[37] ^ x[2];
  assign t[34] = t[38] ^ x[5];
  assign t[35] = t[39] ^ x[8];
  assign t[36] = t[40] ^ x[11];
  assign t[37] = (t[41] & ~t[42]);
  assign t[38] = (t[43] & ~t[44]);
  assign t[39] = (t[45] & ~t[46]);
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (t[47] & ~t[48]);
  assign t[41] = t[49] ^ x[2];
  assign t[42] = t[50] ^ x[1];
  assign t[43] = t[51] ^ x[5];
  assign t[44] = t[52] ^ x[4];
  assign t[45] = t[53] ^ x[8];
  assign t[46] = t[54] ^ x[7];
  assign t[47] = t[55] ^ x[11];
  assign t[48] = t[56] ^ x[10];
  assign t[49] = (x[0]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[0]);
  assign t[51] = (x[3]);
  assign t[52] = (x[3]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[9]);
  assign t[56] = (x[9]);
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[15] ^ t[13];
  assign t[8] = t[16] & t[17];
  assign t[9] = t[29] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind205(x, y);
 input [11:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[15] ^ t[29];
  assign t[12] = t[20] & t[21];
  assign t[13] = ~(t[30]);
  assign t[14] = t[18] ^ t[12];
  assign t[15] = t[31] ^ t[29];
  assign t[16] = ~(t[29]);
  assign t[17] = t[15] ^ t[32];
  assign t[18] = t[22] ^ t[8];
  assign t[19] = t[23] & t[24];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11] ^ t[18]);
  assign t[21] = t[9] ^ t[17];
  assign t[22] = t[25] & t[26];
  assign t[23] = ~(t[22] ^ t[27]);
  assign t[24] = t[7] ^ t[28];
  assign t[25] = ~(t[28]);
  assign t[26] = ~(t[15]);
  assign t[27] = t[9] ^ t[15];
  assign t[28] = t[17] ^ t[29];
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = (t[35]);
  assign t[32] = (t[36]);
  assign t[33] = t[37] ^ x[2];
  assign t[34] = t[38] ^ x[5];
  assign t[35] = t[39] ^ x[8];
  assign t[36] = t[40] ^ x[11];
  assign t[37] = (t[41] & ~t[42]);
  assign t[38] = (t[43] & ~t[44]);
  assign t[39] = (t[45] & ~t[46]);
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (t[47] & ~t[48]);
  assign t[41] = t[49] ^ x[2];
  assign t[42] = t[50] ^ x[1];
  assign t[43] = t[51] ^ x[5];
  assign t[44] = t[52] ^ x[4];
  assign t[45] = t[53] ^ x[8];
  assign t[46] = t[54] ^ x[7];
  assign t[47] = t[55] ^ x[11];
  assign t[48] = t[56] ^ x[10];
  assign t[49] = (x[0]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[0]);
  assign t[51] = (x[3]);
  assign t[52] = (x[3]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[9]);
  assign t[56] = (x[9]);
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[15] ^ t[13];
  assign t[8] = t[16] & t[17];
  assign t[9] = t[29] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind206(x, y);
 input [11:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] ^ t[16];
  assign t[11] = t[17] ^ t[8];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[29] ^ t[28];
  assign t[14] = ~(t[28]);
  assign t[15] = t[13] ^ t[30];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[22] & t[23];
  assign t[18] = ~(t[24] ^ t[11]);
  assign t[19] = t[9] ^ t[15];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[17] ^ t[25]);
  assign t[21] = t[7] ^ t[26];
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[13]);
  assign t[24] = t[13] ^ t[28];
  assign t[25] = t[9] ^ t[13];
  assign t[26] = t[15] ^ t[28];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[2];
  assign t[32] = t[36] ^ x[5];
  assign t[33] = t[37] ^ x[8];
  assign t[34] = t[38] ^ x[11];
  assign t[35] = (t[39] & ~t[40]);
  assign t[36] = (t[41] & ~t[42]);
  assign t[37] = (t[43] & ~t[44]);
  assign t[38] = (t[45] & ~t[46]);
  assign t[39] = t[47] ^ x[2];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[1];
  assign t[41] = t[49] ^ x[5];
  assign t[42] = t[50] ^ x[4];
  assign t[43] = t[51] ^ x[8];
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[11];
  assign t[46] = t[54] ^ x[10];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[5] = ~(t[27]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[13] ^ t[5];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[28] ^ t[5];
  assign y = (t[0]);
endmodule

module R2ind207(x, y);
 input [11:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] ^ t[16];
  assign t[11] = t[17] ^ t[8];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[29] ^ t[28];
  assign t[14] = ~(t[28]);
  assign t[15] = t[13] ^ t[30];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[22] & t[23];
  assign t[18] = ~(t[24] ^ t[11]);
  assign t[19] = t[9] ^ t[15];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[17] ^ t[25]);
  assign t[21] = t[7] ^ t[26];
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[13]);
  assign t[24] = t[13] ^ t[28];
  assign t[25] = t[9] ^ t[13];
  assign t[26] = t[15] ^ t[28];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[2];
  assign t[32] = t[36] ^ x[5];
  assign t[33] = t[37] ^ x[8];
  assign t[34] = t[38] ^ x[11];
  assign t[35] = (t[39] & ~t[40]);
  assign t[36] = (t[41] & ~t[42]);
  assign t[37] = (t[43] & ~t[44]);
  assign t[38] = (t[45] & ~t[46]);
  assign t[39] = t[47] ^ x[2];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[1];
  assign t[41] = t[49] ^ x[5];
  assign t[42] = t[50] ^ x[4];
  assign t[43] = t[51] ^ x[8];
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[11];
  assign t[46] = t[54] ^ x[10];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[5] = ~(t[27]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[13] ^ t[5];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[28] ^ t[5];
  assign y = (t[0]);
endmodule

module R2ind208(x, y);
 input [11:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[7] ^ t[23];
  assign t[11] = t[13] ^ t[4];
  assign t[12] = t[14] & t[15];
  assign t[13] = t[16] & t[17];
  assign t[14] = ~(t[13] ^ t[18]);
  assign t[15] = t[3] ^ t[19];
  assign t[16] = ~(t[19]);
  assign t[17] = ~(t[7]);
  assign t[18] = t[5] ^ t[7];
  assign t[19] = t[10] ^ t[20];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = t[28] ^ x[2];
  assign t[25] = t[29] ^ x[5];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = t[31] ^ x[11];
  assign t[28] = (t[32] & ~t[33]);
  assign t[29] = (t[34] & ~t[35]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[36] & ~t[37]);
  assign t[31] = (t[38] & ~t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[1];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[4];
  assign t[36] = t[44] ^ x[8];
  assign t[37] = t[45] ^ x[7];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[10];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[4] = t[9] & t[10];
  assign t[5] = t[20] ^ t[8];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[21] ^ t[20];
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind209(x, y);
 input [11:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[7] ^ t[23];
  assign t[11] = t[13] ^ t[4];
  assign t[12] = t[14] & t[15];
  assign t[13] = t[16] & t[17];
  assign t[14] = ~(t[13] ^ t[18]);
  assign t[15] = t[3] ^ t[19];
  assign t[16] = ~(t[19]);
  assign t[17] = ~(t[7]);
  assign t[18] = t[5] ^ t[7];
  assign t[19] = t[10] ^ t[20];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = t[28] ^ x[2];
  assign t[25] = t[29] ^ x[5];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = t[31] ^ x[11];
  assign t[28] = (t[32] & ~t[33]);
  assign t[29] = (t[34] & ~t[35]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[36] & ~t[37]);
  assign t[31] = (t[38] & ~t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[1];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[4];
  assign t[36] = t[44] ^ x[8];
  assign t[37] = t[45] ^ x[7];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[10];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[4] = t[9] & t[10];
  assign t[5] = t[20] ^ t[8];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[21] ^ t[20];
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind210(x, y);
 input [11:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[24] ^ t[22];
  assign t[12] = ~(t[22]);
  assign t[13] = t[11] ^ t[25];
  assign t[14] = ~(t[7] ^ t[16]);
  assign t[15] = t[17] ^ t[13];
  assign t[16] = t[18] ^ t[6];
  assign t[17] = t[22] ^ t[9];
  assign t[18] = t[19] & t[20];
  assign t[19] = ~(t[21]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11]);
  assign t[21] = t[13] ^ t[22];
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34] & ~t[35]);
  assign t[31] = (t[36] & ~t[37]);
  assign t[32] = (t[38] & ~t[39]);
  assign t[33] = (t[40] & ~t[41]);
  assign t[34] = t[42] ^ x[2];
  assign t[35] = t[43] ^ x[1];
  assign t[36] = t[44] ^ x[5];
  assign t[37] = t[45] ^ x[4];
  assign t[38] = t[46] ^ x[8];
  assign t[39] = t[47] ^ x[7];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[11];
  assign t[41] = t[49] ^ x[10];
  assign t[42] = (x[0]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[3]);
  assign t[46] = (x[6]);
  assign t[47] = (x[6]);
  assign t[48] = (x[9]);
  assign t[49] = (x[9]);
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[11] ^ t[9];
  assign t[6] = t[12] & t[13];
  assign t[7] = t[11] ^ t[22];
  assign t[8] = t[14] & t[15];
  assign t[9] = ~(t[23]);
  assign y = (t[0]);
endmodule

module R2ind211(x, y);
 input [11:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[24] ^ t[22];
  assign t[12] = ~(t[22]);
  assign t[13] = t[11] ^ t[25];
  assign t[14] = ~(t[7] ^ t[16]);
  assign t[15] = t[17] ^ t[13];
  assign t[16] = t[18] ^ t[6];
  assign t[17] = t[22] ^ t[9];
  assign t[18] = t[19] & t[20];
  assign t[19] = ~(t[21]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11]);
  assign t[21] = t[13] ^ t[22];
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34] & ~t[35]);
  assign t[31] = (t[36] & ~t[37]);
  assign t[32] = (t[38] & ~t[39]);
  assign t[33] = (t[40] & ~t[41]);
  assign t[34] = t[42] ^ x[2];
  assign t[35] = t[43] ^ x[1];
  assign t[36] = t[44] ^ x[5];
  assign t[37] = t[45] ^ x[4];
  assign t[38] = t[46] ^ x[8];
  assign t[39] = t[47] ^ x[7];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[11];
  assign t[41] = t[49] ^ x[10];
  assign t[42] = (x[0]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[3]);
  assign t[46] = (x[6]);
  assign t[47] = (x[6]);
  assign t[48] = (x[9]);
  assign t[49] = (x[9]);
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[11] ^ t[9];
  assign t[6] = t[12] & t[13];
  assign t[7] = t[11] ^ t[22];
  assign t[8] = t[14] & t[15];
  assign t[9] = ~(t[23]);
  assign y = (t[0]);
endmodule

module R2ind212(x, y);
 input [11:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[15] ^ t[29];
  assign t[12] = t[20] & t[21];
  assign t[13] = ~(t[30]);
  assign t[14] = t[18] ^ t[12];
  assign t[15] = t[31] ^ t[29];
  assign t[16] = ~(t[29]);
  assign t[17] = t[15] ^ t[32];
  assign t[18] = t[22] ^ t[8];
  assign t[19] = t[23] & t[24];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11] ^ t[18]);
  assign t[21] = t[9] ^ t[17];
  assign t[22] = t[25] & t[26];
  assign t[23] = ~(t[22] ^ t[27]);
  assign t[24] = t[7] ^ t[28];
  assign t[25] = ~(t[28]);
  assign t[26] = ~(t[15]);
  assign t[27] = t[9] ^ t[15];
  assign t[28] = t[17] ^ t[29];
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = (t[35]);
  assign t[32] = (t[36]);
  assign t[33] = t[37] ^ x[2];
  assign t[34] = t[38] ^ x[5];
  assign t[35] = t[39] ^ x[8];
  assign t[36] = t[40] ^ x[11];
  assign t[37] = (t[41] & ~t[42]);
  assign t[38] = (t[43] & ~t[44]);
  assign t[39] = (t[45] & ~t[46]);
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (t[47] & ~t[48]);
  assign t[41] = t[49] ^ x[2];
  assign t[42] = t[50] ^ x[1];
  assign t[43] = t[51] ^ x[5];
  assign t[44] = t[52] ^ x[4];
  assign t[45] = t[53] ^ x[8];
  assign t[46] = t[54] ^ x[7];
  assign t[47] = t[55] ^ x[11];
  assign t[48] = t[56] ^ x[10];
  assign t[49] = (x[0]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[0]);
  assign t[51] = (x[3]);
  assign t[52] = (x[3]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[9]);
  assign t[56] = (x[9]);
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[15] ^ t[13];
  assign t[8] = t[16] & t[17];
  assign t[9] = t[29] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind213(x, y);
 input [11:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[15] ^ t[29];
  assign t[12] = t[20] & t[21];
  assign t[13] = ~(t[30]);
  assign t[14] = t[18] ^ t[12];
  assign t[15] = t[31] ^ t[29];
  assign t[16] = ~(t[29]);
  assign t[17] = t[15] ^ t[32];
  assign t[18] = t[22] ^ t[8];
  assign t[19] = t[23] & t[24];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11] ^ t[18]);
  assign t[21] = t[9] ^ t[17];
  assign t[22] = t[25] & t[26];
  assign t[23] = ~(t[22] ^ t[27]);
  assign t[24] = t[7] ^ t[28];
  assign t[25] = ~(t[28]);
  assign t[26] = ~(t[15]);
  assign t[27] = t[9] ^ t[15];
  assign t[28] = t[17] ^ t[29];
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = (t[35]);
  assign t[32] = (t[36]);
  assign t[33] = t[37] ^ x[2];
  assign t[34] = t[38] ^ x[5];
  assign t[35] = t[39] ^ x[8];
  assign t[36] = t[40] ^ x[11];
  assign t[37] = (t[41] & ~t[42]);
  assign t[38] = (t[43] & ~t[44]);
  assign t[39] = (t[45] & ~t[46]);
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (t[47] & ~t[48]);
  assign t[41] = t[49] ^ x[2];
  assign t[42] = t[50] ^ x[1];
  assign t[43] = t[51] ^ x[5];
  assign t[44] = t[52] ^ x[4];
  assign t[45] = t[53] ^ x[8];
  assign t[46] = t[54] ^ x[7];
  assign t[47] = t[55] ^ x[11];
  assign t[48] = t[56] ^ x[10];
  assign t[49] = (x[0]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[0]);
  assign t[51] = (x[3]);
  assign t[52] = (x[3]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[9]);
  assign t[56] = (x[9]);
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[15] ^ t[13];
  assign t[8] = t[16] & t[17];
  assign t[9] = t[29] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind214(x, y);
 input [11:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] ^ t[16];
  assign t[11] = t[17] ^ t[8];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[29] ^ t[28];
  assign t[14] = ~(t[28]);
  assign t[15] = t[13] ^ t[30];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[22] & t[23];
  assign t[18] = ~(t[24] ^ t[11]);
  assign t[19] = t[9] ^ t[15];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[17] ^ t[25]);
  assign t[21] = t[7] ^ t[26];
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[13]);
  assign t[24] = t[13] ^ t[28];
  assign t[25] = t[9] ^ t[13];
  assign t[26] = t[15] ^ t[28];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[2];
  assign t[32] = t[36] ^ x[5];
  assign t[33] = t[37] ^ x[8];
  assign t[34] = t[38] ^ x[11];
  assign t[35] = (t[39] & ~t[40]);
  assign t[36] = (t[41] & ~t[42]);
  assign t[37] = (t[43] & ~t[44]);
  assign t[38] = (t[45] & ~t[46]);
  assign t[39] = t[47] ^ x[2];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[1];
  assign t[41] = t[49] ^ x[5];
  assign t[42] = t[50] ^ x[4];
  assign t[43] = t[51] ^ x[8];
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[11];
  assign t[46] = t[54] ^ x[10];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[5] = ~(t[27]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[13] ^ t[5];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[28] ^ t[5];
  assign y = (t[0]);
endmodule

module R2ind215(x, y);
 input [11:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] ^ t[16];
  assign t[11] = t[17] ^ t[8];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[29] ^ t[28];
  assign t[14] = ~(t[28]);
  assign t[15] = t[13] ^ t[30];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[22] & t[23];
  assign t[18] = ~(t[24] ^ t[11]);
  assign t[19] = t[9] ^ t[15];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[17] ^ t[25]);
  assign t[21] = t[7] ^ t[26];
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[13]);
  assign t[24] = t[13] ^ t[28];
  assign t[25] = t[9] ^ t[13];
  assign t[26] = t[15] ^ t[28];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[2];
  assign t[32] = t[36] ^ x[5];
  assign t[33] = t[37] ^ x[8];
  assign t[34] = t[38] ^ x[11];
  assign t[35] = (t[39] & ~t[40]);
  assign t[36] = (t[41] & ~t[42]);
  assign t[37] = (t[43] & ~t[44]);
  assign t[38] = (t[45] & ~t[46]);
  assign t[39] = t[47] ^ x[2];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[1];
  assign t[41] = t[49] ^ x[5];
  assign t[42] = t[50] ^ x[4];
  assign t[43] = t[51] ^ x[8];
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[11];
  assign t[46] = t[54] ^ x[10];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[5] = ~(t[27]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[13] ^ t[5];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[28] ^ t[5];
  assign y = (t[0]);
endmodule

module R2ind216(x, y);
 input [11:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[7] ^ t[23];
  assign t[11] = t[13] ^ t[4];
  assign t[12] = t[14] & t[15];
  assign t[13] = t[16] & t[17];
  assign t[14] = ~(t[13] ^ t[18]);
  assign t[15] = t[3] ^ t[19];
  assign t[16] = ~(t[19]);
  assign t[17] = ~(t[7]);
  assign t[18] = t[5] ^ t[7];
  assign t[19] = t[10] ^ t[20];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = t[28] ^ x[2];
  assign t[25] = t[29] ^ x[5];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = t[31] ^ x[11];
  assign t[28] = (t[32] & ~t[33]);
  assign t[29] = (t[34] & ~t[35]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[36] & ~t[37]);
  assign t[31] = (t[38] & ~t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[1];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[4];
  assign t[36] = t[44] ^ x[8];
  assign t[37] = t[45] ^ x[7];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[10];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[4] = t[9] & t[10];
  assign t[5] = t[20] ^ t[8];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[21] ^ t[20];
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind217(x, y);
 input [11:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[7] ^ t[23];
  assign t[11] = t[13] ^ t[4];
  assign t[12] = t[14] & t[15];
  assign t[13] = t[16] & t[17];
  assign t[14] = ~(t[13] ^ t[18]);
  assign t[15] = t[3] ^ t[19];
  assign t[16] = ~(t[19]);
  assign t[17] = ~(t[7]);
  assign t[18] = t[5] ^ t[7];
  assign t[19] = t[10] ^ t[20];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = t[28] ^ x[2];
  assign t[25] = t[29] ^ x[5];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = t[31] ^ x[11];
  assign t[28] = (t[32] & ~t[33]);
  assign t[29] = (t[34] & ~t[35]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[36] & ~t[37]);
  assign t[31] = (t[38] & ~t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[1];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[4];
  assign t[36] = t[44] ^ x[8];
  assign t[37] = t[45] ^ x[7];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[10];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[4] = t[9] & t[10];
  assign t[5] = t[20] ^ t[8];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[21] ^ t[20];
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind218(x, y);
 input [11:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[24] ^ t[22];
  assign t[12] = ~(t[22]);
  assign t[13] = t[11] ^ t[25];
  assign t[14] = ~(t[7] ^ t[16]);
  assign t[15] = t[17] ^ t[13];
  assign t[16] = t[18] ^ t[6];
  assign t[17] = t[22] ^ t[9];
  assign t[18] = t[19] & t[20];
  assign t[19] = ~(t[21]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11]);
  assign t[21] = t[13] ^ t[22];
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34] & ~t[35]);
  assign t[31] = (t[36] & ~t[37]);
  assign t[32] = (t[38] & ~t[39]);
  assign t[33] = (t[40] & ~t[41]);
  assign t[34] = t[42] ^ x[2];
  assign t[35] = t[43] ^ x[1];
  assign t[36] = t[44] ^ x[5];
  assign t[37] = t[45] ^ x[4];
  assign t[38] = t[46] ^ x[8];
  assign t[39] = t[47] ^ x[7];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[11];
  assign t[41] = t[49] ^ x[10];
  assign t[42] = (x[0]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[3]);
  assign t[46] = (x[6]);
  assign t[47] = (x[6]);
  assign t[48] = (x[9]);
  assign t[49] = (x[9]);
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[11] ^ t[9];
  assign t[6] = t[12] & t[13];
  assign t[7] = t[11] ^ t[22];
  assign t[8] = t[14] & t[15];
  assign t[9] = ~(t[23]);
  assign y = (t[0]);
endmodule

module R2ind219(x, y);
 input [11:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[24] ^ t[22];
  assign t[12] = ~(t[22]);
  assign t[13] = t[11] ^ t[25];
  assign t[14] = ~(t[7] ^ t[16]);
  assign t[15] = t[17] ^ t[13];
  assign t[16] = t[18] ^ t[6];
  assign t[17] = t[22] ^ t[9];
  assign t[18] = t[19] & t[20];
  assign t[19] = ~(t[21]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11]);
  assign t[21] = t[13] ^ t[22];
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34] & ~t[35]);
  assign t[31] = (t[36] & ~t[37]);
  assign t[32] = (t[38] & ~t[39]);
  assign t[33] = (t[40] & ~t[41]);
  assign t[34] = t[42] ^ x[2];
  assign t[35] = t[43] ^ x[1];
  assign t[36] = t[44] ^ x[5];
  assign t[37] = t[45] ^ x[4];
  assign t[38] = t[46] ^ x[8];
  assign t[39] = t[47] ^ x[7];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[11];
  assign t[41] = t[49] ^ x[10];
  assign t[42] = (x[0]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[3]);
  assign t[46] = (x[6]);
  assign t[47] = (x[6]);
  assign t[48] = (x[9]);
  assign t[49] = (x[9]);
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[11] ^ t[9];
  assign t[6] = t[12] & t[13];
  assign t[7] = t[11] ^ t[22];
  assign t[8] = t[14] & t[15];
  assign t[9] = ~(t[23]);
  assign y = (t[0]);
endmodule

module R2ind220(x, y);
 input [11:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[15] ^ t[29];
  assign t[12] = t[20] & t[21];
  assign t[13] = ~(t[30]);
  assign t[14] = t[18] ^ t[12];
  assign t[15] = t[31] ^ t[29];
  assign t[16] = ~(t[29]);
  assign t[17] = t[15] ^ t[32];
  assign t[18] = t[22] ^ t[8];
  assign t[19] = t[23] & t[24];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11] ^ t[18]);
  assign t[21] = t[9] ^ t[17];
  assign t[22] = t[25] & t[26];
  assign t[23] = ~(t[22] ^ t[27]);
  assign t[24] = t[7] ^ t[28];
  assign t[25] = ~(t[28]);
  assign t[26] = ~(t[15]);
  assign t[27] = t[9] ^ t[15];
  assign t[28] = t[17] ^ t[29];
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = (t[35]);
  assign t[32] = (t[36]);
  assign t[33] = t[37] ^ x[2];
  assign t[34] = t[38] ^ x[5];
  assign t[35] = t[39] ^ x[8];
  assign t[36] = t[40] ^ x[11];
  assign t[37] = (t[41] & ~t[42]);
  assign t[38] = (t[43] & ~t[44]);
  assign t[39] = (t[45] & ~t[46]);
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (t[47] & ~t[48]);
  assign t[41] = t[49] ^ x[2];
  assign t[42] = t[50] ^ x[1];
  assign t[43] = t[51] ^ x[5];
  assign t[44] = t[52] ^ x[4];
  assign t[45] = t[53] ^ x[8];
  assign t[46] = t[54] ^ x[7];
  assign t[47] = t[55] ^ x[11];
  assign t[48] = t[56] ^ x[10];
  assign t[49] = (x[0]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[0]);
  assign t[51] = (x[3]);
  assign t[52] = (x[3]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[9]);
  assign t[56] = (x[9]);
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[15] ^ t[13];
  assign t[8] = t[16] & t[17];
  assign t[9] = t[29] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind221(x, y);
 input [11:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[15] ^ t[29];
  assign t[12] = t[20] & t[21];
  assign t[13] = ~(t[30]);
  assign t[14] = t[18] ^ t[12];
  assign t[15] = t[31] ^ t[29];
  assign t[16] = ~(t[29]);
  assign t[17] = t[15] ^ t[32];
  assign t[18] = t[22] ^ t[8];
  assign t[19] = t[23] & t[24];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11] ^ t[18]);
  assign t[21] = t[9] ^ t[17];
  assign t[22] = t[25] & t[26];
  assign t[23] = ~(t[22] ^ t[27]);
  assign t[24] = t[7] ^ t[28];
  assign t[25] = ~(t[28]);
  assign t[26] = ~(t[15]);
  assign t[27] = t[9] ^ t[15];
  assign t[28] = t[17] ^ t[29];
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = (t[35]);
  assign t[32] = (t[36]);
  assign t[33] = t[37] ^ x[2];
  assign t[34] = t[38] ^ x[5];
  assign t[35] = t[39] ^ x[8];
  assign t[36] = t[40] ^ x[11];
  assign t[37] = (t[41] & ~t[42]);
  assign t[38] = (t[43] & ~t[44]);
  assign t[39] = (t[45] & ~t[46]);
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (t[47] & ~t[48]);
  assign t[41] = t[49] ^ x[2];
  assign t[42] = t[50] ^ x[1];
  assign t[43] = t[51] ^ x[5];
  assign t[44] = t[52] ^ x[4];
  assign t[45] = t[53] ^ x[8];
  assign t[46] = t[54] ^ x[7];
  assign t[47] = t[55] ^ x[11];
  assign t[48] = t[56] ^ x[10];
  assign t[49] = (x[0]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[0]);
  assign t[51] = (x[3]);
  assign t[52] = (x[3]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[9]);
  assign t[56] = (x[9]);
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[15] ^ t[13];
  assign t[8] = t[16] & t[17];
  assign t[9] = t[29] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind222(x, y);
 input [11:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] ^ t[16];
  assign t[11] = t[17] ^ t[8];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[29] ^ t[28];
  assign t[14] = ~(t[28]);
  assign t[15] = t[13] ^ t[30];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[22] & t[23];
  assign t[18] = ~(t[24] ^ t[11]);
  assign t[19] = t[9] ^ t[15];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[17] ^ t[25]);
  assign t[21] = t[7] ^ t[26];
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[13]);
  assign t[24] = t[13] ^ t[28];
  assign t[25] = t[9] ^ t[13];
  assign t[26] = t[15] ^ t[28];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[2];
  assign t[32] = t[36] ^ x[5];
  assign t[33] = t[37] ^ x[8];
  assign t[34] = t[38] ^ x[11];
  assign t[35] = (t[39] & ~t[40]);
  assign t[36] = (t[41] & ~t[42]);
  assign t[37] = (t[43] & ~t[44]);
  assign t[38] = (t[45] & ~t[46]);
  assign t[39] = t[47] ^ x[2];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[1];
  assign t[41] = t[49] ^ x[5];
  assign t[42] = t[50] ^ x[4];
  assign t[43] = t[51] ^ x[8];
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[11];
  assign t[46] = t[54] ^ x[10];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[5] = ~(t[27]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[13] ^ t[5];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[28] ^ t[5];
  assign y = (t[0]);
endmodule

module R2ind223(x, y);
 input [11:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] ^ t[16];
  assign t[11] = t[17] ^ t[8];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[29] ^ t[28];
  assign t[14] = ~(t[28]);
  assign t[15] = t[13] ^ t[30];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[22] & t[23];
  assign t[18] = ~(t[24] ^ t[11]);
  assign t[19] = t[9] ^ t[15];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[17] ^ t[25]);
  assign t[21] = t[7] ^ t[26];
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[13]);
  assign t[24] = t[13] ^ t[28];
  assign t[25] = t[9] ^ t[13];
  assign t[26] = t[15] ^ t[28];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[2];
  assign t[32] = t[36] ^ x[5];
  assign t[33] = t[37] ^ x[8];
  assign t[34] = t[38] ^ x[11];
  assign t[35] = (t[39] & ~t[40]);
  assign t[36] = (t[41] & ~t[42]);
  assign t[37] = (t[43] & ~t[44]);
  assign t[38] = (t[45] & ~t[46]);
  assign t[39] = t[47] ^ x[2];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[1];
  assign t[41] = t[49] ^ x[5];
  assign t[42] = t[50] ^ x[4];
  assign t[43] = t[51] ^ x[8];
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[11];
  assign t[46] = t[54] ^ x[10];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[5] = ~(t[27]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[13] ^ t[5];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[28] ^ t[5];
  assign y = (t[0]);
endmodule

module R2ind224(x, y);
 input [11:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[7] ^ t[23];
  assign t[11] = t[13] ^ t[4];
  assign t[12] = t[14] & t[15];
  assign t[13] = t[16] & t[17];
  assign t[14] = ~(t[13] ^ t[18]);
  assign t[15] = t[3] ^ t[19];
  assign t[16] = ~(t[19]);
  assign t[17] = ~(t[7]);
  assign t[18] = t[5] ^ t[7];
  assign t[19] = t[10] ^ t[20];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = t[28] ^ x[2];
  assign t[25] = t[29] ^ x[5];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = t[31] ^ x[11];
  assign t[28] = (t[32] & ~t[33]);
  assign t[29] = (t[34] & ~t[35]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[36] & ~t[37]);
  assign t[31] = (t[38] & ~t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[1];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[4];
  assign t[36] = t[44] ^ x[8];
  assign t[37] = t[45] ^ x[7];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[10];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[4] = t[9] & t[10];
  assign t[5] = t[20] ^ t[8];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[21] ^ t[20];
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind225(x, y);
 input [11:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[7] ^ t[23];
  assign t[11] = t[13] ^ t[4];
  assign t[12] = t[14] & t[15];
  assign t[13] = t[16] & t[17];
  assign t[14] = ~(t[13] ^ t[18]);
  assign t[15] = t[3] ^ t[19];
  assign t[16] = ~(t[19]);
  assign t[17] = ~(t[7]);
  assign t[18] = t[5] ^ t[7];
  assign t[19] = t[10] ^ t[20];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = t[28] ^ x[2];
  assign t[25] = t[29] ^ x[5];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = t[31] ^ x[11];
  assign t[28] = (t[32] & ~t[33]);
  assign t[29] = (t[34] & ~t[35]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[36] & ~t[37]);
  assign t[31] = (t[38] & ~t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[1];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[4];
  assign t[36] = t[44] ^ x[8];
  assign t[37] = t[45] ^ x[7];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[10];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[4] = t[9] & t[10];
  assign t[5] = t[20] ^ t[8];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[21] ^ t[20];
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind226(x, y);
 input [11:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[24] ^ t[22];
  assign t[12] = ~(t[22]);
  assign t[13] = t[11] ^ t[25];
  assign t[14] = ~(t[7] ^ t[16]);
  assign t[15] = t[17] ^ t[13];
  assign t[16] = t[18] ^ t[6];
  assign t[17] = t[22] ^ t[9];
  assign t[18] = t[19] & t[20];
  assign t[19] = ~(t[21]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11]);
  assign t[21] = t[13] ^ t[22];
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34] & ~t[35]);
  assign t[31] = (t[36] & ~t[37]);
  assign t[32] = (t[38] & ~t[39]);
  assign t[33] = (t[40] & ~t[41]);
  assign t[34] = t[42] ^ x[2];
  assign t[35] = t[43] ^ x[1];
  assign t[36] = t[44] ^ x[5];
  assign t[37] = t[45] ^ x[4];
  assign t[38] = t[46] ^ x[8];
  assign t[39] = t[47] ^ x[7];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[11];
  assign t[41] = t[49] ^ x[10];
  assign t[42] = (x[0]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[3]);
  assign t[46] = (x[6]);
  assign t[47] = (x[6]);
  assign t[48] = (x[9]);
  assign t[49] = (x[9]);
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[11] ^ t[9];
  assign t[6] = t[12] & t[13];
  assign t[7] = t[11] ^ t[22];
  assign t[8] = t[14] & t[15];
  assign t[9] = ~(t[23]);
  assign y = (t[0]);
endmodule

module R2ind227(x, y);
 input [11:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[24] ^ t[22];
  assign t[12] = ~(t[22]);
  assign t[13] = t[11] ^ t[25];
  assign t[14] = ~(t[7] ^ t[16]);
  assign t[15] = t[17] ^ t[13];
  assign t[16] = t[18] ^ t[6];
  assign t[17] = t[22] ^ t[9];
  assign t[18] = t[19] & t[20];
  assign t[19] = ~(t[21]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11]);
  assign t[21] = t[13] ^ t[22];
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34] & ~t[35]);
  assign t[31] = (t[36] & ~t[37]);
  assign t[32] = (t[38] & ~t[39]);
  assign t[33] = (t[40] & ~t[41]);
  assign t[34] = t[42] ^ x[2];
  assign t[35] = t[43] ^ x[1];
  assign t[36] = t[44] ^ x[5];
  assign t[37] = t[45] ^ x[4];
  assign t[38] = t[46] ^ x[8];
  assign t[39] = t[47] ^ x[7];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[11];
  assign t[41] = t[49] ^ x[10];
  assign t[42] = (x[0]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[3]);
  assign t[46] = (x[6]);
  assign t[47] = (x[6]);
  assign t[48] = (x[9]);
  assign t[49] = (x[9]);
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[11] ^ t[9];
  assign t[6] = t[12] & t[13];
  assign t[7] = t[11] ^ t[22];
  assign t[8] = t[14] & t[15];
  assign t[9] = ~(t[23]);
  assign y = (t[0]);
endmodule

module R2ind228(x, y);
 input [11:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[15] ^ t[29];
  assign t[12] = t[20] & t[21];
  assign t[13] = ~(t[30]);
  assign t[14] = t[18] ^ t[12];
  assign t[15] = t[31] ^ t[29];
  assign t[16] = ~(t[29]);
  assign t[17] = t[15] ^ t[32];
  assign t[18] = t[22] ^ t[8];
  assign t[19] = t[23] & t[24];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11] ^ t[18]);
  assign t[21] = t[9] ^ t[17];
  assign t[22] = t[25] & t[26];
  assign t[23] = ~(t[22] ^ t[27]);
  assign t[24] = t[7] ^ t[28];
  assign t[25] = ~(t[28]);
  assign t[26] = ~(t[15]);
  assign t[27] = t[9] ^ t[15];
  assign t[28] = t[17] ^ t[29];
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = (t[35]);
  assign t[32] = (t[36]);
  assign t[33] = t[37] ^ x[2];
  assign t[34] = t[38] ^ x[5];
  assign t[35] = t[39] ^ x[8];
  assign t[36] = t[40] ^ x[11];
  assign t[37] = (t[41] & ~t[42]);
  assign t[38] = (t[43] & ~t[44]);
  assign t[39] = (t[45] & ~t[46]);
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (t[47] & ~t[48]);
  assign t[41] = t[49] ^ x[2];
  assign t[42] = t[50] ^ x[1];
  assign t[43] = t[51] ^ x[5];
  assign t[44] = t[52] ^ x[4];
  assign t[45] = t[53] ^ x[8];
  assign t[46] = t[54] ^ x[7];
  assign t[47] = t[55] ^ x[11];
  assign t[48] = t[56] ^ x[10];
  assign t[49] = (x[0]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[0]);
  assign t[51] = (x[3]);
  assign t[52] = (x[3]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[9]);
  assign t[56] = (x[9]);
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[15] ^ t[13];
  assign t[8] = t[16] & t[17];
  assign t[9] = t[29] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind229(x, y);
 input [11:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[15] ^ t[29];
  assign t[12] = t[20] & t[21];
  assign t[13] = ~(t[30]);
  assign t[14] = t[18] ^ t[12];
  assign t[15] = t[31] ^ t[29];
  assign t[16] = ~(t[29]);
  assign t[17] = t[15] ^ t[32];
  assign t[18] = t[22] ^ t[8];
  assign t[19] = t[23] & t[24];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11] ^ t[18]);
  assign t[21] = t[9] ^ t[17];
  assign t[22] = t[25] & t[26];
  assign t[23] = ~(t[22] ^ t[27]);
  assign t[24] = t[7] ^ t[28];
  assign t[25] = ~(t[28]);
  assign t[26] = ~(t[15]);
  assign t[27] = t[9] ^ t[15];
  assign t[28] = t[17] ^ t[29];
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = (t[35]);
  assign t[32] = (t[36]);
  assign t[33] = t[37] ^ x[2];
  assign t[34] = t[38] ^ x[5];
  assign t[35] = t[39] ^ x[8];
  assign t[36] = t[40] ^ x[11];
  assign t[37] = (t[41] & ~t[42]);
  assign t[38] = (t[43] & ~t[44]);
  assign t[39] = (t[45] & ~t[46]);
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (t[47] & ~t[48]);
  assign t[41] = t[49] ^ x[2];
  assign t[42] = t[50] ^ x[1];
  assign t[43] = t[51] ^ x[5];
  assign t[44] = t[52] ^ x[4];
  assign t[45] = t[53] ^ x[8];
  assign t[46] = t[54] ^ x[7];
  assign t[47] = t[55] ^ x[11];
  assign t[48] = t[56] ^ x[10];
  assign t[49] = (x[0]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[0]);
  assign t[51] = (x[3]);
  assign t[52] = (x[3]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[9]);
  assign t[56] = (x[9]);
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[15] ^ t[13];
  assign t[8] = t[16] & t[17];
  assign t[9] = t[29] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind230(x, y);
 input [11:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] ^ t[16];
  assign t[11] = t[17] ^ t[8];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[29] ^ t[28];
  assign t[14] = ~(t[28]);
  assign t[15] = t[13] ^ t[30];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[22] & t[23];
  assign t[18] = ~(t[24] ^ t[11]);
  assign t[19] = t[9] ^ t[15];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[17] ^ t[25]);
  assign t[21] = t[7] ^ t[26];
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[13]);
  assign t[24] = t[13] ^ t[28];
  assign t[25] = t[9] ^ t[13];
  assign t[26] = t[15] ^ t[28];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[2];
  assign t[32] = t[36] ^ x[5];
  assign t[33] = t[37] ^ x[8];
  assign t[34] = t[38] ^ x[11];
  assign t[35] = (t[39] & ~t[40]);
  assign t[36] = (t[41] & ~t[42]);
  assign t[37] = (t[43] & ~t[44]);
  assign t[38] = (t[45] & ~t[46]);
  assign t[39] = t[47] ^ x[2];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[1];
  assign t[41] = t[49] ^ x[5];
  assign t[42] = t[50] ^ x[4];
  assign t[43] = t[51] ^ x[8];
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[11];
  assign t[46] = t[54] ^ x[10];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[5] = ~(t[27]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[13] ^ t[5];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[28] ^ t[5];
  assign y = (t[0]);
endmodule

module R2ind231(x, y);
 input [11:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] ^ t[16];
  assign t[11] = t[17] ^ t[8];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[29] ^ t[28];
  assign t[14] = ~(t[28]);
  assign t[15] = t[13] ^ t[30];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[22] & t[23];
  assign t[18] = ~(t[24] ^ t[11]);
  assign t[19] = t[9] ^ t[15];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[17] ^ t[25]);
  assign t[21] = t[7] ^ t[26];
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[13]);
  assign t[24] = t[13] ^ t[28];
  assign t[25] = t[9] ^ t[13];
  assign t[26] = t[15] ^ t[28];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[2];
  assign t[32] = t[36] ^ x[5];
  assign t[33] = t[37] ^ x[8];
  assign t[34] = t[38] ^ x[11];
  assign t[35] = (t[39] & ~t[40]);
  assign t[36] = (t[41] & ~t[42]);
  assign t[37] = (t[43] & ~t[44]);
  assign t[38] = (t[45] & ~t[46]);
  assign t[39] = t[47] ^ x[2];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[1];
  assign t[41] = t[49] ^ x[5];
  assign t[42] = t[50] ^ x[4];
  assign t[43] = t[51] ^ x[8];
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[11];
  assign t[46] = t[54] ^ x[10];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[5] = ~(t[27]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[13] ^ t[5];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[28] ^ t[5];
  assign y = (t[0]);
endmodule

module R2ind232(x, y);
 input [11:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[7] ^ t[23];
  assign t[11] = t[13] ^ t[4];
  assign t[12] = t[14] & t[15];
  assign t[13] = t[16] & t[17];
  assign t[14] = ~(t[13] ^ t[18]);
  assign t[15] = t[3] ^ t[19];
  assign t[16] = ~(t[19]);
  assign t[17] = ~(t[7]);
  assign t[18] = t[5] ^ t[7];
  assign t[19] = t[10] ^ t[20];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = t[28] ^ x[2];
  assign t[25] = t[29] ^ x[5];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = t[31] ^ x[11];
  assign t[28] = (t[32] & ~t[33]);
  assign t[29] = (t[34] & ~t[35]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[36] & ~t[37]);
  assign t[31] = (t[38] & ~t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[1];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[4];
  assign t[36] = t[44] ^ x[8];
  assign t[37] = t[45] ^ x[7];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[10];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[4] = t[9] & t[10];
  assign t[5] = t[20] ^ t[8];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[21] ^ t[20];
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind233(x, y);
 input [11:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[7] ^ t[23];
  assign t[11] = t[13] ^ t[4];
  assign t[12] = t[14] & t[15];
  assign t[13] = t[16] & t[17];
  assign t[14] = ~(t[13] ^ t[18]);
  assign t[15] = t[3] ^ t[19];
  assign t[16] = ~(t[19]);
  assign t[17] = ~(t[7]);
  assign t[18] = t[5] ^ t[7];
  assign t[19] = t[10] ^ t[20];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = t[28] ^ x[2];
  assign t[25] = t[29] ^ x[5];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = t[31] ^ x[11];
  assign t[28] = (t[32] & ~t[33]);
  assign t[29] = (t[34] & ~t[35]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[36] & ~t[37]);
  assign t[31] = (t[38] & ~t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[1];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[4];
  assign t[36] = t[44] ^ x[8];
  assign t[37] = t[45] ^ x[7];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[10];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[4] = t[9] & t[10];
  assign t[5] = t[20] ^ t[8];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[21] ^ t[20];
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind234(x, y);
 input [11:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[24] ^ t[22];
  assign t[12] = ~(t[22]);
  assign t[13] = t[11] ^ t[25];
  assign t[14] = ~(t[7] ^ t[16]);
  assign t[15] = t[17] ^ t[13];
  assign t[16] = t[18] ^ t[6];
  assign t[17] = t[22] ^ t[9];
  assign t[18] = t[19] & t[20];
  assign t[19] = ~(t[21]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11]);
  assign t[21] = t[13] ^ t[22];
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34] & ~t[35]);
  assign t[31] = (t[36] & ~t[37]);
  assign t[32] = (t[38] & ~t[39]);
  assign t[33] = (t[40] & ~t[41]);
  assign t[34] = t[42] ^ x[2];
  assign t[35] = t[43] ^ x[1];
  assign t[36] = t[44] ^ x[5];
  assign t[37] = t[45] ^ x[4];
  assign t[38] = t[46] ^ x[8];
  assign t[39] = t[47] ^ x[7];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[11];
  assign t[41] = t[49] ^ x[10];
  assign t[42] = (x[0]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[3]);
  assign t[46] = (x[6]);
  assign t[47] = (x[6]);
  assign t[48] = (x[9]);
  assign t[49] = (x[9]);
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[11] ^ t[9];
  assign t[6] = t[12] & t[13];
  assign t[7] = t[11] ^ t[22];
  assign t[8] = t[14] & t[15];
  assign t[9] = ~(t[23]);
  assign y = (t[0]);
endmodule

module R2ind235(x, y);
 input [11:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[24] ^ t[22];
  assign t[12] = ~(t[22]);
  assign t[13] = t[11] ^ t[25];
  assign t[14] = ~(t[7] ^ t[16]);
  assign t[15] = t[17] ^ t[13];
  assign t[16] = t[18] ^ t[6];
  assign t[17] = t[22] ^ t[9];
  assign t[18] = t[19] & t[20];
  assign t[19] = ~(t[21]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11]);
  assign t[21] = t[13] ^ t[22];
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34] & ~t[35]);
  assign t[31] = (t[36] & ~t[37]);
  assign t[32] = (t[38] & ~t[39]);
  assign t[33] = (t[40] & ~t[41]);
  assign t[34] = t[42] ^ x[2];
  assign t[35] = t[43] ^ x[1];
  assign t[36] = t[44] ^ x[5];
  assign t[37] = t[45] ^ x[4];
  assign t[38] = t[46] ^ x[8];
  assign t[39] = t[47] ^ x[7];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[11];
  assign t[41] = t[49] ^ x[10];
  assign t[42] = (x[0]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[3]);
  assign t[46] = (x[6]);
  assign t[47] = (x[6]);
  assign t[48] = (x[9]);
  assign t[49] = (x[9]);
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[11] ^ t[9];
  assign t[6] = t[12] & t[13];
  assign t[7] = t[11] ^ t[22];
  assign t[8] = t[14] & t[15];
  assign t[9] = ~(t[23]);
  assign y = (t[0]);
endmodule

module R2ind236(x, y);
 input [11:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[15] ^ t[29];
  assign t[12] = t[20] & t[21];
  assign t[13] = ~(t[30]);
  assign t[14] = t[18] ^ t[12];
  assign t[15] = t[31] ^ t[29];
  assign t[16] = ~(t[29]);
  assign t[17] = t[15] ^ t[32];
  assign t[18] = t[22] ^ t[8];
  assign t[19] = t[23] & t[24];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11] ^ t[18]);
  assign t[21] = t[9] ^ t[17];
  assign t[22] = t[25] & t[26];
  assign t[23] = ~(t[22] ^ t[27]);
  assign t[24] = t[7] ^ t[28];
  assign t[25] = ~(t[28]);
  assign t[26] = ~(t[15]);
  assign t[27] = t[9] ^ t[15];
  assign t[28] = t[17] ^ t[29];
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = (t[35]);
  assign t[32] = (t[36]);
  assign t[33] = t[37] ^ x[2];
  assign t[34] = t[38] ^ x[5];
  assign t[35] = t[39] ^ x[8];
  assign t[36] = t[40] ^ x[11];
  assign t[37] = (t[41] & ~t[42]);
  assign t[38] = (t[43] & ~t[44]);
  assign t[39] = (t[45] & ~t[46]);
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (t[47] & ~t[48]);
  assign t[41] = t[49] ^ x[2];
  assign t[42] = t[50] ^ x[1];
  assign t[43] = t[51] ^ x[5];
  assign t[44] = t[52] ^ x[4];
  assign t[45] = t[53] ^ x[8];
  assign t[46] = t[54] ^ x[7];
  assign t[47] = t[55] ^ x[11];
  assign t[48] = t[56] ^ x[10];
  assign t[49] = (x[0]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[0]);
  assign t[51] = (x[3]);
  assign t[52] = (x[3]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[9]);
  assign t[56] = (x[9]);
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[15] ^ t[13];
  assign t[8] = t[16] & t[17];
  assign t[9] = t[29] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind237(x, y);
 input [11:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[15] ^ t[29];
  assign t[12] = t[20] & t[21];
  assign t[13] = ~(t[30]);
  assign t[14] = t[18] ^ t[12];
  assign t[15] = t[31] ^ t[29];
  assign t[16] = ~(t[29]);
  assign t[17] = t[15] ^ t[32];
  assign t[18] = t[22] ^ t[8];
  assign t[19] = t[23] & t[24];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11] ^ t[18]);
  assign t[21] = t[9] ^ t[17];
  assign t[22] = t[25] & t[26];
  assign t[23] = ~(t[22] ^ t[27]);
  assign t[24] = t[7] ^ t[28];
  assign t[25] = ~(t[28]);
  assign t[26] = ~(t[15]);
  assign t[27] = t[9] ^ t[15];
  assign t[28] = t[17] ^ t[29];
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = (t[35]);
  assign t[32] = (t[36]);
  assign t[33] = t[37] ^ x[2];
  assign t[34] = t[38] ^ x[5];
  assign t[35] = t[39] ^ x[8];
  assign t[36] = t[40] ^ x[11];
  assign t[37] = (t[41] & ~t[42]);
  assign t[38] = (t[43] & ~t[44]);
  assign t[39] = (t[45] & ~t[46]);
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (t[47] & ~t[48]);
  assign t[41] = t[49] ^ x[2];
  assign t[42] = t[50] ^ x[1];
  assign t[43] = t[51] ^ x[5];
  assign t[44] = t[52] ^ x[4];
  assign t[45] = t[53] ^ x[8];
  assign t[46] = t[54] ^ x[7];
  assign t[47] = t[55] ^ x[11];
  assign t[48] = t[56] ^ x[10];
  assign t[49] = (x[0]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[0]);
  assign t[51] = (x[3]);
  assign t[52] = (x[3]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[9]);
  assign t[56] = (x[9]);
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[15] ^ t[13];
  assign t[8] = t[16] & t[17];
  assign t[9] = t[29] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind238(x, y);
 input [11:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] ^ t[16];
  assign t[11] = t[17] ^ t[8];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[29] ^ t[28];
  assign t[14] = ~(t[28]);
  assign t[15] = t[13] ^ t[30];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[22] & t[23];
  assign t[18] = ~(t[24] ^ t[11]);
  assign t[19] = t[9] ^ t[15];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[17] ^ t[25]);
  assign t[21] = t[7] ^ t[26];
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[13]);
  assign t[24] = t[13] ^ t[28];
  assign t[25] = t[9] ^ t[13];
  assign t[26] = t[15] ^ t[28];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[2];
  assign t[32] = t[36] ^ x[5];
  assign t[33] = t[37] ^ x[8];
  assign t[34] = t[38] ^ x[11];
  assign t[35] = (t[39] & ~t[40]);
  assign t[36] = (t[41] & ~t[42]);
  assign t[37] = (t[43] & ~t[44]);
  assign t[38] = (t[45] & ~t[46]);
  assign t[39] = t[47] ^ x[2];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[1];
  assign t[41] = t[49] ^ x[5];
  assign t[42] = t[50] ^ x[4];
  assign t[43] = t[51] ^ x[8];
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[11];
  assign t[46] = t[54] ^ x[10];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[5] = ~(t[27]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[13] ^ t[5];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[28] ^ t[5];
  assign y = (t[0]);
endmodule

module R2ind239(x, y);
 input [11:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] ^ t[16];
  assign t[11] = t[17] ^ t[8];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[29] ^ t[28];
  assign t[14] = ~(t[28]);
  assign t[15] = t[13] ^ t[30];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[22] & t[23];
  assign t[18] = ~(t[24] ^ t[11]);
  assign t[19] = t[9] ^ t[15];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[17] ^ t[25]);
  assign t[21] = t[7] ^ t[26];
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[13]);
  assign t[24] = t[13] ^ t[28];
  assign t[25] = t[9] ^ t[13];
  assign t[26] = t[15] ^ t[28];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[2];
  assign t[32] = t[36] ^ x[5];
  assign t[33] = t[37] ^ x[8];
  assign t[34] = t[38] ^ x[11];
  assign t[35] = (t[39] & ~t[40]);
  assign t[36] = (t[41] & ~t[42]);
  assign t[37] = (t[43] & ~t[44]);
  assign t[38] = (t[45] & ~t[46]);
  assign t[39] = t[47] ^ x[2];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[1];
  assign t[41] = t[49] ^ x[5];
  assign t[42] = t[50] ^ x[4];
  assign t[43] = t[51] ^ x[8];
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[11];
  assign t[46] = t[54] ^ x[10];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[5] = ~(t[27]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[13] ^ t[5];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[28] ^ t[5];
  assign y = (t[0]);
endmodule

module R2ind240(x, y);
 input [11:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[7] ^ t[23];
  assign t[11] = t[13] ^ t[4];
  assign t[12] = t[14] & t[15];
  assign t[13] = t[16] & t[17];
  assign t[14] = ~(t[13] ^ t[18]);
  assign t[15] = t[3] ^ t[19];
  assign t[16] = ~(t[19]);
  assign t[17] = ~(t[7]);
  assign t[18] = t[5] ^ t[7];
  assign t[19] = t[10] ^ t[20];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = t[28] ^ x[2];
  assign t[25] = t[29] ^ x[5];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = t[31] ^ x[11];
  assign t[28] = (t[32] & ~t[33]);
  assign t[29] = (t[34] & ~t[35]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[36] & ~t[37]);
  assign t[31] = (t[38] & ~t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[1];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[4];
  assign t[36] = t[44] ^ x[8];
  assign t[37] = t[45] ^ x[7];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[10];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[4] = t[9] & t[10];
  assign t[5] = t[20] ^ t[8];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[21] ^ t[20];
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind241(x, y);
 input [11:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[7] ^ t[23];
  assign t[11] = t[13] ^ t[4];
  assign t[12] = t[14] & t[15];
  assign t[13] = t[16] & t[17];
  assign t[14] = ~(t[13] ^ t[18]);
  assign t[15] = t[3] ^ t[19];
  assign t[16] = ~(t[19]);
  assign t[17] = ~(t[7]);
  assign t[18] = t[5] ^ t[7];
  assign t[19] = t[10] ^ t[20];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = t[28] ^ x[2];
  assign t[25] = t[29] ^ x[5];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = t[31] ^ x[11];
  assign t[28] = (t[32] & ~t[33]);
  assign t[29] = (t[34] & ~t[35]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[36] & ~t[37]);
  assign t[31] = (t[38] & ~t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[1];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[4];
  assign t[36] = t[44] ^ x[8];
  assign t[37] = t[45] ^ x[7];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[10];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[4] = t[9] & t[10];
  assign t[5] = t[20] ^ t[8];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[21] ^ t[20];
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind242(x, y);
 input [11:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[24] ^ t[22];
  assign t[12] = ~(t[22]);
  assign t[13] = t[11] ^ t[25];
  assign t[14] = ~(t[7] ^ t[16]);
  assign t[15] = t[17] ^ t[13];
  assign t[16] = t[18] ^ t[6];
  assign t[17] = t[22] ^ t[9];
  assign t[18] = t[19] & t[20];
  assign t[19] = ~(t[21]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11]);
  assign t[21] = t[13] ^ t[22];
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34] & ~t[35]);
  assign t[31] = (t[36] & ~t[37]);
  assign t[32] = (t[38] & ~t[39]);
  assign t[33] = (t[40] & ~t[41]);
  assign t[34] = t[42] ^ x[2];
  assign t[35] = t[43] ^ x[1];
  assign t[36] = t[44] ^ x[5];
  assign t[37] = t[45] ^ x[4];
  assign t[38] = t[46] ^ x[8];
  assign t[39] = t[47] ^ x[7];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[11];
  assign t[41] = t[49] ^ x[10];
  assign t[42] = (x[0]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[3]);
  assign t[46] = (x[6]);
  assign t[47] = (x[6]);
  assign t[48] = (x[9]);
  assign t[49] = (x[9]);
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[11] ^ t[9];
  assign t[6] = t[12] & t[13];
  assign t[7] = t[11] ^ t[22];
  assign t[8] = t[14] & t[15];
  assign t[9] = ~(t[23]);
  assign y = (t[0]);
endmodule

module R2ind243(x, y);
 input [11:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[24] ^ t[22];
  assign t[12] = ~(t[22]);
  assign t[13] = t[11] ^ t[25];
  assign t[14] = ~(t[7] ^ t[16]);
  assign t[15] = t[17] ^ t[13];
  assign t[16] = t[18] ^ t[6];
  assign t[17] = t[22] ^ t[9];
  assign t[18] = t[19] & t[20];
  assign t[19] = ~(t[21]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11]);
  assign t[21] = t[13] ^ t[22];
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34] & ~t[35]);
  assign t[31] = (t[36] & ~t[37]);
  assign t[32] = (t[38] & ~t[39]);
  assign t[33] = (t[40] & ~t[41]);
  assign t[34] = t[42] ^ x[2];
  assign t[35] = t[43] ^ x[1];
  assign t[36] = t[44] ^ x[5];
  assign t[37] = t[45] ^ x[4];
  assign t[38] = t[46] ^ x[8];
  assign t[39] = t[47] ^ x[7];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[11];
  assign t[41] = t[49] ^ x[10];
  assign t[42] = (x[0]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[3]);
  assign t[46] = (x[6]);
  assign t[47] = (x[6]);
  assign t[48] = (x[9]);
  assign t[49] = (x[9]);
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[11] ^ t[9];
  assign t[6] = t[12] & t[13];
  assign t[7] = t[11] ^ t[22];
  assign t[8] = t[14] & t[15];
  assign t[9] = ~(t[23]);
  assign y = (t[0]);
endmodule

module R2ind244(x, y);
 input [11:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[15] ^ t[29];
  assign t[12] = t[20] & t[21];
  assign t[13] = ~(t[30]);
  assign t[14] = t[18] ^ t[12];
  assign t[15] = t[31] ^ t[29];
  assign t[16] = ~(t[29]);
  assign t[17] = t[15] ^ t[32];
  assign t[18] = t[22] ^ t[8];
  assign t[19] = t[23] & t[24];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11] ^ t[18]);
  assign t[21] = t[9] ^ t[17];
  assign t[22] = t[25] & t[26];
  assign t[23] = ~(t[22] ^ t[27]);
  assign t[24] = t[7] ^ t[28];
  assign t[25] = ~(t[28]);
  assign t[26] = ~(t[15]);
  assign t[27] = t[9] ^ t[15];
  assign t[28] = t[17] ^ t[29];
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = (t[35]);
  assign t[32] = (t[36]);
  assign t[33] = t[37] ^ x[2];
  assign t[34] = t[38] ^ x[5];
  assign t[35] = t[39] ^ x[8];
  assign t[36] = t[40] ^ x[11];
  assign t[37] = (t[41] & ~t[42]);
  assign t[38] = (t[43] & ~t[44]);
  assign t[39] = (t[45] & ~t[46]);
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (t[47] & ~t[48]);
  assign t[41] = t[49] ^ x[2];
  assign t[42] = t[50] ^ x[1];
  assign t[43] = t[51] ^ x[5];
  assign t[44] = t[52] ^ x[4];
  assign t[45] = t[53] ^ x[8];
  assign t[46] = t[54] ^ x[7];
  assign t[47] = t[55] ^ x[11];
  assign t[48] = t[56] ^ x[10];
  assign t[49] = (x[0]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[0]);
  assign t[51] = (x[3]);
  assign t[52] = (x[3]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[9]);
  assign t[56] = (x[9]);
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[15] ^ t[13];
  assign t[8] = t[16] & t[17];
  assign t[9] = t[29] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind245(x, y);
 input [11:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[15] ^ t[29];
  assign t[12] = t[20] & t[21];
  assign t[13] = ~(t[30]);
  assign t[14] = t[18] ^ t[12];
  assign t[15] = t[31] ^ t[29];
  assign t[16] = ~(t[29]);
  assign t[17] = t[15] ^ t[32];
  assign t[18] = t[22] ^ t[8];
  assign t[19] = t[23] & t[24];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11] ^ t[18]);
  assign t[21] = t[9] ^ t[17];
  assign t[22] = t[25] & t[26];
  assign t[23] = ~(t[22] ^ t[27]);
  assign t[24] = t[7] ^ t[28];
  assign t[25] = ~(t[28]);
  assign t[26] = ~(t[15]);
  assign t[27] = t[9] ^ t[15];
  assign t[28] = t[17] ^ t[29];
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = (t[35]);
  assign t[32] = (t[36]);
  assign t[33] = t[37] ^ x[2];
  assign t[34] = t[38] ^ x[5];
  assign t[35] = t[39] ^ x[8];
  assign t[36] = t[40] ^ x[11];
  assign t[37] = (t[41] & ~t[42]);
  assign t[38] = (t[43] & ~t[44]);
  assign t[39] = (t[45] & ~t[46]);
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (t[47] & ~t[48]);
  assign t[41] = t[49] ^ x[2];
  assign t[42] = t[50] ^ x[1];
  assign t[43] = t[51] ^ x[5];
  assign t[44] = t[52] ^ x[4];
  assign t[45] = t[53] ^ x[8];
  assign t[46] = t[54] ^ x[7];
  assign t[47] = t[55] ^ x[11];
  assign t[48] = t[56] ^ x[10];
  assign t[49] = (x[0]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[0]);
  assign t[51] = (x[3]);
  assign t[52] = (x[3]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[9]);
  assign t[56] = (x[9]);
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[15] ^ t[13];
  assign t[8] = t[16] & t[17];
  assign t[9] = t[29] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind246(x, y);
 input [11:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] ^ t[16];
  assign t[11] = t[17] ^ t[8];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[29] ^ t[28];
  assign t[14] = ~(t[28]);
  assign t[15] = t[13] ^ t[30];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[22] & t[23];
  assign t[18] = ~(t[24] ^ t[11]);
  assign t[19] = t[9] ^ t[15];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[17] ^ t[25]);
  assign t[21] = t[7] ^ t[26];
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[13]);
  assign t[24] = t[13] ^ t[28];
  assign t[25] = t[9] ^ t[13];
  assign t[26] = t[15] ^ t[28];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[2];
  assign t[32] = t[36] ^ x[5];
  assign t[33] = t[37] ^ x[8];
  assign t[34] = t[38] ^ x[11];
  assign t[35] = (t[39] & ~t[40]);
  assign t[36] = (t[41] & ~t[42]);
  assign t[37] = (t[43] & ~t[44]);
  assign t[38] = (t[45] & ~t[46]);
  assign t[39] = t[47] ^ x[2];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[1];
  assign t[41] = t[49] ^ x[5];
  assign t[42] = t[50] ^ x[4];
  assign t[43] = t[51] ^ x[8];
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[11];
  assign t[46] = t[54] ^ x[10];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[5] = ~(t[27]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[13] ^ t[5];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[28] ^ t[5];
  assign y = (t[0]);
endmodule

module R2ind247(x, y);
 input [11:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] ^ t[16];
  assign t[11] = t[17] ^ t[8];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[29] ^ t[28];
  assign t[14] = ~(t[28]);
  assign t[15] = t[13] ^ t[30];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[22] & t[23];
  assign t[18] = ~(t[24] ^ t[11]);
  assign t[19] = t[9] ^ t[15];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[17] ^ t[25]);
  assign t[21] = t[7] ^ t[26];
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[13]);
  assign t[24] = t[13] ^ t[28];
  assign t[25] = t[9] ^ t[13];
  assign t[26] = t[15] ^ t[28];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[2];
  assign t[32] = t[36] ^ x[5];
  assign t[33] = t[37] ^ x[8];
  assign t[34] = t[38] ^ x[11];
  assign t[35] = (t[39] & ~t[40]);
  assign t[36] = (t[41] & ~t[42]);
  assign t[37] = (t[43] & ~t[44]);
  assign t[38] = (t[45] & ~t[46]);
  assign t[39] = t[47] ^ x[2];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[1];
  assign t[41] = t[49] ^ x[5];
  assign t[42] = t[50] ^ x[4];
  assign t[43] = t[51] ^ x[8];
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[11];
  assign t[46] = t[54] ^ x[10];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[5] = ~(t[27]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[13] ^ t[5];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[28] ^ t[5];
  assign y = (t[0]);
endmodule

module R2ind248(x, y);
 input [11:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[7] ^ t[23];
  assign t[11] = t[13] ^ t[4];
  assign t[12] = t[14] & t[15];
  assign t[13] = t[16] & t[17];
  assign t[14] = ~(t[13] ^ t[18]);
  assign t[15] = t[3] ^ t[19];
  assign t[16] = ~(t[19]);
  assign t[17] = ~(t[7]);
  assign t[18] = t[5] ^ t[7];
  assign t[19] = t[10] ^ t[20];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = t[28] ^ x[2];
  assign t[25] = t[29] ^ x[5];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = t[31] ^ x[11];
  assign t[28] = (t[32] & ~t[33]);
  assign t[29] = (t[34] & ~t[35]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[36] & ~t[37]);
  assign t[31] = (t[38] & ~t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[1];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[4];
  assign t[36] = t[44] ^ x[8];
  assign t[37] = t[45] ^ x[7];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[10];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[4] = t[9] & t[10];
  assign t[5] = t[20] ^ t[8];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[21] ^ t[20];
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind249(x, y);
 input [11:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[7] ^ t[23];
  assign t[11] = t[13] ^ t[4];
  assign t[12] = t[14] & t[15];
  assign t[13] = t[16] & t[17];
  assign t[14] = ~(t[13] ^ t[18]);
  assign t[15] = t[3] ^ t[19];
  assign t[16] = ~(t[19]);
  assign t[17] = ~(t[7]);
  assign t[18] = t[5] ^ t[7];
  assign t[19] = t[10] ^ t[20];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = t[28] ^ x[2];
  assign t[25] = t[29] ^ x[5];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = t[31] ^ x[11];
  assign t[28] = (t[32] & ~t[33]);
  assign t[29] = (t[34] & ~t[35]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[36] & ~t[37]);
  assign t[31] = (t[38] & ~t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[1];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[4];
  assign t[36] = t[44] ^ x[8];
  assign t[37] = t[45] ^ x[7];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[10];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[4] = t[9] & t[10];
  assign t[5] = t[20] ^ t[8];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[21] ^ t[20];
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind250(x, y);
 input [11:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[24] ^ t[22];
  assign t[12] = ~(t[22]);
  assign t[13] = t[11] ^ t[25];
  assign t[14] = ~(t[7] ^ t[16]);
  assign t[15] = t[17] ^ t[13];
  assign t[16] = t[18] ^ t[6];
  assign t[17] = t[22] ^ t[9];
  assign t[18] = t[19] & t[20];
  assign t[19] = ~(t[21]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11]);
  assign t[21] = t[13] ^ t[22];
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34] & ~t[35]);
  assign t[31] = (t[36] & ~t[37]);
  assign t[32] = (t[38] & ~t[39]);
  assign t[33] = (t[40] & ~t[41]);
  assign t[34] = t[42] ^ x[2];
  assign t[35] = t[43] ^ x[1];
  assign t[36] = t[44] ^ x[5];
  assign t[37] = t[45] ^ x[4];
  assign t[38] = t[46] ^ x[8];
  assign t[39] = t[47] ^ x[7];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[11];
  assign t[41] = t[49] ^ x[10];
  assign t[42] = (x[0]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[3]);
  assign t[46] = (x[6]);
  assign t[47] = (x[6]);
  assign t[48] = (x[9]);
  assign t[49] = (x[9]);
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[11] ^ t[9];
  assign t[6] = t[12] & t[13];
  assign t[7] = t[11] ^ t[22];
  assign t[8] = t[14] & t[15];
  assign t[9] = ~(t[23]);
  assign y = (t[0]);
endmodule

module R2ind251(x, y);
 input [11:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[24] ^ t[22];
  assign t[12] = ~(t[22]);
  assign t[13] = t[11] ^ t[25];
  assign t[14] = ~(t[7] ^ t[16]);
  assign t[15] = t[17] ^ t[13];
  assign t[16] = t[18] ^ t[6];
  assign t[17] = t[22] ^ t[9];
  assign t[18] = t[19] & t[20];
  assign t[19] = ~(t[21]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11]);
  assign t[21] = t[13] ^ t[22];
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34] & ~t[35]);
  assign t[31] = (t[36] & ~t[37]);
  assign t[32] = (t[38] & ~t[39]);
  assign t[33] = (t[40] & ~t[41]);
  assign t[34] = t[42] ^ x[2];
  assign t[35] = t[43] ^ x[1];
  assign t[36] = t[44] ^ x[5];
  assign t[37] = t[45] ^ x[4];
  assign t[38] = t[46] ^ x[8];
  assign t[39] = t[47] ^ x[7];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[11];
  assign t[41] = t[49] ^ x[10];
  assign t[42] = (x[0]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[3]);
  assign t[46] = (x[6]);
  assign t[47] = (x[6]);
  assign t[48] = (x[9]);
  assign t[49] = (x[9]);
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[11] ^ t[9];
  assign t[6] = t[12] & t[13];
  assign t[7] = t[11] ^ t[22];
  assign t[8] = t[14] & t[15];
  assign t[9] = ~(t[23]);
  assign y = (t[0]);
endmodule

module R2ind252(x, y);
 input [11:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[15] ^ t[29];
  assign t[12] = t[20] & t[21];
  assign t[13] = ~(t[30]);
  assign t[14] = t[18] ^ t[12];
  assign t[15] = t[31] ^ t[29];
  assign t[16] = ~(t[29]);
  assign t[17] = t[15] ^ t[32];
  assign t[18] = t[22] ^ t[8];
  assign t[19] = t[23] & t[24];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11] ^ t[18]);
  assign t[21] = t[9] ^ t[17];
  assign t[22] = t[25] & t[26];
  assign t[23] = ~(t[22] ^ t[27]);
  assign t[24] = t[7] ^ t[28];
  assign t[25] = ~(t[28]);
  assign t[26] = ~(t[15]);
  assign t[27] = t[9] ^ t[15];
  assign t[28] = t[17] ^ t[29];
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = (t[35]);
  assign t[32] = (t[36]);
  assign t[33] = t[37] ^ x[2];
  assign t[34] = t[38] ^ x[5];
  assign t[35] = t[39] ^ x[8];
  assign t[36] = t[40] ^ x[11];
  assign t[37] = (t[41] & ~t[42]);
  assign t[38] = (t[43] & ~t[44]);
  assign t[39] = (t[45] & ~t[46]);
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (t[47] & ~t[48]);
  assign t[41] = t[49] ^ x[2];
  assign t[42] = t[50] ^ x[1];
  assign t[43] = t[51] ^ x[5];
  assign t[44] = t[52] ^ x[4];
  assign t[45] = t[53] ^ x[8];
  assign t[46] = t[54] ^ x[7];
  assign t[47] = t[55] ^ x[11];
  assign t[48] = t[56] ^ x[10];
  assign t[49] = (x[0]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[0]);
  assign t[51] = (x[3]);
  assign t[52] = (x[3]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[9]);
  assign t[56] = (x[9]);
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[15] ^ t[13];
  assign t[8] = t[16] & t[17];
  assign t[9] = t[29] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind253(x, y);
 input [11:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[15] ^ t[29];
  assign t[12] = t[20] & t[21];
  assign t[13] = ~(t[30]);
  assign t[14] = t[18] ^ t[12];
  assign t[15] = t[31] ^ t[29];
  assign t[16] = ~(t[29]);
  assign t[17] = t[15] ^ t[32];
  assign t[18] = t[22] ^ t[8];
  assign t[19] = t[23] & t[24];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11] ^ t[18]);
  assign t[21] = t[9] ^ t[17];
  assign t[22] = t[25] & t[26];
  assign t[23] = ~(t[22] ^ t[27]);
  assign t[24] = t[7] ^ t[28];
  assign t[25] = ~(t[28]);
  assign t[26] = ~(t[15]);
  assign t[27] = t[9] ^ t[15];
  assign t[28] = t[17] ^ t[29];
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = (t[35]);
  assign t[32] = (t[36]);
  assign t[33] = t[37] ^ x[2];
  assign t[34] = t[38] ^ x[5];
  assign t[35] = t[39] ^ x[8];
  assign t[36] = t[40] ^ x[11];
  assign t[37] = (t[41] & ~t[42]);
  assign t[38] = (t[43] & ~t[44]);
  assign t[39] = (t[45] & ~t[46]);
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (t[47] & ~t[48]);
  assign t[41] = t[49] ^ x[2];
  assign t[42] = t[50] ^ x[1];
  assign t[43] = t[51] ^ x[5];
  assign t[44] = t[52] ^ x[4];
  assign t[45] = t[53] ^ x[8];
  assign t[46] = t[54] ^ x[7];
  assign t[47] = t[55] ^ x[11];
  assign t[48] = t[56] ^ x[10];
  assign t[49] = (x[0]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[0]);
  assign t[51] = (x[3]);
  assign t[52] = (x[3]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[9]);
  assign t[56] = (x[9]);
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[15] ^ t[13];
  assign t[8] = t[16] & t[17];
  assign t[9] = t[29] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind254(x, y);
 input [11:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] ^ t[16];
  assign t[11] = t[17] ^ t[8];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[29] ^ t[28];
  assign t[14] = ~(t[28]);
  assign t[15] = t[13] ^ t[30];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[22] & t[23];
  assign t[18] = ~(t[24] ^ t[11]);
  assign t[19] = t[9] ^ t[15];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[17] ^ t[25]);
  assign t[21] = t[7] ^ t[26];
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[13]);
  assign t[24] = t[13] ^ t[28];
  assign t[25] = t[9] ^ t[13];
  assign t[26] = t[15] ^ t[28];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[2];
  assign t[32] = t[36] ^ x[5];
  assign t[33] = t[37] ^ x[8];
  assign t[34] = t[38] ^ x[11];
  assign t[35] = (t[39] & ~t[40]);
  assign t[36] = (t[41] & ~t[42]);
  assign t[37] = (t[43] & ~t[44]);
  assign t[38] = (t[45] & ~t[46]);
  assign t[39] = t[47] ^ x[2];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[1];
  assign t[41] = t[49] ^ x[5];
  assign t[42] = t[50] ^ x[4];
  assign t[43] = t[51] ^ x[8];
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[11];
  assign t[46] = t[54] ^ x[10];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[5] = ~(t[27]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[13] ^ t[5];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[28] ^ t[5];
  assign y = (t[0]);
endmodule

module R2ind255(x, y);
 input [11:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] ^ t[16];
  assign t[11] = t[17] ^ t[8];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[29] ^ t[28];
  assign t[14] = ~(t[28]);
  assign t[15] = t[13] ^ t[30];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[22] & t[23];
  assign t[18] = ~(t[24] ^ t[11]);
  assign t[19] = t[9] ^ t[15];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[17] ^ t[25]);
  assign t[21] = t[7] ^ t[26];
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[13]);
  assign t[24] = t[13] ^ t[28];
  assign t[25] = t[9] ^ t[13];
  assign t[26] = t[15] ^ t[28];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[2];
  assign t[32] = t[36] ^ x[5];
  assign t[33] = t[37] ^ x[8];
  assign t[34] = t[38] ^ x[11];
  assign t[35] = (t[39] & ~t[40]);
  assign t[36] = (t[41] & ~t[42]);
  assign t[37] = (t[43] & ~t[44]);
  assign t[38] = (t[45] & ~t[46]);
  assign t[39] = t[47] ^ x[2];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[1];
  assign t[41] = t[49] ^ x[5];
  assign t[42] = t[50] ^ x[4];
  assign t[43] = t[51] ^ x[8];
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[11];
  assign t[46] = t[54] ^ x[10];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[5] = ~(t[27]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[13] ^ t[5];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[28] ^ t[5];
  assign y = (t[0]);
endmodule

module R2ind256(x, y);
 input [11:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[7] ^ t[23];
  assign t[11] = t[13] ^ t[4];
  assign t[12] = t[14] & t[15];
  assign t[13] = t[16] & t[17];
  assign t[14] = ~(t[13] ^ t[18]);
  assign t[15] = t[3] ^ t[19];
  assign t[16] = ~(t[19]);
  assign t[17] = ~(t[7]);
  assign t[18] = t[5] ^ t[7];
  assign t[19] = t[10] ^ t[20];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = t[28] ^ x[2];
  assign t[25] = t[29] ^ x[5];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = t[31] ^ x[11];
  assign t[28] = (t[32] & ~t[33]);
  assign t[29] = (t[34] & ~t[35]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[36] & ~t[37]);
  assign t[31] = (t[38] & ~t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[1];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[4];
  assign t[36] = t[44] ^ x[8];
  assign t[37] = t[45] ^ x[7];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[10];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[4] = t[9] & t[10];
  assign t[5] = t[20] ^ t[8];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[21] ^ t[20];
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind257(x, y);
 input [11:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[7] ^ t[23];
  assign t[11] = t[13] ^ t[4];
  assign t[12] = t[14] & t[15];
  assign t[13] = t[16] & t[17];
  assign t[14] = ~(t[13] ^ t[18]);
  assign t[15] = t[3] ^ t[19];
  assign t[16] = ~(t[19]);
  assign t[17] = ~(t[7]);
  assign t[18] = t[5] ^ t[7];
  assign t[19] = t[10] ^ t[20];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = t[28] ^ x[2];
  assign t[25] = t[29] ^ x[5];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = t[31] ^ x[11];
  assign t[28] = (t[32] & ~t[33]);
  assign t[29] = (t[34] & ~t[35]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[36] & ~t[37]);
  assign t[31] = (t[38] & ~t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[1];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[4];
  assign t[36] = t[44] ^ x[8];
  assign t[37] = t[45] ^ x[7];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[10];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[4] = t[9] & t[10];
  assign t[5] = t[20] ^ t[8];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[21] ^ t[20];
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind258(x, y);
 input [11:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[24] ^ t[22];
  assign t[12] = ~(t[22]);
  assign t[13] = t[11] ^ t[25];
  assign t[14] = ~(t[7] ^ t[16]);
  assign t[15] = t[17] ^ t[13];
  assign t[16] = t[18] ^ t[6];
  assign t[17] = t[22] ^ t[9];
  assign t[18] = t[19] & t[20];
  assign t[19] = ~(t[21]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11]);
  assign t[21] = t[13] ^ t[22];
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34] & ~t[35]);
  assign t[31] = (t[36] & ~t[37]);
  assign t[32] = (t[38] & ~t[39]);
  assign t[33] = (t[40] & ~t[41]);
  assign t[34] = t[42] ^ x[2];
  assign t[35] = t[43] ^ x[1];
  assign t[36] = t[44] ^ x[5];
  assign t[37] = t[45] ^ x[4];
  assign t[38] = t[46] ^ x[8];
  assign t[39] = t[47] ^ x[7];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[11];
  assign t[41] = t[49] ^ x[10];
  assign t[42] = (x[0]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[3]);
  assign t[46] = (x[6]);
  assign t[47] = (x[6]);
  assign t[48] = (x[9]);
  assign t[49] = (x[9]);
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[11] ^ t[9];
  assign t[6] = t[12] & t[13];
  assign t[7] = t[11] ^ t[22];
  assign t[8] = t[14] & t[15];
  assign t[9] = ~(t[23]);
  assign y = (t[0]);
endmodule

module R2ind259(x, y);
 input [11:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[24] ^ t[22];
  assign t[12] = ~(t[22]);
  assign t[13] = t[11] ^ t[25];
  assign t[14] = ~(t[7] ^ t[16]);
  assign t[15] = t[17] ^ t[13];
  assign t[16] = t[18] ^ t[6];
  assign t[17] = t[22] ^ t[9];
  assign t[18] = t[19] & t[20];
  assign t[19] = ~(t[21]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11]);
  assign t[21] = t[13] ^ t[22];
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34] & ~t[35]);
  assign t[31] = (t[36] & ~t[37]);
  assign t[32] = (t[38] & ~t[39]);
  assign t[33] = (t[40] & ~t[41]);
  assign t[34] = t[42] ^ x[2];
  assign t[35] = t[43] ^ x[1];
  assign t[36] = t[44] ^ x[5];
  assign t[37] = t[45] ^ x[4];
  assign t[38] = t[46] ^ x[8];
  assign t[39] = t[47] ^ x[7];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[11];
  assign t[41] = t[49] ^ x[10];
  assign t[42] = (x[0]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[3]);
  assign t[46] = (x[6]);
  assign t[47] = (x[6]);
  assign t[48] = (x[9]);
  assign t[49] = (x[9]);
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[11] ^ t[9];
  assign t[6] = t[12] & t[13];
  assign t[7] = t[11] ^ t[22];
  assign t[8] = t[14] & t[15];
  assign t[9] = ~(t[23]);
  assign y = (t[0]);
endmodule

module R2ind260(x, y);
 input [11:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[15] ^ t[29];
  assign t[12] = t[20] & t[21];
  assign t[13] = ~(t[30]);
  assign t[14] = t[18] ^ t[12];
  assign t[15] = t[31] ^ t[29];
  assign t[16] = ~(t[29]);
  assign t[17] = t[15] ^ t[32];
  assign t[18] = t[22] ^ t[8];
  assign t[19] = t[23] & t[24];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11] ^ t[18]);
  assign t[21] = t[9] ^ t[17];
  assign t[22] = t[25] & t[26];
  assign t[23] = ~(t[22] ^ t[27]);
  assign t[24] = t[7] ^ t[28];
  assign t[25] = ~(t[28]);
  assign t[26] = ~(t[15]);
  assign t[27] = t[9] ^ t[15];
  assign t[28] = t[17] ^ t[29];
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = (t[35]);
  assign t[32] = (t[36]);
  assign t[33] = t[37] ^ x[2];
  assign t[34] = t[38] ^ x[5];
  assign t[35] = t[39] ^ x[8];
  assign t[36] = t[40] ^ x[11];
  assign t[37] = (t[41] & ~t[42]);
  assign t[38] = (t[43] & ~t[44]);
  assign t[39] = (t[45] & ~t[46]);
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (t[47] & ~t[48]);
  assign t[41] = t[49] ^ x[2];
  assign t[42] = t[50] ^ x[1];
  assign t[43] = t[51] ^ x[5];
  assign t[44] = t[52] ^ x[4];
  assign t[45] = t[53] ^ x[8];
  assign t[46] = t[54] ^ x[7];
  assign t[47] = t[55] ^ x[11];
  assign t[48] = t[56] ^ x[10];
  assign t[49] = (x[0]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[0]);
  assign t[51] = (x[3]);
  assign t[52] = (x[3]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[9]);
  assign t[56] = (x[9]);
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[15] ^ t[13];
  assign t[8] = t[16] & t[17];
  assign t[9] = t[29] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind261(x, y);
 input [11:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[15] ^ t[29];
  assign t[12] = t[20] & t[21];
  assign t[13] = ~(t[30]);
  assign t[14] = t[18] ^ t[12];
  assign t[15] = t[31] ^ t[29];
  assign t[16] = ~(t[29]);
  assign t[17] = t[15] ^ t[32];
  assign t[18] = t[22] ^ t[8];
  assign t[19] = t[23] & t[24];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11] ^ t[18]);
  assign t[21] = t[9] ^ t[17];
  assign t[22] = t[25] & t[26];
  assign t[23] = ~(t[22] ^ t[27]);
  assign t[24] = t[7] ^ t[28];
  assign t[25] = ~(t[28]);
  assign t[26] = ~(t[15]);
  assign t[27] = t[9] ^ t[15];
  assign t[28] = t[17] ^ t[29];
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = (t[35]);
  assign t[32] = (t[36]);
  assign t[33] = t[37] ^ x[2];
  assign t[34] = t[38] ^ x[5];
  assign t[35] = t[39] ^ x[8];
  assign t[36] = t[40] ^ x[11];
  assign t[37] = (t[41] & ~t[42]);
  assign t[38] = (t[43] & ~t[44]);
  assign t[39] = (t[45] & ~t[46]);
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (t[47] & ~t[48]);
  assign t[41] = t[49] ^ x[2];
  assign t[42] = t[50] ^ x[1];
  assign t[43] = t[51] ^ x[5];
  assign t[44] = t[52] ^ x[4];
  assign t[45] = t[53] ^ x[8];
  assign t[46] = t[54] ^ x[7];
  assign t[47] = t[55] ^ x[11];
  assign t[48] = t[56] ^ x[10];
  assign t[49] = (x[0]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[0]);
  assign t[51] = (x[3]);
  assign t[52] = (x[3]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[9]);
  assign t[56] = (x[9]);
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[15] ^ t[13];
  assign t[8] = t[16] & t[17];
  assign t[9] = t[29] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind262(x, y);
 input [11:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] ^ t[16];
  assign t[11] = t[17] ^ t[8];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[29] ^ t[28];
  assign t[14] = ~(t[28]);
  assign t[15] = t[13] ^ t[30];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[22] & t[23];
  assign t[18] = ~(t[24] ^ t[11]);
  assign t[19] = t[9] ^ t[15];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[17] ^ t[25]);
  assign t[21] = t[7] ^ t[26];
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[13]);
  assign t[24] = t[13] ^ t[28];
  assign t[25] = t[9] ^ t[13];
  assign t[26] = t[15] ^ t[28];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[2];
  assign t[32] = t[36] ^ x[5];
  assign t[33] = t[37] ^ x[8];
  assign t[34] = t[38] ^ x[11];
  assign t[35] = (t[39] & ~t[40]);
  assign t[36] = (t[41] & ~t[42]);
  assign t[37] = (t[43] & ~t[44]);
  assign t[38] = (t[45] & ~t[46]);
  assign t[39] = t[47] ^ x[2];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[1];
  assign t[41] = t[49] ^ x[5];
  assign t[42] = t[50] ^ x[4];
  assign t[43] = t[51] ^ x[8];
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[11];
  assign t[46] = t[54] ^ x[10];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[5] = ~(t[27]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[13] ^ t[5];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[28] ^ t[5];
  assign y = (t[0]);
endmodule

module R2ind263(x, y);
 input [11:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] ^ t[16];
  assign t[11] = t[17] ^ t[8];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[29] ^ t[28];
  assign t[14] = ~(t[28]);
  assign t[15] = t[13] ^ t[30];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[22] & t[23];
  assign t[18] = ~(t[24] ^ t[11]);
  assign t[19] = t[9] ^ t[15];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[17] ^ t[25]);
  assign t[21] = t[7] ^ t[26];
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[13]);
  assign t[24] = t[13] ^ t[28];
  assign t[25] = t[9] ^ t[13];
  assign t[26] = t[15] ^ t[28];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[2];
  assign t[32] = t[36] ^ x[5];
  assign t[33] = t[37] ^ x[8];
  assign t[34] = t[38] ^ x[11];
  assign t[35] = (t[39] & ~t[40]);
  assign t[36] = (t[41] & ~t[42]);
  assign t[37] = (t[43] & ~t[44]);
  assign t[38] = (t[45] & ~t[46]);
  assign t[39] = t[47] ^ x[2];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[1];
  assign t[41] = t[49] ^ x[5];
  assign t[42] = t[50] ^ x[4];
  assign t[43] = t[51] ^ x[8];
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[11];
  assign t[46] = t[54] ^ x[10];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[5] = ~(t[27]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[13] ^ t[5];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[28] ^ t[5];
  assign y = (t[0]);
endmodule

module R2ind264(x, y);
 input [11:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[7] ^ t[23];
  assign t[11] = t[13] ^ t[4];
  assign t[12] = t[14] & t[15];
  assign t[13] = t[16] & t[17];
  assign t[14] = ~(t[13] ^ t[18]);
  assign t[15] = t[3] ^ t[19];
  assign t[16] = ~(t[19]);
  assign t[17] = ~(t[7]);
  assign t[18] = t[5] ^ t[7];
  assign t[19] = t[10] ^ t[20];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = t[28] ^ x[2];
  assign t[25] = t[29] ^ x[5];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = t[31] ^ x[11];
  assign t[28] = (t[32] & ~t[33]);
  assign t[29] = (t[34] & ~t[35]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[36] & ~t[37]);
  assign t[31] = (t[38] & ~t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[1];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[4];
  assign t[36] = t[44] ^ x[8];
  assign t[37] = t[45] ^ x[7];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[10];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[4] = t[9] & t[10];
  assign t[5] = t[20] ^ t[8];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[21] ^ t[20];
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind265(x, y);
 input [11:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[7] ^ t[23];
  assign t[11] = t[13] ^ t[4];
  assign t[12] = t[14] & t[15];
  assign t[13] = t[16] & t[17];
  assign t[14] = ~(t[13] ^ t[18]);
  assign t[15] = t[3] ^ t[19];
  assign t[16] = ~(t[19]);
  assign t[17] = ~(t[7]);
  assign t[18] = t[5] ^ t[7];
  assign t[19] = t[10] ^ t[20];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = t[28] ^ x[2];
  assign t[25] = t[29] ^ x[5];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = t[31] ^ x[11];
  assign t[28] = (t[32] & ~t[33]);
  assign t[29] = (t[34] & ~t[35]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[36] & ~t[37]);
  assign t[31] = (t[38] & ~t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[1];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[4];
  assign t[36] = t[44] ^ x[8];
  assign t[37] = t[45] ^ x[7];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[10];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[4] = t[9] & t[10];
  assign t[5] = t[20] ^ t[8];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[21] ^ t[20];
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind266(x, y);
 input [11:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[24] ^ t[22];
  assign t[12] = ~(t[22]);
  assign t[13] = t[11] ^ t[25];
  assign t[14] = ~(t[7] ^ t[16]);
  assign t[15] = t[17] ^ t[13];
  assign t[16] = t[18] ^ t[6];
  assign t[17] = t[22] ^ t[9];
  assign t[18] = t[19] & t[20];
  assign t[19] = ~(t[21]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11]);
  assign t[21] = t[13] ^ t[22];
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34] & ~t[35]);
  assign t[31] = (t[36] & ~t[37]);
  assign t[32] = (t[38] & ~t[39]);
  assign t[33] = (t[40] & ~t[41]);
  assign t[34] = t[42] ^ x[2];
  assign t[35] = t[43] ^ x[1];
  assign t[36] = t[44] ^ x[5];
  assign t[37] = t[45] ^ x[4];
  assign t[38] = t[46] ^ x[8];
  assign t[39] = t[47] ^ x[7];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[11];
  assign t[41] = t[49] ^ x[10];
  assign t[42] = (x[0]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[3]);
  assign t[46] = (x[6]);
  assign t[47] = (x[6]);
  assign t[48] = (x[9]);
  assign t[49] = (x[9]);
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[11] ^ t[9];
  assign t[6] = t[12] & t[13];
  assign t[7] = t[11] ^ t[22];
  assign t[8] = t[14] & t[15];
  assign t[9] = ~(t[23]);
  assign y = (t[0]);
endmodule

module R2ind267(x, y);
 input [11:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[24] ^ t[22];
  assign t[12] = ~(t[22]);
  assign t[13] = t[11] ^ t[25];
  assign t[14] = ~(t[7] ^ t[16]);
  assign t[15] = t[17] ^ t[13];
  assign t[16] = t[18] ^ t[6];
  assign t[17] = t[22] ^ t[9];
  assign t[18] = t[19] & t[20];
  assign t[19] = ~(t[21]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11]);
  assign t[21] = t[13] ^ t[22];
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34] & ~t[35]);
  assign t[31] = (t[36] & ~t[37]);
  assign t[32] = (t[38] & ~t[39]);
  assign t[33] = (t[40] & ~t[41]);
  assign t[34] = t[42] ^ x[2];
  assign t[35] = t[43] ^ x[1];
  assign t[36] = t[44] ^ x[5];
  assign t[37] = t[45] ^ x[4];
  assign t[38] = t[46] ^ x[8];
  assign t[39] = t[47] ^ x[7];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[11];
  assign t[41] = t[49] ^ x[10];
  assign t[42] = (x[0]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[3]);
  assign t[46] = (x[6]);
  assign t[47] = (x[6]);
  assign t[48] = (x[9]);
  assign t[49] = (x[9]);
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[11] ^ t[9];
  assign t[6] = t[12] & t[13];
  assign t[7] = t[11] ^ t[22];
  assign t[8] = t[14] & t[15];
  assign t[9] = ~(t[23]);
  assign y = (t[0]);
endmodule

module R2ind268(x, y);
 input [11:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[15] ^ t[29];
  assign t[12] = t[20] & t[21];
  assign t[13] = ~(t[30]);
  assign t[14] = t[18] ^ t[12];
  assign t[15] = t[31] ^ t[29];
  assign t[16] = ~(t[29]);
  assign t[17] = t[15] ^ t[32];
  assign t[18] = t[22] ^ t[8];
  assign t[19] = t[23] & t[24];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11] ^ t[18]);
  assign t[21] = t[9] ^ t[17];
  assign t[22] = t[25] & t[26];
  assign t[23] = ~(t[22] ^ t[27]);
  assign t[24] = t[7] ^ t[28];
  assign t[25] = ~(t[28]);
  assign t[26] = ~(t[15]);
  assign t[27] = t[9] ^ t[15];
  assign t[28] = t[17] ^ t[29];
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = (t[35]);
  assign t[32] = (t[36]);
  assign t[33] = t[37] ^ x[2];
  assign t[34] = t[38] ^ x[5];
  assign t[35] = t[39] ^ x[8];
  assign t[36] = t[40] ^ x[11];
  assign t[37] = (t[41] & ~t[42]);
  assign t[38] = (t[43] & ~t[44]);
  assign t[39] = (t[45] & ~t[46]);
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (t[47] & ~t[48]);
  assign t[41] = t[49] ^ x[2];
  assign t[42] = t[50] ^ x[1];
  assign t[43] = t[51] ^ x[5];
  assign t[44] = t[52] ^ x[4];
  assign t[45] = t[53] ^ x[8];
  assign t[46] = t[54] ^ x[7];
  assign t[47] = t[55] ^ x[11];
  assign t[48] = t[56] ^ x[10];
  assign t[49] = (x[0]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[0]);
  assign t[51] = (x[3]);
  assign t[52] = (x[3]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[9]);
  assign t[56] = (x[9]);
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[15] ^ t[13];
  assign t[8] = t[16] & t[17];
  assign t[9] = t[29] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind269(x, y);
 input [11:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[15] ^ t[29];
  assign t[12] = t[20] & t[21];
  assign t[13] = ~(t[30]);
  assign t[14] = t[18] ^ t[12];
  assign t[15] = t[31] ^ t[29];
  assign t[16] = ~(t[29]);
  assign t[17] = t[15] ^ t[32];
  assign t[18] = t[22] ^ t[8];
  assign t[19] = t[23] & t[24];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11] ^ t[18]);
  assign t[21] = t[9] ^ t[17];
  assign t[22] = t[25] & t[26];
  assign t[23] = ~(t[22] ^ t[27]);
  assign t[24] = t[7] ^ t[28];
  assign t[25] = ~(t[28]);
  assign t[26] = ~(t[15]);
  assign t[27] = t[9] ^ t[15];
  assign t[28] = t[17] ^ t[29];
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = (t[35]);
  assign t[32] = (t[36]);
  assign t[33] = t[37] ^ x[2];
  assign t[34] = t[38] ^ x[5];
  assign t[35] = t[39] ^ x[8];
  assign t[36] = t[40] ^ x[11];
  assign t[37] = (t[41] & ~t[42]);
  assign t[38] = (t[43] & ~t[44]);
  assign t[39] = (t[45] & ~t[46]);
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (t[47] & ~t[48]);
  assign t[41] = t[49] ^ x[2];
  assign t[42] = t[50] ^ x[1];
  assign t[43] = t[51] ^ x[5];
  assign t[44] = t[52] ^ x[4];
  assign t[45] = t[53] ^ x[8];
  assign t[46] = t[54] ^ x[7];
  assign t[47] = t[55] ^ x[11];
  assign t[48] = t[56] ^ x[10];
  assign t[49] = (x[0]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[0]);
  assign t[51] = (x[3]);
  assign t[52] = (x[3]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[9]);
  assign t[56] = (x[9]);
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[15] ^ t[13];
  assign t[8] = t[16] & t[17];
  assign t[9] = t[29] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind270(x, y);
 input [11:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] ^ t[16];
  assign t[11] = t[17] ^ t[8];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[29] ^ t[28];
  assign t[14] = ~(t[28]);
  assign t[15] = t[13] ^ t[30];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[22] & t[23];
  assign t[18] = ~(t[24] ^ t[11]);
  assign t[19] = t[9] ^ t[15];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[17] ^ t[25]);
  assign t[21] = t[7] ^ t[26];
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[13]);
  assign t[24] = t[13] ^ t[28];
  assign t[25] = t[9] ^ t[13];
  assign t[26] = t[15] ^ t[28];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[2];
  assign t[32] = t[36] ^ x[5];
  assign t[33] = t[37] ^ x[8];
  assign t[34] = t[38] ^ x[11];
  assign t[35] = (t[39] & ~t[40]);
  assign t[36] = (t[41] & ~t[42]);
  assign t[37] = (t[43] & ~t[44]);
  assign t[38] = (t[45] & ~t[46]);
  assign t[39] = t[47] ^ x[2];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[1];
  assign t[41] = t[49] ^ x[5];
  assign t[42] = t[50] ^ x[4];
  assign t[43] = t[51] ^ x[8];
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[11];
  assign t[46] = t[54] ^ x[10];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[5] = ~(t[27]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[13] ^ t[5];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[28] ^ t[5];
  assign y = (t[0]);
endmodule

module R2ind271(x, y);
 input [11:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] ^ t[16];
  assign t[11] = t[17] ^ t[8];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[29] ^ t[28];
  assign t[14] = ~(t[28]);
  assign t[15] = t[13] ^ t[30];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[22] & t[23];
  assign t[18] = ~(t[24] ^ t[11]);
  assign t[19] = t[9] ^ t[15];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[17] ^ t[25]);
  assign t[21] = t[7] ^ t[26];
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[13]);
  assign t[24] = t[13] ^ t[28];
  assign t[25] = t[9] ^ t[13];
  assign t[26] = t[15] ^ t[28];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[2];
  assign t[32] = t[36] ^ x[5];
  assign t[33] = t[37] ^ x[8];
  assign t[34] = t[38] ^ x[11];
  assign t[35] = (t[39] & ~t[40]);
  assign t[36] = (t[41] & ~t[42]);
  assign t[37] = (t[43] & ~t[44]);
  assign t[38] = (t[45] & ~t[46]);
  assign t[39] = t[47] ^ x[2];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[1];
  assign t[41] = t[49] ^ x[5];
  assign t[42] = t[50] ^ x[4];
  assign t[43] = t[51] ^ x[8];
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[11];
  assign t[46] = t[54] ^ x[10];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[5] = ~(t[27]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[13] ^ t[5];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[28] ^ t[5];
  assign y = (t[0]);
endmodule

module R2ind272(x, y);
 input [11:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[7] ^ t[23];
  assign t[11] = t[13] ^ t[4];
  assign t[12] = t[14] & t[15];
  assign t[13] = t[16] & t[17];
  assign t[14] = ~(t[13] ^ t[18]);
  assign t[15] = t[3] ^ t[19];
  assign t[16] = ~(t[19]);
  assign t[17] = ~(t[7]);
  assign t[18] = t[5] ^ t[7];
  assign t[19] = t[10] ^ t[20];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = t[28] ^ x[2];
  assign t[25] = t[29] ^ x[5];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = t[31] ^ x[11];
  assign t[28] = (t[32] & ~t[33]);
  assign t[29] = (t[34] & ~t[35]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[36] & ~t[37]);
  assign t[31] = (t[38] & ~t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[1];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[4];
  assign t[36] = t[44] ^ x[8];
  assign t[37] = t[45] ^ x[7];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[10];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[4] = t[9] & t[10];
  assign t[5] = t[20] ^ t[8];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[21] ^ t[20];
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind273(x, y);
 input [11:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[7] ^ t[23];
  assign t[11] = t[13] ^ t[4];
  assign t[12] = t[14] & t[15];
  assign t[13] = t[16] & t[17];
  assign t[14] = ~(t[13] ^ t[18]);
  assign t[15] = t[3] ^ t[19];
  assign t[16] = ~(t[19]);
  assign t[17] = ~(t[7]);
  assign t[18] = t[5] ^ t[7];
  assign t[19] = t[10] ^ t[20];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = t[28] ^ x[2];
  assign t[25] = t[29] ^ x[5];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = t[31] ^ x[11];
  assign t[28] = (t[32] & ~t[33]);
  assign t[29] = (t[34] & ~t[35]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[36] & ~t[37]);
  assign t[31] = (t[38] & ~t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[1];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[4];
  assign t[36] = t[44] ^ x[8];
  assign t[37] = t[45] ^ x[7];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[10];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[4] = t[9] & t[10];
  assign t[5] = t[20] ^ t[8];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[21] ^ t[20];
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind274(x, y);
 input [11:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[24] ^ t[22];
  assign t[12] = ~(t[22]);
  assign t[13] = t[11] ^ t[25];
  assign t[14] = ~(t[7] ^ t[16]);
  assign t[15] = t[17] ^ t[13];
  assign t[16] = t[18] ^ t[6];
  assign t[17] = t[22] ^ t[9];
  assign t[18] = t[19] & t[20];
  assign t[19] = ~(t[21]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11]);
  assign t[21] = t[13] ^ t[22];
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34] & ~t[35]);
  assign t[31] = (t[36] & ~t[37]);
  assign t[32] = (t[38] & ~t[39]);
  assign t[33] = (t[40] & ~t[41]);
  assign t[34] = t[42] ^ x[2];
  assign t[35] = t[43] ^ x[1];
  assign t[36] = t[44] ^ x[5];
  assign t[37] = t[45] ^ x[4];
  assign t[38] = t[46] ^ x[8];
  assign t[39] = t[47] ^ x[7];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[11];
  assign t[41] = t[49] ^ x[10];
  assign t[42] = (x[0]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[3]);
  assign t[46] = (x[6]);
  assign t[47] = (x[6]);
  assign t[48] = (x[9]);
  assign t[49] = (x[9]);
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[11] ^ t[9];
  assign t[6] = t[12] & t[13];
  assign t[7] = t[11] ^ t[22];
  assign t[8] = t[14] & t[15];
  assign t[9] = ~(t[23]);
  assign y = (t[0]);
endmodule

module R2ind275(x, y);
 input [11:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[24] ^ t[22];
  assign t[12] = ~(t[22]);
  assign t[13] = t[11] ^ t[25];
  assign t[14] = ~(t[7] ^ t[16]);
  assign t[15] = t[17] ^ t[13];
  assign t[16] = t[18] ^ t[6];
  assign t[17] = t[22] ^ t[9];
  assign t[18] = t[19] & t[20];
  assign t[19] = ~(t[21]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11]);
  assign t[21] = t[13] ^ t[22];
  assign t[22] = (t[26]);
  assign t[23] = (t[27]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = t[30] ^ x[2];
  assign t[27] = t[31] ^ x[5];
  assign t[28] = t[32] ^ x[8];
  assign t[29] = t[33] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34] & ~t[35]);
  assign t[31] = (t[36] & ~t[37]);
  assign t[32] = (t[38] & ~t[39]);
  assign t[33] = (t[40] & ~t[41]);
  assign t[34] = t[42] ^ x[2];
  assign t[35] = t[43] ^ x[1];
  assign t[36] = t[44] ^ x[5];
  assign t[37] = t[45] ^ x[4];
  assign t[38] = t[46] ^ x[8];
  assign t[39] = t[47] ^ x[7];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[11];
  assign t[41] = t[49] ^ x[10];
  assign t[42] = (x[0]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[3]);
  assign t[46] = (x[6]);
  assign t[47] = (x[6]);
  assign t[48] = (x[9]);
  assign t[49] = (x[9]);
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[11] ^ t[9];
  assign t[6] = t[12] & t[13];
  assign t[7] = t[11] ^ t[22];
  assign t[8] = t[14] & t[15];
  assign t[9] = ~(t[23]);
  assign y = (t[0]);
endmodule

module R2ind276(x, y);
 input [11:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[15] ^ t[29];
  assign t[12] = t[20] & t[21];
  assign t[13] = ~(t[30]);
  assign t[14] = t[18] ^ t[12];
  assign t[15] = t[31] ^ t[29];
  assign t[16] = ~(t[29]);
  assign t[17] = t[15] ^ t[32];
  assign t[18] = t[22] ^ t[8];
  assign t[19] = t[23] & t[24];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11] ^ t[18]);
  assign t[21] = t[9] ^ t[17];
  assign t[22] = t[25] & t[26];
  assign t[23] = ~(t[22] ^ t[27]);
  assign t[24] = t[7] ^ t[28];
  assign t[25] = ~(t[28]);
  assign t[26] = ~(t[15]);
  assign t[27] = t[9] ^ t[15];
  assign t[28] = t[17] ^ t[29];
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = (t[35]);
  assign t[32] = (t[36]);
  assign t[33] = t[37] ^ x[2];
  assign t[34] = t[38] ^ x[5];
  assign t[35] = t[39] ^ x[8];
  assign t[36] = t[40] ^ x[11];
  assign t[37] = (t[41] & ~t[42]);
  assign t[38] = (t[43] & ~t[44]);
  assign t[39] = (t[45] & ~t[46]);
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (t[47] & ~t[48]);
  assign t[41] = t[49] ^ x[2];
  assign t[42] = t[50] ^ x[1];
  assign t[43] = t[51] ^ x[5];
  assign t[44] = t[52] ^ x[4];
  assign t[45] = t[53] ^ x[8];
  assign t[46] = t[54] ^ x[7];
  assign t[47] = t[55] ^ x[11];
  assign t[48] = t[56] ^ x[10];
  assign t[49] = (x[0]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[0]);
  assign t[51] = (x[3]);
  assign t[52] = (x[3]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[9]);
  assign t[56] = (x[9]);
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[15] ^ t[13];
  assign t[8] = t[16] & t[17];
  assign t[9] = t[29] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind277(x, y);
 input [11:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[15] ^ t[29];
  assign t[12] = t[20] & t[21];
  assign t[13] = ~(t[30]);
  assign t[14] = t[18] ^ t[12];
  assign t[15] = t[31] ^ t[29];
  assign t[16] = ~(t[29]);
  assign t[17] = t[15] ^ t[32];
  assign t[18] = t[22] ^ t[8];
  assign t[19] = t[23] & t[24];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[11] ^ t[18]);
  assign t[21] = t[9] ^ t[17];
  assign t[22] = t[25] & t[26];
  assign t[23] = ~(t[22] ^ t[27]);
  assign t[24] = t[7] ^ t[28];
  assign t[25] = ~(t[28]);
  assign t[26] = ~(t[15]);
  assign t[27] = t[9] ^ t[15];
  assign t[28] = t[17] ^ t[29];
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = (t[35]);
  assign t[32] = (t[36]);
  assign t[33] = t[37] ^ x[2];
  assign t[34] = t[38] ^ x[5];
  assign t[35] = t[39] ^ x[8];
  assign t[36] = t[40] ^ x[11];
  assign t[37] = (t[41] & ~t[42]);
  assign t[38] = (t[43] & ~t[44]);
  assign t[39] = (t[45] & ~t[46]);
  assign t[3] = t[7] ^ t[8];
  assign t[40] = (t[47] & ~t[48]);
  assign t[41] = t[49] ^ x[2];
  assign t[42] = t[50] ^ x[1];
  assign t[43] = t[51] ^ x[5];
  assign t[44] = t[52] ^ x[4];
  assign t[45] = t[53] ^ x[8];
  assign t[46] = t[54] ^ x[7];
  assign t[47] = t[55] ^ x[11];
  assign t[48] = t[56] ^ x[10];
  assign t[49] = (x[0]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[0]);
  assign t[51] = (x[3]);
  assign t[52] = (x[3]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[9]);
  assign t[56] = (x[9]);
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[15] ^ t[13];
  assign t[8] = t[16] & t[17];
  assign t[9] = t[29] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind278(x, y);
 input [11:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] ^ t[16];
  assign t[11] = t[17] ^ t[8];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[29] ^ t[28];
  assign t[14] = ~(t[28]);
  assign t[15] = t[13] ^ t[30];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[22] & t[23];
  assign t[18] = ~(t[24] ^ t[11]);
  assign t[19] = t[9] ^ t[15];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[17] ^ t[25]);
  assign t[21] = t[7] ^ t[26];
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[13]);
  assign t[24] = t[13] ^ t[28];
  assign t[25] = t[9] ^ t[13];
  assign t[26] = t[15] ^ t[28];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[2];
  assign t[32] = t[36] ^ x[5];
  assign t[33] = t[37] ^ x[8];
  assign t[34] = t[38] ^ x[11];
  assign t[35] = (t[39] & ~t[40]);
  assign t[36] = (t[41] & ~t[42]);
  assign t[37] = (t[43] & ~t[44]);
  assign t[38] = (t[45] & ~t[46]);
  assign t[39] = t[47] ^ x[2];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[1];
  assign t[41] = t[49] ^ x[5];
  assign t[42] = t[50] ^ x[4];
  assign t[43] = t[51] ^ x[8];
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[11];
  assign t[46] = t[54] ^ x[10];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[5] = ~(t[27]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[13] ^ t[5];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[28] ^ t[5];
  assign y = (t[0]);
endmodule

module R2ind279(x, y);
 input [11:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] ^ t[16];
  assign t[11] = t[17] ^ t[8];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[29] ^ t[28];
  assign t[14] = ~(t[28]);
  assign t[15] = t[13] ^ t[30];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[22] & t[23];
  assign t[18] = ~(t[24] ^ t[11]);
  assign t[19] = t[9] ^ t[15];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[17] ^ t[25]);
  assign t[21] = t[7] ^ t[26];
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[13]);
  assign t[24] = t[13] ^ t[28];
  assign t[25] = t[9] ^ t[13];
  assign t[26] = t[15] ^ t[28];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = t[5] ^ t[6];
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[2];
  assign t[32] = t[36] ^ x[5];
  assign t[33] = t[37] ^ x[8];
  assign t[34] = t[38] ^ x[11];
  assign t[35] = (t[39] & ~t[40]);
  assign t[36] = (t[41] & ~t[42]);
  assign t[37] = (t[43] & ~t[44]);
  assign t[38] = (t[45] & ~t[46]);
  assign t[39] = t[47] ^ x[2];
  assign t[3] = t[7] ^ t[8];
  assign t[40] = t[48] ^ x[1];
  assign t[41] = t[49] ^ x[5];
  assign t[42] = t[50] ^ x[4];
  assign t[43] = t[51] ^ x[8];
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[11];
  assign t[46] = t[54] ^ x[10];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = t[9] ^ t[10];
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[5] = ~(t[27]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[13] ^ t[5];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[28] ^ t[5];
  assign y = (t[0]);
endmodule

module R2ind280(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind281(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind282(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind283(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind284(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind285(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind286(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind287(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind288(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind289(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind290(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind291(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind292(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind293(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind294(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind295(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind296(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind297(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind298(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind299(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind300(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind301(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind302(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind303(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind304(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind305(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind306(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind307(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind308(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind309(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind310(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind311(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind312(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind313(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind314(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind315(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind316(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind317(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind318(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind319(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind320(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind321(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind322(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind323(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind324(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind325(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind326(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind327(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind328(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind329(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind330(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind331(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind332(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind333(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind334(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind335(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind336(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind337(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind338(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind339(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind340(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind341(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind342(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind343(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind344(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind345(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind346(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind347(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind348(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind349(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind350(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind351(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind352(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind353(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind354(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind355(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind356(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind357(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind358(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind359(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind360(x, y);
 input [8:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[14] ^ x[1];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[7];
  assign t[13] = (x[0]);
  assign t[14] = (x[0]);
  assign t[15] = (x[6]);
  assign t[16] = (x[6]);
  assign t[1] = t[3] ? x[4] : x[3];
  assign t[2] = ~(~x[5] & ~t[4]);
  assign t[3] = (t[5]);
  assign t[4] = (t[6]);
  assign t[5] = t[7] ^ x[2];
  assign t[6] = t[8] ^ x[8];
  assign t[7] = (t[9] & ~t[10]);
  assign t[8] = (t[11] & ~t[12]);
  assign t[9] = t[13] ^ x[2];
  assign y = (t[0]);
endmodule

module R2ind361(x, y);
 input [8:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[14] ^ x[1];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[7];
  assign t[13] = (x[0]);
  assign t[14] = (x[0]);
  assign t[15] = (x[6]);
  assign t[16] = (x[6]);
  assign t[1] = t[3] ? x[4] : x[3];
  assign t[2] = ~(~x[5] & ~t[4]);
  assign t[3] = (t[5]);
  assign t[4] = (t[6]);
  assign t[5] = t[7] ^ x[2];
  assign t[6] = t[8] ^ x[8];
  assign t[7] = (t[9] & ~t[10]);
  assign t[8] = (t[11] & ~t[12]);
  assign t[9] = t[13] ^ x[2];
  assign y = (t[0]);
endmodule

module R2ind362(x, y);
 input [8:0] x;
 output y;

 wire [18:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = (t[13] & ~t[14]);
  assign t[11] = t[15] ^ x[2];
  assign t[12] = t[16] ^ x[1];
  assign t[13] = t[17] ^ x[8];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = (x[0]);
  assign t[16] = (x[0]);
  assign t[17] = (x[6]);
  assign t[18] = (x[6]);
  assign t[1] = t[5] ? x[4] : x[3];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[4]);
  assign t[4] = ~x[5] & t[6];
  assign t[5] = (t[7]);
  assign t[6] = (t[8]);
  assign t[7] = t[9] ^ x[2];
  assign t[8] = t[10] ^ x[8];
  assign t[9] = (t[11] & ~t[12]);
  assign y = (t[0]);
endmodule

module R2ind363(x, y);
 input [8:0] x;
 output y;

 wire [18:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = (t[13] & ~t[14]);
  assign t[11] = t[15] ^ x[2];
  assign t[12] = t[16] ^ x[1];
  assign t[13] = t[17] ^ x[8];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = (x[0]);
  assign t[16] = (x[0]);
  assign t[17] = (x[6]);
  assign t[18] = (x[6]);
  assign t[1] = t[5] ? x[4] : x[3];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[4]);
  assign t[4] = ~x[5] & t[6];
  assign t[5] = (t[7]);
  assign t[6] = (t[8]);
  assign t[7] = t[9] ^ x[2];
  assign t[8] = t[10] ^ x[8];
  assign t[9] = (t[11] & ~t[12]);
  assign y = (t[0]);
endmodule

module R2ind364(x, y);
 input [8:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[14] ^ x[1];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[7];
  assign t[13] = (x[0]);
  assign t[14] = (x[0]);
  assign t[15] = (x[6]);
  assign t[16] = (x[6]);
  assign t[1] = t[3] ? x[4] : x[3];
  assign t[2] = ~x[5] & t[4];
  assign t[3] = (t[5]);
  assign t[4] = (t[6]);
  assign t[5] = t[7] ^ x[2];
  assign t[6] = t[8] ^ x[8];
  assign t[7] = (t[9] & ~t[10]);
  assign t[8] = (t[11] & ~t[12]);
  assign t[9] = t[13] ^ x[2];
  assign y = (t[0]);
endmodule

module R2ind365(x, y);
 input [8:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[14] ^ x[1];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[7];
  assign t[13] = (x[0]);
  assign t[14] = (x[0]);
  assign t[15] = (x[6]);
  assign t[16] = (x[6]);
  assign t[1] = t[3] ? x[4] : x[3];
  assign t[2] = ~x[5] & t[4];
  assign t[3] = (t[5]);
  assign t[4] = (t[6]);
  assign t[5] = t[7] ^ x[2];
  assign t[6] = t[8] ^ x[8];
  assign t[7] = (t[9] & ~t[10]);
  assign t[8] = (t[11] & ~t[12]);
  assign t[9] = t[13] ^ x[2];
  assign y = (t[0]);
endmodule

module R2ind366(x, y);
 input [4:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = ~t[1];
  assign t[1] = t[2] ? x[4] : x[3];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[2];
  assign t[4] = (t[5] & ~t[6]);
  assign t[5] = t[7] ^ x[2];
  assign t[6] = t[8] ^ x[1];
  assign t[7] = (x[0]);
  assign t[8] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind367(x, y);
 input [4:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = ~t[1];
  assign t[1] = t[2] ? x[4] : x[3];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[2];
  assign t[4] = (t[5] & ~t[6]);
  assign t[5] = t[7] ^ x[2];
  assign t[6] = t[8] ^ x[1];
  assign t[7] = (x[0]);
  assign t[8] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind368(x, y);
 input [8:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[14] ^ x[1];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[7];
  assign t[13] = (x[0]);
  assign t[14] = (x[0]);
  assign t[15] = (x[6]);
  assign t[16] = (x[6]);
  assign t[1] = t[3] ? x[4] : x[3];
  assign t[2] = ~(~x[5] & ~t[4]);
  assign t[3] = (t[5]);
  assign t[4] = (t[6]);
  assign t[5] = t[7] ^ x[2];
  assign t[6] = t[8] ^ x[8];
  assign t[7] = (t[9] & ~t[10]);
  assign t[8] = (t[11] & ~t[12]);
  assign t[9] = t[13] ^ x[2];
  assign y = (t[0]);
endmodule

module R2ind369(x, y);
 input [8:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[14] ^ x[1];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[7];
  assign t[13] = (x[0]);
  assign t[14] = (x[0]);
  assign t[15] = (x[6]);
  assign t[16] = (x[6]);
  assign t[1] = t[3] ? x[4] : x[3];
  assign t[2] = ~(~x[5] & ~t[4]);
  assign t[3] = (t[5]);
  assign t[4] = (t[6]);
  assign t[5] = t[7] ^ x[2];
  assign t[6] = t[8] ^ x[8];
  assign t[7] = (t[9] & ~t[10]);
  assign t[8] = (t[11] & ~t[12]);
  assign t[9] = t[13] ^ x[2];
  assign y = (t[0]);
endmodule

module R2ind370(x, y);
 input [8:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[14] ^ x[1];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[7];
  assign t[13] = (x[0]);
  assign t[14] = (x[0]);
  assign t[15] = (x[6]);
  assign t[16] = (x[6]);
  assign t[1] = t[3] ? x[4] : x[3];
  assign t[2] = ~x[5] & t[4];
  assign t[3] = (t[5]);
  assign t[4] = (t[6]);
  assign t[5] = t[7] ^ x[2];
  assign t[6] = t[8] ^ x[8];
  assign t[7] = (t[9] & ~t[10]);
  assign t[8] = (t[11] & ~t[12]);
  assign t[9] = t[13] ^ x[2];
  assign y = (t[0]);
endmodule

module R2ind371(x, y);
 input [8:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[14] ^ x[1];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[7];
  assign t[13] = (x[0]);
  assign t[14] = (x[0]);
  assign t[15] = (x[6]);
  assign t[16] = (x[6]);
  assign t[1] = t[3] ? x[4] : x[3];
  assign t[2] = ~x[5] & t[4];
  assign t[3] = (t[5]);
  assign t[4] = (t[6]);
  assign t[5] = t[7] ^ x[2];
  assign t[6] = t[8] ^ x[8];
  assign t[7] = (t[9] & ~t[10]);
  assign t[8] = (t[11] & ~t[12]);
  assign t[9] = t[13] ^ x[2];
  assign y = (t[0]);
endmodule

module R2ind372(x, y);
 input [8:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[14] ^ x[1];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[7];
  assign t[13] = (x[0]);
  assign t[14] = (x[0]);
  assign t[15] = (x[6]);
  assign t[16] = (x[6]);
  assign t[1] = t[3] ? x[4] : x[3];
  assign t[2] = ~x[5] & t[4];
  assign t[3] = (t[5]);
  assign t[4] = (t[6]);
  assign t[5] = t[7] ^ x[2];
  assign t[6] = t[8] ^ x[8];
  assign t[7] = (t[9] & ~t[10]);
  assign t[8] = (t[11] & ~t[12]);
  assign t[9] = t[13] ^ x[2];
  assign y = (t[0]);
endmodule

module R2ind373(x, y);
 input [8:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[14] ^ x[1];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[7];
  assign t[13] = (x[0]);
  assign t[14] = (x[0]);
  assign t[15] = (x[6]);
  assign t[16] = (x[6]);
  assign t[1] = t[3] ? x[4] : x[3];
  assign t[2] = ~x[5] & t[4];
  assign t[3] = (t[5]);
  assign t[4] = (t[6]);
  assign t[5] = t[7] ^ x[2];
  assign t[6] = t[8] ^ x[8];
  assign t[7] = (t[9] & ~t[10]);
  assign t[8] = (t[11] & ~t[12]);
  assign t[9] = t[13] ^ x[2];
  assign y = (t[0]);
endmodule

module R2ind374(x, y);
 input [8:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[14] ^ x[1];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[7];
  assign t[13] = (x[0]);
  assign t[14] = (x[0]);
  assign t[15] = (x[6]);
  assign t[16] = (x[6]);
  assign t[1] = t[3] ? x[4] : x[3];
  assign t[2] = ~x[5] & t[4];
  assign t[3] = (t[5]);
  assign t[4] = (t[6]);
  assign t[5] = t[7] ^ x[2];
  assign t[6] = t[8] ^ x[8];
  assign t[7] = (t[9] & ~t[10]);
  assign t[8] = (t[11] & ~t[12]);
  assign t[9] = t[13] ^ x[2];
  assign y = (t[0]);
endmodule

module R2ind375(x, y);
 input [8:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[14] ^ x[1];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[7];
  assign t[13] = (x[0]);
  assign t[14] = (x[0]);
  assign t[15] = (x[6]);
  assign t[16] = (x[6]);
  assign t[1] = t[3] ? x[4] : x[3];
  assign t[2] = ~x[5] & t[4];
  assign t[3] = (t[5]);
  assign t[4] = (t[6]);
  assign t[5] = t[7] ^ x[2];
  assign t[6] = t[8] ^ x[8];
  assign t[7] = (t[9] & ~t[10]);
  assign t[8] = (t[11] & ~t[12]);
  assign t[9] = t[13] ^ x[2];
  assign y = (t[0]);
endmodule

module R2ind376(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind377(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind378(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind379(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind380(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind381(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind382(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind383(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind384(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind385(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind386(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind387(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind388(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind389(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind390(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind391(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind392(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind393(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind394(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind395(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind396(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind397(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind398(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind399(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind400(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind401(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind402(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind403(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind404(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind405(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind406(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind407(x, y);
 input [4:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2_ind(x, y);
 input [737:0] x;
 output [407:0] y;

  R2ind0 R2ind0_inst(.x({x[2], x[1], x[0]}), .y(y[0]));
  R2ind1 R2ind1_inst(.x({x[1], x[2], x[0]}), .y(y[1]));
  R2ind2 R2ind2_inst(.x({x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3]}), .y(y[2]));
  R2ind3 R2ind3_inst(.x({x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3]}), .y(y[3]));
  R2ind4 R2ind4_inst(.x({x[15], x[14], x[13], x[3]}), .y(y[4]));
  R2ind5 R2ind5_inst(.x({x[15], x[14], x[13], x[3]}), .y(y[5]));
  R2ind6 R2ind6_inst(.x({x[12], x[11], x[10], x[3]}), .y(y[6]));
  R2ind7 R2ind7_inst(.x({x[12], x[11], x[10], x[3]}), .y(y[7]));
  R2ind8 R2ind8_inst(.x({x[9], x[8], x[7], x[15], x[14], x[13], x[3]}), .y(y[8]));
  R2ind9 R2ind9_inst(.x({x[9], x[8], x[7], x[15], x[14], x[13], x[3]}), .y(y[9]));
  R2ind10 R2ind10_inst(.x({x[21], x[20], x[19], x[3]}), .y(y[10]));
  R2ind11 R2ind11_inst(.x({x[21], x[20], x[19], x[3]}), .y(y[11]));
  R2ind12 R2ind12_inst(.x({x[24], x[23], x[22], x[3]}), .y(y[12]));
  R2ind13 R2ind13_inst(.x({x[24], x[23], x[22], x[3]}), .y(y[13]));
  R2ind14 R2ind14_inst(.x({x[6], x[5], x[4], x[3]}), .y(y[14]));
  R2ind15 R2ind15_inst(.x({x[6], x[5], x[4], x[3]}), .y(y[15]));
  R2ind16 R2ind16_inst(.x({x[21], x[20], x[19], x[18], x[17], x[16], x[3]}), .y(y[16]));
  R2ind17 R2ind17_inst(.x({x[21], x[20], x[19], x[18], x[17], x[16], x[3]}), .y(y[17]));
  R2ind18 R2ind18_inst(.x({x[27], x[26], x[25]}), .y(y[18]));
  R2ind19 R2ind19_inst(.x({x[27], x[26], x[25]}), .y(y[19]));
  R2ind20 R2ind20_inst(.x({x[30], x[29], x[28], x[3], x[27], x[26], x[25]}), .y(y[20]));
  R2ind21 R2ind21_inst(.x({x[30], x[29], x[28], x[3], x[27], x[26], x[25]}), .y(y[21]));
  R2ind22 R2ind22_inst(.x({x[33], x[32], x[31], x[3]}), .y(y[22]));
  R2ind23 R2ind23_inst(.x({x[33], x[32], x[31], x[3]}), .y(y[23]));
  R2ind24 R2ind24_inst(.x({x[3], x[36], x[35], x[34]}), .y(y[24]));
  R2ind25 R2ind25_inst(.x({x[3], x[39], x[38], x[37]}), .y(y[25]));
  R2ind26 R2ind26_inst(.x({x[3], x[42], x[41], x[40]}), .y(y[26]));
  R2ind27 R2ind27_inst(.x({x[3], x[45], x[44], x[43]}), .y(y[27]));
  R2ind28 R2ind28_inst(.x({x[3], x[48], x[47], x[46]}), .y(y[28]));
  R2ind29 R2ind29_inst(.x({x[3], x[51], x[50], x[49]}), .y(y[29]));
  R2ind30 R2ind30_inst(.x({x[3], x[54], x[53], x[52]}), .y(y[30]));
  R2ind31 R2ind31_inst(.x({x[3], x[57], x[56], x[55]}), .y(y[31]));
  R2ind32 R2ind32_inst(.x({x[3], x[60], x[59], x[58]}), .y(y[32]));
  R2ind33 R2ind33_inst(.x({x[3], x[63], x[62], x[61]}), .y(y[33]));
  R2ind34 R2ind34_inst(.x({x[3], x[66], x[65], x[64]}), .y(y[34]));
  R2ind35 R2ind35_inst(.x({x[3], x[69], x[68], x[67]}), .y(y[35]));
  R2ind36 R2ind36_inst(.x({x[3], x[72], x[71], x[70]}), .y(y[36]));
  R2ind37 R2ind37_inst(.x({x[3], x[75], x[74], x[73]}), .y(y[37]));
  R2ind38 R2ind38_inst(.x({x[3], x[78], x[77], x[76]}), .y(y[38]));
  R2ind39 R2ind39_inst(.x({x[3], x[81], x[80], x[79]}), .y(y[39]));
  R2ind40 R2ind40_inst(.x({x[3], x[84], x[83], x[82]}), .y(y[40]));
  R2ind41 R2ind41_inst(.x({x[3], x[87], x[86], x[85]}), .y(y[41]));
  R2ind42 R2ind42_inst(.x({x[3], x[90], x[89], x[88]}), .y(y[42]));
  R2ind43 R2ind43_inst(.x({x[3], x[93], x[92], x[91]}), .y(y[43]));
  R2ind44 R2ind44_inst(.x({x[3], x[96], x[95], x[94]}), .y(y[44]));
  R2ind45 R2ind45_inst(.x({x[3], x[99], x[98], x[97]}), .y(y[45]));
  R2ind46 R2ind46_inst(.x({x[3], x[102], x[101], x[100]}), .y(y[46]));
  R2ind47 R2ind47_inst(.x({x[3], x[105], x[104], x[103]}), .y(y[47]));
  R2ind48 R2ind48_inst(.x({x[3], x[108], x[107], x[106]}), .y(y[48]));
  R2ind49 R2ind49_inst(.x({x[3], x[111], x[110], x[109]}), .y(y[49]));
  R2ind50 R2ind50_inst(.x({x[3], x[114], x[113], x[112]}), .y(y[50]));
  R2ind51 R2ind51_inst(.x({x[3], x[117], x[116], x[115]}), .y(y[51]));
  R2ind52 R2ind52_inst(.x({x[3], x[120], x[119], x[118]}), .y(y[52]));
  R2ind53 R2ind53_inst(.x({x[3], x[123], x[122], x[121]}), .y(y[53]));
  R2ind54 R2ind54_inst(.x({x[3], x[126], x[125], x[124]}), .y(y[54]));
  R2ind55 R2ind55_inst(.x({x[3], x[129], x[128], x[127]}), .y(y[55]));
  R2ind56 R2ind56_inst(.x({x[3], x[132], x[131], x[130]}), .y(y[56]));
  R2ind57 R2ind57_inst(.x({x[3], x[135], x[134], x[133]}), .y(y[57]));
  R2ind58 R2ind58_inst(.x({x[3], x[138], x[137], x[136]}), .y(y[58]));
  R2ind59 R2ind59_inst(.x({x[3], x[141], x[140], x[139]}), .y(y[59]));
  R2ind60 R2ind60_inst(.x({x[3], x[144], x[143], x[142]}), .y(y[60]));
  R2ind61 R2ind61_inst(.x({x[3], x[147], x[146], x[145]}), .y(y[61]));
  R2ind62 R2ind62_inst(.x({x[3], x[150], x[149], x[148]}), .y(y[62]));
  R2ind63 R2ind63_inst(.x({x[3], x[153], x[152], x[151]}), .y(y[63]));
  R2ind64 R2ind64_inst(.x({x[3], x[156], x[155], x[154]}), .y(y[64]));
  R2ind65 R2ind65_inst(.x({x[3], x[159], x[158], x[157]}), .y(y[65]));
  R2ind66 R2ind66_inst(.x({x[3], x[162], x[161], x[160]}), .y(y[66]));
  R2ind67 R2ind67_inst(.x({x[3], x[165], x[164], x[163]}), .y(y[67]));
  R2ind68 R2ind68_inst(.x({x[3], x[168], x[167], x[166]}), .y(y[68]));
  R2ind69 R2ind69_inst(.x({x[3], x[171], x[170], x[169]}), .y(y[69]));
  R2ind70 R2ind70_inst(.x({x[3], x[174], x[173], x[172]}), .y(y[70]));
  R2ind71 R2ind71_inst(.x({x[3], x[177], x[176], x[175]}), .y(y[71]));
  R2ind72 R2ind72_inst(.x({x[3], x[180], x[179], x[178]}), .y(y[72]));
  R2ind73 R2ind73_inst(.x({x[3], x[183], x[182], x[181]}), .y(y[73]));
  R2ind74 R2ind74_inst(.x({x[3], x[186], x[185], x[184]}), .y(y[74]));
  R2ind75 R2ind75_inst(.x({x[3], x[189], x[188], x[187]}), .y(y[75]));
  R2ind76 R2ind76_inst(.x({x[3], x[192], x[191], x[190]}), .y(y[76]));
  R2ind77 R2ind77_inst(.x({x[3], x[195], x[194], x[193]}), .y(y[77]));
  R2ind78 R2ind78_inst(.x({x[3], x[198], x[197], x[196]}), .y(y[78]));
  R2ind79 R2ind79_inst(.x({x[3], x[201], x[200], x[199]}), .y(y[79]));
  R2ind80 R2ind80_inst(.x({x[3], x[204], x[203], x[202]}), .y(y[80]));
  R2ind81 R2ind81_inst(.x({x[3], x[207], x[206], x[205]}), .y(y[81]));
  R2ind82 R2ind82_inst(.x({x[3], x[210], x[209], x[208]}), .y(y[82]));
  R2ind83 R2ind83_inst(.x({x[3], x[213], x[212], x[211]}), .y(y[83]));
  R2ind84 R2ind84_inst(.x({x[3], x[216], x[215], x[214]}), .y(y[84]));
  R2ind85 R2ind85_inst(.x({x[3], x[219], x[218], x[217]}), .y(y[85]));
  R2ind86 R2ind86_inst(.x({x[3], x[222], x[221], x[220]}), .y(y[86]));
  R2ind87 R2ind87_inst(.x({x[3], x[225], x[224], x[223]}), .y(y[87]));
  R2ind88 R2ind88_inst(.x({x[3], x[228], x[36], x[227], x[226], x[34]}), .y(y[88]));
  R2ind89 R2ind89_inst(.x({x[3], x[231], x[39], x[230], x[229], x[37]}), .y(y[89]));
  R2ind90 R2ind90_inst(.x({x[3], x[234], x[42], x[233], x[232], x[40]}), .y(y[90]));
  R2ind91 R2ind91_inst(.x({x[3], x[237], x[45], x[236], x[235], x[43]}), .y(y[91]));
  R2ind92 R2ind92_inst(.x({x[3], x[240], x[48], x[239], x[238], x[46]}), .y(y[92]));
  R2ind93 R2ind93_inst(.x({x[3], x[243], x[51], x[242], x[241], x[49]}), .y(y[93]));
  R2ind94 R2ind94_inst(.x({x[3], x[54], x[246], x[245], x[52], x[244]}), .y(y[94]));
  R2ind95 R2ind95_inst(.x({x[3], x[57], x[249], x[248], x[55], x[247]}), .y(y[95]));
  R2ind96 R2ind96_inst(.x({x[3], x[60], x[252], x[251], x[58], x[250]}), .y(y[96]));
  R2ind97 R2ind97_inst(.x({x[3], x[63], x[255], x[254], x[61], x[253]}), .y(y[97]));
  R2ind98 R2ind98_inst(.x({x[3], x[66], x[258], x[257], x[64], x[256]}), .y(y[98]));
  R2ind99 R2ind99_inst(.x({x[3], x[69], x[261], x[260], x[67], x[259]}), .y(y[99]));
  R2ind100 R2ind100_inst(.x({x[3], x[72], x[264], x[263], x[70], x[262]}), .y(y[100]));
  R2ind101 R2ind101_inst(.x({x[3], x[75], x[267], x[266], x[73], x[265]}), .y(y[101]));
  R2ind102 R2ind102_inst(.x({x[3], x[78], x[270], x[269], x[76], x[268]}), .y(y[102]));
  R2ind103 R2ind103_inst(.x({x[3], x[81], x[273], x[272], x[79], x[271]}), .y(y[103]));
  R2ind104 R2ind104_inst(.x({x[3], x[84], x[276], x[275], x[82], x[274]}), .y(y[104]));
  R2ind105 R2ind105_inst(.x({x[3], x[87], x[279], x[278], x[85], x[277]}), .y(y[105]));
  R2ind106 R2ind106_inst(.x({x[3], x[90], x[282], x[281], x[88], x[280]}), .y(y[106]));
  R2ind107 R2ind107_inst(.x({x[3], x[93], x[285], x[284], x[91], x[283]}), .y(y[107]));
  R2ind108 R2ind108_inst(.x({x[3], x[288], x[96], x[287], x[286], x[94]}), .y(y[108]));
  R2ind109 R2ind109_inst(.x({x[3], x[291], x[99], x[290], x[289], x[97]}), .y(y[109]));
  R2ind110 R2ind110_inst(.x({x[3], x[294], x[102], x[293], x[292], x[100]}), .y(y[110]));
  R2ind111 R2ind111_inst(.x({x[3], x[297], x[105], x[296], x[295], x[103]}), .y(y[111]));
  R2ind112 R2ind112_inst(.x({x[3], x[300], x[108], x[299], x[298], x[106]}), .y(y[112]));
  R2ind113 R2ind113_inst(.x({x[3], x[303], x[111], x[302], x[301], x[109]}), .y(y[113]));
  R2ind114 R2ind114_inst(.x({x[3], x[306], x[114], x[305], x[304], x[112]}), .y(y[114]));
  R2ind115 R2ind115_inst(.x({x[3], x[309], x[117], x[308], x[307], x[115]}), .y(y[115]));
  R2ind116 R2ind116_inst(.x({x[3], x[312], x[120], x[311], x[310], x[118]}), .y(y[116]));
  R2ind117 R2ind117_inst(.x({x[3], x[315], x[123], x[314], x[313], x[121]}), .y(y[117]));
  R2ind118 R2ind118_inst(.x({x[3], x[318], x[126], x[317], x[316], x[124]}), .y(y[118]));
  R2ind119 R2ind119_inst(.x({x[3], x[321], x[129], x[320], x[319], x[127]}), .y(y[119]));
  R2ind120 R2ind120_inst(.x({x[3], x[324], x[132], x[36], x[323], x[322], x[130], x[34]}), .y(y[120]));
  R2ind121 R2ind121_inst(.x({x[3], x[327], x[135], x[39], x[326], x[325], x[133], x[37]}), .y(y[121]));
  R2ind122 R2ind122_inst(.x({x[3], x[330], x[42], x[138], x[329], x[328], x[40], x[136]}), .y(y[122]));
  R2ind123 R2ind123_inst(.x({x[3], x[333], x[45], x[141], x[332], x[331], x[43], x[139]}), .y(y[123]));
  R2ind124 R2ind124_inst(.x({x[3], x[336], x[48], x[144], x[335], x[334], x[46], x[142]}), .y(y[124]));
  R2ind125 R2ind125_inst(.x({x[3], x[339], x[51], x[147], x[338], x[337], x[49], x[145]}), .y(y[125]));
  R2ind126 R2ind126_inst(.x({x[3], x[342], x[54], x[150], x[341], x[340], x[52], x[148]}), .y(y[126]));
  R2ind127 R2ind127_inst(.x({x[3], x[345], x[57], x[153], x[344], x[343], x[55], x[151]}), .y(y[127]));
  R2ind128 R2ind128_inst(.x({x[3], x[348], x[60], x[156], x[347], x[346], x[58], x[154]}), .y(y[128]));
  R2ind129 R2ind129_inst(.x({x[3], x[351], x[63], x[159], x[350], x[349], x[61], x[157]}), .y(y[129]));
  R2ind130 R2ind130_inst(.x({x[3], x[66], x[354], x[162], x[353], x[64], x[352], x[160]}), .y(y[130]));
  R2ind131 R2ind131_inst(.x({x[3], x[69], x[357], x[165], x[356], x[67], x[355], x[163]}), .y(y[131]));
  R2ind132 R2ind132_inst(.x({x[3], x[72], x[360], x[168], x[359], x[70], x[358], x[166]}), .y(y[132]));
  R2ind133 R2ind133_inst(.x({x[3], x[75], x[363], x[171], x[362], x[73], x[361], x[169]}), .y(y[133]));
  R2ind134 R2ind134_inst(.x({x[3], x[78], x[366], x[174], x[365], x[76], x[364], x[172]}), .y(y[134]));
  R2ind135 R2ind135_inst(.x({x[3], x[81], x[369], x[177], x[368], x[79], x[367], x[175]}), .y(y[135]));
  R2ind136 R2ind136_inst(.x({x[3], x[84], x[372], x[180], x[371], x[82], x[370], x[178]}), .y(y[136]));
  R2ind137 R2ind137_inst(.x({x[3], x[87], x[375], x[183], x[374], x[85], x[373], x[181]}), .y(y[137]));
  R2ind138 R2ind138_inst(.x({x[3], x[90], x[378], x[186], x[377], x[88], x[376], x[184]}), .y(y[138]));
  R2ind139 R2ind139_inst(.x({x[3], x[93], x[381], x[189], x[380], x[91], x[379], x[187]}), .y(y[139]));
  R2ind140 R2ind140_inst(.x({x[3], x[384], x[192], x[96], x[383], x[382], x[190], x[94]}), .y(y[140]));
  R2ind141 R2ind141_inst(.x({x[3], x[387], x[195], x[99], x[386], x[385], x[193], x[97]}), .y(y[141]));
  R2ind142 R2ind142_inst(.x({x[3], x[390], x[198], x[102], x[389], x[388], x[196], x[100]}), .y(y[142]));
  R2ind143 R2ind143_inst(.x({x[3], x[393], x[201], x[105], x[392], x[391], x[199], x[103]}), .y(y[143]));
  R2ind144 R2ind144_inst(.x({x[3], x[396], x[204], x[108], x[395], x[394], x[202], x[106]}), .y(y[144]));
  R2ind145 R2ind145_inst(.x({x[3], x[399], x[207], x[111], x[398], x[397], x[205], x[109]}), .y(y[145]));
  R2ind146 R2ind146_inst(.x({x[3], x[402], x[210], x[114], x[401], x[400], x[208], x[112]}), .y(y[146]));
  R2ind147 R2ind147_inst(.x({x[3], x[405], x[213], x[117], x[404], x[403], x[211], x[115]}), .y(y[147]));
  R2ind148 R2ind148_inst(.x({x[3], x[408], x[216], x[120], x[407], x[406], x[214], x[118]}), .y(y[148]));
  R2ind149 R2ind149_inst(.x({x[3], x[411], x[219], x[123], x[410], x[409], x[217], x[121]}), .y(y[149]));
  R2ind150 R2ind150_inst(.x({x[3], x[414], x[222], x[126], x[413], x[412], x[220], x[124]}), .y(y[150]));
  R2ind151 R2ind151_inst(.x({x[3], x[417], x[225], x[129], x[416], x[415], x[223], x[127]}), .y(y[151]));
  R2ind152 R2ind152_inst(.x({x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[418]}), .y(y[152]));
  R2ind153 R2ind153_inst(.x({x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[418]}), .y(y[153]));
  R2ind154 R2ind154_inst(.x({x[429], x[428], x[427], x[423], x[422], x[421], x[426], x[425], x[424], x[420], x[419], x[418]}), .y(y[154]));
  R2ind155 R2ind155_inst(.x({x[429], x[428], x[427], x[423], x[422], x[421], x[426], x[425], x[424], x[420], x[419], x[418]}), .y(y[155]));
  R2ind156 R2ind156_inst(.x({x[429], x[428], x[427], x[423], x[422], x[421], x[426], x[425], x[424], x[420], x[419], x[418]}), .y(y[156]));
  R2ind157 R2ind157_inst(.x({x[429], x[428], x[427], x[423], x[422], x[421], x[426], x[425], x[424], x[420], x[419], x[418]}), .y(y[157]));
  R2ind158 R2ind158_inst(.x({x[429], x[428], x[427], x[423], x[422], x[421], x[420], x[419], x[418], x[426], x[425], x[424]}), .y(y[158]));
  R2ind159 R2ind159_inst(.x({x[429], x[428], x[427], x[423], x[422], x[421], x[420], x[419], x[418], x[426], x[425], x[424]}), .y(y[159]));
  R2ind160 R2ind160_inst(.x({x[441], x[440], x[439], x[438], x[437], x[436], x[435], x[434], x[433], x[432], x[431], x[430]}), .y(y[160]));
  R2ind161 R2ind161_inst(.x({x[441], x[440], x[439], x[438], x[437], x[436], x[435], x[434], x[433], x[432], x[431], x[430]}), .y(y[161]));
  R2ind162 R2ind162_inst(.x({x[441], x[440], x[439], x[435], x[434], x[433], x[438], x[437], x[436], x[432], x[431], x[430]}), .y(y[162]));
  R2ind163 R2ind163_inst(.x({x[441], x[440], x[439], x[435], x[434], x[433], x[438], x[437], x[436], x[432], x[431], x[430]}), .y(y[163]));
  R2ind164 R2ind164_inst(.x({x[441], x[440], x[439], x[435], x[434], x[433], x[438], x[437], x[436], x[432], x[431], x[430]}), .y(y[164]));
  R2ind165 R2ind165_inst(.x({x[441], x[440], x[439], x[435], x[434], x[433], x[438], x[437], x[436], x[432], x[431], x[430]}), .y(y[165]));
  R2ind166 R2ind166_inst(.x({x[441], x[440], x[439], x[435], x[434], x[433], x[432], x[431], x[430], x[438], x[437], x[436]}), .y(y[166]));
  R2ind167 R2ind167_inst(.x({x[441], x[440], x[439], x[435], x[434], x[433], x[432], x[431], x[430], x[438], x[437], x[436]}), .y(y[167]));
  R2ind168 R2ind168_inst(.x({x[453], x[452], x[451], x[450], x[449], x[448], x[447], x[446], x[445], x[444], x[443], x[442]}), .y(y[168]));
  R2ind169 R2ind169_inst(.x({x[453], x[452], x[451], x[450], x[449], x[448], x[447], x[446], x[445], x[444], x[443], x[442]}), .y(y[169]));
  R2ind170 R2ind170_inst(.x({x[453], x[452], x[451], x[447], x[446], x[445], x[450], x[449], x[448], x[444], x[443], x[442]}), .y(y[170]));
  R2ind171 R2ind171_inst(.x({x[453], x[452], x[451], x[447], x[446], x[445], x[450], x[449], x[448], x[444], x[443], x[442]}), .y(y[171]));
  R2ind172 R2ind172_inst(.x({x[453], x[452], x[451], x[447], x[446], x[445], x[450], x[449], x[448], x[444], x[443], x[442]}), .y(y[172]));
  R2ind173 R2ind173_inst(.x({x[453], x[452], x[451], x[447], x[446], x[445], x[450], x[449], x[448], x[444], x[443], x[442]}), .y(y[173]));
  R2ind174 R2ind174_inst(.x({x[453], x[452], x[451], x[447], x[446], x[445], x[444], x[443], x[442], x[450], x[449], x[448]}), .y(y[174]));
  R2ind175 R2ind175_inst(.x({x[453], x[452], x[451], x[447], x[446], x[445], x[444], x[443], x[442], x[450], x[449], x[448]}), .y(y[175]));
  R2ind176 R2ind176_inst(.x({x[465], x[464], x[463], x[462], x[461], x[460], x[459], x[458], x[457], x[456], x[455], x[454]}), .y(y[176]));
  R2ind177 R2ind177_inst(.x({x[465], x[464], x[463], x[462], x[461], x[460], x[459], x[458], x[457], x[456], x[455], x[454]}), .y(y[177]));
  R2ind178 R2ind178_inst(.x({x[465], x[464], x[463], x[459], x[458], x[457], x[462], x[461], x[460], x[456], x[455], x[454]}), .y(y[178]));
  R2ind179 R2ind179_inst(.x({x[465], x[464], x[463], x[459], x[458], x[457], x[462], x[461], x[460], x[456], x[455], x[454]}), .y(y[179]));
  R2ind180 R2ind180_inst(.x({x[465], x[464], x[463], x[459], x[458], x[457], x[462], x[461], x[460], x[456], x[455], x[454]}), .y(y[180]));
  R2ind181 R2ind181_inst(.x({x[465], x[464], x[463], x[459], x[458], x[457], x[462], x[461], x[460], x[456], x[455], x[454]}), .y(y[181]));
  R2ind182 R2ind182_inst(.x({x[465], x[464], x[463], x[459], x[458], x[457], x[456], x[455], x[454], x[462], x[461], x[460]}), .y(y[182]));
  R2ind183 R2ind183_inst(.x({x[465], x[464], x[463], x[459], x[458], x[457], x[456], x[455], x[454], x[462], x[461], x[460]}), .y(y[183]));
  R2ind184 R2ind184_inst(.x({x[477], x[476], x[475], x[474], x[473], x[472], x[471], x[470], x[469], x[468], x[467], x[466]}), .y(y[184]));
  R2ind185 R2ind185_inst(.x({x[477], x[476], x[475], x[474], x[473], x[472], x[471], x[470], x[469], x[468], x[467], x[466]}), .y(y[185]));
  R2ind186 R2ind186_inst(.x({x[477], x[476], x[475], x[471], x[470], x[469], x[474], x[473], x[472], x[468], x[467], x[466]}), .y(y[186]));
  R2ind187 R2ind187_inst(.x({x[477], x[476], x[475], x[471], x[470], x[469], x[474], x[473], x[472], x[468], x[467], x[466]}), .y(y[187]));
  R2ind188 R2ind188_inst(.x({x[477], x[476], x[475], x[471], x[470], x[469], x[474], x[473], x[472], x[468], x[467], x[466]}), .y(y[188]));
  R2ind189 R2ind189_inst(.x({x[477], x[476], x[475], x[471], x[470], x[469], x[474], x[473], x[472], x[468], x[467], x[466]}), .y(y[189]));
  R2ind190 R2ind190_inst(.x({x[477], x[476], x[475], x[471], x[470], x[469], x[468], x[467], x[466], x[474], x[473], x[472]}), .y(y[190]));
  R2ind191 R2ind191_inst(.x({x[477], x[476], x[475], x[471], x[470], x[469], x[468], x[467], x[466], x[474], x[473], x[472]}), .y(y[191]));
  R2ind192 R2ind192_inst(.x({x[489], x[488], x[487], x[486], x[485], x[484], x[483], x[482], x[481], x[480], x[479], x[478]}), .y(y[192]));
  R2ind193 R2ind193_inst(.x({x[489], x[488], x[487], x[486], x[485], x[484], x[483], x[482], x[481], x[480], x[479], x[478]}), .y(y[193]));
  R2ind194 R2ind194_inst(.x({x[489], x[488], x[487], x[483], x[482], x[481], x[486], x[485], x[484], x[480], x[479], x[478]}), .y(y[194]));
  R2ind195 R2ind195_inst(.x({x[489], x[488], x[487], x[483], x[482], x[481], x[486], x[485], x[484], x[480], x[479], x[478]}), .y(y[195]));
  R2ind196 R2ind196_inst(.x({x[489], x[488], x[487], x[483], x[482], x[481], x[486], x[485], x[484], x[480], x[479], x[478]}), .y(y[196]));
  R2ind197 R2ind197_inst(.x({x[489], x[488], x[487], x[483], x[482], x[481], x[486], x[485], x[484], x[480], x[479], x[478]}), .y(y[197]));
  R2ind198 R2ind198_inst(.x({x[489], x[488], x[487], x[483], x[482], x[481], x[480], x[479], x[478], x[486], x[485], x[484]}), .y(y[198]));
  R2ind199 R2ind199_inst(.x({x[489], x[488], x[487], x[483], x[482], x[481], x[480], x[479], x[478], x[486], x[485], x[484]}), .y(y[199]));
  R2ind200 R2ind200_inst(.x({x[501], x[500], x[499], x[498], x[497], x[496], x[495], x[494], x[493], x[492], x[491], x[490]}), .y(y[200]));
  R2ind201 R2ind201_inst(.x({x[501], x[500], x[499], x[498], x[497], x[496], x[495], x[494], x[493], x[492], x[491], x[490]}), .y(y[201]));
  R2ind202 R2ind202_inst(.x({x[501], x[500], x[499], x[495], x[494], x[493], x[498], x[497], x[496], x[492], x[491], x[490]}), .y(y[202]));
  R2ind203 R2ind203_inst(.x({x[501], x[500], x[499], x[495], x[494], x[493], x[498], x[497], x[496], x[492], x[491], x[490]}), .y(y[203]));
  R2ind204 R2ind204_inst(.x({x[501], x[500], x[499], x[495], x[494], x[493], x[498], x[497], x[496], x[492], x[491], x[490]}), .y(y[204]));
  R2ind205 R2ind205_inst(.x({x[501], x[500], x[499], x[495], x[494], x[493], x[498], x[497], x[496], x[492], x[491], x[490]}), .y(y[205]));
  R2ind206 R2ind206_inst(.x({x[501], x[500], x[499], x[495], x[494], x[493], x[492], x[491], x[490], x[498], x[497], x[496]}), .y(y[206]));
  R2ind207 R2ind207_inst(.x({x[501], x[500], x[499], x[495], x[494], x[493], x[492], x[491], x[490], x[498], x[497], x[496]}), .y(y[207]));
  R2ind208 R2ind208_inst(.x({x[513], x[512], x[511], x[510], x[509], x[508], x[507], x[506], x[505], x[504], x[503], x[502]}), .y(y[208]));
  R2ind209 R2ind209_inst(.x({x[513], x[512], x[511], x[510], x[509], x[508], x[507], x[506], x[505], x[504], x[503], x[502]}), .y(y[209]));
  R2ind210 R2ind210_inst(.x({x[513], x[512], x[511], x[507], x[506], x[505], x[510], x[509], x[508], x[504], x[503], x[502]}), .y(y[210]));
  R2ind211 R2ind211_inst(.x({x[513], x[512], x[511], x[507], x[506], x[505], x[510], x[509], x[508], x[504], x[503], x[502]}), .y(y[211]));
  R2ind212 R2ind212_inst(.x({x[513], x[512], x[511], x[507], x[506], x[505], x[510], x[509], x[508], x[504], x[503], x[502]}), .y(y[212]));
  R2ind213 R2ind213_inst(.x({x[513], x[512], x[511], x[507], x[506], x[505], x[510], x[509], x[508], x[504], x[503], x[502]}), .y(y[213]));
  R2ind214 R2ind214_inst(.x({x[513], x[512], x[511], x[507], x[506], x[505], x[504], x[503], x[502], x[510], x[509], x[508]}), .y(y[214]));
  R2ind215 R2ind215_inst(.x({x[513], x[512], x[511], x[507], x[506], x[505], x[504], x[503], x[502], x[510], x[509], x[508]}), .y(y[215]));
  R2ind216 R2ind216_inst(.x({x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[514]}), .y(y[216]));
  R2ind217 R2ind217_inst(.x({x[525], x[524], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[514]}), .y(y[217]));
  R2ind218 R2ind218_inst(.x({x[525], x[524], x[523], x[519], x[518], x[517], x[522], x[521], x[520], x[516], x[515], x[514]}), .y(y[218]));
  R2ind219 R2ind219_inst(.x({x[525], x[524], x[523], x[519], x[518], x[517], x[522], x[521], x[520], x[516], x[515], x[514]}), .y(y[219]));
  R2ind220 R2ind220_inst(.x({x[525], x[524], x[523], x[519], x[518], x[517], x[522], x[521], x[520], x[516], x[515], x[514]}), .y(y[220]));
  R2ind221 R2ind221_inst(.x({x[525], x[524], x[523], x[519], x[518], x[517], x[522], x[521], x[520], x[516], x[515], x[514]}), .y(y[221]));
  R2ind222 R2ind222_inst(.x({x[525], x[524], x[523], x[519], x[518], x[517], x[516], x[515], x[514], x[522], x[521], x[520]}), .y(y[222]));
  R2ind223 R2ind223_inst(.x({x[525], x[524], x[523], x[519], x[518], x[517], x[516], x[515], x[514], x[522], x[521], x[520]}), .y(y[223]));
  R2ind224 R2ind224_inst(.x({x[537], x[536], x[535], x[534], x[533], x[532], x[531], x[530], x[529], x[528], x[527], x[526]}), .y(y[224]));
  R2ind225 R2ind225_inst(.x({x[537], x[536], x[535], x[534], x[533], x[532], x[531], x[530], x[529], x[528], x[527], x[526]}), .y(y[225]));
  R2ind226 R2ind226_inst(.x({x[537], x[536], x[535], x[531], x[530], x[529], x[534], x[533], x[532], x[528], x[527], x[526]}), .y(y[226]));
  R2ind227 R2ind227_inst(.x({x[537], x[536], x[535], x[531], x[530], x[529], x[534], x[533], x[532], x[528], x[527], x[526]}), .y(y[227]));
  R2ind228 R2ind228_inst(.x({x[537], x[536], x[535], x[531], x[530], x[529], x[534], x[533], x[532], x[528], x[527], x[526]}), .y(y[228]));
  R2ind229 R2ind229_inst(.x({x[537], x[536], x[535], x[531], x[530], x[529], x[534], x[533], x[532], x[528], x[527], x[526]}), .y(y[229]));
  R2ind230 R2ind230_inst(.x({x[537], x[536], x[535], x[531], x[530], x[529], x[528], x[527], x[526], x[534], x[533], x[532]}), .y(y[230]));
  R2ind231 R2ind231_inst(.x({x[537], x[536], x[535], x[531], x[530], x[529], x[528], x[527], x[526], x[534], x[533], x[532]}), .y(y[231]));
  R2ind232 R2ind232_inst(.x({x[549], x[548], x[547], x[546], x[545], x[544], x[543], x[542], x[541], x[540], x[539], x[538]}), .y(y[232]));
  R2ind233 R2ind233_inst(.x({x[549], x[548], x[547], x[546], x[545], x[544], x[543], x[542], x[541], x[540], x[539], x[538]}), .y(y[233]));
  R2ind234 R2ind234_inst(.x({x[549], x[548], x[547], x[543], x[542], x[541], x[546], x[545], x[544], x[540], x[539], x[538]}), .y(y[234]));
  R2ind235 R2ind235_inst(.x({x[549], x[548], x[547], x[543], x[542], x[541], x[546], x[545], x[544], x[540], x[539], x[538]}), .y(y[235]));
  R2ind236 R2ind236_inst(.x({x[549], x[548], x[547], x[543], x[542], x[541], x[546], x[545], x[544], x[540], x[539], x[538]}), .y(y[236]));
  R2ind237 R2ind237_inst(.x({x[549], x[548], x[547], x[543], x[542], x[541], x[546], x[545], x[544], x[540], x[539], x[538]}), .y(y[237]));
  R2ind238 R2ind238_inst(.x({x[549], x[548], x[547], x[543], x[542], x[541], x[540], x[539], x[538], x[546], x[545], x[544]}), .y(y[238]));
  R2ind239 R2ind239_inst(.x({x[549], x[548], x[547], x[543], x[542], x[541], x[540], x[539], x[538], x[546], x[545], x[544]}), .y(y[239]));
  R2ind240 R2ind240_inst(.x({x[561], x[560], x[559], x[558], x[557], x[556], x[555], x[554], x[553], x[552], x[551], x[550]}), .y(y[240]));
  R2ind241 R2ind241_inst(.x({x[561], x[560], x[559], x[558], x[557], x[556], x[555], x[554], x[553], x[552], x[551], x[550]}), .y(y[241]));
  R2ind242 R2ind242_inst(.x({x[561], x[560], x[559], x[555], x[554], x[553], x[558], x[557], x[556], x[552], x[551], x[550]}), .y(y[242]));
  R2ind243 R2ind243_inst(.x({x[561], x[560], x[559], x[555], x[554], x[553], x[558], x[557], x[556], x[552], x[551], x[550]}), .y(y[243]));
  R2ind244 R2ind244_inst(.x({x[561], x[560], x[559], x[555], x[554], x[553], x[558], x[557], x[556], x[552], x[551], x[550]}), .y(y[244]));
  R2ind245 R2ind245_inst(.x({x[561], x[560], x[559], x[555], x[554], x[553], x[558], x[557], x[556], x[552], x[551], x[550]}), .y(y[245]));
  R2ind246 R2ind246_inst(.x({x[561], x[560], x[559], x[555], x[554], x[553], x[552], x[551], x[550], x[558], x[557], x[556]}), .y(y[246]));
  R2ind247 R2ind247_inst(.x({x[561], x[560], x[559], x[555], x[554], x[553], x[552], x[551], x[550], x[558], x[557], x[556]}), .y(y[247]));
  R2ind248 R2ind248_inst(.x({x[573], x[572], x[571], x[570], x[569], x[568], x[567], x[566], x[565], x[564], x[563], x[562]}), .y(y[248]));
  R2ind249 R2ind249_inst(.x({x[573], x[572], x[571], x[570], x[569], x[568], x[567], x[566], x[565], x[564], x[563], x[562]}), .y(y[249]));
  R2ind250 R2ind250_inst(.x({x[573], x[572], x[571], x[567], x[566], x[565], x[570], x[569], x[568], x[564], x[563], x[562]}), .y(y[250]));
  R2ind251 R2ind251_inst(.x({x[573], x[572], x[571], x[567], x[566], x[565], x[570], x[569], x[568], x[564], x[563], x[562]}), .y(y[251]));
  R2ind252 R2ind252_inst(.x({x[573], x[572], x[571], x[567], x[566], x[565], x[570], x[569], x[568], x[564], x[563], x[562]}), .y(y[252]));
  R2ind253 R2ind253_inst(.x({x[573], x[572], x[571], x[567], x[566], x[565], x[570], x[569], x[568], x[564], x[563], x[562]}), .y(y[253]));
  R2ind254 R2ind254_inst(.x({x[573], x[572], x[571], x[567], x[566], x[565], x[564], x[563], x[562], x[570], x[569], x[568]}), .y(y[254]));
  R2ind255 R2ind255_inst(.x({x[573], x[572], x[571], x[567], x[566], x[565], x[564], x[563], x[562], x[570], x[569], x[568]}), .y(y[255]));
  R2ind256 R2ind256_inst(.x({x[585], x[584], x[583], x[582], x[581], x[580], x[579], x[578], x[577], x[576], x[575], x[574]}), .y(y[256]));
  R2ind257 R2ind257_inst(.x({x[585], x[584], x[583], x[582], x[581], x[580], x[579], x[578], x[577], x[576], x[575], x[574]}), .y(y[257]));
  R2ind258 R2ind258_inst(.x({x[585], x[584], x[583], x[579], x[578], x[577], x[582], x[581], x[580], x[576], x[575], x[574]}), .y(y[258]));
  R2ind259 R2ind259_inst(.x({x[585], x[584], x[583], x[579], x[578], x[577], x[582], x[581], x[580], x[576], x[575], x[574]}), .y(y[259]));
  R2ind260 R2ind260_inst(.x({x[585], x[584], x[583], x[579], x[578], x[577], x[582], x[581], x[580], x[576], x[575], x[574]}), .y(y[260]));
  R2ind261 R2ind261_inst(.x({x[585], x[584], x[583], x[579], x[578], x[577], x[582], x[581], x[580], x[576], x[575], x[574]}), .y(y[261]));
  R2ind262 R2ind262_inst(.x({x[585], x[584], x[583], x[579], x[578], x[577], x[576], x[575], x[574], x[582], x[581], x[580]}), .y(y[262]));
  R2ind263 R2ind263_inst(.x({x[585], x[584], x[583], x[579], x[578], x[577], x[576], x[575], x[574], x[582], x[581], x[580]}), .y(y[263]));
  R2ind264 R2ind264_inst(.x({x[597], x[596], x[595], x[594], x[593], x[592], x[591], x[590], x[589], x[588], x[587], x[586]}), .y(y[264]));
  R2ind265 R2ind265_inst(.x({x[597], x[596], x[595], x[594], x[593], x[592], x[591], x[590], x[589], x[588], x[587], x[586]}), .y(y[265]));
  R2ind266 R2ind266_inst(.x({x[597], x[596], x[595], x[591], x[590], x[589], x[594], x[593], x[592], x[588], x[587], x[586]}), .y(y[266]));
  R2ind267 R2ind267_inst(.x({x[597], x[596], x[595], x[591], x[590], x[589], x[594], x[593], x[592], x[588], x[587], x[586]}), .y(y[267]));
  R2ind268 R2ind268_inst(.x({x[597], x[596], x[595], x[591], x[590], x[589], x[594], x[593], x[592], x[588], x[587], x[586]}), .y(y[268]));
  R2ind269 R2ind269_inst(.x({x[597], x[596], x[595], x[591], x[590], x[589], x[594], x[593], x[592], x[588], x[587], x[586]}), .y(y[269]));
  R2ind270 R2ind270_inst(.x({x[597], x[596], x[595], x[591], x[590], x[589], x[588], x[587], x[586], x[594], x[593], x[592]}), .y(y[270]));
  R2ind271 R2ind271_inst(.x({x[597], x[596], x[595], x[591], x[590], x[589], x[588], x[587], x[586], x[594], x[593], x[592]}), .y(y[271]));
  R2ind272 R2ind272_inst(.x({x[609], x[608], x[607], x[606], x[605], x[604], x[603], x[602], x[601], x[600], x[599], x[598]}), .y(y[272]));
  R2ind273 R2ind273_inst(.x({x[609], x[608], x[607], x[606], x[605], x[604], x[603], x[602], x[601], x[600], x[599], x[598]}), .y(y[273]));
  R2ind274 R2ind274_inst(.x({x[609], x[608], x[607], x[603], x[602], x[601], x[606], x[605], x[604], x[600], x[599], x[598]}), .y(y[274]));
  R2ind275 R2ind275_inst(.x({x[609], x[608], x[607], x[603], x[602], x[601], x[606], x[605], x[604], x[600], x[599], x[598]}), .y(y[275]));
  R2ind276 R2ind276_inst(.x({x[609], x[608], x[607], x[603], x[602], x[601], x[606], x[605], x[604], x[600], x[599], x[598]}), .y(y[276]));
  R2ind277 R2ind277_inst(.x({x[609], x[608], x[607], x[603], x[602], x[601], x[606], x[605], x[604], x[600], x[599], x[598]}), .y(y[277]));
  R2ind278 R2ind278_inst(.x({x[609], x[608], x[607], x[603], x[602], x[601], x[600], x[599], x[598], x[606], x[605], x[604]}), .y(y[278]));
  R2ind279 R2ind279_inst(.x({x[609], x[608], x[607], x[603], x[602], x[601], x[600], x[599], x[598], x[606], x[605], x[604]}), .y(y[279]));
  R2ind280 R2ind280_inst(.x({x[611], x[610], x[27], x[26], x[25]}), .y(y[280]));
  R2ind281 R2ind281_inst(.x({x[611], x[610], x[27], x[26], x[25]}), .y(y[281]));
  R2ind282 R2ind282_inst(.x({x[613], x[612], x[27], x[26], x[25]}), .y(y[282]));
  R2ind283 R2ind283_inst(.x({x[613], x[612], x[27], x[26], x[25]}), .y(y[283]));
  R2ind284 R2ind284_inst(.x({x[615], x[614], x[27], x[26], x[25]}), .y(y[284]));
  R2ind285 R2ind285_inst(.x({x[615], x[614], x[27], x[26], x[25]}), .y(y[285]));
  R2ind286 R2ind286_inst(.x({x[617], x[616], x[27], x[26], x[25]}), .y(y[286]));
  R2ind287 R2ind287_inst(.x({x[617], x[616], x[27], x[26], x[25]}), .y(y[287]));
  R2ind288 R2ind288_inst(.x({x[619], x[618], x[27], x[26], x[25]}), .y(y[288]));
  R2ind289 R2ind289_inst(.x({x[619], x[618], x[27], x[26], x[25]}), .y(y[289]));
  R2ind290 R2ind290_inst(.x({x[621], x[620], x[27], x[26], x[25]}), .y(y[290]));
  R2ind291 R2ind291_inst(.x({x[621], x[620], x[27], x[26], x[25]}), .y(y[291]));
  R2ind292 R2ind292_inst(.x({x[623], x[622], x[27], x[26], x[25]}), .y(y[292]));
  R2ind293 R2ind293_inst(.x({x[623], x[622], x[27], x[26], x[25]}), .y(y[293]));
  R2ind294 R2ind294_inst(.x({x[625], x[624], x[27], x[26], x[25]}), .y(y[294]));
  R2ind295 R2ind295_inst(.x({x[625], x[624], x[27], x[26], x[25]}), .y(y[295]));
  R2ind296 R2ind296_inst(.x({x[627], x[626], x[27], x[26], x[25]}), .y(y[296]));
  R2ind297 R2ind297_inst(.x({x[627], x[626], x[27], x[26], x[25]}), .y(y[297]));
  R2ind298 R2ind298_inst(.x({x[629], x[628], x[27], x[26], x[25]}), .y(y[298]));
  R2ind299 R2ind299_inst(.x({x[629], x[628], x[27], x[26], x[25]}), .y(y[299]));
  R2ind300 R2ind300_inst(.x({x[631], x[630], x[27], x[26], x[25]}), .y(y[300]));
  R2ind301 R2ind301_inst(.x({x[631], x[630], x[27], x[26], x[25]}), .y(y[301]));
  R2ind302 R2ind302_inst(.x({x[633], x[632], x[27], x[26], x[25]}), .y(y[302]));
  R2ind303 R2ind303_inst(.x({x[633], x[632], x[27], x[26], x[25]}), .y(y[303]));
  R2ind304 R2ind304_inst(.x({x[635], x[634], x[27], x[26], x[25]}), .y(y[304]));
  R2ind305 R2ind305_inst(.x({x[635], x[634], x[27], x[26], x[25]}), .y(y[305]));
  R2ind306 R2ind306_inst(.x({x[637], x[636], x[27], x[26], x[25]}), .y(y[306]));
  R2ind307 R2ind307_inst(.x({x[637], x[636], x[27], x[26], x[25]}), .y(y[307]));
  R2ind308 R2ind308_inst(.x({x[639], x[638], x[27], x[26], x[25]}), .y(y[308]));
  R2ind309 R2ind309_inst(.x({x[639], x[638], x[27], x[26], x[25]}), .y(y[309]));
  R2ind310 R2ind310_inst(.x({x[641], x[640], x[27], x[26], x[25]}), .y(y[310]));
  R2ind311 R2ind311_inst(.x({x[641], x[640], x[27], x[26], x[25]}), .y(y[311]));
  R2ind312 R2ind312_inst(.x({x[643], x[642], x[27], x[26], x[25]}), .y(y[312]));
  R2ind313 R2ind313_inst(.x({x[643], x[642], x[27], x[26], x[25]}), .y(y[313]));
  R2ind314 R2ind314_inst(.x({x[645], x[644], x[27], x[26], x[25]}), .y(y[314]));
  R2ind315 R2ind315_inst(.x({x[645], x[644], x[27], x[26], x[25]}), .y(y[315]));
  R2ind316 R2ind316_inst(.x({x[647], x[646], x[27], x[26], x[25]}), .y(y[316]));
  R2ind317 R2ind317_inst(.x({x[647], x[646], x[27], x[26], x[25]}), .y(y[317]));
  R2ind318 R2ind318_inst(.x({x[649], x[648], x[27], x[26], x[25]}), .y(y[318]));
  R2ind319 R2ind319_inst(.x({x[649], x[648], x[27], x[26], x[25]}), .y(y[319]));
  R2ind320 R2ind320_inst(.x({x[651], x[650], x[27], x[26], x[25]}), .y(y[320]));
  R2ind321 R2ind321_inst(.x({x[651], x[650], x[27], x[26], x[25]}), .y(y[321]));
  R2ind322 R2ind322_inst(.x({x[653], x[652], x[27], x[26], x[25]}), .y(y[322]));
  R2ind323 R2ind323_inst(.x({x[653], x[652], x[27], x[26], x[25]}), .y(y[323]));
  R2ind324 R2ind324_inst(.x({x[655], x[654], x[27], x[26], x[25]}), .y(y[324]));
  R2ind325 R2ind325_inst(.x({x[655], x[654], x[27], x[26], x[25]}), .y(y[325]));
  R2ind326 R2ind326_inst(.x({x[657], x[656], x[27], x[26], x[25]}), .y(y[326]));
  R2ind327 R2ind327_inst(.x({x[657], x[656], x[27], x[26], x[25]}), .y(y[327]));
  R2ind328 R2ind328_inst(.x({x[659], x[658], x[27], x[26], x[25]}), .y(y[328]));
  R2ind329 R2ind329_inst(.x({x[659], x[658], x[27], x[26], x[25]}), .y(y[329]));
  R2ind330 R2ind330_inst(.x({x[661], x[660], x[27], x[26], x[25]}), .y(y[330]));
  R2ind331 R2ind331_inst(.x({x[661], x[660], x[27], x[26], x[25]}), .y(y[331]));
  R2ind332 R2ind332_inst(.x({x[663], x[662], x[27], x[26], x[25]}), .y(y[332]));
  R2ind333 R2ind333_inst(.x({x[663], x[662], x[27], x[26], x[25]}), .y(y[333]));
  R2ind334 R2ind334_inst(.x({x[665], x[664], x[27], x[26], x[25]}), .y(y[334]));
  R2ind335 R2ind335_inst(.x({x[665], x[664], x[27], x[26], x[25]}), .y(y[335]));
  R2ind336 R2ind336_inst(.x({x[667], x[666], x[27], x[26], x[25]}), .y(y[336]));
  R2ind337 R2ind337_inst(.x({x[667], x[666], x[27], x[26], x[25]}), .y(y[337]));
  R2ind338 R2ind338_inst(.x({x[669], x[668], x[27], x[26], x[25]}), .y(y[338]));
  R2ind339 R2ind339_inst(.x({x[669], x[668], x[27], x[26], x[25]}), .y(y[339]));
  R2ind340 R2ind340_inst(.x({x[671], x[670], x[27], x[26], x[25]}), .y(y[340]));
  R2ind341 R2ind341_inst(.x({x[671], x[670], x[27], x[26], x[25]}), .y(y[341]));
  R2ind342 R2ind342_inst(.x({x[673], x[672], x[27], x[26], x[25]}), .y(y[342]));
  R2ind343 R2ind343_inst(.x({x[673], x[672], x[27], x[26], x[25]}), .y(y[343]));
  R2ind344 R2ind344_inst(.x({x[675], x[674], x[27], x[26], x[25]}), .y(y[344]));
  R2ind345 R2ind345_inst(.x({x[675], x[674], x[27], x[26], x[25]}), .y(y[345]));
  R2ind346 R2ind346_inst(.x({x[677], x[676], x[27], x[26], x[25]}), .y(y[346]));
  R2ind347 R2ind347_inst(.x({x[677], x[676], x[27], x[26], x[25]}), .y(y[347]));
  R2ind348 R2ind348_inst(.x({x[679], x[678], x[27], x[26], x[25]}), .y(y[348]));
  R2ind349 R2ind349_inst(.x({x[679], x[678], x[27], x[26], x[25]}), .y(y[349]));
  R2ind350 R2ind350_inst(.x({x[681], x[680], x[27], x[26], x[25]}), .y(y[350]));
  R2ind351 R2ind351_inst(.x({x[681], x[680], x[27], x[26], x[25]}), .y(y[351]));
  R2ind352 R2ind352_inst(.x({x[683], x[682], x[27], x[26], x[25]}), .y(y[352]));
  R2ind353 R2ind353_inst(.x({x[683], x[682], x[27], x[26], x[25]}), .y(y[353]));
  R2ind354 R2ind354_inst(.x({x[685], x[684], x[27], x[26], x[25]}), .y(y[354]));
  R2ind355 R2ind355_inst(.x({x[685], x[684], x[27], x[26], x[25]}), .y(y[355]));
  R2ind356 R2ind356_inst(.x({x[687], x[686], x[27], x[26], x[25]}), .y(y[356]));
  R2ind357 R2ind357_inst(.x({x[687], x[686], x[27], x[26], x[25]}), .y(y[357]));
  R2ind358 R2ind358_inst(.x({x[689], x[688], x[27], x[26], x[25]}), .y(y[358]));
  R2ind359 R2ind359_inst(.x({x[689], x[688], x[27], x[26], x[25]}), .y(y[359]));
  R2ind360 R2ind360_inst(.x({x[9], x[8], x[7], x[3], x[691], x[690], x[27], x[26], x[25]}), .y(y[360]));
  R2ind361 R2ind361_inst(.x({x[9], x[8], x[7], x[3], x[691], x[690], x[27], x[26], x[25]}), .y(y[361]));
  R2ind362 R2ind362_inst(.x({x[15], x[14], x[13], x[3], x[693], x[692], x[27], x[26], x[25]}), .y(y[362]));
  R2ind363 R2ind363_inst(.x({x[15], x[14], x[13], x[3], x[693], x[692], x[27], x[26], x[25]}), .y(y[363]));
  R2ind364 R2ind364_inst(.x({x[12], x[11], x[10], x[3], x[695], x[694], x[27], x[26], x[25]}), .y(y[364]));
  R2ind365 R2ind365_inst(.x({x[12], x[11], x[10], x[3], x[695], x[694], x[27], x[26], x[25]}), .y(y[365]));
  R2ind366 R2ind366_inst(.x({x[697], x[696], x[27], x[26], x[25]}), .y(y[366]));
  R2ind367 R2ind367_inst(.x({x[697], x[696], x[27], x[26], x[25]}), .y(y[367]));
  R2ind368 R2ind368_inst(.x({x[18], x[17], x[16], x[3], x[699], x[698], x[27], x[26], x[25]}), .y(y[368]));
  R2ind369 R2ind369_inst(.x({x[18], x[17], x[16], x[3], x[699], x[698], x[27], x[26], x[25]}), .y(y[369]));
  R2ind370 R2ind370_inst(.x({x[21], x[20], x[19], x[3], x[701], x[700], x[27], x[26], x[25]}), .y(y[370]));
  R2ind371 R2ind371_inst(.x({x[21], x[20], x[19], x[3], x[701], x[700], x[27], x[26], x[25]}), .y(y[371]));
  R2ind372 R2ind372_inst(.x({x[24], x[23], x[22], x[3], x[703], x[702], x[27], x[26], x[25]}), .y(y[372]));
  R2ind373 R2ind373_inst(.x({x[24], x[23], x[22], x[3], x[703], x[702], x[27], x[26], x[25]}), .y(y[373]));
  R2ind374 R2ind374_inst(.x({x[6], x[5], x[4], x[3], x[705], x[704], x[27], x[26], x[25]}), .y(y[374]));
  R2ind375 R2ind375_inst(.x({x[6], x[5], x[4], x[3], x[705], x[704], x[27], x[26], x[25]}), .y(y[375]));
  R2ind376 R2ind376_inst(.x({x[707], x[706], x[27], x[26], x[25]}), .y(y[376]));
  R2ind377 R2ind377_inst(.x({x[707], x[706], x[27], x[26], x[25]}), .y(y[377]));
  R2ind378 R2ind378_inst(.x({x[709], x[708], x[27], x[26], x[25]}), .y(y[378]));
  R2ind379 R2ind379_inst(.x({x[709], x[708], x[27], x[26], x[25]}), .y(y[379]));
  R2ind380 R2ind380_inst(.x({x[711], x[710], x[27], x[26], x[25]}), .y(y[380]));
  R2ind381 R2ind381_inst(.x({x[711], x[710], x[27], x[26], x[25]}), .y(y[381]));
  R2ind382 R2ind382_inst(.x({x[713], x[712], x[27], x[26], x[25]}), .y(y[382]));
  R2ind383 R2ind383_inst(.x({x[713], x[712], x[27], x[26], x[25]}), .y(y[383]));
  R2ind384 R2ind384_inst(.x({x[715], x[714], x[27], x[26], x[25]}), .y(y[384]));
  R2ind385 R2ind385_inst(.x({x[715], x[714], x[27], x[26], x[25]}), .y(y[385]));
  R2ind386 R2ind386_inst(.x({x[717], x[716], x[27], x[26], x[25]}), .y(y[386]));
  R2ind387 R2ind387_inst(.x({x[717], x[716], x[27], x[26], x[25]}), .y(y[387]));
  R2ind388 R2ind388_inst(.x({x[719], x[718], x[27], x[26], x[25]}), .y(y[388]));
  R2ind389 R2ind389_inst(.x({x[719], x[718], x[27], x[26], x[25]}), .y(y[389]));
  R2ind390 R2ind390_inst(.x({x[721], x[720], x[27], x[26], x[25]}), .y(y[390]));
  R2ind391 R2ind391_inst(.x({x[721], x[720], x[27], x[26], x[25]}), .y(y[391]));
  R2ind392 R2ind392_inst(.x({x[723], x[722], x[27], x[26], x[25]}), .y(y[392]));
  R2ind393 R2ind393_inst(.x({x[723], x[722], x[27], x[26], x[25]}), .y(y[393]));
  R2ind394 R2ind394_inst(.x({x[725], x[724], x[27], x[26], x[25]}), .y(y[394]));
  R2ind395 R2ind395_inst(.x({x[725], x[724], x[27], x[26], x[25]}), .y(y[395]));
  R2ind396 R2ind396_inst(.x({x[727], x[726], x[27], x[26], x[25]}), .y(y[396]));
  R2ind397 R2ind397_inst(.x({x[727], x[726], x[27], x[26], x[25]}), .y(y[397]));
  R2ind398 R2ind398_inst(.x({x[729], x[728], x[27], x[26], x[25]}), .y(y[398]));
  R2ind399 R2ind399_inst(.x({x[729], x[728], x[27], x[26], x[25]}), .y(y[399]));
  R2ind400 R2ind400_inst(.x({x[731], x[730], x[27], x[26], x[25]}), .y(y[400]));
  R2ind401 R2ind401_inst(.x({x[731], x[730], x[27], x[26], x[25]}), .y(y[401]));
  R2ind402 R2ind402_inst(.x({x[733], x[732], x[27], x[26], x[25]}), .y(y[402]));
  R2ind403 R2ind403_inst(.x({x[733], x[732], x[27], x[26], x[25]}), .y(y[403]));
  R2ind404 R2ind404_inst(.x({x[735], x[734], x[27], x[26], x[25]}), .y(y[404]));
  R2ind405 R2ind405_inst(.x({x[735], x[734], x[27], x[26], x[25]}), .y(y[405]));
  R2ind406 R2ind406_inst(.x({x[737], x[736], x[27], x[26], x[25]}), .y(y[406]));
  R2ind407 R2ind407_inst(.x({x[737], x[736], x[27], x[26], x[25]}), .y(y[407]));
endmodule

