/* modified netlist. Source: module PRESENT in file ../CaseStudies/10_PRESENT80_nibble_serial_encryption/netlists/PRESENT.v */
/* 0 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 1 register stage(s) in total */

module PRESENT_LMDPL_Pipeline_d1 (data_in_s0, key_s0, clk, reset, Po_rst, Fresh, data_in_s1, key_s1, data_out_s0, done, data_out_s1);
    input [63:0] data_in_s0 ;
    input [79:0] key_s0 ;
    input clk ;
    input reset ;
    input Po_rst ;
    input [63:0] data_in_s1 ;
    input [79:0] key_s1 ;
    input [3:0] Fresh ;
    output [63:0] data_out_s0 ;
    output done ;
    output [63:0] data_out_s1 ;
    wire selSbox ;
    wire ctrlData_0_ ;
    wire intDone ;
    wire fsm_n15 ;
    wire fsm_n14 ;
    wire fsm_n13 ;
    wire fsm_n12 ;
    wire fsm_n11 ;
    wire fsm_n10 ;
    wire fsm_n9 ;
    wire fsm_n8 ;
    wire fsm_n7 ;
    wire fsm_n6 ;
    wire fsm_n4 ;
    wire fsm_n2 ;
    wire fsm_n5 ;
    wire fsm_n20 ;
    wire fsm_ps_state_0_ ;
    wire fsm_ps_state_1_ ;
    wire fsm_n21 ;
    wire fsm_n3 ;
    wire fsm_rst_countSerial ;
    wire fsm_en_countRound ;
    wire fsm_cnt_rnd_n33 ;
    wire fsm_cnt_rnd_n32 ;
    wire fsm_cnt_rnd_n31 ;
    wire fsm_cnt_rnd_n30 ;
    wire fsm_cnt_rnd_n29 ;
    wire fsm_cnt_rnd_n28 ;
    wire fsm_cnt_rnd_n27 ;
    wire fsm_cnt_rnd_n26 ;
    wire fsm_cnt_rnd_n23 ;
    wire fsm_cnt_rnd_n22 ;
    wire fsm_cnt_rnd_n21 ;
    wire fsm_cnt_rnd_n20 ;
    wire fsm_cnt_rnd_n19 ;
    wire fsm_cnt_rnd_n17 ;
    wire fsm_cnt_rnd_n15 ;
    wire fsm_cnt_rnd_n13 ;
    wire fsm_cnt_rnd_n12 ;
    wire fsm_cnt_rnd_n11 ;
    wire fsm_cnt_rnd_n10 ;
    wire fsm_cnt_rnd_n9 ;
    wire fsm_cnt_rnd_n8 ;
    wire fsm_cnt_rnd_n7 ;
    wire fsm_cnt_rnd_n6 ;
    wire fsm_cnt_rnd_n5 ;
    wire fsm_cnt_rnd_n3 ;
    wire fsm_cnt_rnd_n24 ;
    wire fsm_cnt_rnd_n41 ;
    wire fsm_cnt_rnd_n25 ;
    wire fsm_cnt_rnd_n1 ;
    wire fsm_cnt_rnd_n18 ;
    wire fsm_cnt_rnd_n16 ;
    wire fsm_cnt_rnd_n14 ;
    wire fsm_cnt_ser_n10 ;
    wire fsm_cnt_ser_n9 ;
    wire fsm_cnt_ser_n8 ;
    wire fsm_cnt_ser_n7 ;
    wire fsm_cnt_ser_n6 ;
    wire fsm_cnt_ser_n5 ;
    wire fsm_cnt_ser_n4 ;
    wire fsm_cnt_ser_n2 ;
    wire fsm_cnt_ser_n20 ;
    wire fsm_cnt_ser_n28 ;
    wire fsm_cnt_ser_n26 ;
    wire fsm_cnt_ser_n3 ;
    wire fsm_cnt_ser_n1 ;
    wire stateFF_state_n7 ;
    wire stateFF_state_n6 ;
    wire stateFF_state_n5 ;
    wire keyFF_keystate_n8 ;
    wire keyFF_keystate_n7 ;
    wire keyFF_keystate_n6 ;
    wire sboxInst_n3 ;
    wire sboxInst_n2 ;
    wire sboxInst_n1 ;
    wire sboxInst_L8 ;
    wire sboxInst_L7 ;
    wire sboxInst_T3 ;
    wire sboxInst_T1 ;
    wire sboxInst_Q7 ;
    wire sboxInst_Q6 ;
    wire sboxInst_L5 ;
    wire sboxInst_T2 ;
    wire sboxInst_L4 ;
    wire sboxInst_Q3 ;
    wire sboxInst_L3 ;
    wire sboxInst_Q2 ;
    wire sboxInst_T0 ;
    wire sboxInst_L2 ;
    wire sboxInst_L1 ;
    wire sboxInst_L0 ;
    wire [4:0] counter ;
    wire [3:0] serialIn ;
    wire [3:0] sboxOut ;
    wire [3:0] roundkey ;
    wire [3:1] keyRegKS ;
    wire [3:0] sboxIn ;
    wire [3:0] stateXORroundkey ;
    wire [3:0] fsm_countSerial ;
    wire [63:0] stateFF_inputPar ;
    wire [3:0] stateFF_state_gff_1_s_next_state ;
    wire [3:0] stateFF_state_gff_2_s_next_state ;
    wire [3:0] stateFF_state_gff_3_s_next_state ;
    wire [3:0] stateFF_state_gff_4_s_next_state ;
    wire [3:0] stateFF_state_gff_5_s_next_state ;
    wire [3:0] stateFF_state_gff_6_s_next_state ;
    wire [3:0] stateFF_state_gff_7_s_next_state ;
    wire [3:0] stateFF_state_gff_8_s_next_state ;
    wire [3:0] stateFF_state_gff_9_s_next_state ;
    wire [3:0] stateFF_state_gff_10_s_next_state ;
    wire [3:0] stateFF_state_gff_11_s_next_state ;
    wire [3:0] stateFF_state_gff_12_s_next_state ;
    wire [3:0] stateFF_state_gff_13_s_next_state ;
    wire [3:0] stateFF_state_gff_14_s_next_state ;
    wire [3:0] stateFF_state_gff_15_s_next_state ;
    wire [3:0] stateFF_state_gff_16_s_next_state ;
    wire [4:0] keyFF_counterAdd ;
    wire [75:3] keyFF_outputPar ;
    wire [79:0] keyFF_inputPar ;
    wire [3:0] keyFF_keystate_gff_1_s_next_state ;
    wire [3:0] keyFF_keystate_gff_2_s_next_state ;
    wire [3:0] keyFF_keystate_gff_3_s_next_state ;
    wire [3:0] keyFF_keystate_gff_4_s_next_state ;
    wire [3:0] keyFF_keystate_gff_5_s_next_state ;
    wire [3:0] keyFF_keystate_gff_6_s_next_state ;
    wire [3:0] keyFF_keystate_gff_7_s_next_state ;
    wire [3:0] keyFF_keystate_gff_8_s_next_state ;
    wire [3:0] keyFF_keystate_gff_9_s_next_state ;
    wire [3:0] keyFF_keystate_gff_10_s_next_state ;
    wire [3:0] keyFF_keystate_gff_11_s_next_state ;
    wire [3:0] keyFF_keystate_gff_12_s_next_state ;
    wire [3:0] keyFF_keystate_gff_13_s_next_state ;
    wire [3:0] keyFF_keystate_gff_14_s_next_state ;
    wire [3:0] keyFF_keystate_gff_15_s_next_state ;
    wire [3:0] keyFF_keystate_gff_16_s_next_state ;
    wire [3:0] keyFF_keystate_gff_17_s_next_state ;
    wire [3:0] keyFF_keystate_gff_18_s_next_state ;
    wire [3:0] keyFF_keystate_gff_19_s_next_state ;
    wire [3:0] keyFF_keystate_gff_20_s_next_state ;
    wire LMDPL_pre1 ;
    wire LMDPL_pre2 ;
    wire mid_rst ;
    wire new_AGEMA_signal_860 ;
    wire new_AGEMA_signal_861 ;
    wire new_AGEMA_signal_863 ;
    wire new_AGEMA_signal_864 ;
    wire new_AGEMA_signal_865 ;
    wire new_AGEMA_signal_866 ;
    wire new_AGEMA_signal_867 ;
    wire new_AGEMA_signal_869 ;
    wire new_AGEMA_signal_870 ;
    wire new_AGEMA_signal_871 ;
    wire new_AGEMA_signal_872 ;
    wire new_AGEMA_signal_873 ;
    wire new_AGEMA_signal_875 ;
    wire new_AGEMA_signal_876 ;
    wire new_AGEMA_signal_877 ;
    wire new_AGEMA_signal_878 ;
    wire new_AGEMA_signal_879 ;
    wire new_AGEMA_signal_881 ;
    wire new_AGEMA_signal_882 ;
    wire new_AGEMA_signal_883 ;
    wire new_AGEMA_signal_884 ;
    wire new_AGEMA_signal_885 ;
    wire new_AGEMA_signal_887 ;
    wire new_AGEMA_signal_888 ;
    wire new_AGEMA_signal_889 ;
    wire new_AGEMA_signal_890 ;
    wire new_AGEMA_signal_891 ;
    wire new_AGEMA_signal_893 ;
    wire new_AGEMA_signal_894 ;
    wire new_AGEMA_signal_895 ;
    wire new_AGEMA_signal_896 ;
    wire new_AGEMA_signal_897 ;
    wire new_AGEMA_signal_899 ;
    wire new_AGEMA_signal_900 ;
    wire new_AGEMA_signal_901 ;
    wire new_AGEMA_signal_902 ;
    wire new_AGEMA_signal_903 ;
    wire new_AGEMA_signal_905 ;
    wire new_AGEMA_signal_906 ;
    wire new_AGEMA_signal_907 ;
    wire new_AGEMA_signal_908 ;
    wire new_AGEMA_signal_909 ;
    wire new_AGEMA_signal_911 ;
    wire new_AGEMA_signal_912 ;
    wire new_AGEMA_signal_913 ;
    wire new_AGEMA_signal_914 ;
    wire new_AGEMA_signal_915 ;
    wire new_AGEMA_signal_917 ;
    wire new_AGEMA_signal_918 ;
    wire new_AGEMA_signal_919 ;
    wire new_AGEMA_signal_920 ;
    wire new_AGEMA_signal_921 ;
    wire new_AGEMA_signal_923 ;
    wire new_AGEMA_signal_924 ;
    wire new_AGEMA_signal_925 ;
    wire new_AGEMA_signal_926 ;
    wire new_AGEMA_signal_927 ;
    wire new_AGEMA_signal_929 ;
    wire new_AGEMA_signal_930 ;
    wire new_AGEMA_signal_931 ;
    wire new_AGEMA_signal_932 ;
    wire new_AGEMA_signal_933 ;
    wire new_AGEMA_signal_935 ;
    wire new_AGEMA_signal_936 ;
    wire new_AGEMA_signal_937 ;
    wire new_AGEMA_signal_938 ;
    wire new_AGEMA_signal_939 ;
    wire new_AGEMA_signal_941 ;
    wire new_AGEMA_signal_942 ;
    wire new_AGEMA_signal_943 ;
    wire new_AGEMA_signal_944 ;
    wire new_AGEMA_signal_945 ;
    wire new_AGEMA_signal_947 ;
    wire new_AGEMA_signal_948 ;
    wire new_AGEMA_signal_949 ;
    wire new_AGEMA_signal_950 ;
    wire new_AGEMA_signal_951 ;
    wire new_AGEMA_signal_953 ;
    wire new_AGEMA_signal_954 ;
    wire new_AGEMA_signal_955 ;
    wire new_AGEMA_signal_956 ;
    wire new_AGEMA_signal_957 ;
    wire new_AGEMA_signal_959 ;
    wire new_AGEMA_signal_960 ;
    wire new_AGEMA_signal_961 ;
    wire new_AGEMA_signal_962 ;
    wire new_AGEMA_signal_963 ;
    wire new_AGEMA_signal_965 ;
    wire new_AGEMA_signal_966 ;
    wire new_AGEMA_signal_967 ;
    wire new_AGEMA_signal_968 ;
    wire new_AGEMA_signal_969 ;
    wire new_AGEMA_signal_971 ;
    wire new_AGEMA_signal_972 ;
    wire new_AGEMA_signal_973 ;
    wire new_AGEMA_signal_974 ;
    wire new_AGEMA_signal_975 ;
    wire new_AGEMA_signal_976 ;
    wire new_AGEMA_signal_977 ;
    wire new_AGEMA_signal_978 ;
    wire new_AGEMA_signal_979 ;
    wire new_AGEMA_signal_981 ;
    wire new_AGEMA_signal_982 ;
    wire new_AGEMA_signal_983 ;
    wire new_AGEMA_signal_984 ;
    wire new_AGEMA_signal_985 ;
    wire new_AGEMA_signal_987 ;
    wire new_AGEMA_signal_988 ;
    wire new_AGEMA_signal_989 ;
    wire new_AGEMA_signal_990 ;
    wire new_AGEMA_signal_991 ;
    wire new_AGEMA_signal_993 ;
    wire new_AGEMA_signal_994 ;
    wire new_AGEMA_signal_995 ;
    wire new_AGEMA_signal_996 ;
    wire new_AGEMA_signal_997 ;
    wire new_AGEMA_signal_999 ;
    wire new_AGEMA_signal_1000 ;
    wire new_AGEMA_signal_1001 ;
    wire new_AGEMA_signal_1002 ;
    wire new_AGEMA_signal_1003 ;
    wire new_AGEMA_signal_1005 ;
    wire new_AGEMA_signal_1006 ;
    wire new_AGEMA_signal_1007 ;
    wire new_AGEMA_signal_1008 ;
    wire new_AGEMA_signal_1009 ;
    wire new_AGEMA_signal_1011 ;
    wire new_AGEMA_signal_1012 ;
    wire new_AGEMA_signal_1013 ;
    wire new_AGEMA_signal_1014 ;
    wire new_AGEMA_signal_1015 ;
    wire new_AGEMA_signal_1017 ;
    wire new_AGEMA_signal_1018 ;
    wire new_AGEMA_signal_1019 ;
    wire new_AGEMA_signal_1020 ;
    wire new_AGEMA_signal_1021 ;
    wire new_AGEMA_signal_1023 ;
    wire new_AGEMA_signal_1024 ;
    wire new_AGEMA_signal_1025 ;
    wire new_AGEMA_signal_1026 ;
    wire new_AGEMA_signal_1027 ;
    wire new_AGEMA_signal_1029 ;
    wire new_AGEMA_signal_1030 ;
    wire new_AGEMA_signal_1031 ;
    wire new_AGEMA_signal_1032 ;
    wire new_AGEMA_signal_1033 ;
    wire new_AGEMA_signal_1035 ;
    wire new_AGEMA_signal_1036 ;
    wire new_AGEMA_signal_1037 ;
    wire new_AGEMA_signal_1038 ;
    wire new_AGEMA_signal_1039 ;
    wire new_AGEMA_signal_1041 ;
    wire new_AGEMA_signal_1042 ;
    wire new_AGEMA_signal_1043 ;
    wire new_AGEMA_signal_1044 ;
    wire new_AGEMA_signal_1045 ;
    wire new_AGEMA_signal_1047 ;
    wire new_AGEMA_signal_1048 ;
    wire new_AGEMA_signal_1049 ;
    wire new_AGEMA_signal_1050 ;
    wire new_AGEMA_signal_1051 ;
    wire new_AGEMA_signal_1053 ;
    wire new_AGEMA_signal_1054 ;
    wire new_AGEMA_signal_1055 ;
    wire new_AGEMA_signal_1056 ;
    wire new_AGEMA_signal_1057 ;
    wire new_AGEMA_signal_1059 ;
    wire new_AGEMA_signal_1060 ;
    wire new_AGEMA_signal_1061 ;
    wire new_AGEMA_signal_1062 ;
    wire new_AGEMA_signal_1063 ;
    wire new_AGEMA_signal_1065 ;
    wire new_AGEMA_signal_1066 ;
    wire new_AGEMA_signal_1067 ;
    wire new_AGEMA_signal_1068 ;
    wire new_AGEMA_signal_1069 ;
    wire new_AGEMA_signal_1070 ;
    wire new_AGEMA_signal_1071 ;
    wire new_AGEMA_signal_1072 ;
    wire new_AGEMA_signal_1073 ;
    wire new_AGEMA_signal_1075 ;
    wire new_AGEMA_signal_1076 ;
    wire new_AGEMA_signal_1077 ;
    wire new_AGEMA_signal_1078 ;
    wire new_AGEMA_signal_1079 ;
    wire new_AGEMA_signal_1081 ;
    wire new_AGEMA_signal_1082 ;
    wire new_AGEMA_signal_1083 ;
    wire new_AGEMA_signal_1084 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1087 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1089 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1091 ;
    wire new_AGEMA_signal_1093 ;
    wire new_AGEMA_signal_1094 ;
    wire new_AGEMA_signal_1095 ;
    wire new_AGEMA_signal_1096 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1099 ;
    wire new_AGEMA_signal_1100 ;
    wire new_AGEMA_signal_1101 ;
    wire new_AGEMA_signal_1102 ;
    wire new_AGEMA_signal_1103 ;
    wire new_AGEMA_signal_1105 ;
    wire new_AGEMA_signal_1106 ;
    wire new_AGEMA_signal_1107 ;
    wire new_AGEMA_signal_1108 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1111 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1113 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1115 ;
    wire new_AGEMA_signal_1117 ;
    wire new_AGEMA_signal_1118 ;
    wire new_AGEMA_signal_1119 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1121 ;
    wire new_AGEMA_signal_1123 ;
    wire new_AGEMA_signal_1124 ;
    wire new_AGEMA_signal_1125 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1127 ;
    wire new_AGEMA_signal_1129 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1131 ;
    wire new_AGEMA_signal_1132 ;
    wire new_AGEMA_signal_1133 ;
    wire new_AGEMA_signal_1135 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1137 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1139 ;
    wire new_AGEMA_signal_1141 ;
    wire new_AGEMA_signal_1142 ;
    wire new_AGEMA_signal_1143 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1147 ;
    wire new_AGEMA_signal_1148 ;
    wire new_AGEMA_signal_1149 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1153 ;
    wire new_AGEMA_signal_1154 ;
    wire new_AGEMA_signal_1155 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1159 ;
    wire new_AGEMA_signal_1160 ;
    wire new_AGEMA_signal_1161 ;
    wire new_AGEMA_signal_1162 ;
    wire new_AGEMA_signal_1163 ;
    wire new_AGEMA_signal_1164 ;
    wire new_AGEMA_signal_1165 ;
    wire new_AGEMA_signal_1166 ;
    wire new_AGEMA_signal_1167 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1170 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1172 ;
    wire new_AGEMA_signal_1173 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1176 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1179 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1182 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1184 ;
    wire new_AGEMA_signal_1185 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1188 ;
    wire new_AGEMA_signal_1189 ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1193 ;
    wire new_AGEMA_signal_1194 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1196 ;
    wire new_AGEMA_signal_1197 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1200 ;
    wire new_AGEMA_signal_1201 ;
    wire new_AGEMA_signal_1202 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1206 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1208 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1211 ;
    wire new_AGEMA_signal_1212 ;
    wire new_AGEMA_signal_1213 ;
    wire new_AGEMA_signal_1214 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1217 ;
    wire new_AGEMA_signal_1218 ;
    wire new_AGEMA_signal_1219 ;
    wire new_AGEMA_signal_1220 ;
    wire new_AGEMA_signal_1221 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1224 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1227 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1230 ;
    wire new_AGEMA_signal_1231 ;
    wire new_AGEMA_signal_1232 ;
    wire new_AGEMA_signal_1233 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1236 ;
    wire new_AGEMA_signal_1237 ;
    wire new_AGEMA_signal_1238 ;
    wire new_AGEMA_signal_1239 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1242 ;
    wire new_AGEMA_signal_1243 ;
    wire new_AGEMA_signal_1244 ;
    wire new_AGEMA_signal_1245 ;
    wire new_AGEMA_signal_1247 ;
    wire new_AGEMA_signal_1248 ;
    wire new_AGEMA_signal_1249 ;
    wire new_AGEMA_signal_1250 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1253 ;
    wire new_AGEMA_signal_1254 ;
    wire new_AGEMA_signal_1255 ;
    wire new_AGEMA_signal_1256 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1259 ;
    wire new_AGEMA_signal_1260 ;
    wire new_AGEMA_signal_1261 ;
    wire new_AGEMA_signal_1262 ;
    wire new_AGEMA_signal_1263 ;
    wire new_AGEMA_signal_1264 ;
    wire new_AGEMA_signal_1265 ;
    wire new_AGEMA_signal_1266 ;
    wire new_AGEMA_signal_1267 ;
    wire new_AGEMA_signal_1268 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1270 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1272 ;
    wire new_AGEMA_signal_1273 ;
    wire new_AGEMA_signal_1274 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1276 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1278 ;
    wire new_AGEMA_signal_1279 ;
    wire new_AGEMA_signal_1280 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1282 ;
    wire new_AGEMA_signal_1283 ;
    wire new_AGEMA_signal_1284 ;
    wire new_AGEMA_signal_1285 ;
    wire new_AGEMA_signal_1286 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1288 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1291 ;
    wire new_AGEMA_signal_1292 ;
    wire new_AGEMA_signal_1293 ;
    wire new_AGEMA_signal_1294 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1296 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1300 ;
    wire new_AGEMA_signal_1301 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1304 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1308 ;
    wire new_AGEMA_signal_1309 ;
    wire new_AGEMA_signal_1310 ;
    wire new_AGEMA_signal_1311 ;
    wire new_AGEMA_signal_1312 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1316 ;
    wire new_AGEMA_signal_1317 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1320 ;
    wire new_AGEMA_signal_1321 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1326 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1344 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1352 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1364 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1381 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1400 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1412 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1441 ;
    wire new_AGEMA_signal_1442 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1444 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1456 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1459 ;
    wire new_AGEMA_signal_1460 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1465 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1471 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1474 ;
    wire new_AGEMA_signal_1475 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1483 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1492 ;
    wire new_AGEMA_signal_1493 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1501 ;
    wire new_AGEMA_signal_1502 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1510 ;
    wire new_AGEMA_signal_1511 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1519 ;
    wire new_AGEMA_signal_1520 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1522 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1528 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1547 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1555 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1559 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1563 ;
    wire new_AGEMA_signal_1564 ;
    wire new_AGEMA_signal_1565 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1573 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1579 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1581 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1583 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1591 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1593 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1599 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1609 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1619 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1627 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1645 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1653 ;
    wire new_AGEMA_signal_1654 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1663 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1699 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1701 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1789 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1799 ;
    wire new_AGEMA_signal_1800 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1835 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1870 ;
    wire new_AGEMA_signal_1871 ;
    wire new_AGEMA_signal_1872 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1880 ;
    wire new_AGEMA_signal_1881 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1888 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1896 ;
    wire new_AGEMA_signal_1897 ;
    wire new_AGEMA_signal_1898 ;
    wire new_AGEMA_signal_1899 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1906 ;
    wire new_AGEMA_signal_1907 ;
    wire new_AGEMA_signal_1908 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1914 ;
    wire new_AGEMA_signal_1915 ;
    wire new_AGEMA_signal_1916 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1923 ;
    wire new_AGEMA_signal_1924 ;
    wire new_AGEMA_signal_1925 ;
    wire new_AGEMA_signal_1926 ;
    wire new_AGEMA_signal_1927 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1931 ;
    wire new_AGEMA_signal_1932 ;
    wire new_AGEMA_signal_1933 ;
    wire new_AGEMA_signal_1934 ;
    wire new_AGEMA_signal_1935 ;
    wire new_AGEMA_signal_1936 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1938 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1940 ;
    wire new_AGEMA_signal_1941 ;
    wire new_AGEMA_signal_1942 ;
    wire new_AGEMA_signal_1943 ;
    wire new_AGEMA_signal_1944 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1947 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1949 ;
    wire new_AGEMA_signal_1950 ;
    wire new_AGEMA_signal_1951 ;
    wire new_AGEMA_signal_1952 ;
    wire new_AGEMA_signal_1953 ;
    wire new_AGEMA_signal_1954 ;
    wire new_AGEMA_signal_1955 ;
    wire new_AGEMA_signal_1956 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1958 ;
    wire new_AGEMA_signal_1959 ;
    wire new_AGEMA_signal_1960 ;
    wire new_AGEMA_signal_1961 ;
    wire new_AGEMA_signal_1962 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1967 ;
    wire new_AGEMA_signal_1968 ;
    wire new_AGEMA_signal_1969 ;
    wire new_AGEMA_signal_1970 ;
    wire new_AGEMA_signal_1971 ;
    wire new_AGEMA_signal_1972 ;
    wire new_AGEMA_signal_1973 ;
    wire new_AGEMA_signal_1974 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1976 ;
    wire new_AGEMA_signal_1977 ;
    wire new_AGEMA_signal_1978 ;
    wire new_AGEMA_signal_1979 ;
    wire new_AGEMA_signal_1980 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1985 ;
    wire new_AGEMA_signal_1986 ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1988 ;
    wire new_AGEMA_signal_1989 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1995 ;
    wire new_AGEMA_signal_1996 ;
    wire new_AGEMA_signal_1997 ;
    wire new_AGEMA_signal_1998 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2003 ;
    wire new_AGEMA_signal_2004 ;
    wire new_AGEMA_signal_2005 ;
    wire new_AGEMA_signal_2006 ;
    wire new_AGEMA_signal_2007 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2014 ;
    wire new_AGEMA_signal_2015 ;
    wire new_AGEMA_signal_2016 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2022 ;
    wire new_AGEMA_signal_2023 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2025 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2032 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2034 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2041 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2043 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2050 ;
    wire new_AGEMA_signal_2051 ;
    wire new_AGEMA_signal_2052 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2059 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2061 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2086 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2097 ;
    wire new_AGEMA_signal_2098 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2102 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2104 ;
    wire new_AGEMA_signal_2105 ;
    wire new_AGEMA_signal_2106 ;
    wire new_AGEMA_signal_2107 ;

    /* cells in depth 0 */
    linear_LMDPL #(.CONF(1'b0)) U9 ( .a ({new_AGEMA_signal_861, new_AGEMA_signal_860, roundkey[0]}), .b ({new_AGEMA_signal_863, data_out_s1[60], data_out_s0[60]}), .c ({new_AGEMA_signal_865, new_AGEMA_signal_864, stateXORroundkey[0]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) U10 ( .a ({new_AGEMA_signal_867, new_AGEMA_signal_866, roundkey[1]}), .b ({new_AGEMA_signal_869, data_out_s1[61], data_out_s0[61]}), .c ({new_AGEMA_signal_871, new_AGEMA_signal_870, stateXORroundkey[1]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) U11 ( .a ({new_AGEMA_signal_873, new_AGEMA_signal_872, roundkey[2]}), .b ({new_AGEMA_signal_875, data_out_s1[62], data_out_s0[62]}), .c ({new_AGEMA_signal_877, new_AGEMA_signal_876, stateXORroundkey[2]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) U12 ( .a ({new_AGEMA_signal_879, new_AGEMA_signal_878, roundkey[3]}), .b ({new_AGEMA_signal_881, data_out_s1[63], data_out_s0[63]}), .c ({new_AGEMA_signal_883, new_AGEMA_signal_882, stateXORroundkey[3]}) ) ;
    NOR2_X1 fsm_U20 ( .A1 (reset), .A2 (fsm_n15), .ZN (fsm_n21) ) ;
    NOR2_X1 fsm_U19 ( .A1 (fsm_n14), .A2 (done), .ZN (fsm_n15) ) ;
    NOR2_X1 fsm_U18 ( .A1 (reset), .A2 (fsm_n13), .ZN (fsm_n20) ) ;
    NOR2_X1 fsm_U17 ( .A1 (fsm_ps_state_1_), .A2 (fsm_n12), .ZN (fsm_n13) ) ;
    NOR2_X1 fsm_U16 ( .A1 (fsm_n11), .A2 (fsm_n10), .ZN (fsm_n12) ) ;
    NAND2_X1 fsm_U15 ( .A1 (counter[3]), .A2 (counter[1]), .ZN (fsm_n10) ) ;
    OR2_X1 fsm_U14 ( .A1 (fsm_n9), .A2 (fsm_n8), .ZN (fsm_n11) ) ;
    NAND2_X1 fsm_U13 ( .A1 (counter[0]), .A2 (counter[4]), .ZN (fsm_n8) ) ;
    NAND2_X1 fsm_U12 ( .A1 (counter[2]), .A2 (fsm_ps_state_0_), .ZN (fsm_n9) ) ;
    NOR2_X1 fsm_U11 ( .A1 (fsm_n3), .A2 (fsm_n5), .ZN (done) ) ;
    AND2_X1 fsm_U10 ( .A1 (fsm_n14), .A2 (fsm_n5), .ZN (fsm_en_countRound) ) ;
    AND2_X1 fsm_U9 ( .A1 (fsm_countSerial[2]), .A2 (fsm_n7), .ZN (fsm_n14) ) ;
    NOR2_X1 fsm_U8 ( .A1 (fsm_n6), .A2 (fsm_n4), .ZN (fsm_n7) ) ;
    NAND2_X1 fsm_U7 ( .A1 (fsm_countSerial[1]), .A2 (fsm_countSerial[0]), .ZN (fsm_n4) ) ;
    NAND2_X1 fsm_U6 ( .A1 (fsm_n3), .A2 (fsm_countSerial[3]), .ZN (fsm_n6) ) ;
    NOR2_X1 fsm_U5 ( .A1 (fsm_ps_state_0_), .A2 (fsm_n5), .ZN (intDone) ) ;
    NOR2_X1 fsm_U4 ( .A1 (fsm_ps_state_1_), .A2 (fsm_n3), .ZN (selSbox) ) ;
    NOR2_X1 fsm_U3 ( .A1 (reset), .A2 (selSbox), .ZN (fsm_rst_countSerial) ) ;
    INV_X1 fsm_U2 ( .A (reset), .ZN (fsm_n2) ) ;
    INV_X1 fsm_U1 ( .A (fsm_rst_countSerial), .ZN (ctrlData_0_) ) ;
    NAND2_X1 fsm_cnt_rnd_U28 ( .A1 (fsm_cnt_rnd_n33), .A2 (fsm_cnt_rnd_n32), .ZN (fsm_cnt_rnd_n41) ) ;
    NAND2_X1 fsm_cnt_rnd_U27 ( .A1 (fsm_cnt_rnd_n31), .A2 (counter[1]), .ZN (fsm_cnt_rnd_n32) ) ;
    NAND2_X1 fsm_cnt_rnd_U26 ( .A1 (fsm_cnt_rnd_n30), .A2 (fsm_cnt_rnd_n24), .ZN (fsm_cnt_rnd_n33) ) ;
    NAND2_X1 fsm_cnt_rnd_U25 ( .A1 (fsm_cnt_rnd_n29), .A2 (counter[0]), .ZN (fsm_cnt_rnd_n30) ) ;
    NAND2_X1 fsm_cnt_rnd_U24 ( .A1 (fsm_cnt_rnd_n28), .A2 (fsm_cnt_rnd_n27), .ZN (fsm_cnt_rnd_n18) ) ;
    NAND2_X1 fsm_cnt_rnd_U23 ( .A1 (fsm_cnt_rnd_n26), .A2 (counter[0]), .ZN (fsm_cnt_rnd_n27) ) ;
    MUX2_X1 fsm_cnt_rnd_U22 ( .S (fsm_cnt_rnd_n5), .A (fsm_cnt_rnd_n23), .B (fsm_cnt_rnd_n22), .Z (fsm_cnt_rnd_n16) ) ;
    NAND2_X1 fsm_cnt_rnd_U21 ( .A1 (fsm_cnt_rnd_n31), .A2 (fsm_cnt_rnd_n21), .ZN (fsm_cnt_rnd_n23) ) ;
    NAND2_X1 fsm_cnt_rnd_U20 ( .A1 (fsm_cnt_rnd_n29), .A2 (fsm_cnt_rnd_n24), .ZN (fsm_cnt_rnd_n21) ) ;
    NOR2_X1 fsm_cnt_rnd_U19 ( .A1 (fsm_cnt_rnd_n20), .A2 (fsm_cnt_rnd_n26), .ZN (fsm_cnt_rnd_n31) ) ;
    NOR2_X1 fsm_cnt_rnd_U18 ( .A1 (fsm_en_countRound), .A2 (fsm_cnt_rnd_n6), .ZN (fsm_cnt_rnd_n26) ) ;
    INV_X1 fsm_cnt_rnd_U17 ( .A (fsm_cnt_rnd_n28), .ZN (fsm_cnt_rnd_n20) ) ;
    NAND2_X1 fsm_cnt_rnd_U16 ( .A1 (fsm_cnt_rnd_n29), .A2 (fsm_cnt_rnd_n3), .ZN (fsm_cnt_rnd_n28) ) ;
    MUX2_X1 fsm_cnt_rnd_U15 ( .S (counter[4]), .A (fsm_cnt_rnd_n19), .B (fsm_cnt_rnd_n17), .Z (fsm_cnt_rnd_n14) ) ;
    NAND2_X1 fsm_cnt_rnd_U14 ( .A1 (fsm_cnt_rnd_n15), .A2 (fsm_cnt_rnd_n13), .ZN (fsm_cnt_rnd_n17) ) ;
    NAND2_X1 fsm_cnt_rnd_U13 ( .A1 (fsm_cnt_rnd_n29), .A2 (fsm_cnt_rnd_n25), .ZN (fsm_cnt_rnd_n15) ) ;
    INV_X1 fsm_cnt_rnd_U12 ( .A (fsm_cnt_rnd_n12), .ZN (fsm_cnt_rnd_n29) ) ;
    NOR2_X1 fsm_cnt_rnd_U11 ( .A1 (fsm_cnt_rnd_n25), .A2 (fsm_cnt_rnd_n11), .ZN (fsm_cnt_rnd_n19) ) ;
    INV_X1 fsm_cnt_rnd_U10 ( .A (fsm_cnt_rnd_n10), .ZN (fsm_cnt_rnd_n1) ) ;
    MUX2_X1 fsm_cnt_rnd_U9 ( .S (fsm_cnt_rnd_n25), .A (fsm_cnt_rnd_n13), .B (fsm_cnt_rnd_n11), .Z (fsm_cnt_rnd_n10) ) ;
    NAND2_X1 fsm_cnt_rnd_U8 ( .A1 (counter[2]), .A2 (fsm_cnt_rnd_n22), .ZN (fsm_cnt_rnd_n11) ) ;
    NOR2_X1 fsm_cnt_rnd_U7 ( .A1 (fsm_cnt_rnd_n12), .A2 (fsm_cnt_rnd_n9), .ZN (fsm_cnt_rnd_n22) ) ;
    NAND2_X1 fsm_cnt_rnd_U6 ( .A1 (fsm_en_countRound), .A2 (fsm_n2), .ZN (fsm_cnt_rnd_n12) ) ;
    NAND2_X1 fsm_cnt_rnd_U5 ( .A1 (fsm_n2), .A2 (fsm_cnt_rnd_n8), .ZN (fsm_cnt_rnd_n13) ) ;
    NAND2_X1 fsm_cnt_rnd_U4 ( .A1 (fsm_en_countRound), .A2 (fsm_cnt_rnd_n7), .ZN (fsm_cnt_rnd_n8) ) ;
    NOR2_X1 fsm_cnt_rnd_U3 ( .A1 (fsm_cnt_rnd_n5), .A2 (fsm_cnt_rnd_n9), .ZN (fsm_cnt_rnd_n7) ) ;
    OR2_X1 fsm_cnt_rnd_U2 ( .A1 (fsm_cnt_rnd_n24), .A2 (fsm_cnt_rnd_n3), .ZN (fsm_cnt_rnd_n9) ) ;
    INV_X1 fsm_cnt_rnd_U1 ( .A (fsm_n2), .ZN (fsm_cnt_rnd_n6) ) ;
    INV_X1 fsm_cnt_rnd_count_reg_reg_2__U1 ( .A (counter[2]), .ZN (fsm_cnt_rnd_n5) ) ;
    INV_X1 fsm_cnt_rnd_count_reg_reg_0__U1 ( .A (counter[0]), .ZN (fsm_cnt_rnd_n3) ) ;
    INV_X1 fsm_cnt_rnd_count_reg_reg_3__U1 ( .A (counter[3]), .ZN (fsm_cnt_rnd_n25) ) ;
    INV_X1 fsm_cnt_rnd_count_reg_reg_1__U1 ( .A (fsm_cnt_rnd_n24), .ZN (counter[1]) ) ;
    NOR2_X1 fsm_cnt_ser_U12 ( .A1 (fsm_cnt_ser_n10), .A2 (fsm_cnt_ser_n9), .ZN (fsm_cnt_ser_n3) ) ;
    XNOR2_X1 fsm_cnt_ser_U11 ( .A (fsm_n3), .B (fsm_countSerial[0]), .ZN (fsm_cnt_ser_n10) ) ;
    NOR2_X1 fsm_cnt_ser_U10 ( .A1 (fsm_cnt_ser_n9), .A2 (fsm_cnt_ser_n8), .ZN (fsm_cnt_ser_n28) ) ;
    XOR2_X1 fsm_cnt_ser_U9 ( .A (fsm_countSerial[1]), .B (fsm_cnt_ser_n7), .Z (fsm_cnt_ser_n8) ) ;
    NOR2_X1 fsm_cnt_ser_U8 ( .A1 (fsm_cnt_ser_n9), .A2 (fsm_cnt_ser_n6), .ZN (fsm_cnt_ser_n26) ) ;
    XOR2_X1 fsm_cnt_ser_U7 ( .A (fsm_countSerial[3]), .B (fsm_cnt_ser_n5), .Z (fsm_cnt_ser_n6) ) ;
    NAND2_X1 fsm_cnt_ser_U6 ( .A1 (fsm_cnt_ser_n4), .A2 (fsm_countSerial[2]), .ZN (fsm_cnt_ser_n5) ) ;
    NOR2_X1 fsm_cnt_ser_U5 ( .A1 (fsm_cnt_ser_n2), .A2 (fsm_cnt_ser_n9), .ZN (fsm_cnt_ser_n1) ) ;
    INV_X1 fsm_cnt_ser_U4 ( .A (fsm_rst_countSerial), .ZN (fsm_cnt_ser_n9) ) ;
    XNOR2_X1 fsm_cnt_ser_U3 ( .A (fsm_cnt_ser_n4), .B (fsm_countSerial[2]), .ZN (fsm_cnt_ser_n2) ) ;
    NOR2_X1 fsm_cnt_ser_U2 ( .A1 (fsm_cnt_ser_n20), .A2 (fsm_cnt_ser_n7), .ZN (fsm_cnt_ser_n4) ) ;
    NAND2_X1 fsm_cnt_ser_U1 ( .A1 (fsm_n3), .A2 (fsm_countSerial[0]), .ZN (fsm_cnt_ser_n7) ) ;
    INV_X1 fsm_cnt_ser_count_reg_reg_1__U1 ( .A (fsm_countSerial[1]), .ZN (fsm_cnt_ser_n20) ) ;
    INV_X1 fsm_ps_state_reg_0__U1 ( .A (fsm_ps_state_0_), .ZN (fsm_n3) ) ;
    INV_X1 fsm_ps_state_reg_1__U1 ( .A (fsm_ps_state_1_), .ZN (fsm_n5) ) ;
    INV_X1 stateFF_state_U3 ( .A (stateFF_state_n7), .ZN (stateFF_state_n6) ) ;
    INV_X1 stateFF_state_U2 ( .A (stateFF_state_n7), .ZN (stateFF_state_n5) ) ;
    INV_X1 stateFF_state_U1 ( .A (ctrlData_0_), .ZN (stateFF_state_n7) ) ;
    mux2_masked_LMDPL stateFF_state_gff_1_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, ctrlData_0_}), .b ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, serialIn[0]}), .a ({new_AGEMA_signal_891, new_AGEMA_signal_890, stateFF_inputPar[0]}), .c ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, stateFF_state_gff_1_s_next_state[0]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_1_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, ctrlData_0_}), .b ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, serialIn[1]}), .a ({new_AGEMA_signal_897, new_AGEMA_signal_896, stateFF_inputPar[1]}), .c ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, stateFF_state_gff_1_s_next_state[1]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_1_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, ctrlData_0_}), .b ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, serialIn[2]}), .a ({new_AGEMA_signal_903, new_AGEMA_signal_902, stateFF_inputPar[2]}), .c ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, stateFF_state_gff_1_s_next_state[2]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_1_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, ctrlData_0_}), .b ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, serialIn[3]}), .a ({new_AGEMA_signal_909, new_AGEMA_signal_908, stateFF_inputPar[3]}), .c ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, stateFF_state_gff_1_s_next_state[3]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_2_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, ctrlData_0_}), .b ({new_AGEMA_signal_887, data_out_s1[0], data_out_s0[0]}), .a ({new_AGEMA_signal_915, new_AGEMA_signal_914, stateFF_inputPar[4]}), .c ({new_AGEMA_signal_1753, new_AGEMA_signal_1752, stateFF_state_gff_2_s_next_state[0]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_2_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, ctrlData_0_}), .b ({new_AGEMA_signal_981, data_out_s1[1], data_out_s0[1]}), .a ({new_AGEMA_signal_921, new_AGEMA_signal_920, stateFF_inputPar[5]}), .c ({new_AGEMA_signal_1755, new_AGEMA_signal_1754, stateFF_state_gff_2_s_next_state[1]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_2_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, ctrlData_0_}), .b ({new_AGEMA_signal_1075, data_out_s1[2], data_out_s0[2]}), .a ({new_AGEMA_signal_927, new_AGEMA_signal_926, stateFF_inputPar[6]}), .c ({new_AGEMA_signal_1757, new_AGEMA_signal_1756, stateFF_state_gff_2_s_next_state[2]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_2_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, ctrlData_0_}), .b ({new_AGEMA_signal_1169, data_out_s1[3], data_out_s0[3]}), .a ({new_AGEMA_signal_933, new_AGEMA_signal_932, stateFF_inputPar[7]}), .c ({new_AGEMA_signal_1759, new_AGEMA_signal_1758, stateFF_state_gff_2_s_next_state[3]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_3_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, stateFF_state_n6}), .b ({new_AGEMA_signal_893, data_out_s1[4], data_out_s0[4]}), .a ({new_AGEMA_signal_939, new_AGEMA_signal_938, stateFF_inputPar[8]}), .c ({new_AGEMA_signal_1793, new_AGEMA_signal_1792, stateFF_state_gff_3_s_next_state[0]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_3_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, stateFF_state_n6}), .b ({new_AGEMA_signal_987, data_out_s1[5], data_out_s0[5]}), .a ({new_AGEMA_signal_945, new_AGEMA_signal_944, stateFF_inputPar[9]}), .c ({new_AGEMA_signal_1795, new_AGEMA_signal_1794, stateFF_state_gff_3_s_next_state[1]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_3_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, stateFF_state_n6}), .b ({new_AGEMA_signal_1081, data_out_s1[6], data_out_s0[6]}), .a ({new_AGEMA_signal_951, new_AGEMA_signal_950, stateFF_inputPar[10]}), .c ({new_AGEMA_signal_1797, new_AGEMA_signal_1796, stateFF_state_gff_3_s_next_state[2]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_3_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, stateFF_state_n6}), .b ({new_AGEMA_signal_1175, data_out_s1[7], data_out_s0[7]}), .a ({new_AGEMA_signal_957, new_AGEMA_signal_956, stateFF_inputPar[11]}), .c ({new_AGEMA_signal_1799, new_AGEMA_signal_1798, stateFF_state_gff_3_s_next_state[3]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_4_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, stateFF_state_n6}), .b ({new_AGEMA_signal_899, data_out_s1[8], data_out_s0[8]}), .a ({new_AGEMA_signal_963, new_AGEMA_signal_962, stateFF_inputPar[12]}), .c ({new_AGEMA_signal_1801, new_AGEMA_signal_1800, stateFF_state_gff_4_s_next_state[0]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_4_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, stateFF_state_n6}), .b ({new_AGEMA_signal_993, data_out_s1[9], data_out_s0[9]}), .a ({new_AGEMA_signal_969, new_AGEMA_signal_968, stateFF_inputPar[13]}), .c ({new_AGEMA_signal_1803, new_AGEMA_signal_1802, stateFF_state_gff_4_s_next_state[1]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_4_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, stateFF_state_n6}), .b ({new_AGEMA_signal_1087, data_out_s1[10], data_out_s0[10]}), .a ({new_AGEMA_signal_975, new_AGEMA_signal_974, stateFF_inputPar[14]}), .c ({new_AGEMA_signal_1805, new_AGEMA_signal_1804, stateFF_state_gff_4_s_next_state[2]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_4_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, stateFF_state_n6}), .b ({new_AGEMA_signal_1181, data_out_s1[11], data_out_s0[11]}), .a ({new_AGEMA_signal_979, new_AGEMA_signal_978, stateFF_inputPar[15]}), .c ({new_AGEMA_signal_1807, new_AGEMA_signal_1806, stateFF_state_gff_4_s_next_state[3]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_5_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, stateFF_state_n6}), .b ({new_AGEMA_signal_905, data_out_s1[12], data_out_s0[12]}), .a ({new_AGEMA_signal_985, new_AGEMA_signal_984, stateFF_inputPar[16]}), .c ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, stateFF_state_gff_5_s_next_state[0]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_5_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, stateFF_state_n6}), .b ({new_AGEMA_signal_999, data_out_s1[13], data_out_s0[13]}), .a ({new_AGEMA_signal_991, new_AGEMA_signal_990, stateFF_inputPar[17]}), .c ({new_AGEMA_signal_1811, new_AGEMA_signal_1810, stateFF_state_gff_5_s_next_state[1]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_5_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, stateFF_state_n6}), .b ({new_AGEMA_signal_1093, data_out_s1[14], data_out_s0[14]}), .a ({new_AGEMA_signal_997, new_AGEMA_signal_996, stateFF_inputPar[18]}), .c ({new_AGEMA_signal_1813, new_AGEMA_signal_1812, stateFF_state_gff_5_s_next_state[2]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_5_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, stateFF_state_n6}), .b ({new_AGEMA_signal_1187, data_out_s1[15], data_out_s0[15]}), .a ({new_AGEMA_signal_1003, new_AGEMA_signal_1002, stateFF_inputPar[19]}), .c ({new_AGEMA_signal_1815, new_AGEMA_signal_1814, stateFF_state_gff_5_s_next_state[3]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_6_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, stateFF_state_n6}), .b ({new_AGEMA_signal_911, data_out_s1[16], data_out_s0[16]}), .a ({new_AGEMA_signal_1009, new_AGEMA_signal_1008, stateFF_inputPar[20]}), .c ({new_AGEMA_signal_1817, new_AGEMA_signal_1816, stateFF_state_gff_6_s_next_state[0]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_6_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, stateFF_state_n6}), .b ({new_AGEMA_signal_1005, data_out_s1[17], data_out_s0[17]}), .a ({new_AGEMA_signal_1015, new_AGEMA_signal_1014, stateFF_inputPar[21]}), .c ({new_AGEMA_signal_1819, new_AGEMA_signal_1818, stateFF_state_gff_6_s_next_state[1]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_6_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, stateFF_state_n6}), .b ({new_AGEMA_signal_1099, data_out_s1[18], data_out_s0[18]}), .a ({new_AGEMA_signal_1021, new_AGEMA_signal_1020, stateFF_inputPar[22]}), .c ({new_AGEMA_signal_1821, new_AGEMA_signal_1820, stateFF_state_gff_6_s_next_state[2]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_6_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, stateFF_state_n6}), .b ({new_AGEMA_signal_1193, data_out_s1[19], data_out_s0[19]}), .a ({new_AGEMA_signal_1027, new_AGEMA_signal_1026, stateFF_inputPar[23]}), .c ({new_AGEMA_signal_1823, new_AGEMA_signal_1822, stateFF_state_gff_6_s_next_state[3]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_7_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, stateFF_state_n6}), .b ({new_AGEMA_signal_917, data_out_s1[20], data_out_s0[20]}), .a ({new_AGEMA_signal_1033, new_AGEMA_signal_1032, stateFF_inputPar[24]}), .c ({new_AGEMA_signal_1825, new_AGEMA_signal_1824, stateFF_state_gff_7_s_next_state[0]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_7_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, stateFF_state_n6}), .b ({new_AGEMA_signal_1011, data_out_s1[21], data_out_s0[21]}), .a ({new_AGEMA_signal_1039, new_AGEMA_signal_1038, stateFF_inputPar[25]}), .c ({new_AGEMA_signal_1827, new_AGEMA_signal_1826, stateFF_state_gff_7_s_next_state[1]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_7_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, stateFF_state_n6}), .b ({new_AGEMA_signal_1105, data_out_s1[22], data_out_s0[22]}), .a ({new_AGEMA_signal_1045, new_AGEMA_signal_1044, stateFF_inputPar[26]}), .c ({new_AGEMA_signal_1829, new_AGEMA_signal_1828, stateFF_state_gff_7_s_next_state[2]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_7_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, stateFF_state_n6}), .b ({new_AGEMA_signal_1199, data_out_s1[23], data_out_s0[23]}), .a ({new_AGEMA_signal_1051, new_AGEMA_signal_1050, stateFF_inputPar[27]}), .c ({new_AGEMA_signal_1831, new_AGEMA_signal_1830, stateFF_state_gff_7_s_next_state[3]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_8_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, stateFF_state_n6}), .b ({new_AGEMA_signal_923, data_out_s1[24], data_out_s0[24]}), .a ({new_AGEMA_signal_1057, new_AGEMA_signal_1056, stateFF_inputPar[28]}), .c ({new_AGEMA_signal_1833, new_AGEMA_signal_1832, stateFF_state_gff_8_s_next_state[0]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_8_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, stateFF_state_n6}), .b ({new_AGEMA_signal_1017, data_out_s1[25], data_out_s0[25]}), .a ({new_AGEMA_signal_1063, new_AGEMA_signal_1062, stateFF_inputPar[29]}), .c ({new_AGEMA_signal_1835, new_AGEMA_signal_1834, stateFF_state_gff_8_s_next_state[1]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_8_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, stateFF_state_n6}), .b ({new_AGEMA_signal_1111, data_out_s1[26], data_out_s0[26]}), .a ({new_AGEMA_signal_1069, new_AGEMA_signal_1068, stateFF_inputPar[30]}), .c ({new_AGEMA_signal_1837, new_AGEMA_signal_1836, stateFF_state_gff_8_s_next_state[2]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_8_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, stateFF_state_n6}), .b ({new_AGEMA_signal_1205, data_out_s1[27], data_out_s0[27]}), .a ({new_AGEMA_signal_1073, new_AGEMA_signal_1072, stateFF_inputPar[31]}), .c ({new_AGEMA_signal_1839, new_AGEMA_signal_1838, stateFF_state_gff_8_s_next_state[3]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_9_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, stateFF_state_n6}), .b ({new_AGEMA_signal_929, data_out_s1[28], data_out_s0[28]}), .a ({new_AGEMA_signal_1079, new_AGEMA_signal_1078, stateFF_inputPar[32]}), .c ({new_AGEMA_signal_1841, new_AGEMA_signal_1840, stateFF_state_gff_9_s_next_state[0]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_9_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, stateFF_state_n6}), .b ({new_AGEMA_signal_1023, data_out_s1[29], data_out_s0[29]}), .a ({new_AGEMA_signal_1085, new_AGEMA_signal_1084, stateFF_inputPar[33]}), .c ({new_AGEMA_signal_1843, new_AGEMA_signal_1842, stateFF_state_gff_9_s_next_state[1]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_9_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, stateFF_state_n6}), .b ({new_AGEMA_signal_1117, data_out_s1[30], data_out_s0[30]}), .a ({new_AGEMA_signal_1091, new_AGEMA_signal_1090, stateFF_inputPar[34]}), .c ({new_AGEMA_signal_1845, new_AGEMA_signal_1844, stateFF_state_gff_9_s_next_state[2]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_9_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, stateFF_state_n6}), .b ({new_AGEMA_signal_1211, data_out_s1[31], data_out_s0[31]}), .a ({new_AGEMA_signal_1097, new_AGEMA_signal_1096, stateFF_inputPar[35]}), .c ({new_AGEMA_signal_1847, new_AGEMA_signal_1846, stateFF_state_gff_9_s_next_state[3]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_10_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, stateFF_state_n5}), .b ({new_AGEMA_signal_935, data_out_s1[32], data_out_s0[32]}), .a ({new_AGEMA_signal_1103, new_AGEMA_signal_1102, stateFF_inputPar[36]}), .c ({new_AGEMA_signal_1851, new_AGEMA_signal_1850, stateFF_state_gff_10_s_next_state[0]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_10_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, stateFF_state_n5}), .b ({new_AGEMA_signal_1029, data_out_s1[33], data_out_s0[33]}), .a ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, stateFF_inputPar[37]}), .c ({new_AGEMA_signal_1853, new_AGEMA_signal_1852, stateFF_state_gff_10_s_next_state[1]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_10_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, stateFF_state_n5}), .b ({new_AGEMA_signal_1123, data_out_s1[34], data_out_s0[34]}), .a ({new_AGEMA_signal_1115, new_AGEMA_signal_1114, stateFF_inputPar[38]}), .c ({new_AGEMA_signal_1855, new_AGEMA_signal_1854, stateFF_state_gff_10_s_next_state[2]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_10_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, stateFF_state_n5}), .b ({new_AGEMA_signal_1217, data_out_s1[35], data_out_s0[35]}), .a ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, stateFF_inputPar[39]}), .c ({new_AGEMA_signal_1857, new_AGEMA_signal_1856, stateFF_state_gff_10_s_next_state[3]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_11_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, stateFF_state_n5}), .b ({new_AGEMA_signal_941, data_out_s1[36], data_out_s0[36]}), .a ({new_AGEMA_signal_1127, new_AGEMA_signal_1126, stateFF_inputPar[40]}), .c ({new_AGEMA_signal_1859, new_AGEMA_signal_1858, stateFF_state_gff_11_s_next_state[0]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_11_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, stateFF_state_n5}), .b ({new_AGEMA_signal_1035, data_out_s1[37], data_out_s0[37]}), .a ({new_AGEMA_signal_1133, new_AGEMA_signal_1132, stateFF_inputPar[41]}), .c ({new_AGEMA_signal_1861, new_AGEMA_signal_1860, stateFF_state_gff_11_s_next_state[1]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_11_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, stateFF_state_n5}), .b ({new_AGEMA_signal_1129, data_out_s1[38], data_out_s0[38]}), .a ({new_AGEMA_signal_1139, new_AGEMA_signal_1138, stateFF_inputPar[42]}), .c ({new_AGEMA_signal_1863, new_AGEMA_signal_1862, stateFF_state_gff_11_s_next_state[2]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_11_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, stateFF_state_n5}), .b ({new_AGEMA_signal_1223, data_out_s1[39], data_out_s0[39]}), .a ({new_AGEMA_signal_1145, new_AGEMA_signal_1144, stateFF_inputPar[43]}), .c ({new_AGEMA_signal_1865, new_AGEMA_signal_1864, stateFF_state_gff_11_s_next_state[3]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_12_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, stateFF_state_n5}), .b ({new_AGEMA_signal_947, data_out_s1[40], data_out_s0[40]}), .a ({new_AGEMA_signal_1151, new_AGEMA_signal_1150, stateFF_inputPar[44]}), .c ({new_AGEMA_signal_1867, new_AGEMA_signal_1866, stateFF_state_gff_12_s_next_state[0]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_12_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, stateFF_state_n5}), .b ({new_AGEMA_signal_1041, data_out_s1[41], data_out_s0[41]}), .a ({new_AGEMA_signal_1157, new_AGEMA_signal_1156, stateFF_inputPar[45]}), .c ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, stateFF_state_gff_12_s_next_state[1]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_12_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, stateFF_state_n5}), .b ({new_AGEMA_signal_1135, data_out_s1[42], data_out_s0[42]}), .a ({new_AGEMA_signal_1163, new_AGEMA_signal_1162, stateFF_inputPar[46]}), .c ({new_AGEMA_signal_1871, new_AGEMA_signal_1870, stateFF_state_gff_12_s_next_state[2]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_12_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, stateFF_state_n5}), .b ({new_AGEMA_signal_1229, data_out_s1[43], data_out_s0[43]}), .a ({new_AGEMA_signal_1167, new_AGEMA_signal_1166, stateFF_inputPar[47]}), .c ({new_AGEMA_signal_1873, new_AGEMA_signal_1872, stateFF_state_gff_12_s_next_state[3]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_13_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, stateFF_state_n5}), .b ({new_AGEMA_signal_953, data_out_s1[44], data_out_s0[44]}), .a ({new_AGEMA_signal_1173, new_AGEMA_signal_1172, stateFF_inputPar[48]}), .c ({new_AGEMA_signal_1875, new_AGEMA_signal_1874, stateFF_state_gff_13_s_next_state[0]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_13_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, stateFF_state_n5}), .b ({new_AGEMA_signal_1047, data_out_s1[45], data_out_s0[45]}), .a ({new_AGEMA_signal_1179, new_AGEMA_signal_1178, stateFF_inputPar[49]}), .c ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, stateFF_state_gff_13_s_next_state[1]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_13_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, stateFF_state_n5}), .b ({new_AGEMA_signal_1141, data_out_s1[46], data_out_s0[46]}), .a ({new_AGEMA_signal_1185, new_AGEMA_signal_1184, stateFF_inputPar[50]}), .c ({new_AGEMA_signal_1879, new_AGEMA_signal_1878, stateFF_state_gff_13_s_next_state[2]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_13_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, stateFF_state_n5}), .b ({new_AGEMA_signal_1235, data_out_s1[47], data_out_s0[47]}), .a ({new_AGEMA_signal_1191, new_AGEMA_signal_1190, stateFF_inputPar[51]}), .c ({new_AGEMA_signal_1881, new_AGEMA_signal_1880, stateFF_state_gff_13_s_next_state[3]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_14_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, stateFF_state_n5}), .b ({new_AGEMA_signal_959, data_out_s1[48], data_out_s0[48]}), .a ({new_AGEMA_signal_1197, new_AGEMA_signal_1196, stateFF_inputPar[52]}), .c ({new_AGEMA_signal_1883, new_AGEMA_signal_1882, stateFF_state_gff_14_s_next_state[0]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_14_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, stateFF_state_n5}), .b ({new_AGEMA_signal_1053, data_out_s1[49], data_out_s0[49]}), .a ({new_AGEMA_signal_1203, new_AGEMA_signal_1202, stateFF_inputPar[53]}), .c ({new_AGEMA_signal_1885, new_AGEMA_signal_1884, stateFF_state_gff_14_s_next_state[1]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_14_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, stateFF_state_n5}), .b ({new_AGEMA_signal_1147, data_out_s1[50], data_out_s0[50]}), .a ({new_AGEMA_signal_1209, new_AGEMA_signal_1208, stateFF_inputPar[54]}), .c ({new_AGEMA_signal_1887, new_AGEMA_signal_1886, stateFF_state_gff_14_s_next_state[2]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_14_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, stateFF_state_n5}), .b ({new_AGEMA_signal_1241, data_out_s1[51], data_out_s0[51]}), .a ({new_AGEMA_signal_1215, new_AGEMA_signal_1214, stateFF_inputPar[55]}), .c ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, stateFF_state_gff_14_s_next_state[3]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_15_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, stateFF_state_n5}), .b ({new_AGEMA_signal_965, data_out_s1[52], data_out_s0[52]}), .a ({new_AGEMA_signal_1221, new_AGEMA_signal_1220, stateFF_inputPar[56]}), .c ({new_AGEMA_signal_1891, new_AGEMA_signal_1890, stateFF_state_gff_15_s_next_state[0]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_15_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, stateFF_state_n5}), .b ({new_AGEMA_signal_1059, data_out_s1[53], data_out_s0[53]}), .a ({new_AGEMA_signal_1227, new_AGEMA_signal_1226, stateFF_inputPar[57]}), .c ({new_AGEMA_signal_1893, new_AGEMA_signal_1892, stateFF_state_gff_15_s_next_state[1]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_15_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, stateFF_state_n5}), .b ({new_AGEMA_signal_1153, data_out_s1[54], data_out_s0[54]}), .a ({new_AGEMA_signal_1233, new_AGEMA_signal_1232, stateFF_inputPar[58]}), .c ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, stateFF_state_gff_15_s_next_state[2]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_15_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, stateFF_state_n5}), .b ({new_AGEMA_signal_1247, data_out_s1[55], data_out_s0[55]}), .a ({new_AGEMA_signal_1239, new_AGEMA_signal_1238, stateFF_inputPar[59]}), .c ({new_AGEMA_signal_1897, new_AGEMA_signal_1896, stateFF_state_gff_15_s_next_state[3]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_16_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, stateFF_state_n5}), .b ({new_AGEMA_signal_971, data_out_s1[56], data_out_s0[56]}), .a ({new_AGEMA_signal_1245, new_AGEMA_signal_1244, stateFF_inputPar[60]}), .c ({new_AGEMA_signal_1899, new_AGEMA_signal_1898, stateFF_state_gff_16_s_next_state[0]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_16_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, stateFF_state_n5}), .b ({new_AGEMA_signal_1065, data_out_s1[57], data_out_s0[57]}), .a ({new_AGEMA_signal_1251, new_AGEMA_signal_1250, stateFF_inputPar[61]}), .c ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, stateFF_state_gff_16_s_next_state[1]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_16_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, stateFF_state_n5}), .b ({new_AGEMA_signal_1159, data_out_s1[58], data_out_s0[58]}), .a ({new_AGEMA_signal_1257, new_AGEMA_signal_1256, stateFF_inputPar[62]}), .c ({new_AGEMA_signal_1903, new_AGEMA_signal_1902, stateFF_state_gff_16_s_next_state[2]}) ) ;
    mux2_masked_LMDPL stateFF_state_gff_16_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, stateFF_state_n5}), .b ({new_AGEMA_signal_1253, data_out_s1[59], data_out_s0[59]}), .a ({new_AGEMA_signal_1261, new_AGEMA_signal_1260, stateFF_inputPar[63]}), .c ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, stateFF_state_gff_16_s_next_state[3]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_0_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_887, data_out_s1[0], data_out_s0[0]}), .a ({new_AGEMA_signal_889, new_AGEMA_signal_888, data_in_s0[0]}), .c ({new_AGEMA_signal_891, new_AGEMA_signal_890, stateFF_inputPar[0]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_1_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_893, data_out_s1[4], data_out_s0[4]}), .a ({new_AGEMA_signal_895, new_AGEMA_signal_894, data_in_s0[1]}), .c ({new_AGEMA_signal_897, new_AGEMA_signal_896, stateFF_inputPar[1]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_2_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_899, data_out_s1[8], data_out_s0[8]}), .a ({new_AGEMA_signal_901, new_AGEMA_signal_900, data_in_s0[2]}), .c ({new_AGEMA_signal_903, new_AGEMA_signal_902, stateFF_inputPar[2]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_3_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_905, data_out_s1[12], data_out_s0[12]}), .a ({new_AGEMA_signal_907, new_AGEMA_signal_906, data_in_s0[3]}), .c ({new_AGEMA_signal_909, new_AGEMA_signal_908, stateFF_inputPar[3]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_4_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_911, data_out_s1[16], data_out_s0[16]}), .a ({new_AGEMA_signal_913, new_AGEMA_signal_912, data_in_s0[4]}), .c ({new_AGEMA_signal_915, new_AGEMA_signal_914, stateFF_inputPar[4]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_5_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_917, data_out_s1[20], data_out_s0[20]}), .a ({new_AGEMA_signal_919, new_AGEMA_signal_918, data_in_s0[5]}), .c ({new_AGEMA_signal_921, new_AGEMA_signal_920, stateFF_inputPar[5]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_6_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_923, data_out_s1[24], data_out_s0[24]}), .a ({new_AGEMA_signal_925, new_AGEMA_signal_924, data_in_s0[6]}), .c ({new_AGEMA_signal_927, new_AGEMA_signal_926, stateFF_inputPar[6]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_7_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_929, data_out_s1[28], data_out_s0[28]}), .a ({new_AGEMA_signal_931, new_AGEMA_signal_930, data_in_s0[7]}), .c ({new_AGEMA_signal_933, new_AGEMA_signal_932, stateFF_inputPar[7]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_8_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_935, data_out_s1[32], data_out_s0[32]}), .a ({new_AGEMA_signal_937, new_AGEMA_signal_936, data_in_s0[8]}), .c ({new_AGEMA_signal_939, new_AGEMA_signal_938, stateFF_inputPar[8]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_9_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_941, data_out_s1[36], data_out_s0[36]}), .a ({new_AGEMA_signal_943, new_AGEMA_signal_942, data_in_s0[9]}), .c ({new_AGEMA_signal_945, new_AGEMA_signal_944, stateFF_inputPar[9]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_10_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_947, data_out_s1[40], data_out_s0[40]}), .a ({new_AGEMA_signal_949, new_AGEMA_signal_948, data_in_s0[10]}), .c ({new_AGEMA_signal_951, new_AGEMA_signal_950, stateFF_inputPar[10]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_11_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_953, data_out_s1[44], data_out_s0[44]}), .a ({new_AGEMA_signal_955, new_AGEMA_signal_954, data_in_s0[11]}), .c ({new_AGEMA_signal_957, new_AGEMA_signal_956, stateFF_inputPar[11]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_12_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_959, data_out_s1[48], data_out_s0[48]}), .a ({new_AGEMA_signal_961, new_AGEMA_signal_960, data_in_s0[12]}), .c ({new_AGEMA_signal_963, new_AGEMA_signal_962, stateFF_inputPar[12]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_13_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_965, data_out_s1[52], data_out_s0[52]}), .a ({new_AGEMA_signal_967, new_AGEMA_signal_966, data_in_s0[13]}), .c ({new_AGEMA_signal_969, new_AGEMA_signal_968, stateFF_inputPar[13]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_14_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_971, data_out_s1[56], data_out_s0[56]}), .a ({new_AGEMA_signal_973, new_AGEMA_signal_972, data_in_s0[14]}), .c ({new_AGEMA_signal_975, new_AGEMA_signal_974, stateFF_inputPar[14]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_15_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_863, data_out_s1[60], data_out_s0[60]}), .a ({new_AGEMA_signal_977, new_AGEMA_signal_976, data_in_s0[15]}), .c ({new_AGEMA_signal_979, new_AGEMA_signal_978, stateFF_inputPar[15]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_16_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_981, data_out_s1[1], data_out_s0[1]}), .a ({new_AGEMA_signal_983, new_AGEMA_signal_982, data_in_s0[16]}), .c ({new_AGEMA_signal_985, new_AGEMA_signal_984, stateFF_inputPar[16]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_17_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_987, data_out_s1[5], data_out_s0[5]}), .a ({new_AGEMA_signal_989, new_AGEMA_signal_988, data_in_s0[17]}), .c ({new_AGEMA_signal_991, new_AGEMA_signal_990, stateFF_inputPar[17]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_18_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_993, data_out_s1[9], data_out_s0[9]}), .a ({new_AGEMA_signal_995, new_AGEMA_signal_994, data_in_s0[18]}), .c ({new_AGEMA_signal_997, new_AGEMA_signal_996, stateFF_inputPar[18]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_19_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_999, data_out_s1[13], data_out_s0[13]}), .a ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, data_in_s0[19]}), .c ({new_AGEMA_signal_1003, new_AGEMA_signal_1002, stateFF_inputPar[19]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_20_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1005, data_out_s1[17], data_out_s0[17]}), .a ({new_AGEMA_signal_1007, new_AGEMA_signal_1006, data_in_s0[20]}), .c ({new_AGEMA_signal_1009, new_AGEMA_signal_1008, stateFF_inputPar[20]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_21_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1011, data_out_s1[21], data_out_s0[21]}), .a ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, data_in_s0[21]}), .c ({new_AGEMA_signal_1015, new_AGEMA_signal_1014, stateFF_inputPar[21]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_22_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1017, data_out_s1[25], data_out_s0[25]}), .a ({new_AGEMA_signal_1019, new_AGEMA_signal_1018, data_in_s0[22]}), .c ({new_AGEMA_signal_1021, new_AGEMA_signal_1020, stateFF_inputPar[22]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_23_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1023, data_out_s1[29], data_out_s0[29]}), .a ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, data_in_s0[23]}), .c ({new_AGEMA_signal_1027, new_AGEMA_signal_1026, stateFF_inputPar[23]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_24_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1029, data_out_s1[33], data_out_s0[33]}), .a ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, data_in_s0[24]}), .c ({new_AGEMA_signal_1033, new_AGEMA_signal_1032, stateFF_inputPar[24]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_25_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1035, data_out_s1[37], data_out_s0[37]}), .a ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, data_in_s0[25]}), .c ({new_AGEMA_signal_1039, new_AGEMA_signal_1038, stateFF_inputPar[25]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_26_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1041, data_out_s1[41], data_out_s0[41]}), .a ({new_AGEMA_signal_1043, new_AGEMA_signal_1042, data_in_s0[26]}), .c ({new_AGEMA_signal_1045, new_AGEMA_signal_1044, stateFF_inputPar[26]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_27_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1047, data_out_s1[45], data_out_s0[45]}), .a ({new_AGEMA_signal_1049, new_AGEMA_signal_1048, data_in_s0[27]}), .c ({new_AGEMA_signal_1051, new_AGEMA_signal_1050, stateFF_inputPar[27]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_28_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1053, data_out_s1[49], data_out_s0[49]}), .a ({new_AGEMA_signal_1055, new_AGEMA_signal_1054, data_in_s0[28]}), .c ({new_AGEMA_signal_1057, new_AGEMA_signal_1056, stateFF_inputPar[28]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_29_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1059, data_out_s1[53], data_out_s0[53]}), .a ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, data_in_s0[29]}), .c ({new_AGEMA_signal_1063, new_AGEMA_signal_1062, stateFF_inputPar[29]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_30_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1065, data_out_s1[57], data_out_s0[57]}), .a ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, data_in_s0[30]}), .c ({new_AGEMA_signal_1069, new_AGEMA_signal_1068, stateFF_inputPar[30]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_31_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_869, data_out_s1[61], data_out_s0[61]}), .a ({new_AGEMA_signal_1071, new_AGEMA_signal_1070, data_in_s0[31]}), .c ({new_AGEMA_signal_1073, new_AGEMA_signal_1072, stateFF_inputPar[31]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_32_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1075, data_out_s1[2], data_out_s0[2]}), .a ({new_AGEMA_signal_1077, new_AGEMA_signal_1076, data_in_s0[32]}), .c ({new_AGEMA_signal_1079, new_AGEMA_signal_1078, stateFF_inputPar[32]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_33_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1081, data_out_s1[6], data_out_s0[6]}), .a ({new_AGEMA_signal_1083, new_AGEMA_signal_1082, data_in_s0[33]}), .c ({new_AGEMA_signal_1085, new_AGEMA_signal_1084, stateFF_inputPar[33]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_34_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1087, data_out_s1[10], data_out_s0[10]}), .a ({new_AGEMA_signal_1089, new_AGEMA_signal_1088, data_in_s0[34]}), .c ({new_AGEMA_signal_1091, new_AGEMA_signal_1090, stateFF_inputPar[34]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_35_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1093, data_out_s1[14], data_out_s0[14]}), .a ({new_AGEMA_signal_1095, new_AGEMA_signal_1094, data_in_s0[35]}), .c ({new_AGEMA_signal_1097, new_AGEMA_signal_1096, stateFF_inputPar[35]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_36_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1099, data_out_s1[18], data_out_s0[18]}), .a ({new_AGEMA_signal_1101, new_AGEMA_signal_1100, data_in_s0[36]}), .c ({new_AGEMA_signal_1103, new_AGEMA_signal_1102, stateFF_inputPar[36]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_37_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1105, data_out_s1[22], data_out_s0[22]}), .a ({new_AGEMA_signal_1107, new_AGEMA_signal_1106, data_in_s0[37]}), .c ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, stateFF_inputPar[37]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_38_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1111, data_out_s1[26], data_out_s0[26]}), .a ({new_AGEMA_signal_1113, new_AGEMA_signal_1112, data_in_s0[38]}), .c ({new_AGEMA_signal_1115, new_AGEMA_signal_1114, stateFF_inputPar[38]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_39_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1117, data_out_s1[30], data_out_s0[30]}), .a ({new_AGEMA_signal_1119, new_AGEMA_signal_1118, data_in_s0[39]}), .c ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, stateFF_inputPar[39]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_40_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1123, data_out_s1[34], data_out_s0[34]}), .a ({new_AGEMA_signal_1125, new_AGEMA_signal_1124, data_in_s0[40]}), .c ({new_AGEMA_signal_1127, new_AGEMA_signal_1126, stateFF_inputPar[40]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_41_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1129, data_out_s1[38], data_out_s0[38]}), .a ({new_AGEMA_signal_1131, new_AGEMA_signal_1130, data_in_s0[41]}), .c ({new_AGEMA_signal_1133, new_AGEMA_signal_1132, stateFF_inputPar[41]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_42_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1135, data_out_s1[42], data_out_s0[42]}), .a ({new_AGEMA_signal_1137, new_AGEMA_signal_1136, data_in_s0[42]}), .c ({new_AGEMA_signal_1139, new_AGEMA_signal_1138, stateFF_inputPar[42]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_43_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1141, data_out_s1[46], data_out_s0[46]}), .a ({new_AGEMA_signal_1143, new_AGEMA_signal_1142, data_in_s0[43]}), .c ({new_AGEMA_signal_1145, new_AGEMA_signal_1144, stateFF_inputPar[43]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_44_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1147, data_out_s1[50], data_out_s0[50]}), .a ({new_AGEMA_signal_1149, new_AGEMA_signal_1148, data_in_s0[44]}), .c ({new_AGEMA_signal_1151, new_AGEMA_signal_1150, stateFF_inputPar[44]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_45_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1153, data_out_s1[54], data_out_s0[54]}), .a ({new_AGEMA_signal_1155, new_AGEMA_signal_1154, data_in_s0[45]}), .c ({new_AGEMA_signal_1157, new_AGEMA_signal_1156, stateFF_inputPar[45]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_46_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1159, data_out_s1[58], data_out_s0[58]}), .a ({new_AGEMA_signal_1161, new_AGEMA_signal_1160, data_in_s0[46]}), .c ({new_AGEMA_signal_1163, new_AGEMA_signal_1162, stateFF_inputPar[46]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_47_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_875, data_out_s1[62], data_out_s0[62]}), .a ({new_AGEMA_signal_1165, new_AGEMA_signal_1164, data_in_s0[47]}), .c ({new_AGEMA_signal_1167, new_AGEMA_signal_1166, stateFF_inputPar[47]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_48_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1169, data_out_s1[3], data_out_s0[3]}), .a ({new_AGEMA_signal_1171, new_AGEMA_signal_1170, data_in_s0[48]}), .c ({new_AGEMA_signal_1173, new_AGEMA_signal_1172, stateFF_inputPar[48]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_49_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1175, data_out_s1[7], data_out_s0[7]}), .a ({new_AGEMA_signal_1177, new_AGEMA_signal_1176, data_in_s0[49]}), .c ({new_AGEMA_signal_1179, new_AGEMA_signal_1178, stateFF_inputPar[49]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_50_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1181, data_out_s1[11], data_out_s0[11]}), .a ({new_AGEMA_signal_1183, new_AGEMA_signal_1182, data_in_s0[50]}), .c ({new_AGEMA_signal_1185, new_AGEMA_signal_1184, stateFF_inputPar[50]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_51_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1187, data_out_s1[15], data_out_s0[15]}), .a ({new_AGEMA_signal_1189, new_AGEMA_signal_1188, data_in_s0[51]}), .c ({new_AGEMA_signal_1191, new_AGEMA_signal_1190, stateFF_inputPar[51]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_52_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1193, data_out_s1[19], data_out_s0[19]}), .a ({new_AGEMA_signal_1195, new_AGEMA_signal_1194, data_in_s0[52]}), .c ({new_AGEMA_signal_1197, new_AGEMA_signal_1196, stateFF_inputPar[52]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_53_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1199, data_out_s1[23], data_out_s0[23]}), .a ({new_AGEMA_signal_1201, new_AGEMA_signal_1200, data_in_s0[53]}), .c ({new_AGEMA_signal_1203, new_AGEMA_signal_1202, stateFF_inputPar[53]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_54_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1205, data_out_s1[27], data_out_s0[27]}), .a ({new_AGEMA_signal_1207, new_AGEMA_signal_1206, data_in_s0[54]}), .c ({new_AGEMA_signal_1209, new_AGEMA_signal_1208, stateFF_inputPar[54]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_55_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1211, data_out_s1[31], data_out_s0[31]}), .a ({new_AGEMA_signal_1213, new_AGEMA_signal_1212, data_in_s0[55]}), .c ({new_AGEMA_signal_1215, new_AGEMA_signal_1214, stateFF_inputPar[55]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_56_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1217, data_out_s1[35], data_out_s0[35]}), .a ({new_AGEMA_signal_1219, new_AGEMA_signal_1218, data_in_s0[56]}), .c ({new_AGEMA_signal_1221, new_AGEMA_signal_1220, stateFF_inputPar[56]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_57_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1223, data_out_s1[39], data_out_s0[39]}), .a ({new_AGEMA_signal_1225, new_AGEMA_signal_1224, data_in_s0[57]}), .c ({new_AGEMA_signal_1227, new_AGEMA_signal_1226, stateFF_inputPar[57]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_58_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1229, data_out_s1[43], data_out_s0[43]}), .a ({new_AGEMA_signal_1231, new_AGEMA_signal_1230, data_in_s0[58]}), .c ({new_AGEMA_signal_1233, new_AGEMA_signal_1232, stateFF_inputPar[58]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_59_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1235, data_out_s1[47], data_out_s0[47]}), .a ({new_AGEMA_signal_1237, new_AGEMA_signal_1236, data_in_s0[59]}), .c ({new_AGEMA_signal_1239, new_AGEMA_signal_1238, stateFF_inputPar[59]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_60_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1241, data_out_s1[51], data_out_s0[51]}), .a ({new_AGEMA_signal_1243, new_AGEMA_signal_1242, data_in_s0[60]}), .c ({new_AGEMA_signal_1245, new_AGEMA_signal_1244, stateFF_inputPar[60]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_61_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1247, data_out_s1[55], data_out_s0[55]}), .a ({new_AGEMA_signal_1249, new_AGEMA_signal_1248, data_in_s0[61]}), .c ({new_AGEMA_signal_1251, new_AGEMA_signal_1250, stateFF_inputPar[61]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_62_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1253, data_out_s1[59], data_out_s0[59]}), .a ({new_AGEMA_signal_1255, new_AGEMA_signal_1254, data_in_s0[62]}), .c ({new_AGEMA_signal_1257, new_AGEMA_signal_1256, stateFF_inputPar[62]}) ) ;
    mux2_masked_LMDPL stateFF_MUX_inputPar_mux_inst_63_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_881, data_out_s1[63], data_out_s0[63]}), .a ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, data_in_s0[63]}), .c ({new_AGEMA_signal_1261, new_AGEMA_signal_1260, stateFF_inputPar[63]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) keyFF_U5 ( .a ({LMDPL_pre1, 1'b0, counter[4]}), .b ({new_AGEMA_signal_1263, new_AGEMA_signal_1262, keyFF_outputPar[22]}), .c ({new_AGEMA_signal_1265, new_AGEMA_signal_1264, keyFF_counterAdd[4]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) keyFF_U4 ( .a ({LMDPL_pre1, 1'b0, counter[3]}), .b ({new_AGEMA_signal_1267, new_AGEMA_signal_1266, keyFF_outputPar[21]}), .c ({new_AGEMA_signal_1269, new_AGEMA_signal_1268, keyFF_counterAdd[3]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) keyFF_U3 ( .a ({LMDPL_pre1, 1'b0, counter[2]}), .b ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, keyFF_outputPar[20]}), .c ({new_AGEMA_signal_1273, new_AGEMA_signal_1272, keyFF_counterAdd[2]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) keyFF_U2 ( .a ({LMDPL_pre1, 1'b0, counter[1]}), .b ({new_AGEMA_signal_1699, new_AGEMA_signal_1698, keyFF_outputPar[19]}), .c ({new_AGEMA_signal_1701, new_AGEMA_signal_1700, keyFF_counterAdd[1]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) keyFF_U1 ( .a ({LMDPL_pre1, 1'b0, counter[0]}), .b ({new_AGEMA_signal_1275, new_AGEMA_signal_1274, keyFF_outputPar[18]}), .c ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, keyFF_counterAdd[0]}) ) ;
    INV_X1 keyFF_keystate_U3 ( .A (keyFF_keystate_n8), .ZN (keyFF_keystate_n6) ) ;
    INV_X1 keyFF_keystate_U2 ( .A (keyFF_keystate_n8), .ZN (keyFF_keystate_n7) ) ;
    INV_X1 keyFF_keystate_U1 ( .A (ctrlData_0_), .ZN (keyFF_keystate_n8) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_1_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_861, new_AGEMA_signal_860, roundkey[0]}), .a ({new_AGEMA_signal_1283, new_AGEMA_signal_1282, keyFF_inputPar[0]}), .c ({new_AGEMA_signal_1909, new_AGEMA_signal_1908, keyFF_keystate_gff_1_s_next_state[0]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_1_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_867, new_AGEMA_signal_866, roundkey[1]}), .a ({new_AGEMA_signal_1289, new_AGEMA_signal_1288, keyFF_inputPar[1]}), .c ({new_AGEMA_signal_1911, new_AGEMA_signal_1910, keyFF_keystate_gff_1_s_next_state[1]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_1_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_873, new_AGEMA_signal_872, roundkey[2]}), .a ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, keyFF_inputPar[2]}), .c ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, keyFF_keystate_gff_1_s_next_state[2]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_1_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_879, new_AGEMA_signal_878, roundkey[3]}), .a ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, keyFF_inputPar[3]}), .c ({new_AGEMA_signal_1915, new_AGEMA_signal_1914, keyFF_keystate_gff_1_s_next_state[3]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_2_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_1727, new_AGEMA_signal_1726, keyRegKS[1]}), .a ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, keyFF_inputPar[4]}), .c ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, keyFF_keystate_gff_2_s_next_state[0]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_2_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_1731, new_AGEMA_signal_1730, keyRegKS[2]}), .a ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, keyFF_inputPar[5]}), .c ({new_AGEMA_signal_1919, new_AGEMA_signal_1918, keyFF_keystate_gff_2_s_next_state[1]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_2_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_1735, new_AGEMA_signal_1734, keyRegKS[3]}), .a ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, keyFF_inputPar[6]}), .c ({new_AGEMA_signal_1921, new_AGEMA_signal_1920, keyFF_keystate_gff_2_s_next_state[2]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_2_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_1279, new_AGEMA_signal_1278, keyFF_outputPar[3]}), .a ({new_AGEMA_signal_1325, new_AGEMA_signal_1324, keyFF_inputPar[7]}), .c ({new_AGEMA_signal_1923, new_AGEMA_signal_1922, keyFF_keystate_gff_2_s_next_state[3]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_3_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1285, new_AGEMA_signal_1284, keyFF_outputPar[4]}), .a ({new_AGEMA_signal_1331, new_AGEMA_signal_1330, keyFF_inputPar[8]}), .c ({new_AGEMA_signal_1927, new_AGEMA_signal_1926, keyFF_keystate_gff_3_s_next_state[0]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_3_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1291, new_AGEMA_signal_1290, keyFF_outputPar[5]}), .a ({new_AGEMA_signal_1337, new_AGEMA_signal_1336, keyFF_inputPar[9]}), .c ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, keyFF_keystate_gff_3_s_next_state[1]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_3_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1297, new_AGEMA_signal_1296, keyFF_outputPar[6]}), .a ({new_AGEMA_signal_1343, new_AGEMA_signal_1342, keyFF_inputPar[10]}), .c ({new_AGEMA_signal_1931, new_AGEMA_signal_1930, keyFF_keystate_gff_3_s_next_state[2]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_3_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1303, new_AGEMA_signal_1302, keyFF_outputPar[7]}), .a ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, keyFF_inputPar[11]}), .c ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, keyFF_keystate_gff_3_s_next_state[3]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_4_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1309, new_AGEMA_signal_1308, keyFF_outputPar[8]}), .a ({new_AGEMA_signal_1355, new_AGEMA_signal_1354, keyFF_inputPar[12]}), .c ({new_AGEMA_signal_1935, new_AGEMA_signal_1934, keyFF_keystate_gff_4_s_next_state[0]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_4_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1315, new_AGEMA_signal_1314, keyFF_outputPar[9]}), .a ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, keyFF_inputPar[13]}), .c ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, keyFF_keystate_gff_4_s_next_state[1]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_4_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1321, new_AGEMA_signal_1320, keyFF_outputPar[10]}), .a ({new_AGEMA_signal_1367, new_AGEMA_signal_1366, keyFF_inputPar[14]}), .c ({new_AGEMA_signal_1939, new_AGEMA_signal_1938, keyFF_keystate_gff_4_s_next_state[2]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_4_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1327, new_AGEMA_signal_1326, keyFF_outputPar[11]}), .a ({new_AGEMA_signal_1705, new_AGEMA_signal_1704, keyFF_inputPar[15]}), .c ({new_AGEMA_signal_1941, new_AGEMA_signal_1940, keyFF_keystate_gff_4_s_next_state[3]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_5_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, ctrlData_0_}), .b ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, keyFF_outputPar[12]}), .a ({new_AGEMA_signal_1721, new_AGEMA_signal_1720, keyFF_inputPar[16]}), .c ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, keyFF_keystate_gff_5_s_next_state[0]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_5_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, ctrlData_0_}), .b ({new_AGEMA_signal_1339, new_AGEMA_signal_1338, keyFF_outputPar[13]}), .a ({new_AGEMA_signal_1709, new_AGEMA_signal_1708, keyFF_inputPar[17]}), .c ({new_AGEMA_signal_1763, new_AGEMA_signal_1762, keyFF_keystate_gff_5_s_next_state[1]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_5_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, ctrlData_0_}), .b ({new_AGEMA_signal_1345, new_AGEMA_signal_1344, keyFF_outputPar[14]}), .a ({new_AGEMA_signal_1713, new_AGEMA_signal_1712, keyFF_inputPar[18]}), .c ({new_AGEMA_signal_1765, new_AGEMA_signal_1764, keyFF_keystate_gff_5_s_next_state[2]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_5_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, ctrlData_0_}), .b ({new_AGEMA_signal_1351, new_AGEMA_signal_1350, keyFF_outputPar[15]}), .a ({new_AGEMA_signal_1717, new_AGEMA_signal_1716, keyFF_inputPar[19]}), .c ({new_AGEMA_signal_1767, new_AGEMA_signal_1766, keyFF_keystate_gff_5_s_next_state[3]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_6_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, ctrlData_0_}), .b ({new_AGEMA_signal_1357, new_AGEMA_signal_1356, keyFF_outputPar[16]}), .a ({new_AGEMA_signal_1373, new_AGEMA_signal_1372, keyFF_inputPar[20]}), .c ({new_AGEMA_signal_1769, new_AGEMA_signal_1768, keyFF_keystate_gff_6_s_next_state[0]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_6_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, ctrlData_0_}), .b ({new_AGEMA_signal_1363, new_AGEMA_signal_1362, keyFF_outputPar[17]}), .a ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, keyFF_inputPar[21]}), .c ({new_AGEMA_signal_1771, new_AGEMA_signal_1770, keyFF_keystate_gff_6_s_next_state[1]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_6_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, ctrlData_0_}), .b ({new_AGEMA_signal_1275, new_AGEMA_signal_1274, keyFF_outputPar[18]}), .a ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, keyFF_inputPar[22]}), .c ({new_AGEMA_signal_1773, new_AGEMA_signal_1772, keyFF_keystate_gff_6_s_next_state[2]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_6_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, ctrlData_0_}), .b ({new_AGEMA_signal_1699, new_AGEMA_signal_1698, keyFF_outputPar[19]}), .a ({new_AGEMA_signal_1391, new_AGEMA_signal_1390, keyFF_inputPar[23]}), .c ({new_AGEMA_signal_1775, new_AGEMA_signal_1774, keyFF_keystate_gff_6_s_next_state[3]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_7_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, keyFF_outputPar[20]}), .a ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, keyFF_inputPar[24]}), .c ({new_AGEMA_signal_1943, new_AGEMA_signal_1942, keyFF_keystate_gff_7_s_next_state[0]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_7_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_1267, new_AGEMA_signal_1266, keyFF_outputPar[21]}), .a ({new_AGEMA_signal_1403, new_AGEMA_signal_1402, keyFF_inputPar[25]}), .c ({new_AGEMA_signal_1945, new_AGEMA_signal_1944, keyFF_keystate_gff_7_s_next_state[1]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_7_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_1263, new_AGEMA_signal_1262, keyFF_outputPar[22]}), .a ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, keyFF_inputPar[26]}), .c ({new_AGEMA_signal_1947, new_AGEMA_signal_1946, keyFF_keystate_gff_7_s_next_state[2]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_7_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_1369, new_AGEMA_signal_1368, keyFF_outputPar[23]}), .a ({new_AGEMA_signal_1415, new_AGEMA_signal_1414, keyFF_inputPar[27]}), .c ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, keyFF_keystate_gff_7_s_next_state[3]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_8_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_1375, new_AGEMA_signal_1374, keyFF_outputPar[24]}), .a ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, keyFF_inputPar[28]}), .c ({new_AGEMA_signal_1951, new_AGEMA_signal_1950, keyFF_keystate_gff_8_s_next_state[0]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_8_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_1381, new_AGEMA_signal_1380, keyFF_outputPar[25]}), .a ({new_AGEMA_signal_1427, new_AGEMA_signal_1426, keyFF_inputPar[29]}), .c ({new_AGEMA_signal_1953, new_AGEMA_signal_1952, keyFF_keystate_gff_8_s_next_state[1]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_8_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_1387, new_AGEMA_signal_1386, keyFF_outputPar[26]}), .a ({new_AGEMA_signal_1433, new_AGEMA_signal_1432, keyFF_inputPar[30]}), .c ({new_AGEMA_signal_1955, new_AGEMA_signal_1954, keyFF_keystate_gff_8_s_next_state[2]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_8_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_1393, new_AGEMA_signal_1392, keyFF_outputPar[27]}), .a ({new_AGEMA_signal_1439, new_AGEMA_signal_1438, keyFF_inputPar[31]}), .c ({new_AGEMA_signal_1957, new_AGEMA_signal_1956, keyFF_keystate_gff_8_s_next_state[3]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_9_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_1399, new_AGEMA_signal_1398, keyFF_outputPar[28]}), .a ({new_AGEMA_signal_1445, new_AGEMA_signal_1444, keyFF_inputPar[32]}), .c ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, keyFF_keystate_gff_9_s_next_state[0]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_9_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_1405, new_AGEMA_signal_1404, keyFF_outputPar[29]}), .a ({new_AGEMA_signal_1451, new_AGEMA_signal_1450, keyFF_inputPar[33]}), .c ({new_AGEMA_signal_1961, new_AGEMA_signal_1960, keyFF_keystate_gff_9_s_next_state[1]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_9_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_1411, new_AGEMA_signal_1410, keyFF_outputPar[30]}), .a ({new_AGEMA_signal_1457, new_AGEMA_signal_1456, keyFF_inputPar[34]}), .c ({new_AGEMA_signal_1963, new_AGEMA_signal_1962, keyFF_keystate_gff_9_s_next_state[2]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_9_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_1417, new_AGEMA_signal_1416, keyFF_outputPar[31]}), .a ({new_AGEMA_signal_1463, new_AGEMA_signal_1462, keyFF_inputPar[35]}), .c ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, keyFF_keystate_gff_9_s_next_state[3]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_10_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_1423, new_AGEMA_signal_1422, keyFF_outputPar[32]}), .a ({new_AGEMA_signal_1469, new_AGEMA_signal_1468, keyFF_inputPar[36]}), .c ({new_AGEMA_signal_1967, new_AGEMA_signal_1966, keyFF_keystate_gff_10_s_next_state[0]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_10_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_1429, new_AGEMA_signal_1428, keyFF_outputPar[33]}), .a ({new_AGEMA_signal_1475, new_AGEMA_signal_1474, keyFF_inputPar[37]}), .c ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, keyFF_keystate_gff_10_s_next_state[1]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_10_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_1435, new_AGEMA_signal_1434, keyFF_outputPar[34]}), .a ({new_AGEMA_signal_1481, new_AGEMA_signal_1480, keyFF_inputPar[38]}), .c ({new_AGEMA_signal_1971, new_AGEMA_signal_1970, keyFF_keystate_gff_10_s_next_state[2]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_10_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_1441, new_AGEMA_signal_1440, keyFF_outputPar[35]}), .a ({new_AGEMA_signal_1487, new_AGEMA_signal_1486, keyFF_inputPar[39]}), .c ({new_AGEMA_signal_1973, new_AGEMA_signal_1972, keyFF_keystate_gff_10_s_next_state[3]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_11_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_1447, new_AGEMA_signal_1446, keyFF_outputPar[36]}), .a ({new_AGEMA_signal_1493, new_AGEMA_signal_1492, keyFF_inputPar[40]}), .c ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, keyFF_keystate_gff_11_s_next_state[0]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_11_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_1453, new_AGEMA_signal_1452, keyFF_outputPar[37]}), .a ({new_AGEMA_signal_1499, new_AGEMA_signal_1498, keyFF_inputPar[41]}), .c ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, keyFF_keystate_gff_11_s_next_state[1]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_11_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_1459, new_AGEMA_signal_1458, keyFF_outputPar[38]}), .a ({new_AGEMA_signal_1505, new_AGEMA_signal_1504, keyFF_inputPar[42]}), .c ({new_AGEMA_signal_1979, new_AGEMA_signal_1978, keyFF_keystate_gff_11_s_next_state[2]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_11_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, keyFF_outputPar[39]}), .a ({new_AGEMA_signal_1511, new_AGEMA_signal_1510, keyFF_inputPar[43]}), .c ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, keyFF_keystate_gff_11_s_next_state[3]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_12_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_1471, new_AGEMA_signal_1470, keyFF_outputPar[40]}), .a ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, keyFF_inputPar[44]}), .c ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, keyFF_keystate_gff_12_s_next_state[0]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_12_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_1477, new_AGEMA_signal_1476, keyFF_outputPar[41]}), .a ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, keyFF_inputPar[45]}), .c ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, keyFF_keystate_gff_12_s_next_state[1]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_12_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_1483, new_AGEMA_signal_1482, keyFF_outputPar[42]}), .a ({new_AGEMA_signal_1529, new_AGEMA_signal_1528, keyFF_inputPar[46]}), .c ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, keyFF_keystate_gff_12_s_next_state[2]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_12_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_1489, new_AGEMA_signal_1488, keyFF_outputPar[43]}), .a ({new_AGEMA_signal_1535, new_AGEMA_signal_1534, keyFF_inputPar[47]}), .c ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, keyFF_keystate_gff_12_s_next_state[3]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_13_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_1495, new_AGEMA_signal_1494, keyFF_outputPar[44]}), .a ({new_AGEMA_signal_1541, new_AGEMA_signal_1540, keyFF_inputPar[48]}), .c ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, keyFF_keystate_gff_13_s_next_state[0]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_13_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_1501, new_AGEMA_signal_1500, keyFF_outputPar[45]}), .a ({new_AGEMA_signal_1547, new_AGEMA_signal_1546, keyFF_inputPar[49]}), .c ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, keyFF_keystate_gff_13_s_next_state[1]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_13_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_1507, new_AGEMA_signal_1506, keyFF_outputPar[46]}), .a ({new_AGEMA_signal_1553, new_AGEMA_signal_1552, keyFF_inputPar[50]}), .c ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, keyFF_keystate_gff_13_s_next_state[2]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_13_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, keyFF_keystate_n7}), .b ({new_AGEMA_signal_1513, new_AGEMA_signal_1512, keyFF_outputPar[47]}), .a ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, keyFF_inputPar[51]}), .c ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, keyFF_keystate_gff_13_s_next_state[3]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_14_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1519, new_AGEMA_signal_1518, keyFF_outputPar[48]}), .a ({new_AGEMA_signal_1565, new_AGEMA_signal_1564, keyFF_inputPar[52]}), .c ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, keyFF_keystate_gff_14_s_next_state[0]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_14_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1525, new_AGEMA_signal_1524, keyFF_outputPar[49]}), .a ({new_AGEMA_signal_1571, new_AGEMA_signal_1570, keyFF_inputPar[53]}), .c ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, keyFF_keystate_gff_14_s_next_state[1]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_14_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1531, new_AGEMA_signal_1530, keyFF_outputPar[50]}), .a ({new_AGEMA_signal_1577, new_AGEMA_signal_1576, keyFF_inputPar[54]}), .c ({new_AGEMA_signal_2003, new_AGEMA_signal_2002, keyFF_keystate_gff_14_s_next_state[2]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_14_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1537, new_AGEMA_signal_1536, keyFF_outputPar[51]}), .a ({new_AGEMA_signal_1583, new_AGEMA_signal_1582, keyFF_inputPar[55]}), .c ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, keyFF_keystate_gff_14_s_next_state[3]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_15_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1543, new_AGEMA_signal_1542, keyFF_outputPar[52]}), .a ({new_AGEMA_signal_1589, new_AGEMA_signal_1588, keyFF_inputPar[56]}), .c ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, keyFF_keystate_gff_15_s_next_state[0]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_15_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1549, new_AGEMA_signal_1548, keyFF_outputPar[53]}), .a ({new_AGEMA_signal_1595, new_AGEMA_signal_1594, keyFF_inputPar[57]}), .c ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, keyFF_keystate_gff_15_s_next_state[1]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_15_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1555, new_AGEMA_signal_1554, keyFF_outputPar[54]}), .a ({new_AGEMA_signal_1601, new_AGEMA_signal_1600, keyFF_inputPar[58]}), .c ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, keyFF_keystate_gff_15_s_next_state[2]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_15_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1561, new_AGEMA_signal_1560, keyFF_outputPar[55]}), .a ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, keyFF_inputPar[59]}), .c ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, keyFF_keystate_gff_15_s_next_state[3]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_16_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1567, new_AGEMA_signal_1566, keyFF_outputPar[56]}), .a ({new_AGEMA_signal_1613, new_AGEMA_signal_1612, keyFF_inputPar[60]}), .c ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, keyFF_keystate_gff_16_s_next_state[0]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_16_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1573, new_AGEMA_signal_1572, keyFF_outputPar[57]}), .a ({new_AGEMA_signal_1619, new_AGEMA_signal_1618, keyFF_inputPar[61]}), .c ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, keyFF_keystate_gff_16_s_next_state[1]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_16_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1579, new_AGEMA_signal_1578, keyFF_outputPar[58]}), .a ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, keyFF_inputPar[62]}), .c ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, keyFF_keystate_gff_16_s_next_state[2]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_16_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1585, new_AGEMA_signal_1584, keyFF_outputPar[59]}), .a ({new_AGEMA_signal_1631, new_AGEMA_signal_1630, keyFF_inputPar[63]}), .c ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, keyFF_keystate_gff_16_s_next_state[3]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_17_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1591, new_AGEMA_signal_1590, keyFF_outputPar[60]}), .a ({new_AGEMA_signal_1637, new_AGEMA_signal_1636, keyFF_inputPar[64]}), .c ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, keyFF_keystate_gff_17_s_next_state[0]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_17_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1597, new_AGEMA_signal_1596, keyFF_outputPar[61]}), .a ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, keyFF_inputPar[65]}), .c ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, keyFF_keystate_gff_17_s_next_state[1]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_17_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1603, new_AGEMA_signal_1602, keyFF_outputPar[62]}), .a ({new_AGEMA_signal_1649, new_AGEMA_signal_1648, keyFF_inputPar[66]}), .c ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, keyFF_keystate_gff_17_s_next_state[2]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_17_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1609, new_AGEMA_signal_1608, keyFF_outputPar[63]}), .a ({new_AGEMA_signal_1655, new_AGEMA_signal_1654, keyFF_inputPar[67]}), .c ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, keyFF_keystate_gff_17_s_next_state[3]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_18_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1615, new_AGEMA_signal_1614, keyFF_outputPar[64]}), .a ({new_AGEMA_signal_1661, new_AGEMA_signal_1660, keyFF_inputPar[68]}), .c ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, keyFF_keystate_gff_18_s_next_state[0]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_18_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1621, new_AGEMA_signal_1620, keyFF_outputPar[65]}), .a ({new_AGEMA_signal_1667, new_AGEMA_signal_1666, keyFF_inputPar[69]}), .c ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, keyFF_keystate_gff_18_s_next_state[1]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_18_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1627, new_AGEMA_signal_1626, keyFF_outputPar[66]}), .a ({new_AGEMA_signal_1673, new_AGEMA_signal_1672, keyFF_inputPar[70]}), .c ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, keyFF_keystate_gff_18_s_next_state[2]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_18_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1633, new_AGEMA_signal_1632, keyFF_outputPar[67]}), .a ({new_AGEMA_signal_1679, new_AGEMA_signal_1678, keyFF_inputPar[71]}), .c ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, keyFF_keystate_gff_18_s_next_state[3]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_19_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1639, new_AGEMA_signal_1638, keyFF_outputPar[68]}), .a ({new_AGEMA_signal_1685, new_AGEMA_signal_1684, keyFF_inputPar[72]}), .c ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, keyFF_keystate_gff_19_s_next_state[0]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_19_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1645, new_AGEMA_signal_1644, keyFF_outputPar[69]}), .a ({new_AGEMA_signal_1689, new_AGEMA_signal_1688, keyFF_inputPar[73]}), .c ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, keyFF_keystate_gff_19_s_next_state[1]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_19_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1651, new_AGEMA_signal_1650, keyFF_outputPar[70]}), .a ({new_AGEMA_signal_1693, new_AGEMA_signal_1692, keyFF_inputPar[74]}), .c ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, keyFF_keystate_gff_19_s_next_state[2]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_19_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1657, new_AGEMA_signal_1656, keyFF_outputPar[71]}), .a ({new_AGEMA_signal_1697, new_AGEMA_signal_1696, keyFF_inputPar[75]}), .c ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, keyFF_keystate_gff_19_s_next_state[3]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_20_MUX_inst1_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1663, new_AGEMA_signal_1662, keyFF_outputPar[72]}), .a ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, keyFF_inputPar[76]}), .c ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, keyFF_keystate_gff_20_s_next_state[0]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_20_MUX_inst1_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1669, new_AGEMA_signal_1668, keyFF_outputPar[73]}), .a ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, keyFF_inputPar[77]}), .c ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, keyFF_keystate_gff_20_s_next_state[1]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_20_MUX_inst1_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1675, new_AGEMA_signal_1674, keyFF_outputPar[74]}), .a ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, keyFF_inputPar[78]}), .c ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, keyFF_keystate_gff_20_s_next_state[2]}) ) ;
    mux2_masked_LMDPL keyFF_keystate_gff_20_MUX_inst1_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, keyFF_keystate_n6}), .b ({new_AGEMA_signal_1681, new_AGEMA_signal_1680, keyFF_outputPar[75]}), .a ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, keyFF_inputPar[79]}), .c ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, keyFF_keystate_gff_20_s_next_state[3]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_0_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1279, new_AGEMA_signal_1278, keyFF_outputPar[3]}), .a ({new_AGEMA_signal_1281, new_AGEMA_signal_1280, key_s0[0]}), .c ({new_AGEMA_signal_1283, new_AGEMA_signal_1282, keyFF_inputPar[0]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_1_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1285, new_AGEMA_signal_1284, keyFF_outputPar[4]}), .a ({new_AGEMA_signal_1287, new_AGEMA_signal_1286, key_s0[1]}), .c ({new_AGEMA_signal_1289, new_AGEMA_signal_1288, keyFF_inputPar[1]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_2_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1291, new_AGEMA_signal_1290, keyFF_outputPar[5]}), .a ({new_AGEMA_signal_1293, new_AGEMA_signal_1292, key_s0[2]}), .c ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, keyFF_inputPar[2]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_3_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1297, new_AGEMA_signal_1296, keyFF_outputPar[6]}), .a ({new_AGEMA_signal_1299, new_AGEMA_signal_1298, key_s0[3]}), .c ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, keyFF_inputPar[3]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_4_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1303, new_AGEMA_signal_1302, keyFF_outputPar[7]}), .a ({new_AGEMA_signal_1305, new_AGEMA_signal_1304, key_s0[4]}), .c ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, keyFF_inputPar[4]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_5_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1309, new_AGEMA_signal_1308, keyFF_outputPar[8]}), .a ({new_AGEMA_signal_1311, new_AGEMA_signal_1310, key_s0[5]}), .c ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, keyFF_inputPar[5]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_6_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1315, new_AGEMA_signal_1314, keyFF_outputPar[9]}), .a ({new_AGEMA_signal_1317, new_AGEMA_signal_1316, key_s0[6]}), .c ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, keyFF_inputPar[6]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_7_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1321, new_AGEMA_signal_1320, keyFF_outputPar[10]}), .a ({new_AGEMA_signal_1323, new_AGEMA_signal_1322, key_s0[7]}), .c ({new_AGEMA_signal_1325, new_AGEMA_signal_1324, keyFF_inputPar[7]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_8_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1327, new_AGEMA_signal_1326, keyFF_outputPar[11]}), .a ({new_AGEMA_signal_1329, new_AGEMA_signal_1328, key_s0[8]}), .c ({new_AGEMA_signal_1331, new_AGEMA_signal_1330, keyFF_inputPar[8]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_9_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, keyFF_outputPar[12]}), .a ({new_AGEMA_signal_1335, new_AGEMA_signal_1334, key_s0[9]}), .c ({new_AGEMA_signal_1337, new_AGEMA_signal_1336, keyFF_inputPar[9]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_10_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1339, new_AGEMA_signal_1338, keyFF_outputPar[13]}), .a ({new_AGEMA_signal_1341, new_AGEMA_signal_1340, key_s0[10]}), .c ({new_AGEMA_signal_1343, new_AGEMA_signal_1342, keyFF_inputPar[10]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_11_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1345, new_AGEMA_signal_1344, keyFF_outputPar[14]}), .a ({new_AGEMA_signal_1347, new_AGEMA_signal_1346, key_s0[11]}), .c ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, keyFF_inputPar[11]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_12_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1351, new_AGEMA_signal_1350, keyFF_outputPar[15]}), .a ({new_AGEMA_signal_1353, new_AGEMA_signal_1352, key_s0[12]}), .c ({new_AGEMA_signal_1355, new_AGEMA_signal_1354, keyFF_inputPar[12]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_13_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1357, new_AGEMA_signal_1356, keyFF_outputPar[16]}), .a ({new_AGEMA_signal_1359, new_AGEMA_signal_1358, key_s0[13]}), .c ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, keyFF_inputPar[13]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_14_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1363, new_AGEMA_signal_1362, keyFF_outputPar[17]}), .a ({new_AGEMA_signal_1365, new_AGEMA_signal_1364, key_s0[14]}), .c ({new_AGEMA_signal_1367, new_AGEMA_signal_1366, keyFF_inputPar[14]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_15_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, keyFF_counterAdd[0]}), .a ({new_AGEMA_signal_1703, new_AGEMA_signal_1702, key_s0[15]}), .c ({new_AGEMA_signal_1705, new_AGEMA_signal_1704, keyFF_inputPar[15]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_16_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1701, new_AGEMA_signal_1700, keyFF_counterAdd[1]}), .a ({new_AGEMA_signal_1719, new_AGEMA_signal_1718, key_s0[16]}), .c ({new_AGEMA_signal_1721, new_AGEMA_signal_1720, keyFF_inputPar[16]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_17_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1273, new_AGEMA_signal_1272, keyFF_counterAdd[2]}), .a ({new_AGEMA_signal_1707, new_AGEMA_signal_1706, key_s0[17]}), .c ({new_AGEMA_signal_1709, new_AGEMA_signal_1708, keyFF_inputPar[17]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_18_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1269, new_AGEMA_signal_1268, keyFF_counterAdd[3]}), .a ({new_AGEMA_signal_1711, new_AGEMA_signal_1710, key_s0[18]}), .c ({new_AGEMA_signal_1713, new_AGEMA_signal_1712, keyFF_inputPar[18]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_19_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1265, new_AGEMA_signal_1264, keyFF_counterAdd[4]}), .a ({new_AGEMA_signal_1715, new_AGEMA_signal_1714, key_s0[19]}), .c ({new_AGEMA_signal_1717, new_AGEMA_signal_1716, keyFF_inputPar[19]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_20_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1369, new_AGEMA_signal_1368, keyFF_outputPar[23]}), .a ({new_AGEMA_signal_1371, new_AGEMA_signal_1370, key_s0[20]}), .c ({new_AGEMA_signal_1373, new_AGEMA_signal_1372, keyFF_inputPar[20]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_21_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1375, new_AGEMA_signal_1374, keyFF_outputPar[24]}), .a ({new_AGEMA_signal_1377, new_AGEMA_signal_1376, key_s0[21]}), .c ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, keyFF_inputPar[21]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_22_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1381, new_AGEMA_signal_1380, keyFF_outputPar[25]}), .a ({new_AGEMA_signal_1383, new_AGEMA_signal_1382, key_s0[22]}), .c ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, keyFF_inputPar[22]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_23_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1387, new_AGEMA_signal_1386, keyFF_outputPar[26]}), .a ({new_AGEMA_signal_1389, new_AGEMA_signal_1388, key_s0[23]}), .c ({new_AGEMA_signal_1391, new_AGEMA_signal_1390, keyFF_inputPar[23]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_24_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1393, new_AGEMA_signal_1392, keyFF_outputPar[27]}), .a ({new_AGEMA_signal_1395, new_AGEMA_signal_1394, key_s0[24]}), .c ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, keyFF_inputPar[24]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_25_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1399, new_AGEMA_signal_1398, keyFF_outputPar[28]}), .a ({new_AGEMA_signal_1401, new_AGEMA_signal_1400, key_s0[25]}), .c ({new_AGEMA_signal_1403, new_AGEMA_signal_1402, keyFF_inputPar[25]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_26_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1405, new_AGEMA_signal_1404, keyFF_outputPar[29]}), .a ({new_AGEMA_signal_1407, new_AGEMA_signal_1406, key_s0[26]}), .c ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, keyFF_inputPar[26]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_27_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1411, new_AGEMA_signal_1410, keyFF_outputPar[30]}), .a ({new_AGEMA_signal_1413, new_AGEMA_signal_1412, key_s0[27]}), .c ({new_AGEMA_signal_1415, new_AGEMA_signal_1414, keyFF_inputPar[27]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_28_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1417, new_AGEMA_signal_1416, keyFF_outputPar[31]}), .a ({new_AGEMA_signal_1419, new_AGEMA_signal_1418, key_s0[28]}), .c ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, keyFF_inputPar[28]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_29_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1423, new_AGEMA_signal_1422, keyFF_outputPar[32]}), .a ({new_AGEMA_signal_1425, new_AGEMA_signal_1424, key_s0[29]}), .c ({new_AGEMA_signal_1427, new_AGEMA_signal_1426, keyFF_inputPar[29]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_30_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1429, new_AGEMA_signal_1428, keyFF_outputPar[33]}), .a ({new_AGEMA_signal_1431, new_AGEMA_signal_1430, key_s0[30]}), .c ({new_AGEMA_signal_1433, new_AGEMA_signal_1432, keyFF_inputPar[30]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_31_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1435, new_AGEMA_signal_1434, keyFF_outputPar[34]}), .a ({new_AGEMA_signal_1437, new_AGEMA_signal_1436, key_s0[31]}), .c ({new_AGEMA_signal_1439, new_AGEMA_signal_1438, keyFF_inputPar[31]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_32_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1441, new_AGEMA_signal_1440, keyFF_outputPar[35]}), .a ({new_AGEMA_signal_1443, new_AGEMA_signal_1442, key_s0[32]}), .c ({new_AGEMA_signal_1445, new_AGEMA_signal_1444, keyFF_inputPar[32]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_33_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1447, new_AGEMA_signal_1446, keyFF_outputPar[36]}), .a ({new_AGEMA_signal_1449, new_AGEMA_signal_1448, key_s0[33]}), .c ({new_AGEMA_signal_1451, new_AGEMA_signal_1450, keyFF_inputPar[33]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_34_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1453, new_AGEMA_signal_1452, keyFF_outputPar[37]}), .a ({new_AGEMA_signal_1455, new_AGEMA_signal_1454, key_s0[34]}), .c ({new_AGEMA_signal_1457, new_AGEMA_signal_1456, keyFF_inputPar[34]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_35_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1459, new_AGEMA_signal_1458, keyFF_outputPar[38]}), .a ({new_AGEMA_signal_1461, new_AGEMA_signal_1460, key_s0[35]}), .c ({new_AGEMA_signal_1463, new_AGEMA_signal_1462, keyFF_inputPar[35]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_36_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, keyFF_outputPar[39]}), .a ({new_AGEMA_signal_1467, new_AGEMA_signal_1466, key_s0[36]}), .c ({new_AGEMA_signal_1469, new_AGEMA_signal_1468, keyFF_inputPar[36]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_37_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1471, new_AGEMA_signal_1470, keyFF_outputPar[40]}), .a ({new_AGEMA_signal_1473, new_AGEMA_signal_1472, key_s0[37]}), .c ({new_AGEMA_signal_1475, new_AGEMA_signal_1474, keyFF_inputPar[37]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_38_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1477, new_AGEMA_signal_1476, keyFF_outputPar[41]}), .a ({new_AGEMA_signal_1479, new_AGEMA_signal_1478, key_s0[38]}), .c ({new_AGEMA_signal_1481, new_AGEMA_signal_1480, keyFF_inputPar[38]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_39_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1483, new_AGEMA_signal_1482, keyFF_outputPar[42]}), .a ({new_AGEMA_signal_1485, new_AGEMA_signal_1484, key_s0[39]}), .c ({new_AGEMA_signal_1487, new_AGEMA_signal_1486, keyFF_inputPar[39]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_40_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1489, new_AGEMA_signal_1488, keyFF_outputPar[43]}), .a ({new_AGEMA_signal_1491, new_AGEMA_signal_1490, key_s0[40]}), .c ({new_AGEMA_signal_1493, new_AGEMA_signal_1492, keyFF_inputPar[40]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_41_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1495, new_AGEMA_signal_1494, keyFF_outputPar[44]}), .a ({new_AGEMA_signal_1497, new_AGEMA_signal_1496, key_s0[41]}), .c ({new_AGEMA_signal_1499, new_AGEMA_signal_1498, keyFF_inputPar[41]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_42_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1501, new_AGEMA_signal_1500, keyFF_outputPar[45]}), .a ({new_AGEMA_signal_1503, new_AGEMA_signal_1502, key_s0[42]}), .c ({new_AGEMA_signal_1505, new_AGEMA_signal_1504, keyFF_inputPar[42]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_43_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1507, new_AGEMA_signal_1506, keyFF_outputPar[46]}), .a ({new_AGEMA_signal_1509, new_AGEMA_signal_1508, key_s0[43]}), .c ({new_AGEMA_signal_1511, new_AGEMA_signal_1510, keyFF_inputPar[43]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_44_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1513, new_AGEMA_signal_1512, keyFF_outputPar[47]}), .a ({new_AGEMA_signal_1515, new_AGEMA_signal_1514, key_s0[44]}), .c ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, keyFF_inputPar[44]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_45_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1519, new_AGEMA_signal_1518, keyFF_outputPar[48]}), .a ({new_AGEMA_signal_1521, new_AGEMA_signal_1520, key_s0[45]}), .c ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, keyFF_inputPar[45]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_46_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1525, new_AGEMA_signal_1524, keyFF_outputPar[49]}), .a ({new_AGEMA_signal_1527, new_AGEMA_signal_1526, key_s0[46]}), .c ({new_AGEMA_signal_1529, new_AGEMA_signal_1528, keyFF_inputPar[46]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_47_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1531, new_AGEMA_signal_1530, keyFF_outputPar[50]}), .a ({new_AGEMA_signal_1533, new_AGEMA_signal_1532, key_s0[47]}), .c ({new_AGEMA_signal_1535, new_AGEMA_signal_1534, keyFF_inputPar[47]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_48_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1537, new_AGEMA_signal_1536, keyFF_outputPar[51]}), .a ({new_AGEMA_signal_1539, new_AGEMA_signal_1538, key_s0[48]}), .c ({new_AGEMA_signal_1541, new_AGEMA_signal_1540, keyFF_inputPar[48]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_49_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1543, new_AGEMA_signal_1542, keyFF_outputPar[52]}), .a ({new_AGEMA_signal_1545, new_AGEMA_signal_1544, key_s0[49]}), .c ({new_AGEMA_signal_1547, new_AGEMA_signal_1546, keyFF_inputPar[49]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_50_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1549, new_AGEMA_signal_1548, keyFF_outputPar[53]}), .a ({new_AGEMA_signal_1551, new_AGEMA_signal_1550, key_s0[50]}), .c ({new_AGEMA_signal_1553, new_AGEMA_signal_1552, keyFF_inputPar[50]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_51_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1555, new_AGEMA_signal_1554, keyFF_outputPar[54]}), .a ({new_AGEMA_signal_1557, new_AGEMA_signal_1556, key_s0[51]}), .c ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, keyFF_inputPar[51]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_52_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1561, new_AGEMA_signal_1560, keyFF_outputPar[55]}), .a ({new_AGEMA_signal_1563, new_AGEMA_signal_1562, key_s0[52]}), .c ({new_AGEMA_signal_1565, new_AGEMA_signal_1564, keyFF_inputPar[52]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_53_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1567, new_AGEMA_signal_1566, keyFF_outputPar[56]}), .a ({new_AGEMA_signal_1569, new_AGEMA_signal_1568, key_s0[53]}), .c ({new_AGEMA_signal_1571, new_AGEMA_signal_1570, keyFF_inputPar[53]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_54_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1573, new_AGEMA_signal_1572, keyFF_outputPar[57]}), .a ({new_AGEMA_signal_1575, new_AGEMA_signal_1574, key_s0[54]}), .c ({new_AGEMA_signal_1577, new_AGEMA_signal_1576, keyFF_inputPar[54]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_55_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1579, new_AGEMA_signal_1578, keyFF_outputPar[58]}), .a ({new_AGEMA_signal_1581, new_AGEMA_signal_1580, key_s0[55]}), .c ({new_AGEMA_signal_1583, new_AGEMA_signal_1582, keyFF_inputPar[55]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_56_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1585, new_AGEMA_signal_1584, keyFF_outputPar[59]}), .a ({new_AGEMA_signal_1587, new_AGEMA_signal_1586, key_s0[56]}), .c ({new_AGEMA_signal_1589, new_AGEMA_signal_1588, keyFF_inputPar[56]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_57_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1591, new_AGEMA_signal_1590, keyFF_outputPar[60]}), .a ({new_AGEMA_signal_1593, new_AGEMA_signal_1592, key_s0[57]}), .c ({new_AGEMA_signal_1595, new_AGEMA_signal_1594, keyFF_inputPar[57]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_58_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1597, new_AGEMA_signal_1596, keyFF_outputPar[61]}), .a ({new_AGEMA_signal_1599, new_AGEMA_signal_1598, key_s0[58]}), .c ({new_AGEMA_signal_1601, new_AGEMA_signal_1600, keyFF_inputPar[58]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_59_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1603, new_AGEMA_signal_1602, keyFF_outputPar[62]}), .a ({new_AGEMA_signal_1605, new_AGEMA_signal_1604, key_s0[59]}), .c ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, keyFF_inputPar[59]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_60_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1609, new_AGEMA_signal_1608, keyFF_outputPar[63]}), .a ({new_AGEMA_signal_1611, new_AGEMA_signal_1610, key_s0[60]}), .c ({new_AGEMA_signal_1613, new_AGEMA_signal_1612, keyFF_inputPar[60]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_61_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1615, new_AGEMA_signal_1614, keyFF_outputPar[64]}), .a ({new_AGEMA_signal_1617, new_AGEMA_signal_1616, key_s0[61]}), .c ({new_AGEMA_signal_1619, new_AGEMA_signal_1618, keyFF_inputPar[61]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_62_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1621, new_AGEMA_signal_1620, keyFF_outputPar[65]}), .a ({new_AGEMA_signal_1623, new_AGEMA_signal_1622, key_s0[62]}), .c ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, keyFF_inputPar[62]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_63_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1627, new_AGEMA_signal_1626, keyFF_outputPar[66]}), .a ({new_AGEMA_signal_1629, new_AGEMA_signal_1628, key_s0[63]}), .c ({new_AGEMA_signal_1631, new_AGEMA_signal_1630, keyFF_inputPar[63]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_64_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1633, new_AGEMA_signal_1632, keyFF_outputPar[67]}), .a ({new_AGEMA_signal_1635, new_AGEMA_signal_1634, key_s0[64]}), .c ({new_AGEMA_signal_1637, new_AGEMA_signal_1636, keyFF_inputPar[64]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_65_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1639, new_AGEMA_signal_1638, keyFF_outputPar[68]}), .a ({new_AGEMA_signal_1641, new_AGEMA_signal_1640, key_s0[65]}), .c ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, keyFF_inputPar[65]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_66_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1645, new_AGEMA_signal_1644, keyFF_outputPar[69]}), .a ({new_AGEMA_signal_1647, new_AGEMA_signal_1646, key_s0[66]}), .c ({new_AGEMA_signal_1649, new_AGEMA_signal_1648, keyFF_inputPar[66]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_67_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1651, new_AGEMA_signal_1650, keyFF_outputPar[70]}), .a ({new_AGEMA_signal_1653, new_AGEMA_signal_1652, key_s0[67]}), .c ({new_AGEMA_signal_1655, new_AGEMA_signal_1654, keyFF_inputPar[67]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_68_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1657, new_AGEMA_signal_1656, keyFF_outputPar[71]}), .a ({new_AGEMA_signal_1659, new_AGEMA_signal_1658, key_s0[68]}), .c ({new_AGEMA_signal_1661, new_AGEMA_signal_1660, keyFF_inputPar[68]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_69_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1663, new_AGEMA_signal_1662, keyFF_outputPar[72]}), .a ({new_AGEMA_signal_1665, new_AGEMA_signal_1664, key_s0[69]}), .c ({new_AGEMA_signal_1667, new_AGEMA_signal_1666, keyFF_inputPar[69]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_70_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1669, new_AGEMA_signal_1668, keyFF_outputPar[73]}), .a ({new_AGEMA_signal_1671, new_AGEMA_signal_1670, key_s0[70]}), .c ({new_AGEMA_signal_1673, new_AGEMA_signal_1672, keyFF_inputPar[70]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_71_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1675, new_AGEMA_signal_1674, keyFF_outputPar[74]}), .a ({new_AGEMA_signal_1677, new_AGEMA_signal_1676, key_s0[71]}), .c ({new_AGEMA_signal_1679, new_AGEMA_signal_1678, keyFF_inputPar[71]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_72_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1681, new_AGEMA_signal_1680, keyFF_outputPar[75]}), .a ({new_AGEMA_signal_1683, new_AGEMA_signal_1682, key_s0[72]}), .c ({new_AGEMA_signal_1685, new_AGEMA_signal_1684, keyFF_inputPar[72]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_73_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_861, new_AGEMA_signal_860, roundkey[0]}), .a ({new_AGEMA_signal_1687, new_AGEMA_signal_1686, key_s0[73]}), .c ({new_AGEMA_signal_1689, new_AGEMA_signal_1688, keyFF_inputPar[73]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_74_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_867, new_AGEMA_signal_866, roundkey[1]}), .a ({new_AGEMA_signal_1691, new_AGEMA_signal_1690, key_s0[74]}), .c ({new_AGEMA_signal_1693, new_AGEMA_signal_1692, keyFF_inputPar[74]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_75_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_873, new_AGEMA_signal_872, roundkey[2]}), .a ({new_AGEMA_signal_1695, new_AGEMA_signal_1694, key_s0[75]}), .c ({new_AGEMA_signal_1697, new_AGEMA_signal_1696, keyFF_inputPar[75]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_76_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_1789, new_AGEMA_signal_1788, sboxOut[0]}), .a ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, key_s0[76]}), .c ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, keyFF_inputPar[76]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_77_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, sboxOut[1]}), .a ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, key_s0[77]}), .c ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, keyFF_inputPar[77]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_78_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, sboxOut[2]}), .a ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, key_s0[78]}), .c ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, keyFF_inputPar[78]}) ) ;
    mux2_masked_LMDPL keyFF_MUX_inputPar_mux_inst_79_U1 ( .s ({new_AGEMA_signal_885, new_AGEMA_signal_884, reset}), .b ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, sboxOut[3]}), .a ({new_AGEMA_signal_2099, new_AGEMA_signal_2098, key_s0[79]}), .c ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, keyFF_inputPar[79]}) ) ;
    not_LMDPL sboxInst_U3 ( .x ({new_AGEMA_signal_1743, new_AGEMA_signal_1742, sboxInst_L0}), .y ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, sboxInst_n1}) ) ;
    not_LMDPL sboxInst_U2 ( .x ({new_AGEMA_signal_1737, new_AGEMA_signal_1736, sboxIn[3]}), .y ({new_AGEMA_signal_1739, new_AGEMA_signal_1738, sboxInst_n2}) ) ;
    not_LMDPL sboxInst_U1 ( .x ({new_AGEMA_signal_1729, new_AGEMA_signal_1728, sboxIn[1]}), .y ({new_AGEMA_signal_1741, new_AGEMA_signal_1740, sboxInst_n3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) sboxInst_XOR1_U1 ( .a ({new_AGEMA_signal_1733, new_AGEMA_signal_1732, sboxIn[2]}), .b ({new_AGEMA_signal_1729, new_AGEMA_signal_1728, sboxIn[1]}), .c ({new_AGEMA_signal_1743, new_AGEMA_signal_1742, sboxInst_L0}) ) ;
    linear_LMDPL #(.CONF(1'b0)) sboxInst_XOR2_U1 ( .a ({new_AGEMA_signal_1729, new_AGEMA_signal_1728, sboxIn[1]}), .b ({new_AGEMA_signal_1725, new_AGEMA_signal_1724, sboxIn[0]}), .c ({new_AGEMA_signal_1745, new_AGEMA_signal_1744, sboxInst_L1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) sboxInst_XOR3_U1 ( .a ({new_AGEMA_signal_1745, new_AGEMA_signal_1744, sboxInst_L1}), .b ({new_AGEMA_signal_1737, new_AGEMA_signal_1736, sboxIn[3]}), .c ({new_AGEMA_signal_1779, new_AGEMA_signal_1778, sboxInst_L2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) sboxInst_XOR16_U1 ( .a ({new_AGEMA_signal_1787, new_AGEMA_signal_1786, sboxInst_T0}), .b ({new_AGEMA_signal_1779, new_AGEMA_signal_1778, sboxInst_L2}), .c ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, sboxInst_Q2}) ) ;
    linear_LMDPL #(.CONF(1'b0)) sboxInst_XOR4_U1 ( .a ({new_AGEMA_signal_1737, new_AGEMA_signal_1736, sboxIn[3]}), .b ({new_AGEMA_signal_1725, new_AGEMA_signal_1724, sboxIn[0]}), .c ({new_AGEMA_signal_1747, new_AGEMA_signal_1746, sboxInst_L3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) sboxInst_XOR5_U1 ( .a ({new_AGEMA_signal_1747, new_AGEMA_signal_1746, sboxInst_L3}), .b ({new_AGEMA_signal_1743, new_AGEMA_signal_1742, sboxInst_L0}), .c ({new_AGEMA_signal_1781, new_AGEMA_signal_1780, sboxInst_Q3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) sboxInst_XOR6_U1 ( .a ({new_AGEMA_signal_1737, new_AGEMA_signal_1736, sboxIn[3]}), .b ({new_AGEMA_signal_1729, new_AGEMA_signal_1728, sboxIn[1]}), .c ({new_AGEMA_signal_1749, new_AGEMA_signal_1748, sboxInst_L4}) ) ;
    linear_LMDPL #(.CONF(1'b0)) sboxInst_XOR7_U1 ( .a ({new_AGEMA_signal_1787, new_AGEMA_signal_1786, sboxInst_T0}), .b ({new_AGEMA_signal_1785, new_AGEMA_signal_1784, sboxInst_T2}), .c ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, sboxInst_L5}) ) ;
    linear_LMDPL #(.CONF(1'b1)) sboxInst_XOR8_U1 ( .a ({new_AGEMA_signal_1749, new_AGEMA_signal_1748, sboxInst_L4}), .b ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, sboxInst_L5}), .c ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, sboxInst_Q6}) ) ;
    linear_LMDPL #(.CONF(1'b0)) sboxInst_XOR9_U1 ( .a ({new_AGEMA_signal_1745, new_AGEMA_signal_1744, sboxInst_L1}), .b ({new_AGEMA_signal_1733, new_AGEMA_signal_1732, sboxIn[2]}), .c ({new_AGEMA_signal_1783, new_AGEMA_signal_1782, sboxInst_Q7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) sboxInst_AND1_U1 ( .a ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, sboxInst_n1}), .b ({new_AGEMA_signal_1739, new_AGEMA_signal_1738, sboxInst_n2}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[0]), .c ({new_AGEMA_signal_1787, new_AGEMA_signal_1786, sboxInst_T0}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) sboxInst_AND2_U1 ( .a ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, sboxInst_Q2}), .b ({new_AGEMA_signal_1781, new_AGEMA_signal_1780, sboxInst_Q3}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[1]), .c ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, sboxInst_T1}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) sboxInst_AND3_U1 ( .a ({new_AGEMA_signal_1741, new_AGEMA_signal_1740, sboxInst_n3}), .b ({new_AGEMA_signal_1733, new_AGEMA_signal_1732, sboxIn[2]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[2]), .c ({new_AGEMA_signal_1785, new_AGEMA_signal_1784, sboxInst_T2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) sboxInst_AND4_U1 ( .a ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, sboxInst_Q6}), .b ({new_AGEMA_signal_1783, new_AGEMA_signal_1782, sboxInst_Q7}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[3]), .c ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, sboxInst_T3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) sboxInst_XOR10_U1 ( .a ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, sboxInst_L5}), .b ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, sboxInst_T3}), .c ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, sboxInst_L7}) ) ;
    linear_LMDPL #(.CONF(1'b0)) sboxInst_XOR11_U1 ( .a ({new_AGEMA_signal_1725, new_AGEMA_signal_1724, sboxIn[0]}), .b ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, sboxInst_L7}), .c ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, sboxOut[3]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) sboxInst_XOR12_U1 ( .a ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, sboxInst_L5}), .b ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, sboxInst_T1}), .c ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, sboxInst_L8}) ) ;
    linear_LMDPL #(.CONF(1'b0)) sboxInst_XOR13_U1 ( .a ({new_AGEMA_signal_1745, new_AGEMA_signal_1744, sboxInst_L1}), .b ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, sboxInst_L8}), .c ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, sboxOut[2]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) sboxInst_XOR14_U1 ( .a ({new_AGEMA_signal_1749, new_AGEMA_signal_1748, sboxInst_L4}), .b ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, sboxInst_T3}), .c ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, sboxOut[1]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) sboxInst_XOR15_U1 ( .a ({new_AGEMA_signal_1747, new_AGEMA_signal_1746, sboxInst_L3}), .b ({new_AGEMA_signal_1785, new_AGEMA_signal_1784, sboxInst_T2}), .c ({new_AGEMA_signal_1789, new_AGEMA_signal_1788, sboxOut[0]}) ) ;
    mux2_masked_LMDPL MUX_sboxin_mux_inst_0_U1 ( .s ({new_AGEMA_signal_1723, new_AGEMA_signal_1722, selSbox}), .b ({new_AGEMA_signal_865, new_AGEMA_signal_864, stateXORroundkey[0]}), .a ({new_AGEMA_signal_879, new_AGEMA_signal_878, roundkey[3]}), .c ({new_AGEMA_signal_1725, new_AGEMA_signal_1724, sboxIn[0]}) ) ;
    mux2_masked_LMDPL MUX_sboxin_mux_inst_1_U1 ( .s ({new_AGEMA_signal_1723, new_AGEMA_signal_1722, selSbox}), .b ({new_AGEMA_signal_871, new_AGEMA_signal_870, stateXORroundkey[1]}), .a ({new_AGEMA_signal_1727, new_AGEMA_signal_1726, keyRegKS[1]}), .c ({new_AGEMA_signal_1729, new_AGEMA_signal_1728, sboxIn[1]}) ) ;
    mux2_masked_LMDPL MUX_sboxin_mux_inst_2_U1 ( .s ({new_AGEMA_signal_1723, new_AGEMA_signal_1722, selSbox}), .b ({new_AGEMA_signal_877, new_AGEMA_signal_876, stateXORroundkey[2]}), .a ({new_AGEMA_signal_1731, new_AGEMA_signal_1730, keyRegKS[2]}), .c ({new_AGEMA_signal_1733, new_AGEMA_signal_1732, sboxIn[2]}) ) ;
    mux2_masked_LMDPL MUX_sboxin_mux_inst_3_U1 ( .s ({new_AGEMA_signal_1723, new_AGEMA_signal_1722, selSbox}), .b ({new_AGEMA_signal_883, new_AGEMA_signal_882, stateXORroundkey[3]}), .a ({new_AGEMA_signal_1735, new_AGEMA_signal_1734, keyRegKS[3]}), .c ({new_AGEMA_signal_1737, new_AGEMA_signal_1736, sboxIn[3]}) ) ;
    mux2_masked_LMDPL MUX_serialIn_mux_inst_0_U1 ( .s ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, intDone}), .b ({new_AGEMA_signal_1789, new_AGEMA_signal_1788, sboxOut[0]}), .a ({new_AGEMA_signal_865, new_AGEMA_signal_864, stateXORroundkey[0]}), .c ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, serialIn[0]}) ) ;
    mux2_masked_LMDPL MUX_serialIn_mux_inst_1_U1 ( .s ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, intDone}), .b ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, sboxOut[1]}), .a ({new_AGEMA_signal_871, new_AGEMA_signal_870, stateXORroundkey[1]}), .c ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, serialIn[1]}) ) ;
    mux2_masked_LMDPL MUX_serialIn_mux_inst_2_U1 ( .s ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, intDone}), .b ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, sboxOut[2]}), .a ({new_AGEMA_signal_877, new_AGEMA_signal_876, stateXORroundkey[2]}), .c ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, serialIn[2]}) ) ;
    mux2_masked_LMDPL MUX_serialIn_mux_inst_3_U1 ( .s ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, intDone}), .b ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, sboxOut[3]}), .a ({new_AGEMA_signal_883, new_AGEMA_signal_882, stateXORroundkey[3]}), .c ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, serialIn[3]}) ) ;
    Precharger_reg new_AGEMA_gate_704 ( .D (reset), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_885, new_AGEMA_signal_884}) ) ;
    Precharger_reg new_AGEMA_gate_705 ( .D (selSbox), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_1723, new_AGEMA_signal_1722}) ) ;
    Precharger_reg new_AGEMA_gate_706 ( .D (ctrlData_0_), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_1751, new_AGEMA_signal_1750}) ) ;
    Precharger_reg new_AGEMA_gate_707 ( .D (stateFF_state_n6), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_1791, new_AGEMA_signal_1790}) ) ;
    Precharger_reg new_AGEMA_gate_708 ( .D (stateFF_state_n5), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_1849, new_AGEMA_signal_1848}) ) ;
    Precharger_reg new_AGEMA_gate_709 ( .D (keyFF_keystate_n7), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_1907, new_AGEMA_signal_1906}) ) ;
    Precharger_reg new_AGEMA_gate_710 ( .D (keyFF_keystate_n6), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_1925, new_AGEMA_signal_1924}) ) ;
    Precharger_reg new_AGEMA_gate_711 ( .D (intDone), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_2055, new_AGEMA_signal_2054}) ) ;
    ClockController_LMDPL ClockControllerInst ( .clk (clk), .Po_rst (Po_rst), .pre1 (LMDPL_pre1), .pre2 (LMDPL_pre2), .mid_rst (mid_rst) ) ;
    Precharger PrechargeCell_0 ( .D (data_in_s1[63]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1259, new_AGEMA_signal_1258}) ) ;
    Precharger PrechargeCell_1 ( .D (data_in_s1[62]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1255, new_AGEMA_signal_1254}) ) ;
    Precharger PrechargeCell_2 ( .D (data_in_s1[61]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1249, new_AGEMA_signal_1248}) ) ;
    Precharger PrechargeCell_3 ( .D (data_in_s1[60]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1243, new_AGEMA_signal_1242}) ) ;
    Precharger PrechargeCell_4 ( .D (data_in_s1[59]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1237, new_AGEMA_signal_1236}) ) ;
    Precharger PrechargeCell_5 ( .D (data_in_s1[58]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1231, new_AGEMA_signal_1230}) ) ;
    Precharger PrechargeCell_6 ( .D (data_in_s1[57]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1225, new_AGEMA_signal_1224}) ) ;
    Precharger PrechargeCell_7 ( .D (data_in_s1[56]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1219, new_AGEMA_signal_1218}) ) ;
    Precharger PrechargeCell_8 ( .D (data_in_s1[55]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1213, new_AGEMA_signal_1212}) ) ;
    Precharger PrechargeCell_9 ( .D (data_in_s1[54]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1207, new_AGEMA_signal_1206}) ) ;
    Precharger PrechargeCell_10 ( .D (data_in_s1[53]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1201, new_AGEMA_signal_1200}) ) ;
    Precharger PrechargeCell_11 ( .D (data_in_s1[52]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1195, new_AGEMA_signal_1194}) ) ;
    Precharger PrechargeCell_12 ( .D (data_in_s1[51]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1189, new_AGEMA_signal_1188}) ) ;
    Precharger PrechargeCell_13 ( .D (data_in_s1[50]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1183, new_AGEMA_signal_1182}) ) ;
    Precharger PrechargeCell_14 ( .D (data_in_s1[49]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1177, new_AGEMA_signal_1176}) ) ;
    Precharger PrechargeCell_15 ( .D (data_in_s1[48]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1171, new_AGEMA_signal_1170}) ) ;
    Precharger PrechargeCell_16 ( .D (data_in_s1[47]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1165, new_AGEMA_signal_1164}) ) ;
    Precharger PrechargeCell_17 ( .D (data_in_s1[46]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1161, new_AGEMA_signal_1160}) ) ;
    Precharger PrechargeCell_18 ( .D (data_in_s1[45]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1155, new_AGEMA_signal_1154}) ) ;
    Precharger PrechargeCell_19 ( .D (data_in_s1[44]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1149, new_AGEMA_signal_1148}) ) ;
    Precharger PrechargeCell_20 ( .D (data_in_s1[43]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1143, new_AGEMA_signal_1142}) ) ;
    Precharger PrechargeCell_21 ( .D (data_in_s1[42]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1137, new_AGEMA_signal_1136}) ) ;
    Precharger PrechargeCell_22 ( .D (data_in_s1[41]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1131, new_AGEMA_signal_1130}) ) ;
    Precharger PrechargeCell_23 ( .D (data_in_s1[40]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1125, new_AGEMA_signal_1124}) ) ;
    Precharger PrechargeCell_24 ( .D (data_in_s1[39]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1119, new_AGEMA_signal_1118}) ) ;
    Precharger PrechargeCell_25 ( .D (data_in_s1[38]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1113, new_AGEMA_signal_1112}) ) ;
    Precharger PrechargeCell_26 ( .D (data_in_s1[37]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1107, new_AGEMA_signal_1106}) ) ;
    Precharger PrechargeCell_27 ( .D (data_in_s1[36]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1101, new_AGEMA_signal_1100}) ) ;
    Precharger PrechargeCell_28 ( .D (data_in_s1[35]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1095, new_AGEMA_signal_1094}) ) ;
    Precharger PrechargeCell_29 ( .D (data_in_s1[34]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1089, new_AGEMA_signal_1088}) ) ;
    Precharger PrechargeCell_30 ( .D (data_in_s1[33]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1083, new_AGEMA_signal_1082}) ) ;
    Precharger PrechargeCell_31 ( .D (data_in_s1[32]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1077, new_AGEMA_signal_1076}) ) ;
    Precharger PrechargeCell_32 ( .D (data_in_s1[31]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1071, new_AGEMA_signal_1070}) ) ;
    Precharger PrechargeCell_33 ( .D (data_in_s1[30]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1067, new_AGEMA_signal_1066}) ) ;
    Precharger PrechargeCell_34 ( .D (data_in_s1[29]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1061, new_AGEMA_signal_1060}) ) ;
    Precharger PrechargeCell_35 ( .D (data_in_s1[28]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1055, new_AGEMA_signal_1054}) ) ;
    Precharger PrechargeCell_36 ( .D (data_in_s1[27]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1049, new_AGEMA_signal_1048}) ) ;
    Precharger PrechargeCell_37 ( .D (data_in_s1[26]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1043, new_AGEMA_signal_1042}) ) ;
    Precharger PrechargeCell_38 ( .D (data_in_s1[25]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1037, new_AGEMA_signal_1036}) ) ;
    Precharger PrechargeCell_39 ( .D (data_in_s1[24]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1031, new_AGEMA_signal_1030}) ) ;
    Precharger PrechargeCell_40 ( .D (data_in_s1[23]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1025, new_AGEMA_signal_1024}) ) ;
    Precharger PrechargeCell_41 ( .D (data_in_s1[22]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1019, new_AGEMA_signal_1018}) ) ;
    Precharger PrechargeCell_42 ( .D (data_in_s1[21]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1013, new_AGEMA_signal_1012}) ) ;
    Precharger PrechargeCell_43 ( .D (data_in_s1[20]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1007, new_AGEMA_signal_1006}) ) ;
    Precharger PrechargeCell_44 ( .D (data_in_s1[19]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1001, new_AGEMA_signal_1000}) ) ;
    Precharger PrechargeCell_45 ( .D (data_in_s1[18]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_995, new_AGEMA_signal_994}) ) ;
    Precharger PrechargeCell_46 ( .D (data_in_s1[17]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_989, new_AGEMA_signal_988}) ) ;
    Precharger PrechargeCell_47 ( .D (data_in_s1[16]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_983, new_AGEMA_signal_982}) ) ;
    Precharger PrechargeCell_48 ( .D (data_in_s1[15]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_977, new_AGEMA_signal_976}) ) ;
    Precharger PrechargeCell_49 ( .D (data_in_s1[14]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_973, new_AGEMA_signal_972}) ) ;
    Precharger PrechargeCell_50 ( .D (data_in_s1[13]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_967, new_AGEMA_signal_966}) ) ;
    Precharger PrechargeCell_51 ( .D (data_in_s1[12]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_961, new_AGEMA_signal_960}) ) ;
    Precharger PrechargeCell_52 ( .D (data_in_s1[11]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_955, new_AGEMA_signal_954}) ) ;
    Precharger PrechargeCell_53 ( .D (data_in_s1[10]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_949, new_AGEMA_signal_948}) ) ;
    Precharger PrechargeCell_54 ( .D (data_in_s1[9]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_943, new_AGEMA_signal_942}) ) ;
    Precharger PrechargeCell_55 ( .D (data_in_s1[8]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_937, new_AGEMA_signal_936}) ) ;
    Precharger PrechargeCell_56 ( .D (data_in_s1[7]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_931, new_AGEMA_signal_930}) ) ;
    Precharger PrechargeCell_57 ( .D (data_in_s1[6]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_925, new_AGEMA_signal_924}) ) ;
    Precharger PrechargeCell_58 ( .D (data_in_s1[5]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_919, new_AGEMA_signal_918}) ) ;
    Precharger PrechargeCell_59 ( .D (data_in_s1[4]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_913, new_AGEMA_signal_912}) ) ;
    Precharger PrechargeCell_60 ( .D (data_in_s1[3]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_907, new_AGEMA_signal_906}) ) ;
    Precharger PrechargeCell_61 ( .D (data_in_s1[2]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_901, new_AGEMA_signal_900}) ) ;
    Precharger PrechargeCell_62 ( .D (data_in_s1[1]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_895, new_AGEMA_signal_894}) ) ;
    Precharger PrechargeCell_63 ( .D (data_in_s1[0]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_889, new_AGEMA_signal_888}) ) ;
    Precharger PrechargeCell_64 ( .D (key_s1[79]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2099, new_AGEMA_signal_2098}) ) ;
    Precharger PrechargeCell_65 ( .D (key_s1[78]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2081, new_AGEMA_signal_2080}) ) ;
    Precharger PrechargeCell_66 ( .D (key_s1[77]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2077, new_AGEMA_signal_2076}) ) ;
    Precharger PrechargeCell_67 ( .D (key_s1[76]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2047, new_AGEMA_signal_2046}) ) ;
    Precharger PrechargeCell_68 ( .D (key_s1[75]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1695, new_AGEMA_signal_1694}) ) ;
    Precharger PrechargeCell_69 ( .D (key_s1[74]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1691, new_AGEMA_signal_1690}) ) ;
    Precharger PrechargeCell_70 ( .D (key_s1[73]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1687, new_AGEMA_signal_1686}) ) ;
    Precharger PrechargeCell_71 ( .D (key_s1[72]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1683, new_AGEMA_signal_1682}) ) ;
    Precharger PrechargeCell_72 ( .D (key_s1[71]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1677, new_AGEMA_signal_1676}) ) ;
    Precharger PrechargeCell_73 ( .D (key_s1[70]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1671, new_AGEMA_signal_1670}) ) ;
    Precharger PrechargeCell_74 ( .D (key_s1[69]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1665, new_AGEMA_signal_1664}) ) ;
    Precharger PrechargeCell_75 ( .D (key_s1[68]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1659, new_AGEMA_signal_1658}) ) ;
    Precharger PrechargeCell_76 ( .D (key_s1[67]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1653, new_AGEMA_signal_1652}) ) ;
    Precharger PrechargeCell_77 ( .D (key_s1[66]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1647, new_AGEMA_signal_1646}) ) ;
    Precharger PrechargeCell_78 ( .D (key_s1[65]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1641, new_AGEMA_signal_1640}) ) ;
    Precharger PrechargeCell_79 ( .D (key_s1[64]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1635, new_AGEMA_signal_1634}) ) ;
    Precharger PrechargeCell_80 ( .D (key_s1[63]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1629, new_AGEMA_signal_1628}) ) ;
    Precharger PrechargeCell_81 ( .D (key_s1[62]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1623, new_AGEMA_signal_1622}) ) ;
    Precharger PrechargeCell_82 ( .D (key_s1[61]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1617, new_AGEMA_signal_1616}) ) ;
    Precharger PrechargeCell_83 ( .D (key_s1[60]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1611, new_AGEMA_signal_1610}) ) ;
    Precharger PrechargeCell_84 ( .D (key_s1[59]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1605, new_AGEMA_signal_1604}) ) ;
    Precharger PrechargeCell_85 ( .D (key_s1[58]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1599, new_AGEMA_signal_1598}) ) ;
    Precharger PrechargeCell_86 ( .D (key_s1[57]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1593, new_AGEMA_signal_1592}) ) ;
    Precharger PrechargeCell_87 ( .D (key_s1[56]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1587, new_AGEMA_signal_1586}) ) ;
    Precharger PrechargeCell_88 ( .D (key_s1[55]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1581, new_AGEMA_signal_1580}) ) ;
    Precharger PrechargeCell_89 ( .D (key_s1[54]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1575, new_AGEMA_signal_1574}) ) ;
    Precharger PrechargeCell_90 ( .D (key_s1[53]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1569, new_AGEMA_signal_1568}) ) ;
    Precharger PrechargeCell_91 ( .D (key_s1[52]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1563, new_AGEMA_signal_1562}) ) ;
    Precharger PrechargeCell_92 ( .D (key_s1[51]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1557, new_AGEMA_signal_1556}) ) ;
    Precharger PrechargeCell_93 ( .D (key_s1[50]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1551, new_AGEMA_signal_1550}) ) ;
    Precharger PrechargeCell_94 ( .D (key_s1[49]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1545, new_AGEMA_signal_1544}) ) ;
    Precharger PrechargeCell_95 ( .D (key_s1[48]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1539, new_AGEMA_signal_1538}) ) ;
    Precharger PrechargeCell_96 ( .D (key_s1[47]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1533, new_AGEMA_signal_1532}) ) ;
    Precharger PrechargeCell_97 ( .D (key_s1[46]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1527, new_AGEMA_signal_1526}) ) ;
    Precharger PrechargeCell_98 ( .D (key_s1[45]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1521, new_AGEMA_signal_1520}) ) ;
    Precharger PrechargeCell_99 ( .D (key_s1[44]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1515, new_AGEMA_signal_1514}) ) ;
    Precharger PrechargeCell_100 ( .D (key_s1[43]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1509, new_AGEMA_signal_1508}) ) ;
    Precharger PrechargeCell_101 ( .D (key_s1[42]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1503, new_AGEMA_signal_1502}) ) ;
    Precharger PrechargeCell_102 ( .D (key_s1[41]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1497, new_AGEMA_signal_1496}) ) ;
    Precharger PrechargeCell_103 ( .D (key_s1[40]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1491, new_AGEMA_signal_1490}) ) ;
    Precharger PrechargeCell_104 ( .D (key_s1[39]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1485, new_AGEMA_signal_1484}) ) ;
    Precharger PrechargeCell_105 ( .D (key_s1[38]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1479, new_AGEMA_signal_1478}) ) ;
    Precharger PrechargeCell_106 ( .D (key_s1[37]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1473, new_AGEMA_signal_1472}) ) ;
    Precharger PrechargeCell_107 ( .D (key_s1[36]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1467, new_AGEMA_signal_1466}) ) ;
    Precharger PrechargeCell_108 ( .D (key_s1[35]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1461, new_AGEMA_signal_1460}) ) ;
    Precharger PrechargeCell_109 ( .D (key_s1[34]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1455, new_AGEMA_signal_1454}) ) ;
    Precharger PrechargeCell_110 ( .D (key_s1[33]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1449, new_AGEMA_signal_1448}) ) ;
    Precharger PrechargeCell_111 ( .D (key_s1[32]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1443, new_AGEMA_signal_1442}) ) ;
    Precharger PrechargeCell_112 ( .D (key_s1[31]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1437, new_AGEMA_signal_1436}) ) ;
    Precharger PrechargeCell_113 ( .D (key_s1[30]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1431, new_AGEMA_signal_1430}) ) ;
    Precharger PrechargeCell_114 ( .D (key_s1[29]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1425, new_AGEMA_signal_1424}) ) ;
    Precharger PrechargeCell_115 ( .D (key_s1[28]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1419, new_AGEMA_signal_1418}) ) ;
    Precharger PrechargeCell_116 ( .D (key_s1[27]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1413, new_AGEMA_signal_1412}) ) ;
    Precharger PrechargeCell_117 ( .D (key_s1[26]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1407, new_AGEMA_signal_1406}) ) ;
    Precharger PrechargeCell_118 ( .D (key_s1[25]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1401, new_AGEMA_signal_1400}) ) ;
    Precharger PrechargeCell_119 ( .D (key_s1[24]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1395, new_AGEMA_signal_1394}) ) ;
    Precharger PrechargeCell_120 ( .D (key_s1[23]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1389, new_AGEMA_signal_1388}) ) ;
    Precharger PrechargeCell_121 ( .D (key_s1[22]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1383, new_AGEMA_signal_1382}) ) ;
    Precharger PrechargeCell_122 ( .D (key_s1[21]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1377, new_AGEMA_signal_1376}) ) ;
    Precharger PrechargeCell_123 ( .D (key_s1[20]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1371, new_AGEMA_signal_1370}) ) ;
    Precharger PrechargeCell_124 ( .D (key_s1[19]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1715, new_AGEMA_signal_1714}) ) ;
    Precharger PrechargeCell_125 ( .D (key_s1[18]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1711, new_AGEMA_signal_1710}) ) ;
    Precharger PrechargeCell_126 ( .D (key_s1[17]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1707, new_AGEMA_signal_1706}) ) ;
    Precharger PrechargeCell_127 ( .D (key_s1[16]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1719, new_AGEMA_signal_1718}) ) ;
    Precharger PrechargeCell_128 ( .D (key_s1[15]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1703, new_AGEMA_signal_1702}) ) ;
    Precharger PrechargeCell_129 ( .D (key_s1[14]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1365, new_AGEMA_signal_1364}) ) ;
    Precharger PrechargeCell_130 ( .D (key_s1[13]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1359, new_AGEMA_signal_1358}) ) ;
    Precharger PrechargeCell_131 ( .D (key_s1[12]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1353, new_AGEMA_signal_1352}) ) ;
    Precharger PrechargeCell_132 ( .D (key_s1[11]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1347, new_AGEMA_signal_1346}) ) ;
    Precharger PrechargeCell_133 ( .D (key_s1[10]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1341, new_AGEMA_signal_1340}) ) ;
    Precharger PrechargeCell_134 ( .D (key_s1[9]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1335, new_AGEMA_signal_1334}) ) ;
    Precharger PrechargeCell_135 ( .D (key_s1[8]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1329, new_AGEMA_signal_1328}) ) ;
    Precharger PrechargeCell_136 ( .D (key_s1[7]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1323, new_AGEMA_signal_1322}) ) ;
    Precharger PrechargeCell_137 ( .D (key_s1[6]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1317, new_AGEMA_signal_1316}) ) ;
    Precharger PrechargeCell_138 ( .D (key_s1[5]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1311, new_AGEMA_signal_1310}) ) ;
    Precharger PrechargeCell_139 ( .D (key_s1[4]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1305, new_AGEMA_signal_1304}) ) ;
    Precharger PrechargeCell_140 ( .D (key_s1[3]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1299, new_AGEMA_signal_1298}) ) ;
    Precharger PrechargeCell_141 ( .D (key_s1[2]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1293, new_AGEMA_signal_1292}) ) ;
    Precharger PrechargeCell_142 ( .D (key_s1[1]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1287, new_AGEMA_signal_1286}) ) ;
    Precharger PrechargeCell_143 ( .D (key_s1[0]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1281, new_AGEMA_signal_1280}) ) ;

    /* register cells */
    reg_sr_LMDPL fsm_cnt_rnd_count_reg_reg_4__FF_FF ( .D (fsm_cnt_rnd_n14), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (counter[4]), .QN () ) ;
    reg_sr_LMDPL fsm_cnt_rnd_count_reg_reg_2__FF_FF ( .D (fsm_cnt_rnd_n16), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (counter[2]), .QN () ) ;
    reg_sr_LMDPL fsm_cnt_rnd_count_reg_reg_0__FF_FF ( .D (fsm_cnt_rnd_n18), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (counter[0]), .QN () ) ;
    reg_sr_LMDPL fsm_cnt_rnd_count_reg_reg_3__FF_FF ( .D (fsm_cnt_rnd_n1), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (counter[3]), .QN () ) ;
    reg_sr_LMDPL fsm_cnt_rnd_count_reg_reg_1__FF_FF ( .D (fsm_cnt_rnd_n41), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (fsm_cnt_rnd_n24), .QN () ) ;
    reg_sr_LMDPL fsm_cnt_ser_count_reg_reg_2__FF_FF ( .D (fsm_cnt_ser_n1), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (fsm_countSerial[2]), .QN () ) ;
    reg_sr_LMDPL fsm_cnt_ser_count_reg_reg_0__FF_FF ( .D (fsm_cnt_ser_n3), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (fsm_countSerial[0]), .QN () ) ;
    reg_sr_LMDPL fsm_cnt_ser_count_reg_reg_3__FF_FF ( .D (fsm_cnt_ser_n26), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (fsm_countSerial[3]), .QN () ) ;
    reg_sr_LMDPL fsm_cnt_ser_count_reg_reg_1__FF_FF ( .D (fsm_cnt_ser_n28), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (fsm_countSerial[1]), .QN () ) ;
    reg_sr_LMDPL fsm_ps_state_reg_0__FF_FF ( .D (fsm_n21), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (fsm_ps_state_0_), .QN () ) ;
    reg_sr_LMDPL fsm_ps_state_reg_1__FF_FF ( .D (fsm_n20), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (fsm_ps_state_1_), .QN () ) ;
    reg_LMDPL stateFF_state_gff_1_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, stateFF_state_gff_1_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_887, data_out_s1[0], data_out_s0[0]}) ) ;
    reg_LMDPL stateFF_state_gff_1_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, stateFF_state_gff_1_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1075, data_out_s1[2], data_out_s0[2]}) ) ;
    reg_LMDPL stateFF_state_gff_1_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, stateFF_state_gff_1_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_981, data_out_s1[1], data_out_s0[1]}) ) ;
    reg_LMDPL stateFF_state_gff_1_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, stateFF_state_gff_1_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1169, data_out_s1[3], data_out_s0[3]}) ) ;
    reg_LMDPL stateFF_state_gff_2_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_1759, new_AGEMA_signal_1758, stateFF_state_gff_2_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1175, data_out_s1[7], data_out_s0[7]}) ) ;
    reg_LMDPL stateFF_state_gff_2_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_1757, new_AGEMA_signal_1756, stateFF_state_gff_2_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1081, data_out_s1[6], data_out_s0[6]}) ) ;
    reg_LMDPL stateFF_state_gff_2_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_1755, new_AGEMA_signal_1754, stateFF_state_gff_2_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_987, data_out_s1[5], data_out_s0[5]}) ) ;
    reg_LMDPL stateFF_state_gff_2_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_1753, new_AGEMA_signal_1752, stateFF_state_gff_2_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_893, data_out_s1[4], data_out_s0[4]}) ) ;
    reg_LMDPL stateFF_state_gff_3_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_1799, new_AGEMA_signal_1798, stateFF_state_gff_3_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1181, data_out_s1[11], data_out_s0[11]}) ) ;
    reg_LMDPL stateFF_state_gff_3_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_1797, new_AGEMA_signal_1796, stateFF_state_gff_3_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1087, data_out_s1[10], data_out_s0[10]}) ) ;
    reg_LMDPL stateFF_state_gff_3_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_1795, new_AGEMA_signal_1794, stateFF_state_gff_3_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_993, data_out_s1[9], data_out_s0[9]}) ) ;
    reg_LMDPL stateFF_state_gff_3_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_1793, new_AGEMA_signal_1792, stateFF_state_gff_3_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_899, data_out_s1[8], data_out_s0[8]}) ) ;
    reg_LMDPL stateFF_state_gff_4_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_1807, new_AGEMA_signal_1806, stateFF_state_gff_4_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1187, data_out_s1[15], data_out_s0[15]}) ) ;
    reg_LMDPL stateFF_state_gff_4_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_1805, new_AGEMA_signal_1804, stateFF_state_gff_4_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1093, data_out_s1[14], data_out_s0[14]}) ) ;
    reg_LMDPL stateFF_state_gff_4_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_1803, new_AGEMA_signal_1802, stateFF_state_gff_4_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_999, data_out_s1[13], data_out_s0[13]}) ) ;
    reg_LMDPL stateFF_state_gff_4_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_1801, new_AGEMA_signal_1800, stateFF_state_gff_4_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_905, data_out_s1[12], data_out_s0[12]}) ) ;
    reg_LMDPL stateFF_state_gff_5_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_1815, new_AGEMA_signal_1814, stateFF_state_gff_5_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1193, data_out_s1[19], data_out_s0[19]}) ) ;
    reg_LMDPL stateFF_state_gff_5_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_1813, new_AGEMA_signal_1812, stateFF_state_gff_5_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1099, data_out_s1[18], data_out_s0[18]}) ) ;
    reg_LMDPL stateFF_state_gff_5_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_1811, new_AGEMA_signal_1810, stateFF_state_gff_5_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1005, data_out_s1[17], data_out_s0[17]}) ) ;
    reg_LMDPL stateFF_state_gff_5_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, stateFF_state_gff_5_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_911, data_out_s1[16], data_out_s0[16]}) ) ;
    reg_LMDPL stateFF_state_gff_6_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_1823, new_AGEMA_signal_1822, stateFF_state_gff_6_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1199, data_out_s1[23], data_out_s0[23]}) ) ;
    reg_LMDPL stateFF_state_gff_6_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_1821, new_AGEMA_signal_1820, stateFF_state_gff_6_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1105, data_out_s1[22], data_out_s0[22]}) ) ;
    reg_LMDPL stateFF_state_gff_6_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_1819, new_AGEMA_signal_1818, stateFF_state_gff_6_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1011, data_out_s1[21], data_out_s0[21]}) ) ;
    reg_LMDPL stateFF_state_gff_6_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_1817, new_AGEMA_signal_1816, stateFF_state_gff_6_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_917, data_out_s1[20], data_out_s0[20]}) ) ;
    reg_LMDPL stateFF_state_gff_7_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_1831, new_AGEMA_signal_1830, stateFF_state_gff_7_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1205, data_out_s1[27], data_out_s0[27]}) ) ;
    reg_LMDPL stateFF_state_gff_7_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_1829, new_AGEMA_signal_1828, stateFF_state_gff_7_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1111, data_out_s1[26], data_out_s0[26]}) ) ;
    reg_LMDPL stateFF_state_gff_7_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_1827, new_AGEMA_signal_1826, stateFF_state_gff_7_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1017, data_out_s1[25], data_out_s0[25]}) ) ;
    reg_LMDPL stateFF_state_gff_7_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_1825, new_AGEMA_signal_1824, stateFF_state_gff_7_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_923, data_out_s1[24], data_out_s0[24]}) ) ;
    reg_LMDPL stateFF_state_gff_8_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_1839, new_AGEMA_signal_1838, stateFF_state_gff_8_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1211, data_out_s1[31], data_out_s0[31]}) ) ;
    reg_LMDPL stateFF_state_gff_8_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_1837, new_AGEMA_signal_1836, stateFF_state_gff_8_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1117, data_out_s1[30], data_out_s0[30]}) ) ;
    reg_LMDPL stateFF_state_gff_8_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_1835, new_AGEMA_signal_1834, stateFF_state_gff_8_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1023, data_out_s1[29], data_out_s0[29]}) ) ;
    reg_LMDPL stateFF_state_gff_8_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_1833, new_AGEMA_signal_1832, stateFF_state_gff_8_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_929, data_out_s1[28], data_out_s0[28]}) ) ;
    reg_LMDPL stateFF_state_gff_9_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_1847, new_AGEMA_signal_1846, stateFF_state_gff_9_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1217, data_out_s1[35], data_out_s0[35]}) ) ;
    reg_LMDPL stateFF_state_gff_9_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_1845, new_AGEMA_signal_1844, stateFF_state_gff_9_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1123, data_out_s1[34], data_out_s0[34]}) ) ;
    reg_LMDPL stateFF_state_gff_9_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_1843, new_AGEMA_signal_1842, stateFF_state_gff_9_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1029, data_out_s1[33], data_out_s0[33]}) ) ;
    reg_LMDPL stateFF_state_gff_9_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_1841, new_AGEMA_signal_1840, stateFF_state_gff_9_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_935, data_out_s1[32], data_out_s0[32]}) ) ;
    reg_LMDPL stateFF_state_gff_10_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_1857, new_AGEMA_signal_1856, stateFF_state_gff_10_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1223, data_out_s1[39], data_out_s0[39]}) ) ;
    reg_LMDPL stateFF_state_gff_10_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_1855, new_AGEMA_signal_1854, stateFF_state_gff_10_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1129, data_out_s1[38], data_out_s0[38]}) ) ;
    reg_LMDPL stateFF_state_gff_10_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_1853, new_AGEMA_signal_1852, stateFF_state_gff_10_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1035, data_out_s1[37], data_out_s0[37]}) ) ;
    reg_LMDPL stateFF_state_gff_10_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_1851, new_AGEMA_signal_1850, stateFF_state_gff_10_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_941, data_out_s1[36], data_out_s0[36]}) ) ;
    reg_LMDPL stateFF_state_gff_11_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_1865, new_AGEMA_signal_1864, stateFF_state_gff_11_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1229, data_out_s1[43], data_out_s0[43]}) ) ;
    reg_LMDPL stateFF_state_gff_11_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_1863, new_AGEMA_signal_1862, stateFF_state_gff_11_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1135, data_out_s1[42], data_out_s0[42]}) ) ;
    reg_LMDPL stateFF_state_gff_11_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_1861, new_AGEMA_signal_1860, stateFF_state_gff_11_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1041, data_out_s1[41], data_out_s0[41]}) ) ;
    reg_LMDPL stateFF_state_gff_11_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_1859, new_AGEMA_signal_1858, stateFF_state_gff_11_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_947, data_out_s1[40], data_out_s0[40]}) ) ;
    reg_LMDPL stateFF_state_gff_12_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_1873, new_AGEMA_signal_1872, stateFF_state_gff_12_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1235, data_out_s1[47], data_out_s0[47]}) ) ;
    reg_LMDPL stateFF_state_gff_12_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_1871, new_AGEMA_signal_1870, stateFF_state_gff_12_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1141, data_out_s1[46], data_out_s0[46]}) ) ;
    reg_LMDPL stateFF_state_gff_12_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, stateFF_state_gff_12_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1047, data_out_s1[45], data_out_s0[45]}) ) ;
    reg_LMDPL stateFF_state_gff_12_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_1867, new_AGEMA_signal_1866, stateFF_state_gff_12_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_953, data_out_s1[44], data_out_s0[44]}) ) ;
    reg_LMDPL stateFF_state_gff_13_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_1881, new_AGEMA_signal_1880, stateFF_state_gff_13_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1241, data_out_s1[51], data_out_s0[51]}) ) ;
    reg_LMDPL stateFF_state_gff_13_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_1879, new_AGEMA_signal_1878, stateFF_state_gff_13_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1147, data_out_s1[50], data_out_s0[50]}) ) ;
    reg_LMDPL stateFF_state_gff_13_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, stateFF_state_gff_13_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1053, data_out_s1[49], data_out_s0[49]}) ) ;
    reg_LMDPL stateFF_state_gff_13_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_1875, new_AGEMA_signal_1874, stateFF_state_gff_13_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_959, data_out_s1[48], data_out_s0[48]}) ) ;
    reg_LMDPL stateFF_state_gff_14_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, stateFF_state_gff_14_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1247, data_out_s1[55], data_out_s0[55]}) ) ;
    reg_LMDPL stateFF_state_gff_14_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_1887, new_AGEMA_signal_1886, stateFF_state_gff_14_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1153, data_out_s1[54], data_out_s0[54]}) ) ;
    reg_LMDPL stateFF_state_gff_14_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_1885, new_AGEMA_signal_1884, stateFF_state_gff_14_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1059, data_out_s1[53], data_out_s0[53]}) ) ;
    reg_LMDPL stateFF_state_gff_14_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_1883, new_AGEMA_signal_1882, stateFF_state_gff_14_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_965, data_out_s1[52], data_out_s0[52]}) ) ;
    reg_LMDPL stateFF_state_gff_15_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_1897, new_AGEMA_signal_1896, stateFF_state_gff_15_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1253, data_out_s1[59], data_out_s0[59]}) ) ;
    reg_LMDPL stateFF_state_gff_15_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, stateFF_state_gff_15_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1159, data_out_s1[58], data_out_s0[58]}) ) ;
    reg_LMDPL stateFF_state_gff_15_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_1893, new_AGEMA_signal_1892, stateFF_state_gff_15_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1065, data_out_s1[57], data_out_s0[57]}) ) ;
    reg_LMDPL stateFF_state_gff_15_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_1891, new_AGEMA_signal_1890, stateFF_state_gff_15_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_971, data_out_s1[56], data_out_s0[56]}) ) ;
    reg_LMDPL stateFF_state_gff_16_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, stateFF_state_gff_16_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_881, data_out_s1[63], data_out_s0[63]}) ) ;
    reg_LMDPL stateFF_state_gff_16_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_1903, new_AGEMA_signal_1902, stateFF_state_gff_16_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_875, data_out_s1[62], data_out_s0[62]}) ) ;
    reg_LMDPL stateFF_state_gff_16_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, stateFF_state_gff_16_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_869, data_out_s1[61], data_out_s0[61]}) ) ;
    reg_LMDPL stateFF_state_gff_16_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_1899, new_AGEMA_signal_1898, stateFF_state_gff_16_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_863, data_out_s1[60], data_out_s0[60]}) ) ;
    reg_LMDPL keyFF_keystate_gff_1_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_1915, new_AGEMA_signal_1914, keyFF_keystate_gff_1_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1279, new_AGEMA_signal_1278, keyFF_outputPar[3]}) ) ;
    reg_LMDPL keyFF_keystate_gff_1_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, keyFF_keystate_gff_1_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1735, new_AGEMA_signal_1734, keyRegKS[3]}) ) ;
    reg_LMDPL keyFF_keystate_gff_1_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_1911, new_AGEMA_signal_1910, keyFF_keystate_gff_1_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1731, new_AGEMA_signal_1730, keyRegKS[2]}) ) ;
    reg_LMDPL keyFF_keystate_gff_1_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_1909, new_AGEMA_signal_1908, keyFF_keystate_gff_1_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1727, new_AGEMA_signal_1726, keyRegKS[1]}) ) ;
    reg_LMDPL keyFF_keystate_gff_2_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_1923, new_AGEMA_signal_1922, keyFF_keystate_gff_2_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1303, new_AGEMA_signal_1302, keyFF_outputPar[7]}) ) ;
    reg_LMDPL keyFF_keystate_gff_2_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_1921, new_AGEMA_signal_1920, keyFF_keystate_gff_2_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1297, new_AGEMA_signal_1296, keyFF_outputPar[6]}) ) ;
    reg_LMDPL keyFF_keystate_gff_2_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_1919, new_AGEMA_signal_1918, keyFF_keystate_gff_2_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1291, new_AGEMA_signal_1290, keyFF_outputPar[5]}) ) ;
    reg_LMDPL keyFF_keystate_gff_2_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, keyFF_keystate_gff_2_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1285, new_AGEMA_signal_1284, keyFF_outputPar[4]}) ) ;
    reg_LMDPL keyFF_keystate_gff_3_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, keyFF_keystate_gff_3_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1327, new_AGEMA_signal_1326, keyFF_outputPar[11]}) ) ;
    reg_LMDPL keyFF_keystate_gff_3_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_1931, new_AGEMA_signal_1930, keyFF_keystate_gff_3_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1321, new_AGEMA_signal_1320, keyFF_outputPar[10]}) ) ;
    reg_LMDPL keyFF_keystate_gff_3_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, keyFF_keystate_gff_3_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1315, new_AGEMA_signal_1314, keyFF_outputPar[9]}) ) ;
    reg_LMDPL keyFF_keystate_gff_3_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_1927, new_AGEMA_signal_1926, keyFF_keystate_gff_3_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1309, new_AGEMA_signal_1308, keyFF_outputPar[8]}) ) ;
    reg_LMDPL keyFF_keystate_gff_4_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_1941, new_AGEMA_signal_1940, keyFF_keystate_gff_4_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1351, new_AGEMA_signal_1350, keyFF_outputPar[15]}) ) ;
    reg_LMDPL keyFF_keystate_gff_4_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_1939, new_AGEMA_signal_1938, keyFF_keystate_gff_4_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1345, new_AGEMA_signal_1344, keyFF_outputPar[14]}) ) ;
    reg_LMDPL keyFF_keystate_gff_4_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, keyFF_keystate_gff_4_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1339, new_AGEMA_signal_1338, keyFF_outputPar[13]}) ) ;
    reg_LMDPL keyFF_keystate_gff_4_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_1935, new_AGEMA_signal_1934, keyFF_keystate_gff_4_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, keyFF_outputPar[12]}) ) ;
    reg_LMDPL keyFF_keystate_gff_5_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_1767, new_AGEMA_signal_1766, keyFF_keystate_gff_5_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1699, new_AGEMA_signal_1698, keyFF_outputPar[19]}) ) ;
    reg_LMDPL keyFF_keystate_gff_5_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_1765, new_AGEMA_signal_1764, keyFF_keystate_gff_5_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1275, new_AGEMA_signal_1274, keyFF_outputPar[18]}) ) ;
    reg_LMDPL keyFF_keystate_gff_5_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_1763, new_AGEMA_signal_1762, keyFF_keystate_gff_5_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1363, new_AGEMA_signal_1362, keyFF_outputPar[17]}) ) ;
    reg_LMDPL keyFF_keystate_gff_5_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, keyFF_keystate_gff_5_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1357, new_AGEMA_signal_1356, keyFF_outputPar[16]}) ) ;
    reg_LMDPL keyFF_keystate_gff_6_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_1775, new_AGEMA_signal_1774, keyFF_keystate_gff_6_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1369, new_AGEMA_signal_1368, keyFF_outputPar[23]}) ) ;
    reg_LMDPL keyFF_keystate_gff_6_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_1773, new_AGEMA_signal_1772, keyFF_keystate_gff_6_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1263, new_AGEMA_signal_1262, keyFF_outputPar[22]}) ) ;
    reg_LMDPL keyFF_keystate_gff_6_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_1771, new_AGEMA_signal_1770, keyFF_keystate_gff_6_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1267, new_AGEMA_signal_1266, keyFF_outputPar[21]}) ) ;
    reg_LMDPL keyFF_keystate_gff_6_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_1769, new_AGEMA_signal_1768, keyFF_keystate_gff_6_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, keyFF_outputPar[20]}) ) ;
    reg_LMDPL keyFF_keystate_gff_7_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, keyFF_keystate_gff_7_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1393, new_AGEMA_signal_1392, keyFF_outputPar[27]}) ) ;
    reg_LMDPL keyFF_keystate_gff_7_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_1947, new_AGEMA_signal_1946, keyFF_keystate_gff_7_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1387, new_AGEMA_signal_1386, keyFF_outputPar[26]}) ) ;
    reg_LMDPL keyFF_keystate_gff_7_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_1945, new_AGEMA_signal_1944, keyFF_keystate_gff_7_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1381, new_AGEMA_signal_1380, keyFF_outputPar[25]}) ) ;
    reg_LMDPL keyFF_keystate_gff_7_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_1943, new_AGEMA_signal_1942, keyFF_keystate_gff_7_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1375, new_AGEMA_signal_1374, keyFF_outputPar[24]}) ) ;
    reg_LMDPL keyFF_keystate_gff_8_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_1957, new_AGEMA_signal_1956, keyFF_keystate_gff_8_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1417, new_AGEMA_signal_1416, keyFF_outputPar[31]}) ) ;
    reg_LMDPL keyFF_keystate_gff_8_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_1955, new_AGEMA_signal_1954, keyFF_keystate_gff_8_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1411, new_AGEMA_signal_1410, keyFF_outputPar[30]}) ) ;
    reg_LMDPL keyFF_keystate_gff_8_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_1953, new_AGEMA_signal_1952, keyFF_keystate_gff_8_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1405, new_AGEMA_signal_1404, keyFF_outputPar[29]}) ) ;
    reg_LMDPL keyFF_keystate_gff_8_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_1951, new_AGEMA_signal_1950, keyFF_keystate_gff_8_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1399, new_AGEMA_signal_1398, keyFF_outputPar[28]}) ) ;
    reg_LMDPL keyFF_keystate_gff_9_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, keyFF_keystate_gff_9_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1441, new_AGEMA_signal_1440, keyFF_outputPar[35]}) ) ;
    reg_LMDPL keyFF_keystate_gff_9_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_1963, new_AGEMA_signal_1962, keyFF_keystate_gff_9_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1435, new_AGEMA_signal_1434, keyFF_outputPar[34]}) ) ;
    reg_LMDPL keyFF_keystate_gff_9_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_1961, new_AGEMA_signal_1960, keyFF_keystate_gff_9_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1429, new_AGEMA_signal_1428, keyFF_outputPar[33]}) ) ;
    reg_LMDPL keyFF_keystate_gff_9_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, keyFF_keystate_gff_9_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1423, new_AGEMA_signal_1422, keyFF_outputPar[32]}) ) ;
    reg_LMDPL keyFF_keystate_gff_10_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_1973, new_AGEMA_signal_1972, keyFF_keystate_gff_10_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, keyFF_outputPar[39]}) ) ;
    reg_LMDPL keyFF_keystate_gff_10_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_1971, new_AGEMA_signal_1970, keyFF_keystate_gff_10_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1459, new_AGEMA_signal_1458, keyFF_outputPar[38]}) ) ;
    reg_LMDPL keyFF_keystate_gff_10_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, keyFF_keystate_gff_10_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1453, new_AGEMA_signal_1452, keyFF_outputPar[37]}) ) ;
    reg_LMDPL keyFF_keystate_gff_10_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_1967, new_AGEMA_signal_1966, keyFF_keystate_gff_10_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1447, new_AGEMA_signal_1446, keyFF_outputPar[36]}) ) ;
    reg_LMDPL keyFF_keystate_gff_11_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, keyFF_keystate_gff_11_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1489, new_AGEMA_signal_1488, keyFF_outputPar[43]}) ) ;
    reg_LMDPL keyFF_keystate_gff_11_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_1979, new_AGEMA_signal_1978, keyFF_keystate_gff_11_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1483, new_AGEMA_signal_1482, keyFF_outputPar[42]}) ) ;
    reg_LMDPL keyFF_keystate_gff_11_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, keyFF_keystate_gff_11_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1477, new_AGEMA_signal_1476, keyFF_outputPar[41]}) ) ;
    reg_LMDPL keyFF_keystate_gff_11_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, keyFF_keystate_gff_11_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1471, new_AGEMA_signal_1470, keyFF_outputPar[40]}) ) ;
    reg_LMDPL keyFF_keystate_gff_12_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, keyFF_keystate_gff_12_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1513, new_AGEMA_signal_1512, keyFF_outputPar[47]}) ) ;
    reg_LMDPL keyFF_keystate_gff_12_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, keyFF_keystate_gff_12_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1507, new_AGEMA_signal_1506, keyFF_outputPar[46]}) ) ;
    reg_LMDPL keyFF_keystate_gff_12_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, keyFF_keystate_gff_12_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1501, new_AGEMA_signal_1500, keyFF_outputPar[45]}) ) ;
    reg_LMDPL keyFF_keystate_gff_12_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, keyFF_keystate_gff_12_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1495, new_AGEMA_signal_1494, keyFF_outputPar[44]}) ) ;
    reg_LMDPL keyFF_keystate_gff_13_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, keyFF_keystate_gff_13_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1537, new_AGEMA_signal_1536, keyFF_outputPar[51]}) ) ;
    reg_LMDPL keyFF_keystate_gff_13_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, keyFF_keystate_gff_13_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1531, new_AGEMA_signal_1530, keyFF_outputPar[50]}) ) ;
    reg_LMDPL keyFF_keystate_gff_13_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, keyFF_keystate_gff_13_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1525, new_AGEMA_signal_1524, keyFF_outputPar[49]}) ) ;
    reg_LMDPL keyFF_keystate_gff_13_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, keyFF_keystate_gff_13_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1519, new_AGEMA_signal_1518, keyFF_outputPar[48]}) ) ;
    reg_LMDPL keyFF_keystate_gff_14_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, keyFF_keystate_gff_14_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1561, new_AGEMA_signal_1560, keyFF_outputPar[55]}) ) ;
    reg_LMDPL keyFF_keystate_gff_14_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_2003, new_AGEMA_signal_2002, keyFF_keystate_gff_14_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1555, new_AGEMA_signal_1554, keyFF_outputPar[54]}) ) ;
    reg_LMDPL keyFF_keystate_gff_14_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, keyFF_keystate_gff_14_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1549, new_AGEMA_signal_1548, keyFF_outputPar[53]}) ) ;
    reg_LMDPL keyFF_keystate_gff_14_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, keyFF_keystate_gff_14_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1543, new_AGEMA_signal_1542, keyFF_outputPar[52]}) ) ;
    reg_LMDPL keyFF_keystate_gff_15_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, keyFF_keystate_gff_15_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1585, new_AGEMA_signal_1584, keyFF_outputPar[59]}) ) ;
    reg_LMDPL keyFF_keystate_gff_15_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, keyFF_keystate_gff_15_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1579, new_AGEMA_signal_1578, keyFF_outputPar[58]}) ) ;
    reg_LMDPL keyFF_keystate_gff_15_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, keyFF_keystate_gff_15_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1573, new_AGEMA_signal_1572, keyFF_outputPar[57]}) ) ;
    reg_LMDPL keyFF_keystate_gff_15_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, keyFF_keystate_gff_15_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1567, new_AGEMA_signal_1566, keyFF_outputPar[56]}) ) ;
    reg_LMDPL keyFF_keystate_gff_16_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, keyFF_keystate_gff_16_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1609, new_AGEMA_signal_1608, keyFF_outputPar[63]}) ) ;
    reg_LMDPL keyFF_keystate_gff_16_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, keyFF_keystate_gff_16_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1603, new_AGEMA_signal_1602, keyFF_outputPar[62]}) ) ;
    reg_LMDPL keyFF_keystate_gff_16_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, keyFF_keystate_gff_16_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1597, new_AGEMA_signal_1596, keyFF_outputPar[61]}) ) ;
    reg_LMDPL keyFF_keystate_gff_16_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, keyFF_keystate_gff_16_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1591, new_AGEMA_signal_1590, keyFF_outputPar[60]}) ) ;
    reg_LMDPL keyFF_keystate_gff_17_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, keyFF_keystate_gff_17_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1633, new_AGEMA_signal_1632, keyFF_outputPar[67]}) ) ;
    reg_LMDPL keyFF_keystate_gff_17_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, keyFF_keystate_gff_17_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1627, new_AGEMA_signal_1626, keyFF_outputPar[66]}) ) ;
    reg_LMDPL keyFF_keystate_gff_17_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, keyFF_keystate_gff_17_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1621, new_AGEMA_signal_1620, keyFF_outputPar[65]}) ) ;
    reg_LMDPL keyFF_keystate_gff_17_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, keyFF_keystate_gff_17_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1615, new_AGEMA_signal_1614, keyFF_outputPar[64]}) ) ;
    reg_LMDPL keyFF_keystate_gff_18_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, keyFF_keystate_gff_18_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1657, new_AGEMA_signal_1656, keyFF_outputPar[71]}) ) ;
    reg_LMDPL keyFF_keystate_gff_18_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, keyFF_keystate_gff_18_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1651, new_AGEMA_signal_1650, keyFF_outputPar[70]}) ) ;
    reg_LMDPL keyFF_keystate_gff_18_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, keyFF_keystate_gff_18_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1645, new_AGEMA_signal_1644, keyFF_outputPar[69]}) ) ;
    reg_LMDPL keyFF_keystate_gff_18_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, keyFF_keystate_gff_18_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1639, new_AGEMA_signal_1638, keyFF_outputPar[68]}) ) ;
    reg_LMDPL keyFF_keystate_gff_19_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, keyFF_keystate_gff_19_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1681, new_AGEMA_signal_1680, keyFF_outputPar[75]}) ) ;
    reg_LMDPL keyFF_keystate_gff_19_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, keyFF_keystate_gff_19_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1675, new_AGEMA_signal_1674, keyFF_outputPar[74]}) ) ;
    reg_LMDPL keyFF_keystate_gff_19_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, keyFF_keystate_gff_19_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1669, new_AGEMA_signal_1668, keyFF_outputPar[73]}) ) ;
    reg_LMDPL keyFF_keystate_gff_19_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, keyFF_keystate_gff_19_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1663, new_AGEMA_signal_1662, keyFF_outputPar[72]}) ) ;
    reg_LMDPL keyFF_keystate_gff_20_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, keyFF_keystate_gff_20_s_next_state[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_879, new_AGEMA_signal_878, roundkey[3]}) ) ;
    reg_LMDPL keyFF_keystate_gff_20_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, keyFF_keystate_gff_20_s_next_state[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_873, new_AGEMA_signal_872, roundkey[2]}) ) ;
    reg_LMDPL keyFF_keystate_gff_20_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, keyFF_keystate_gff_20_s_next_state[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_867, new_AGEMA_signal_866, roundkey[1]}) ) ;
    reg_LMDPL keyFF_keystate_gff_20_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, keyFF_keystate_gff_20_s_next_state[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_861, new_AGEMA_signal_860, roundkey[0]}) ) ;
endmodule
