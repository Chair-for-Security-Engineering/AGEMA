/* modified netlist. Source: module SkinnyTop in file Designs/Skinny64_64_round-based/AGEMA/SkinnyTop.v */
/* clock gating is added to the circuit, the latency increased 4 time(s)  */

module SkinnyTop_HPC2_AIG_ClockGating_d1 (Plaintext_s0, Key_s0, clk, rst, Key_s1, Plaintext_s1, Fresh, Ciphertext_s0, done, Ciphertext_s1, Synch);
    input [63:0] Plaintext_s0 ;
    input [63:0] Key_s0 ;
    input clk ;
    input rst ;
    input [63:0] Key_s1 ;
    input [63:0] Plaintext_s1 ;
    input [63:0] Fresh ;
    output [63:0] Ciphertext_s0 ;
    output done ;
    output [63:0] Ciphertext_s1 ;
    output Synch ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_768 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_771 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_774 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_777 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_780 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_783 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_786 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_789 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_792 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_809 ;
    wire signal_810 ;
    wire signal_811 ;
    wire signal_812 ;
    wire signal_813 ;
    wire signal_814 ;
    wire signal_815 ;
    wire signal_816 ;
    wire signal_817 ;
    wire signal_818 ;
    wire signal_819 ;
    wire signal_820 ;
    wire signal_821 ;
    wire signal_822 ;
    wire signal_823 ;
    wire signal_824 ;
    wire signal_825 ;
    wire signal_826 ;
    wire signal_827 ;
    wire signal_828 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_831 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_834 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_837 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_840 ;
    wire signal_841 ;
    wire signal_842 ;
    wire signal_843 ;
    wire signal_844 ;
    wire signal_845 ;
    wire signal_846 ;
    wire signal_847 ;
    wire signal_848 ;
    wire signal_849 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_852 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_855 ;
    wire signal_856 ;
    wire signal_857 ;
    wire signal_858 ;
    wire signal_859 ;
    wire signal_860 ;
    wire signal_861 ;
    wire signal_862 ;
    wire signal_863 ;
    wire signal_864 ;
    wire signal_865 ;
    wire signal_866 ;
    wire signal_867 ;
    wire signal_868 ;
    wire signal_869 ;
    wire signal_870 ;
    wire signal_871 ;
    wire signal_872 ;
    wire signal_873 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_879 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_885 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_888 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_891 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_894 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_897 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_900 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_903 ;
    wire signal_939 ;
    wire signal_940 ;
    wire signal_943 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1276 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1279 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1282 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1285 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1288 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1294 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1297 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1300 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1303 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1309 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1494 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1499 ;
    wire signal_1500 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1503 ;
    wire signal_1504 ;
    wire signal_1505 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1509 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1512 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1518 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1521 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1527 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1530 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1536 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1539 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1564 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1623 ;
    wire signal_1624 ;
    wire signal_1625 ;
    wire signal_1626 ;
    wire signal_1627 ;
    wire signal_1628 ;
    wire signal_1629 ;
    wire signal_1630 ;
    wire signal_1631 ;
    wire signal_1632 ;
    wire signal_1633 ;
    wire signal_1634 ;
    wire signal_1635 ;
    wire signal_1636 ;
    wire signal_1637 ;
    wire signal_1638 ;
    wire signal_1639 ;
    wire signal_1640 ;
    wire signal_1641 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1661 ;
    wire signal_1662 ;
    wire signal_1664 ;
    wire signal_1665 ;
    wire signal_1667 ;
    wire signal_1668 ;
    wire signal_1670 ;
    wire signal_1671 ;
    wire signal_1673 ;
    wire signal_1674 ;
    wire signal_1676 ;
    wire signal_1677 ;
    wire signal_1679 ;
    wire signal_1680 ;
    wire signal_1682 ;
    wire signal_1683 ;
    wire signal_1685 ;
    wire signal_1686 ;
    wire signal_1688 ;
    wire signal_1689 ;
    wire signal_1691 ;
    wire signal_1692 ;
    wire signal_1694 ;
    wire signal_1695 ;
    wire signal_1697 ;
    wire signal_1698 ;
    wire signal_1700 ;
    wire signal_1701 ;
    wire signal_1703 ;
    wire signal_1704 ;
    wire signal_1706 ;
    wire signal_1707 ;
    wire signal_1709 ;
    wire signal_1710 ;
    wire signal_1712 ;
    wire signal_1713 ;
    wire signal_1715 ;
    wire signal_1716 ;
    wire signal_1718 ;
    wire signal_1719 ;
    wire signal_1721 ;
    wire signal_1722 ;
    wire signal_1724 ;
    wire signal_1725 ;
    wire signal_1727 ;
    wire signal_1728 ;
    wire signal_1730 ;
    wire signal_1731 ;
    wire signal_1733 ;
    wire signal_1734 ;
    wire signal_1736 ;
    wire signal_1737 ;
    wire signal_1739 ;
    wire signal_1740 ;
    wire signal_1742 ;
    wire signal_1743 ;
    wire signal_1745 ;
    wire signal_1746 ;
    wire signal_1748 ;
    wire signal_1749 ;
    wire signal_1751 ;
    wire signal_1752 ;
    wire signal_1754 ;
    wire signal_1755 ;
    wire signal_1757 ;
    wire signal_1758 ;
    wire signal_1760 ;
    wire signal_1761 ;
    wire signal_1763 ;
    wire signal_1764 ;
    wire signal_1766 ;
    wire signal_1767 ;
    wire signal_1769 ;
    wire signal_1770 ;
    wire signal_1772 ;
    wire signal_1773 ;
    wire signal_1775 ;
    wire signal_1776 ;
    wire signal_1778 ;
    wire signal_1779 ;
    wire signal_1781 ;
    wire signal_1782 ;
    wire signal_1784 ;
    wire signal_1785 ;
    wire signal_1787 ;
    wire signal_1788 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1838 ;
    wire signal_1840 ;
    wire signal_1842 ;
    wire signal_1844 ;
    wire signal_1846 ;
    wire signal_1848 ;
    wire signal_1850 ;
    wire signal_1852 ;
    wire signal_1854 ;
    wire signal_1856 ;
    wire signal_1858 ;
    wire signal_1860 ;
    wire signal_1862 ;
    wire signal_1864 ;
    wire signal_1866 ;
    wire signal_1868 ;
    wire signal_1870 ;
    wire signal_1872 ;
    wire signal_1874 ;
    wire signal_1876 ;
    wire signal_1878 ;
    wire signal_1880 ;
    wire signal_1882 ;
    wire signal_1884 ;
    wire signal_1886 ;
    wire signal_1888 ;
    wire signal_1890 ;
    wire signal_1892 ;
    wire signal_1894 ;
    wire signal_1896 ;
    wire signal_1898 ;
    wire signal_1900 ;
    wire signal_1902 ;
    wire signal_1904 ;
    wire signal_1906 ;
    wire signal_1908 ;
    wire signal_1910 ;
    wire signal_1912 ;
    wire signal_1914 ;
    wire signal_1916 ;
    wire signal_1918 ;
    wire signal_1920 ;
    wire signal_1922 ;
    wire signal_1924 ;
    wire signal_1926 ;
    wire signal_1928 ;
    wire signal_1930 ;
    wire signal_1932 ;
    wire signal_1934 ;
    wire signal_1936 ;
    wire signal_1938 ;
    wire signal_1940 ;
    wire signal_1942 ;
    wire signal_1944 ;
    wire signal_1946 ;
    wire signal_1948 ;
    wire signal_1950 ;
    wire signal_1952 ;
    wire signal_1954 ;
    wire signal_1956 ;
    wire signal_1958 ;
    wire signal_1960 ;
    wire signal_1962 ;
    wire signal_1964 ;
    wire signal_1966 ;
    wire signal_1967 ;
    wire signal_1968 ;
    wire signal_1969 ;
    wire signal_1970 ;
    wire signal_1971 ;
    wire signal_1972 ;
    wire signal_1973 ;
    wire signal_1974 ;
    wire signal_1975 ;
    wire signal_1976 ;
    wire signal_1977 ;
    wire signal_1978 ;
    wire signal_1979 ;
    wire signal_1980 ;
    wire signal_1981 ;
    wire signal_1982 ;
    wire signal_1983 ;
    wire signal_1984 ;
    wire signal_1985 ;
    wire signal_1986 ;
    wire signal_1987 ;
    wire signal_1988 ;
    wire signal_1989 ;
    wire signal_1990 ;
    wire signal_1991 ;
    wire signal_1992 ;
    wire signal_1993 ;
    wire signal_1994 ;
    wire signal_1995 ;
    wire signal_1996 ;
    wire signal_1997 ;
    wire signal_1998 ;
    wire signal_1999 ;
    wire signal_2000 ;
    wire signal_2001 ;
    wire signal_2002 ;
    wire signal_2003 ;
    wire signal_2004 ;
    wire signal_2005 ;
    wire signal_2006 ;
    wire signal_2007 ;
    wire signal_2008 ;
    wire signal_2009 ;
    wire signal_2010 ;
    wire signal_2011 ;
    wire signal_2012 ;
    wire signal_2013 ;
    wire signal_2014 ;
    wire signal_2015 ;
    wire signal_2016 ;
    wire signal_2017 ;
    wire signal_2018 ;
    wire signal_2019 ;
    wire signal_2020 ;
    wire signal_2021 ;
    wire signal_2022 ;
    wire signal_2023 ;
    wire signal_2024 ;
    wire signal_2025 ;
    wire signal_2026 ;
    wire signal_2027 ;
    wire signal_2028 ;
    wire signal_2029 ;
    wire signal_2030 ;
    wire signal_2031 ;
    wire signal_2032 ;
    wire signal_2033 ;
    wire signal_2034 ;
    wire signal_2035 ;
    wire signal_2036 ;
    wire signal_2037 ;
    wire signal_2038 ;
    wire signal_2039 ;
    wire signal_2040 ;
    wire signal_2041 ;
    wire signal_2042 ;
    wire signal_2043 ;
    wire signal_2044 ;
    wire signal_2045 ;
    wire signal_2046 ;
    wire signal_2047 ;
    wire signal_2048 ;
    wire signal_2049 ;
    wire signal_2050 ;
    wire signal_2051 ;
    wire signal_2052 ;
    wire signal_2053 ;
    wire signal_2054 ;
    wire signal_2055 ;
    wire signal_2056 ;
    wire signal_2057 ;
    wire signal_2058 ;
    wire signal_2059 ;
    wire signal_2060 ;
    wire signal_2061 ;
    wire signal_2062 ;
    wire signal_2063 ;
    wire signal_2064 ;
    wire signal_2065 ;
    wire signal_2066 ;
    wire signal_2067 ;
    wire signal_2068 ;
    wire signal_2069 ;
    wire signal_2070 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2079 ;
    wire signal_2080 ;
    wire signal_2081 ;
    wire signal_2082 ;
    wire signal_2083 ;
    wire signal_2084 ;
    wire signal_2085 ;
    wire signal_2086 ;
    wire signal_2087 ;
    wire signal_2088 ;
    wire signal_2089 ;
    wire signal_2090 ;
    wire signal_2091 ;
    wire signal_2092 ;
    wire signal_2093 ;
    wire signal_2094 ;
    wire signal_2095 ;
    wire signal_2096 ;
    wire signal_2097 ;
    wire signal_2098 ;
    wire signal_2099 ;
    wire signal_2100 ;
    wire signal_2101 ;
    wire signal_2102 ;
    wire signal_2103 ;
    wire signal_2104 ;
    wire signal_2105 ;
    wire signal_2106 ;
    wire signal_2107 ;
    wire signal_2108 ;
    wire signal_2109 ;
    wire signal_2110 ;
    wire signal_2111 ;
    wire signal_2112 ;
    wire signal_2113 ;
    wire signal_2114 ;
    wire signal_2115 ;
    wire signal_2116 ;
    wire signal_2117 ;
    wire signal_2118 ;
    wire signal_2119 ;
    wire signal_2120 ;
    wire signal_2121 ;
    wire signal_2122 ;
    wire signal_2123 ;
    wire signal_2124 ;
    wire signal_2125 ;
    wire signal_2126 ;
    wire signal_2127 ;
    wire signal_2128 ;
    wire signal_2129 ;
    wire signal_2130 ;
    wire signal_2131 ;
    wire signal_2132 ;
    wire signal_2133 ;
    wire signal_2134 ;
    wire signal_2135 ;
    wire signal_2136 ;
    wire signal_2137 ;
    wire signal_2138 ;
    wire signal_2139 ;
    wire signal_2140 ;
    wire signal_2141 ;
    wire signal_2142 ;
    wire signal_2143 ;
    wire signal_2144 ;
    wire signal_2145 ;
    wire signal_2146 ;
    wire signal_2147 ;
    wire signal_2148 ;
    wire signal_2149 ;
    wire signal_2150 ;
    wire signal_2151 ;
    wire signal_2152 ;
    wire signal_2153 ;
    wire signal_2154 ;
    wire signal_2155 ;
    wire signal_2156 ;
    wire signal_2157 ;
    wire signal_2158 ;
    wire signal_2159 ;
    wire signal_2160 ;
    wire signal_2161 ;
    wire signal_2162 ;
    wire signal_2163 ;
    wire signal_2164 ;
    wire signal_2165 ;
    wire signal_2166 ;
    wire signal_2167 ;
    wire signal_2168 ;
    wire signal_2169 ;
    wire signal_2170 ;
    wire signal_2171 ;
    wire signal_2172 ;
    wire signal_2173 ;
    wire signal_2174 ;
    wire signal_2175 ;
    wire signal_2176 ;
    wire signal_2177 ;
    wire signal_2178 ;
    wire signal_2179 ;
    wire signal_2180 ;
    wire signal_2181 ;
    wire signal_2182 ;
    wire signal_2183 ;
    wire signal_2184 ;
    wire signal_2185 ;
    wire signal_2186 ;
    wire signal_2187 ;
    wire signal_2188 ;
    wire signal_2189 ;
    wire signal_2190 ;
    wire signal_2191 ;
    wire signal_2192 ;
    wire signal_2193 ;
    wire signal_2194 ;
    wire signal_2195 ;
    wire signal_2196 ;
    wire signal_2197 ;
    wire signal_2198 ;
    wire signal_2199 ;
    wire signal_2200 ;
    wire signal_2201 ;
    wire signal_2202 ;
    wire signal_2203 ;
    wire signal_2204 ;
    wire signal_2205 ;
    wire signal_2206 ;
    wire signal_2207 ;
    wire signal_2208 ;
    wire signal_2209 ;
    wire signal_2210 ;
    wire signal_2211 ;
    wire signal_2212 ;
    wire signal_2213 ;
    wire signal_2214 ;
    wire signal_2215 ;
    wire signal_2216 ;
    wire signal_2217 ;
    wire signal_2218 ;
    wire signal_2219 ;
    wire signal_2220 ;
    wire signal_2221 ;
    wire signal_2222 ;
    wire signal_2223 ;
    wire signal_2224 ;
    wire signal_2225 ;
    wire signal_2226 ;
    wire signal_2227 ;
    wire signal_2228 ;
    wire signal_2229 ;
    wire signal_2230 ;
    wire signal_2231 ;
    wire signal_2232 ;
    wire signal_2233 ;
    wire signal_2234 ;
    wire signal_2235 ;
    wire signal_2236 ;
    wire signal_2237 ;
    wire signal_2238 ;
    wire signal_2239 ;
    wire signal_2240 ;
    wire signal_2241 ;
    wire signal_2242 ;
    wire signal_2243 ;
    wire signal_2244 ;
    wire signal_2245 ;
    wire signal_2246 ;
    wire signal_2247 ;
    wire signal_2248 ;
    wire signal_2249 ;
    wire signal_2251 ;
    wire signal_2253 ;
    wire signal_2255 ;
    wire signal_2256 ;
    wire signal_2257 ;
    wire signal_2258 ;
    wire signal_2259 ;
    wire signal_2260 ;
    wire signal_2261 ;
    wire signal_2262 ;
    wire signal_2263 ;
    wire signal_2264 ;
    wire signal_2265 ;
    wire signal_2266 ;
    wire signal_2267 ;
    wire signal_2268 ;
    wire signal_2269 ;
    wire signal_2270 ;
    wire signal_2271 ;
    wire signal_2272 ;
    wire signal_2273 ;
    wire signal_2274 ;
    wire signal_2275 ;
    wire signal_2276 ;
    wire signal_2277 ;
    wire signal_2278 ;
    wire signal_2279 ;
    wire signal_2280 ;
    wire signal_2281 ;
    wire signal_2282 ;
    wire signal_2283 ;
    wire signal_2284 ;
    wire signal_2285 ;
    wire signal_2286 ;
    wire signal_2287 ;
    wire signal_2288 ;
    wire signal_2289 ;
    wire signal_2290 ;
    wire signal_2291 ;
    wire signal_2292 ;
    wire signal_2293 ;
    wire signal_2294 ;
    wire signal_2295 ;
    wire signal_2296 ;
    wire signal_2297 ;
    wire signal_2298 ;
    wire signal_2299 ;
    wire signal_2300 ;
    wire signal_2301 ;
    wire signal_2302 ;
    wire signal_2303 ;
    wire signal_2304 ;
    wire signal_2305 ;
    wire signal_2306 ;
    wire signal_2308 ;
    wire signal_2310 ;
    wire signal_2312 ;
    wire signal_2314 ;
    wire signal_2316 ;
    wire signal_2318 ;
    wire signal_2319 ;
    wire signal_2320 ;
    wire signal_2321 ;
    wire signal_2322 ;
    wire signal_2323 ;
    wire signal_2324 ;
    wire signal_2325 ;
    wire signal_2326 ;
    wire signal_2327 ;
    wire signal_2328 ;
    wire signal_2329 ;
    wire signal_2330 ;
    wire signal_2331 ;
    wire signal_2332 ;
    wire signal_2333 ;
    wire signal_2334 ;
    wire signal_2335 ;
    wire signal_2336 ;
    wire signal_2337 ;
    wire signal_2338 ;
    wire signal_2339 ;
    wire signal_2340 ;
    wire signal_2341 ;
    wire signal_2342 ;
    wire signal_2343 ;
    wire signal_2344 ;
    wire signal_2345 ;
    wire signal_2346 ;
    wire signal_2347 ;
    wire signal_2348 ;
    wire signal_2349 ;
    wire signal_2350 ;
    wire signal_2351 ;
    wire signal_2352 ;
    wire signal_2353 ;
    wire signal_2354 ;
    wire signal_2355 ;
    wire signal_2356 ;
    wire signal_2357 ;
    wire signal_2358 ;
    wire signal_2359 ;
    wire signal_2360 ;
    wire signal_2361 ;
    wire signal_2362 ;
    wire signal_2363 ;
    wire signal_2365 ;
    wire signal_2367 ;
    wire signal_2369 ;
    wire signal_2371 ;
    wire signal_2373 ;
    wire signal_2375 ;
    wire signal_2377 ;
    wire signal_2378 ;
    wire signal_2379 ;
    wire signal_2380 ;
    wire signal_2381 ;
    wire signal_2382 ;
    wire signal_2383 ;
    wire signal_2384 ;
    wire signal_2385 ;
    wire signal_2386 ;
    wire signal_2387 ;
    wire signal_2388 ;
    wire signal_2389 ;
    wire signal_2390 ;
    wire signal_2391 ;
    wire signal_2392 ;
    wire signal_2393 ;
    wire signal_2394 ;
    wire signal_2395 ;
    wire signal_2396 ;
    wire signal_2397 ;
    wire signal_2398 ;
    wire signal_2399 ;
    wire signal_2400 ;
    wire signal_2401 ;
    wire signal_2402 ;
    wire signal_2403 ;
    wire signal_2404 ;
    wire signal_2405 ;
    wire signal_2406 ;
    wire signal_2407 ;
    wire signal_2408 ;
    wire signal_2409 ;
    wire signal_2410 ;
    wire signal_2411 ;
    wire signal_2413 ;
    wire signal_2415 ;
    wire signal_2417 ;
    wire signal_2419 ;
    wire signal_2421 ;
    wire signal_2423 ;
    wire signal_2425 ;
    wire signal_2427 ;
    wire signal_2429 ;
    wire signal_2431 ;
    wire signal_2433 ;
    wire signal_2434 ;
    wire signal_2435 ;
    wire signal_2436 ;
    wire signal_2437 ;
    wire signal_2438 ;
    wire signal_2439 ;
    wire signal_2440 ;
    wire signal_2441 ;
    wire signal_2442 ;
    wire signal_2443 ;
    wire signal_2444 ;
    wire signal_2445 ;
    wire signal_2446 ;
    wire signal_2447 ;
    wire signal_2448 ;
    wire signal_2449 ;
    wire signal_2450 ;
    wire signal_2451 ;
    wire signal_2452 ;
    wire signal_2453 ;
    wire signal_2454 ;
    wire signal_2455 ;
    wire signal_2456 ;
    wire signal_2458 ;
    wire signal_2460 ;
    wire signal_2462 ;
    wire signal_2464 ;
    wire signal_2466 ;
    wire signal_2468 ;
    wire signal_2470 ;
    wire signal_2472 ;
    wire signal_2473 ;
    wire signal_2474 ;
    wire signal_2475 ;
    wire signal_2476 ;
    wire signal_2477 ;
    wire signal_2478 ;
    wire signal_2479 ;
    wire signal_2480 ;
    wire signal_2481 ;
    wire signal_2482 ;
    wire signal_2483 ;
    wire signal_2484 ;
    wire signal_2485 ;
    wire signal_2486 ;
    wire signal_2487 ;
    wire signal_2488 ;
    wire signal_2489 ;
    wire signal_2490 ;
    wire signal_2491 ;
    wire signal_2492 ;
    wire signal_2493 ;
    wire signal_2494 ;
    wire signal_2496 ;
    wire signal_2498 ;
    wire signal_2500 ;
    wire signal_2502 ;
    wire signal_2504 ;
    wire signal_2506 ;
    wire signal_2508 ;
    wire signal_2510 ;
    wire signal_2512 ;
    wire signal_2514 ;
    wire signal_2516 ;
    wire signal_2518 ;
    wire signal_2519 ;
    wire signal_2520 ;
    wire signal_2521 ;
    wire signal_2522 ;
    wire signal_2523 ;
    wire signal_2524 ;
    wire signal_2525 ;
    wire signal_2526 ;
    wire signal_2527 ;
    wire signal_2528 ;
    wire signal_2529 ;
    wire signal_2530 ;
    wire signal_2531 ;
    wire signal_2532 ;
    wire signal_2534 ;
    wire signal_2536 ;
    wire signal_2538 ;
    wire signal_2540 ;
    wire signal_2542 ;
    wire signal_2544 ;
    wire signal_2546 ;
    wire signal_2548 ;
    wire signal_2549 ;
    wire signal_2550 ;
    wire signal_2551 ;
    wire signal_2552 ;
    wire signal_2553 ;
    wire signal_2554 ;
    wire signal_2555 ;
    wire signal_2556 ;
    wire signal_2558 ;
    wire signal_2560 ;
    wire signal_2562 ;
    wire signal_2564 ;
    wire signal_2566 ;
    wire signal_2568 ;
    wire signal_2569 ;
    wire signal_2570 ;
    wire signal_2571 ;
    wire signal_2573 ;
    wire signal_2575 ;
    wire signal_2577 ;
    wire signal_2642 ;

    /* cells in depth 0 */
    mux2_masked #(.security_order(1), .pipeline(0)) cell_769 ( .s (rst), .b ({signal_1647, signal_1163}), .a ({Key_s1[0], Key_s0[0]}), .c ({signal_1649, signal_1099}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_770 ( .s (rst), .b ({signal_1650, signal_1162}), .a ({Key_s1[1], Key_s0[1]}), .c ({signal_1652, signal_1098}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_771 ( .s (rst), .b ({signal_1653, signal_1161}), .a ({Key_s1[2], Key_s0[2]}), .c ({signal_1655, signal_1097}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_772 ( .s (rst), .b ({signal_1656, signal_1160}), .a ({Key_s1[3], Key_s0[3]}), .c ({signal_1658, signal_1096}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_773 ( .s (rst), .b ({signal_1659, signal_1159}), .a ({Key_s1[4], Key_s0[4]}), .c ({signal_1661, signal_1095}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_774 ( .s (rst), .b ({signal_1662, signal_1158}), .a ({Key_s1[5], Key_s0[5]}), .c ({signal_1664, signal_1094}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_775 ( .s (rst), .b ({signal_1665, signal_1157}), .a ({Key_s1[6], Key_s0[6]}), .c ({signal_1667, signal_1093}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_776 ( .s (rst), .b ({signal_1668, signal_1156}), .a ({Key_s1[7], Key_s0[7]}), .c ({signal_1670, signal_1092}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_777 ( .s (rst), .b ({signal_1671, signal_1155}), .a ({Key_s1[8], Key_s0[8]}), .c ({signal_1673, signal_1091}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_778 ( .s (rst), .b ({signal_1674, signal_1154}), .a ({Key_s1[9], Key_s0[9]}), .c ({signal_1676, signal_1090}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_779 ( .s (rst), .b ({signal_1677, signal_1153}), .a ({Key_s1[10], Key_s0[10]}), .c ({signal_1679, signal_1089}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_780 ( .s (rst), .b ({signal_1680, signal_1152}), .a ({Key_s1[11], Key_s0[11]}), .c ({signal_1682, signal_1088}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_781 ( .s (rst), .b ({signal_1683, signal_1151}), .a ({Key_s1[12], Key_s0[12]}), .c ({signal_1685, signal_1087}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_782 ( .s (rst), .b ({signal_1686, signal_1150}), .a ({Key_s1[13], Key_s0[13]}), .c ({signal_1688, signal_1086}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_783 ( .s (rst), .b ({signal_1689, signal_1149}), .a ({Key_s1[14], Key_s0[14]}), .c ({signal_1691, signal_1085}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_784 ( .s (rst), .b ({signal_1692, signal_1148}), .a ({Key_s1[15], Key_s0[15]}), .c ({signal_1694, signal_1084}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_785 ( .s (rst), .b ({signal_1695, signal_1147}), .a ({Key_s1[16], Key_s0[16]}), .c ({signal_1697, signal_1083}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_786 ( .s (rst), .b ({signal_1698, signal_1146}), .a ({Key_s1[17], Key_s0[17]}), .c ({signal_1700, signal_1082}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_787 ( .s (rst), .b ({signal_1701, signal_1145}), .a ({Key_s1[18], Key_s0[18]}), .c ({signal_1703, signal_1081}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_788 ( .s (rst), .b ({signal_1704, signal_1144}), .a ({Key_s1[19], Key_s0[19]}), .c ({signal_1706, signal_1080}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_789 ( .s (rst), .b ({signal_1707, signal_1143}), .a ({Key_s1[20], Key_s0[20]}), .c ({signal_1709, signal_1079}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_790 ( .s (rst), .b ({signal_1710, signal_1142}), .a ({Key_s1[21], Key_s0[21]}), .c ({signal_1712, signal_1078}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_791 ( .s (rst), .b ({signal_1713, signal_1141}), .a ({Key_s1[22], Key_s0[22]}), .c ({signal_1715, signal_1077}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_792 ( .s (rst), .b ({signal_1716, signal_1140}), .a ({Key_s1[23], Key_s0[23]}), .c ({signal_1718, signal_1076}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_793 ( .s (rst), .b ({signal_1719, signal_1139}), .a ({Key_s1[24], Key_s0[24]}), .c ({signal_1721, signal_1075}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_794 ( .s (rst), .b ({signal_1722, signal_1138}), .a ({Key_s1[25], Key_s0[25]}), .c ({signal_1724, signal_1074}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_795 ( .s (rst), .b ({signal_1725, signal_1137}), .a ({Key_s1[26], Key_s0[26]}), .c ({signal_1727, signal_1073}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_796 ( .s (rst), .b ({signal_1728, signal_1136}), .a ({Key_s1[27], Key_s0[27]}), .c ({signal_1730, signal_1072}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_797 ( .s (rst), .b ({signal_1731, signal_1135}), .a ({Key_s1[28], Key_s0[28]}), .c ({signal_1733, signal_1071}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_798 ( .s (rst), .b ({signal_1734, signal_1134}), .a ({Key_s1[29], Key_s0[29]}), .c ({signal_1736, signal_1070}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_799 ( .s (rst), .b ({signal_1737, signal_1133}), .a ({Key_s1[30], Key_s0[30]}), .c ({signal_1739, signal_1069}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_800 ( .s (rst), .b ({signal_1740, signal_1132}), .a ({Key_s1[31], Key_s0[31]}), .c ({signal_1742, signal_1068}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_801 ( .s (rst), .b ({signal_1743, signal_1131}), .a ({Key_s1[32], Key_s0[32]}), .c ({signal_1745, signal_1067}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_802 ( .s (rst), .b ({signal_1746, signal_1130}), .a ({Key_s1[33], Key_s0[33]}), .c ({signal_1748, signal_1066}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_803 ( .s (rst), .b ({signal_1749, signal_1129}), .a ({Key_s1[34], Key_s0[34]}), .c ({signal_1751, signal_1065}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_804 ( .s (rst), .b ({signal_1752, signal_1128}), .a ({Key_s1[35], Key_s0[35]}), .c ({signal_1754, signal_1064}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_805 ( .s (rst), .b ({signal_1755, signal_1127}), .a ({Key_s1[36], Key_s0[36]}), .c ({signal_1757, signal_1063}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_806 ( .s (rst), .b ({signal_1758, signal_1126}), .a ({Key_s1[37], Key_s0[37]}), .c ({signal_1760, signal_1062}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_807 ( .s (rst), .b ({signal_1761, signal_1125}), .a ({Key_s1[38], Key_s0[38]}), .c ({signal_1763, signal_1061}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_808 ( .s (rst), .b ({signal_1764, signal_1124}), .a ({Key_s1[39], Key_s0[39]}), .c ({signal_1766, signal_1060}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_809 ( .s (rst), .b ({signal_1767, signal_1123}), .a ({Key_s1[40], Key_s0[40]}), .c ({signal_1769, signal_1059}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_810 ( .s (rst), .b ({signal_1770, signal_1122}), .a ({Key_s1[41], Key_s0[41]}), .c ({signal_1772, signal_1058}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_811 ( .s (rst), .b ({signal_1773, signal_1121}), .a ({Key_s1[42], Key_s0[42]}), .c ({signal_1775, signal_1057}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_812 ( .s (rst), .b ({signal_1776, signal_1120}), .a ({Key_s1[43], Key_s0[43]}), .c ({signal_1778, signal_1056}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_813 ( .s (rst), .b ({signal_1779, signal_1119}), .a ({Key_s1[44], Key_s0[44]}), .c ({signal_1781, signal_1055}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_814 ( .s (rst), .b ({signal_1782, signal_1118}), .a ({Key_s1[45], Key_s0[45]}), .c ({signal_1784, signal_1054}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_815 ( .s (rst), .b ({signal_1785, signal_1117}), .a ({Key_s1[46], Key_s0[46]}), .c ({signal_1787, signal_1053}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_816 ( .s (rst), .b ({signal_1788, signal_1116}), .a ({Key_s1[47], Key_s0[47]}), .c ({signal_1790, signal_1052}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_817 ( .s (rst), .b ({signal_1791, signal_1115}), .a ({Key_s1[48], Key_s0[48]}), .c ({signal_1793, signal_1051}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_818 ( .s (rst), .b ({signal_1794, signal_1114}), .a ({Key_s1[49], Key_s0[49]}), .c ({signal_1796, signal_1050}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_819 ( .s (rst), .b ({signal_1797, signal_1113}), .a ({Key_s1[50], Key_s0[50]}), .c ({signal_1799, signal_1049}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_820 ( .s (rst), .b ({signal_1800, signal_1112}), .a ({Key_s1[51], Key_s0[51]}), .c ({signal_1802, signal_1048}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_821 ( .s (rst), .b ({signal_1803, signal_1111}), .a ({Key_s1[52], Key_s0[52]}), .c ({signal_1805, signal_1047}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_822 ( .s (rst), .b ({signal_1806, signal_1110}), .a ({Key_s1[53], Key_s0[53]}), .c ({signal_1808, signal_1046}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_823 ( .s (rst), .b ({signal_1809, signal_1109}), .a ({Key_s1[54], Key_s0[54]}), .c ({signal_1811, signal_1045}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_824 ( .s (rst), .b ({signal_1812, signal_1108}), .a ({Key_s1[55], Key_s0[55]}), .c ({signal_1814, signal_1044}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_825 ( .s (rst), .b ({signal_1815, signal_1107}), .a ({Key_s1[56], Key_s0[56]}), .c ({signal_1817, signal_1043}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_826 ( .s (rst), .b ({signal_1818, signal_1106}), .a ({Key_s1[57], Key_s0[57]}), .c ({signal_1820, signal_1042}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_827 ( .s (rst), .b ({signal_1821, signal_1105}), .a ({Key_s1[58], Key_s0[58]}), .c ({signal_1823, signal_1041}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_828 ( .s (rst), .b ({signal_1824, signal_1104}), .a ({Key_s1[59], Key_s0[59]}), .c ({signal_1826, signal_1040}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_829 ( .s (rst), .b ({signal_1827, signal_1103}), .a ({Key_s1[60], Key_s0[60]}), .c ({signal_1829, signal_1039}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_830 ( .s (rst), .b ({signal_1830, signal_1102}), .a ({Key_s1[61], Key_s0[61]}), .c ({signal_1832, signal_1038}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_831 ( .s (rst), .b ({signal_1833, signal_1101}), .a ({Key_s1[62], Key_s0[62]}), .c ({signal_1835, signal_1037}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_832 ( .s (rst), .b ({signal_1836, signal_1100}), .a ({Key_s1[63], Key_s0[63]}), .c ({signal_1838, signal_1036}) ) ;
    MUX2_X1 cell_961 ( .S (rst), .A (signal_1029), .B (1'b1), .Z (signal_1035) ) ;
    MUX2_X1 cell_962 ( .S (rst), .A (signal_1028), .B (1'b0), .Z (signal_1034) ) ;
    MUX2_X1 cell_963 ( .S (rst), .A (signal_1027), .B (1'b0), .Z (signal_1033) ) ;
    MUX2_X1 cell_964 ( .S (rst), .A (signal_1026), .B (1'b0), .Z (signal_1032) ) ;
    MUX2_X1 cell_965 ( .S (rst), .A (signal_1025), .B (1'b0), .Z (signal_1031) ) ;
    MUX2_X1 cell_966 ( .S (rst), .A (signal_1024), .B (1'b0), .Z (signal_1030) ) ;
    MUX2_X1 cell_979 ( .S (signal_940), .A (signal_759), .B (signal_939), .Z (signal_1029) ) ;
    NAND2_X1 cell_980 ( .A1 (signal_939), .A2 (signal_760), .ZN (signal_759) ) ;
    NAND2_X1 cell_981 ( .A1 (signal_761), .A2 (signal_762), .ZN (signal_760) ) ;
    NOR2_X1 cell_982 ( .A1 (signal_1026), .A2 (signal_1025), .ZN (signal_762) ) ;
    AND2_X1 cell_983 ( .A1 (signal_1028), .A2 (signal_943), .ZN (signal_761) ) ;
    AND2_X1 cell_984 ( .A1 (signal_763), .A2 (signal_943), .ZN (signal_1027) ) ;
    NAND2_X1 cell_985 ( .A1 (signal_764), .A2 (signal_939), .ZN (signal_763) ) ;
    NOR2_X1 cell_986 ( .A1 (signal_940), .A2 (signal_765), .ZN (signal_764) ) ;
    NAND2_X1 cell_987 ( .A1 (signal_1028), .A2 (signal_766), .ZN (signal_765) ) ;
    NOR2_X1 cell_988 ( .A1 (signal_1026), .A2 (signal_1025), .ZN (signal_766) ) ;
    OR2_X1 cell_989 ( .A1 (signal_940), .A2 (signal_767), .ZN (signal_1024) ) ;
    NOR2_X1 cell_990 ( .A1 (signal_1025), .A2 (signal_768), .ZN (signal_767) ) ;
    NAND2_X1 cell_991 ( .A1 (signal_939), .A2 (signal_769), .ZN (signal_768) ) ;
    NOR2_X1 cell_992 ( .A1 (signal_1026), .A2 (signal_770), .ZN (signal_769) ) ;
    NAND2_X1 cell_993 ( .A1 (signal_1028), .A2 (signal_943), .ZN (signal_770) ) ;
    NOR2_X1 cell_994 ( .A1 (signal_771), .A2 (signal_772), .ZN (done) ) ;
    NAND2_X1 cell_995 ( .A1 (signal_940), .A2 (signal_939), .ZN (signal_772) ) ;
    NAND2_X1 cell_996 ( .A1 (signal_773), .A2 (signal_774), .ZN (signal_771) ) ;
    NOR2_X1 cell_997 ( .A1 (signal_1025), .A2 (signal_775), .ZN (signal_774) ) ;
    INV_X1 cell_998 ( .A (signal_1028), .ZN (signal_775) ) ;
    NOR2_X1 cell_999 ( .A1 (signal_943), .A2 (signal_1026), .ZN (signal_773) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1000 ( .a ({Ciphertext_s1[2], Ciphertext_s0[2]}), .b ({signal_1840, signal_1164}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1001 ( .a ({Ciphertext_s1[6], Ciphertext_s0[6]}), .b ({signal_1842, signal_1165}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1002 ( .a ({Ciphertext_s1[10], Ciphertext_s0[10]}), .b ({signal_1844, signal_1166}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1003 ( .a ({Ciphertext_s1[14], Ciphertext_s0[14]}), .b ({signal_1846, signal_1167}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1004 ( .a ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({signal_1848, signal_1168}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1005 ( .a ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({signal_1850, signal_1169}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1006 ( .a ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({signal_1852, signal_1170}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1007 ( .a ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({signal_1854, signal_1171}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1008 ( .a ({Ciphertext_s1[34], Ciphertext_s0[34]}), .b ({signal_1856, signal_1172}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1009 ( .a ({Ciphertext_s1[38], Ciphertext_s0[38]}), .b ({signal_1858, signal_1173}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1010 ( .a ({Ciphertext_s1[42], Ciphertext_s0[42]}), .b ({signal_1860, signal_1174}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1011 ( .a ({Ciphertext_s1[46], Ciphertext_s0[46]}), .b ({signal_1862, signal_1175}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1012 ( .a ({Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({signal_1864, signal_1176}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1013 ( .a ({Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({signal_1866, signal_1177}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1014 ( .a ({Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({signal_1868, signal_1178}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1015 ( .a ({Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({signal_1870, signal_1179}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1016 ( .a ({Ciphertext_s1[2], Ciphertext_s0[2]}), .b ({Ciphertext_s1[3], Ciphertext_s0[3]}), .c ({signal_1872, signal_1180}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1017 ( .a ({Ciphertext_s1[0], Ciphertext_s0[0]}), .b ({Ciphertext_s1[2], Ciphertext_s0[2]}), .c ({signal_1874, signal_1181}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1018 ( .a ({Ciphertext_s1[6], Ciphertext_s0[6]}), .b ({Ciphertext_s1[7], Ciphertext_s0[7]}), .c ({signal_1876, signal_1182}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1019 ( .a ({Ciphertext_s1[4], Ciphertext_s0[4]}), .b ({Ciphertext_s1[6], Ciphertext_s0[6]}), .c ({signal_1878, signal_1183}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1020 ( .a ({Ciphertext_s1[10], Ciphertext_s0[10]}), .b ({Ciphertext_s1[11], Ciphertext_s0[11]}), .c ({signal_1880, signal_1184}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1021 ( .a ({Ciphertext_s1[8], Ciphertext_s0[8]}), .b ({Ciphertext_s1[10], Ciphertext_s0[10]}), .c ({signal_1882, signal_1185}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1022 ( .a ({Ciphertext_s1[14], Ciphertext_s0[14]}), .b ({Ciphertext_s1[15], Ciphertext_s0[15]}), .c ({signal_1884, signal_1186}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1023 ( .a ({Ciphertext_s1[12], Ciphertext_s0[12]}), .b ({Ciphertext_s1[14], Ciphertext_s0[14]}), .c ({signal_1886, signal_1187}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1024 ( .a ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({Ciphertext_s1[19], Ciphertext_s0[19]}), .c ({signal_1888, signal_1188}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1025 ( .a ({Ciphertext_s1[16], Ciphertext_s0[16]}), .b ({Ciphertext_s1[18], Ciphertext_s0[18]}), .c ({signal_1890, signal_1189}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1026 ( .a ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({Ciphertext_s1[23], Ciphertext_s0[23]}), .c ({signal_1892, signal_1190}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1027 ( .a ({Ciphertext_s1[20], Ciphertext_s0[20]}), .b ({Ciphertext_s1[22], Ciphertext_s0[22]}), .c ({signal_1894, signal_1191}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1028 ( .a ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({Ciphertext_s1[27], Ciphertext_s0[27]}), .c ({signal_1896, signal_1192}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1029 ( .a ({Ciphertext_s1[24], Ciphertext_s0[24]}), .b ({Ciphertext_s1[26], Ciphertext_s0[26]}), .c ({signal_1898, signal_1193}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1030 ( .a ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({Ciphertext_s1[31], Ciphertext_s0[31]}), .c ({signal_1900, signal_1194}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1031 ( .a ({Ciphertext_s1[28], Ciphertext_s0[28]}), .b ({Ciphertext_s1[30], Ciphertext_s0[30]}), .c ({signal_1902, signal_1195}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1032 ( .a ({Ciphertext_s1[34], Ciphertext_s0[34]}), .b ({Ciphertext_s1[35], Ciphertext_s0[35]}), .c ({signal_1904, signal_1196}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1033 ( .a ({Ciphertext_s1[32], Ciphertext_s0[32]}), .b ({Ciphertext_s1[34], Ciphertext_s0[34]}), .c ({signal_1906, signal_1197}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1034 ( .a ({Ciphertext_s1[38], Ciphertext_s0[38]}), .b ({Ciphertext_s1[39], Ciphertext_s0[39]}), .c ({signal_1908, signal_1198}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1035 ( .a ({Ciphertext_s1[36], Ciphertext_s0[36]}), .b ({Ciphertext_s1[38], Ciphertext_s0[38]}), .c ({signal_1910, signal_1199}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1036 ( .a ({Ciphertext_s1[42], Ciphertext_s0[42]}), .b ({Ciphertext_s1[43], Ciphertext_s0[43]}), .c ({signal_1912, signal_1200}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1037 ( .a ({Ciphertext_s1[40], Ciphertext_s0[40]}), .b ({Ciphertext_s1[42], Ciphertext_s0[42]}), .c ({signal_1914, signal_1201}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1038 ( .a ({Ciphertext_s1[46], Ciphertext_s0[46]}), .b ({Ciphertext_s1[47], Ciphertext_s0[47]}), .c ({signal_1916, signal_1202}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1039 ( .a ({Ciphertext_s1[44], Ciphertext_s0[44]}), .b ({Ciphertext_s1[46], Ciphertext_s0[46]}), .c ({signal_1918, signal_1203}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1040 ( .a ({Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({Ciphertext_s1[51], Ciphertext_s0[51]}), .c ({signal_1920, signal_1204}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1041 ( .a ({Ciphertext_s1[48], Ciphertext_s0[48]}), .b ({Ciphertext_s1[50], Ciphertext_s0[50]}), .c ({signal_1922, signal_1205}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1042 ( .a ({Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({Ciphertext_s1[55], Ciphertext_s0[55]}), .c ({signal_1924, signal_1206}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1043 ( .a ({Ciphertext_s1[52], Ciphertext_s0[52]}), .b ({Ciphertext_s1[54], Ciphertext_s0[54]}), .c ({signal_1926, signal_1207}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1044 ( .a ({Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({Ciphertext_s1[59], Ciphertext_s0[59]}), .c ({signal_1928, signal_1208}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1045 ( .a ({Ciphertext_s1[56], Ciphertext_s0[56]}), .b ({Ciphertext_s1[58], Ciphertext_s0[58]}), .c ({signal_1930, signal_1209}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1046 ( .a ({Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({Ciphertext_s1[63], Ciphertext_s0[63]}), .c ({signal_1932, signal_1210}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1047 ( .a ({Ciphertext_s1[60], Ciphertext_s0[60]}), .b ({Ciphertext_s1[62], Ciphertext_s0[62]}), .c ({signal_1934, signal_1211}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1048 ( .a ({Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({Ciphertext_s1[2], Ciphertext_s0[2]}), .c ({signal_1936, signal_1212}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1049 ( .a ({Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({Ciphertext_s1[6], Ciphertext_s0[6]}), .c ({signal_1938, signal_1213}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1050 ( .a ({Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({Ciphertext_s1[10], Ciphertext_s0[10]}), .c ({signal_1940, signal_1214}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1051 ( .a ({Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({Ciphertext_s1[14], Ciphertext_s0[14]}), .c ({signal_1942, signal_1215}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1052 ( .a ({Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({Ciphertext_s1[18], Ciphertext_s0[18]}), .c ({signal_1944, signal_1216}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1053 ( .a ({Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({Ciphertext_s1[22], Ciphertext_s0[22]}), .c ({signal_1946, signal_1217}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1054 ( .a ({Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({Ciphertext_s1[26], Ciphertext_s0[26]}), .c ({signal_1948, signal_1218}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1055 ( .a ({Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({Ciphertext_s1[30], Ciphertext_s0[30]}), .c ({signal_1950, signal_1219}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1056 ( .a ({Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({Ciphertext_s1[34], Ciphertext_s0[34]}), .c ({signal_1952, signal_1220}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1057 ( .a ({Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({Ciphertext_s1[38], Ciphertext_s0[38]}), .c ({signal_1954, signal_1221}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1058 ( .a ({Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({Ciphertext_s1[42], Ciphertext_s0[42]}), .c ({signal_1956, signal_1222}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1059 ( .a ({Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({Ciphertext_s1[46], Ciphertext_s0[46]}), .c ({signal_1958, signal_1223}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1060 ( .a ({Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({Ciphertext_s1[50], Ciphertext_s0[50]}), .c ({signal_1960, signal_1224}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1061 ( .a ({Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({Ciphertext_s1[54], Ciphertext_s0[54]}), .c ({signal_1962, signal_1225}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1062 ( .a ({Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({Ciphertext_s1[58], Ciphertext_s0[58]}), .c ({signal_1964, signal_1226}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1063 ( .a ({Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({Ciphertext_s1[62], Ciphertext_s0[62]}), .c ({signal_1966, signal_1227}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1080 ( .a ({Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({signal_1874, signal_1181}), .c ({signal_1983, signal_1244}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1081 ( .a ({Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({signal_1872, signal_1180}), .c ({signal_1984, signal_1245}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1082 ( .a ({Ciphertext_s1[2], Ciphertext_s0[2]}), .b ({signal_1874, signal_1181}), .c ({signal_1985, signal_1246}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1083 ( .a ({Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({signal_1878, signal_1183}), .c ({signal_1986, signal_1247}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1084 ( .a ({Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({signal_1876, signal_1182}), .c ({signal_1987, signal_1248}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1085 ( .a ({Ciphertext_s1[6], Ciphertext_s0[6]}), .b ({signal_1878, signal_1183}), .c ({signal_1988, signal_1249}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1086 ( .a ({Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({signal_1882, signal_1185}), .c ({signal_1989, signal_1250}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1087 ( .a ({Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({signal_1880, signal_1184}), .c ({signal_1990, signal_1251}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1088 ( .a ({Ciphertext_s1[10], Ciphertext_s0[10]}), .b ({signal_1882, signal_1185}), .c ({signal_1991, signal_1252}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1089 ( .a ({Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({signal_1886, signal_1187}), .c ({signal_1992, signal_1253}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1090 ( .a ({Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({signal_1884, signal_1186}), .c ({signal_1993, signal_1254}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1091 ( .a ({Ciphertext_s1[14], Ciphertext_s0[14]}), .b ({signal_1886, signal_1187}), .c ({signal_1994, signal_1255}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1092 ( .a ({Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({signal_1890, signal_1189}), .c ({signal_1995, signal_1256}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1093 ( .a ({Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({signal_1888, signal_1188}), .c ({signal_1996, signal_1257}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1094 ( .a ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({signal_1890, signal_1189}), .c ({signal_1997, signal_1258}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1095 ( .a ({Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({signal_1894, signal_1191}), .c ({signal_1998, signal_1259}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1096 ( .a ({Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({signal_1892, signal_1190}), .c ({signal_1999, signal_1260}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1097 ( .a ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({signal_1894, signal_1191}), .c ({signal_2000, signal_1261}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1098 ( .a ({Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({signal_1898, signal_1193}), .c ({signal_2001, signal_1262}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1099 ( .a ({Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({signal_1896, signal_1192}), .c ({signal_2002, signal_1263}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1100 ( .a ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({signal_1898, signal_1193}), .c ({signal_2003, signal_1264}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1101 ( .a ({Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({signal_1902, signal_1195}), .c ({signal_2004, signal_1265}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1102 ( .a ({Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({signal_1900, signal_1194}), .c ({signal_2005, signal_1266}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1103 ( .a ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({signal_1902, signal_1195}), .c ({signal_2006, signal_1267}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1104 ( .a ({Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({signal_1906, signal_1197}), .c ({signal_2007, signal_1268}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1105 ( .a ({Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({signal_1904, signal_1196}), .c ({signal_2008, signal_1269}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1106 ( .a ({Ciphertext_s1[34], Ciphertext_s0[34]}), .b ({signal_1906, signal_1197}), .c ({signal_2009, signal_1270}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1107 ( .a ({Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({signal_1910, signal_1199}), .c ({signal_2010, signal_1271}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1108 ( .a ({Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({signal_1908, signal_1198}), .c ({signal_2011, signal_1272}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1109 ( .a ({Ciphertext_s1[38], Ciphertext_s0[38]}), .b ({signal_1910, signal_1199}), .c ({signal_2012, signal_1273}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1110 ( .a ({Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({signal_1914, signal_1201}), .c ({signal_2013, signal_1274}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1111 ( .a ({Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({signal_1912, signal_1200}), .c ({signal_2014, signal_1275}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1112 ( .a ({Ciphertext_s1[42], Ciphertext_s0[42]}), .b ({signal_1914, signal_1201}), .c ({signal_2015, signal_1276}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1113 ( .a ({Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({signal_1918, signal_1203}), .c ({signal_2016, signal_1277}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1114 ( .a ({Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({signal_1916, signal_1202}), .c ({signal_2017, signal_1278}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1115 ( .a ({Ciphertext_s1[46], Ciphertext_s0[46]}), .b ({signal_1918, signal_1203}), .c ({signal_2018, signal_1279}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1116 ( .a ({Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({signal_1922, signal_1205}), .c ({signal_2019, signal_1280}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1117 ( .a ({Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({signal_1920, signal_1204}), .c ({signal_2020, signal_1281}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1118 ( .a ({Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({signal_1922, signal_1205}), .c ({signal_2021, signal_1282}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1119 ( .a ({Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({signal_1926, signal_1207}), .c ({signal_2022, signal_1283}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1120 ( .a ({Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({signal_1924, signal_1206}), .c ({signal_2023, signal_1284}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1121 ( .a ({Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({signal_1926, signal_1207}), .c ({signal_2024, signal_1285}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1122 ( .a ({Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({signal_1930, signal_1209}), .c ({signal_2025, signal_1286}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1123 ( .a ({Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({signal_1928, signal_1208}), .c ({signal_2026, signal_1287}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1124 ( .a ({Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({signal_1930, signal_1209}), .c ({signal_2027, signal_1288}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1125 ( .a ({Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({signal_1934, signal_1211}), .c ({signal_2028, signal_1289}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1126 ( .a ({Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({signal_1932, signal_1210}), .c ({signal_2029, signal_1290}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1127 ( .a ({Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({signal_1934, signal_1211}), .c ({signal_2030, signal_1291}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1128 ( .a ({signal_1985, signal_1246}), .b ({signal_2031, signal_1292}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1129 ( .a ({signal_1988, signal_1249}), .b ({signal_2032, signal_1293}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1130 ( .a ({signal_1991, signal_1252}), .b ({signal_2033, signal_1294}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1131 ( .a ({signal_1994, signal_1255}), .b ({signal_2034, signal_1295}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1132 ( .a ({signal_1997, signal_1258}), .b ({signal_2035, signal_1296}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1133 ( .a ({signal_2000, signal_1261}), .b ({signal_2036, signal_1297}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1134 ( .a ({signal_2003, signal_1264}), .b ({signal_2037, signal_1298}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1135 ( .a ({signal_2006, signal_1267}), .b ({signal_2038, signal_1299}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1136 ( .a ({signal_2009, signal_1270}), .b ({signal_2039, signal_1300}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1137 ( .a ({signal_2012, signal_1273}), .b ({signal_2040, signal_1301}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1138 ( .a ({signal_2015, signal_1276}), .b ({signal_2041, signal_1302}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1139 ( .a ({signal_2018, signal_1279}), .b ({signal_2042, signal_1303}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1140 ( .a ({signal_2021, signal_1282}), .b ({signal_2043, signal_1304}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1141 ( .a ({signal_2024, signal_1285}), .b ({signal_2044, signal_1305}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1142 ( .a ({signal_2027, signal_1288}), .b ({signal_2045, signal_1306}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1143 ( .a ({signal_2030, signal_1291}), .b ({signal_2046, signal_1307}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1160 ( .a ({signal_1984, signal_1245}), .b ({signal_1985, signal_1246}), .c ({signal_2063, signal_1324}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1161 ( .a ({signal_1987, signal_1248}), .b ({signal_1988, signal_1249}), .c ({signal_2064, signal_1325}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1162 ( .a ({signal_1990, signal_1251}), .b ({signal_1991, signal_1252}), .c ({signal_2065, signal_1326}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1163 ( .a ({signal_1993, signal_1254}), .b ({signal_1994, signal_1255}), .c ({signal_2066, signal_1327}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1164 ( .a ({signal_1996, signal_1257}), .b ({signal_1997, signal_1258}), .c ({signal_2067, signal_1328}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1165 ( .a ({signal_1999, signal_1260}), .b ({signal_2000, signal_1261}), .c ({signal_2068, signal_1329}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1166 ( .a ({signal_2002, signal_1263}), .b ({signal_2003, signal_1264}), .c ({signal_2069, signal_1330}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1167 ( .a ({signal_2005, signal_1266}), .b ({signal_2006, signal_1267}), .c ({signal_2070, signal_1331}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1168 ( .a ({signal_2008, signal_1269}), .b ({signal_2009, signal_1270}), .c ({signal_2071, signal_1332}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1169 ( .a ({signal_2011, signal_1272}), .b ({signal_2012, signal_1273}), .c ({signal_2072, signal_1333}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1170 ( .a ({signal_2014, signal_1275}), .b ({signal_2015, signal_1276}), .c ({signal_2073, signal_1334}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1171 ( .a ({signal_2017, signal_1278}), .b ({signal_2018, signal_1279}), .c ({signal_2074, signal_1335}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1172 ( .a ({signal_2020, signal_1281}), .b ({signal_2021, signal_1282}), .c ({signal_2075, signal_1336}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1173 ( .a ({signal_2023, signal_1284}), .b ({signal_2024, signal_1285}), .c ({signal_2076, signal_1337}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1174 ( .a ({signal_2026, signal_1287}), .b ({signal_2027, signal_1288}), .c ({signal_2077, signal_1338}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1175 ( .a ({signal_2029, signal_1290}), .b ({signal_2030, signal_1291}), .c ({signal_2078, signal_1339}) ) ;
    ClockGatingController #(5) cell_1547 ( .clk (clk), .rst (rst), .GatedClk (signal_2642), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    mux2_masked #(.security_order(1), .pipeline(0)) cell_2 ( .s (rst), .b ({signal_2304, signal_837}), .a ({Plaintext_s1[2], Plaintext_s0[2]}), .c ({signal_2308, signal_901}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3 ( .s (rst), .b ({signal_2406, signal_836}), .a ({Plaintext_s1[3], Plaintext_s0[3]}), .c ({signal_2413, signal_900}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_6 ( .s (rst), .b ({signal_2305, signal_833}), .a ({Plaintext_s1[6], Plaintext_s0[6]}), .c ({signal_2310, signal_897}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_7 ( .s (rst), .b ({signal_2407, signal_832}), .a ({Plaintext_s1[7], Plaintext_s0[7]}), .c ({signal_2415, signal_896}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_10 ( .s (rst), .b ({signal_2306, signal_829}), .a ({Plaintext_s1[10], Plaintext_s0[10]}), .c ({signal_2312, signal_893}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_11 ( .s (rst), .b ({signal_2408, signal_828}), .a ({Plaintext_s1[11], Plaintext_s0[11]}), .c ({signal_2417, signal_892}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_14 ( .s (rst), .b ({signal_2411, signal_825}), .a ({Plaintext_s1[14], Plaintext_s0[14]}), .c ({signal_2419, signal_889}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_15 ( .s (rst), .b ({signal_2494, signal_824}), .a ({Plaintext_s1[15], Plaintext_s0[15]}), .c ({signal_2502, signal_888}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_18 ( .s (rst), .b ({signal_2301, signal_821}), .a ({Plaintext_s1[18], Plaintext_s0[18]}), .c ({signal_2314, signal_885}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_19 ( .s (rst), .b ({signal_2403, signal_820}), .a ({Plaintext_s1[19], Plaintext_s0[19]}), .c ({signal_2421, signal_884}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_22 ( .s (rst), .b ({signal_2302, signal_817}), .a ({Plaintext_s1[22], Plaintext_s0[22]}), .c ({signal_2316, signal_881}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_23 ( .s (rst), .b ({signal_2404, signal_816}), .a ({Plaintext_s1[23], Plaintext_s0[23]}), .c ({signal_2423, signal_880}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_26 ( .s (rst), .b ({signal_2410, signal_813}), .a ({Plaintext_s1[26], Plaintext_s0[26]}), .c ({signal_2425, signal_877}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_27 ( .s (rst), .b ({signal_2493, signal_812}), .a ({Plaintext_s1[27], Plaintext_s0[27]}), .c ({signal_2508, signal_876}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_30 ( .s (rst), .b ({signal_2303, signal_809}), .a ({Plaintext_s1[30], Plaintext_s0[30]}), .c ({signal_2318, signal_873}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_31 ( .s (rst), .b ({signal_2405, signal_808}), .a ({Plaintext_s1[31], Plaintext_s0[31]}), .c ({signal_2427, signal_872}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_34 ( .s (rst), .b ({signal_2211, signal_805}), .a ({Plaintext_s1[34], Plaintext_s0[34]}), .c ({signal_2251, signal_869}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_35 ( .s (rst), .b ({signal_2319, signal_804}), .a ({Plaintext_s1[35], Plaintext_s0[35]}), .c ({signal_2365, signal_868}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_38 ( .s (rst), .b ({signal_2212, signal_801}), .a ({Plaintext_s1[38], Plaintext_s0[38]}), .c ({signal_2253, signal_865}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_39 ( .s (rst), .b ({signal_2320, signal_800}), .a ({Plaintext_s1[39], Plaintext_s0[39]}), .c ({signal_2367, signal_864}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_42 ( .s (rst), .b ({signal_2213, signal_797}), .a ({Plaintext_s1[42], Plaintext_s0[42]}), .c ({signal_2255, signal_861}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_43 ( .s (rst), .b ({signal_2321, signal_796}), .a ({Plaintext_s1[43], Plaintext_s0[43]}), .c ({signal_2369, signal_860}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_46 ( .s (rst), .b ({signal_2322, signal_793}), .a ({Plaintext_s1[46], Plaintext_s0[46]}), .c ({signal_2371, signal_857}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_47 ( .s (rst), .b ({signal_2434, signal_792}), .a ({Plaintext_s1[47], Plaintext_s0[47]}), .c ({signal_2464, signal_856}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_50 ( .s (rst), .b ({signal_2323, signal_789}), .a ({Plaintext_s1[50], Plaintext_s0[50]}), .c ({signal_2373, signal_853}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_51 ( .s (rst), .b ({signal_2435, signal_788}), .a ({Plaintext_s1[51], Plaintext_s0[51]}), .c ({signal_2466, signal_852}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_54 ( .s (rst), .b ({signal_2324, signal_785}), .a ({Plaintext_s1[54], Plaintext_s0[54]}), .c ({signal_2375, signal_849}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_55 ( .s (rst), .b ({signal_2436, signal_784}), .a ({Plaintext_s1[55], Plaintext_s0[55]}), .c ({signal_2468, signal_848}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_58 ( .s (rst), .b ({signal_2325, signal_781}), .a ({Plaintext_s1[58], Plaintext_s0[58]}), .c ({signal_2377, signal_845}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_59 ( .s (rst), .b ({signal_2437, signal_780}), .a ({Plaintext_s1[59], Plaintext_s0[59]}), .c ({signal_2470, signal_844}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_62 ( .s (rst), .b ({signal_2438, signal_777}), .a ({Plaintext_s1[62], Plaintext_s0[62]}), .c ({signal_2472, signal_841}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_63 ( .s (rst), .b ({signal_2519, signal_776}), .a ({Plaintext_s1[63], Plaintext_s0[63]}), .c ({signal_2548, signal_840}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1064 ( .a ({signal_1840, signal_1164}), .b ({signal_1936, signal_1212}), .clk (clk), .r (Fresh[0]), .c ({signal_1967, signal_1228}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1065 ( .a ({signal_1842, signal_1165}), .b ({signal_1938, signal_1213}), .clk (clk), .r (Fresh[1]), .c ({signal_1968, signal_1229}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1066 ( .a ({signal_1844, signal_1166}), .b ({signal_1940, signal_1214}), .clk (clk), .r (Fresh[2]), .c ({signal_1969, signal_1230}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1067 ( .a ({signal_1846, signal_1167}), .b ({signal_1942, signal_1215}), .clk (clk), .r (Fresh[3]), .c ({signal_1970, signal_1231}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1068 ( .a ({signal_1848, signal_1168}), .b ({signal_1944, signal_1216}), .clk (clk), .r (Fresh[4]), .c ({signal_1971, signal_1232}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1069 ( .a ({signal_1850, signal_1169}), .b ({signal_1946, signal_1217}), .clk (clk), .r (Fresh[5]), .c ({signal_1972, signal_1233}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1070 ( .a ({signal_1852, signal_1170}), .b ({signal_1948, signal_1218}), .clk (clk), .r (Fresh[6]), .c ({signal_1973, signal_1234}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1071 ( .a ({signal_1854, signal_1171}), .b ({signal_1950, signal_1219}), .clk (clk), .r (Fresh[7]), .c ({signal_1974, signal_1235}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1072 ( .a ({signal_1856, signal_1172}), .b ({signal_1952, signal_1220}), .clk (clk), .r (Fresh[8]), .c ({signal_1975, signal_1236}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1073 ( .a ({signal_1858, signal_1173}), .b ({signal_1954, signal_1221}), .clk (clk), .r (Fresh[9]), .c ({signal_1976, signal_1237}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1074 ( .a ({signal_1860, signal_1174}), .b ({signal_1956, signal_1222}), .clk (clk), .r (Fresh[10]), .c ({signal_1977, signal_1238}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1075 ( .a ({signal_1862, signal_1175}), .b ({signal_1958, signal_1223}), .clk (clk), .r (Fresh[11]), .c ({signal_1978, signal_1239}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1076 ( .a ({signal_1864, signal_1176}), .b ({signal_1960, signal_1224}), .clk (clk), .r (Fresh[12]), .c ({signal_1979, signal_1240}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1077 ( .a ({signal_1866, signal_1177}), .b ({signal_1962, signal_1225}), .clk (clk), .r (Fresh[13]), .c ({signal_1980, signal_1241}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1078 ( .a ({signal_1868, signal_1178}), .b ({signal_1964, signal_1226}), .clk (clk), .r (Fresh[14]), .c ({signal_1981, signal_1242}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1079 ( .a ({signal_1870, signal_1179}), .b ({signal_1966, signal_1227}), .clk (clk), .r (Fresh[15]), .c ({signal_1982, signal_1243}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1144 ( .a ({signal_1840, signal_1164}), .b ({signal_1984, signal_1245}), .clk (clk), .r (Fresh[16]), .c ({signal_2047, signal_1308}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1145 ( .a ({signal_1842, signal_1165}), .b ({signal_1987, signal_1248}), .clk (clk), .r (Fresh[17]), .c ({signal_2048, signal_1309}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1146 ( .a ({signal_1844, signal_1166}), .b ({signal_1990, signal_1251}), .clk (clk), .r (Fresh[18]), .c ({signal_2049, signal_1310}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1147 ( .a ({signal_1846, signal_1167}), .b ({signal_1993, signal_1254}), .clk (clk), .r (Fresh[19]), .c ({signal_2050, signal_1311}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1148 ( .a ({signal_1848, signal_1168}), .b ({signal_1996, signal_1257}), .clk (clk), .r (Fresh[20]), .c ({signal_2051, signal_1312}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1149 ( .a ({signal_1850, signal_1169}), .b ({signal_1999, signal_1260}), .clk (clk), .r (Fresh[21]), .c ({signal_2052, signal_1313}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1150 ( .a ({signal_1852, signal_1170}), .b ({signal_2002, signal_1263}), .clk (clk), .r (Fresh[22]), .c ({signal_2053, signal_1314}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1151 ( .a ({signal_1854, signal_1171}), .b ({signal_2005, signal_1266}), .clk (clk), .r (Fresh[23]), .c ({signal_2054, signal_1315}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1152 ( .a ({signal_1856, signal_1172}), .b ({signal_2008, signal_1269}), .clk (clk), .r (Fresh[24]), .c ({signal_2055, signal_1316}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1153 ( .a ({signal_1858, signal_1173}), .b ({signal_2011, signal_1272}), .clk (clk), .r (Fresh[25]), .c ({signal_2056, signal_1317}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1154 ( .a ({signal_1860, signal_1174}), .b ({signal_2014, signal_1275}), .clk (clk), .r (Fresh[26]), .c ({signal_2057, signal_1318}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1155 ( .a ({signal_1862, signal_1175}), .b ({signal_2017, signal_1278}), .clk (clk), .r (Fresh[27]), .c ({signal_2058, signal_1319}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1156 ( .a ({signal_1864, signal_1176}), .b ({signal_2020, signal_1281}), .clk (clk), .r (Fresh[28]), .c ({signal_2059, signal_1320}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1157 ( .a ({signal_1866, signal_1177}), .b ({signal_2023, signal_1284}), .clk (clk), .r (Fresh[29]), .c ({signal_2060, signal_1321}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1158 ( .a ({signal_1868, signal_1178}), .b ({signal_2026, signal_1287}), .clk (clk), .r (Fresh[30]), .c ({signal_2061, signal_1322}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1159 ( .a ({signal_1870, signal_1179}), .b ({signal_2029, signal_1290}), .clk (clk), .r (Fresh[31]), .c ({signal_2062, signal_1323}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1176 ( .a ({signal_1872, signal_1180}), .b ({signal_1967, signal_1228}), .c ({signal_2079, signal_1340}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1177 ( .a ({signal_1876, signal_1182}), .b ({signal_1968, signal_1229}), .c ({signal_2080, signal_1341}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1178 ( .a ({signal_1880, signal_1184}), .b ({signal_1969, signal_1230}), .c ({signal_2081, signal_1342}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1179 ( .a ({signal_1884, signal_1186}), .b ({signal_1970, signal_1231}), .c ({signal_2082, signal_1343}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1180 ( .a ({signal_1888, signal_1188}), .b ({signal_1971, signal_1232}), .c ({signal_2083, signal_1344}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1181 ( .a ({signal_1892, signal_1190}), .b ({signal_1972, signal_1233}), .c ({signal_2084, signal_1345}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1182 ( .a ({signal_1896, signal_1192}), .b ({signal_1973, signal_1234}), .c ({signal_2085, signal_1346}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1183 ( .a ({signal_1900, signal_1194}), .b ({signal_1974, signal_1235}), .c ({signal_2086, signal_1347}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1184 ( .a ({signal_1904, signal_1196}), .b ({signal_1975, signal_1236}), .c ({signal_2087, signal_1348}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1185 ( .a ({signal_1908, signal_1198}), .b ({signal_1976, signal_1237}), .c ({signal_2088, signal_1349}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1186 ( .a ({signal_1912, signal_1200}), .b ({signal_1977, signal_1238}), .c ({signal_2089, signal_1350}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1187 ( .a ({signal_1916, signal_1202}), .b ({signal_1978, signal_1239}), .c ({signal_2090, signal_1351}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1188 ( .a ({signal_1920, signal_1204}), .b ({signal_1979, signal_1240}), .c ({signal_2091, signal_1352}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1189 ( .a ({signal_1924, signal_1206}), .b ({signal_1980, signal_1241}), .c ({signal_2092, signal_1353}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1190 ( .a ({signal_1928, signal_1208}), .b ({signal_1981, signal_1242}), .c ({signal_2093, signal_1354}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1191 ( .a ({signal_1932, signal_1210}), .b ({signal_1982, signal_1243}), .c ({signal_2094, signal_1355}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1192 ( .a ({signal_1983, signal_1244}), .b ({signal_2047, signal_1308}), .c ({signal_2095, signal_1356}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1193 ( .a ({signal_1967, signal_1228}), .b ({signal_2063, signal_1324}), .c ({signal_2096, signal_1357}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1194 ( .a ({signal_1874, signal_1181}), .b ({signal_2047, signal_1308}), .c ({signal_2097, signal_1358}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1195 ( .a ({signal_1986, signal_1247}), .b ({signal_2048, signal_1309}), .c ({signal_2098, signal_1359}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1196 ( .a ({signal_1968, signal_1229}), .b ({signal_2064, signal_1325}), .c ({signal_2099, signal_1360}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1197 ( .a ({signal_1878, signal_1183}), .b ({signal_2048, signal_1309}), .c ({signal_2100, signal_1361}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1198 ( .a ({signal_1989, signal_1250}), .b ({signal_2049, signal_1310}), .c ({signal_2101, signal_1362}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1199 ( .a ({signal_1969, signal_1230}), .b ({signal_2065, signal_1326}), .c ({signal_2102, signal_1363}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1200 ( .a ({signal_1882, signal_1185}), .b ({signal_2049, signal_1310}), .c ({signal_2103, signal_1364}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1201 ( .a ({signal_1992, signal_1253}), .b ({signal_2050, signal_1311}), .c ({signal_2104, signal_1365}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1202 ( .a ({signal_1970, signal_1231}), .b ({signal_2066, signal_1327}), .c ({signal_2105, signal_1366}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1203 ( .a ({signal_1886, signal_1187}), .b ({signal_2050, signal_1311}), .c ({signal_2106, signal_1367}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1204 ( .a ({signal_1995, signal_1256}), .b ({signal_2051, signal_1312}), .c ({signal_2107, signal_1368}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1205 ( .a ({signal_1971, signal_1232}), .b ({signal_2067, signal_1328}), .c ({signal_2108, signal_1369}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1206 ( .a ({signal_1890, signal_1189}), .b ({signal_2051, signal_1312}), .c ({signal_2109, signal_1370}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1207 ( .a ({signal_1998, signal_1259}), .b ({signal_2052, signal_1313}), .c ({signal_2110, signal_1371}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1208 ( .a ({signal_1972, signal_1233}), .b ({signal_2068, signal_1329}), .c ({signal_2111, signal_1372}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1209 ( .a ({signal_1894, signal_1191}), .b ({signal_2052, signal_1313}), .c ({signal_2112, signal_1373}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1210 ( .a ({signal_2001, signal_1262}), .b ({signal_2053, signal_1314}), .c ({signal_2113, signal_1374}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1211 ( .a ({signal_1973, signal_1234}), .b ({signal_2069, signal_1330}), .c ({signal_2114, signal_1375}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1212 ( .a ({signal_1898, signal_1193}), .b ({signal_2053, signal_1314}), .c ({signal_2115, signal_1376}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1213 ( .a ({signal_2004, signal_1265}), .b ({signal_2054, signal_1315}), .c ({signal_2116, signal_1377}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1214 ( .a ({signal_1974, signal_1235}), .b ({signal_2070, signal_1331}), .c ({signal_2117, signal_1378}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1215 ( .a ({signal_1902, signal_1195}), .b ({signal_2054, signal_1315}), .c ({signal_2118, signal_1379}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1216 ( .a ({signal_2007, signal_1268}), .b ({signal_2055, signal_1316}), .c ({signal_2119, signal_1380}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1217 ( .a ({signal_1975, signal_1236}), .b ({signal_2071, signal_1332}), .c ({signal_2120, signal_1381}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1218 ( .a ({signal_1906, signal_1197}), .b ({signal_2055, signal_1316}), .c ({signal_2121, signal_1382}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1219 ( .a ({signal_2010, signal_1271}), .b ({signal_2056, signal_1317}), .c ({signal_2122, signal_1383}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1220 ( .a ({signal_1976, signal_1237}), .b ({signal_2072, signal_1333}), .c ({signal_2123, signal_1384}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1221 ( .a ({signal_1910, signal_1199}), .b ({signal_2056, signal_1317}), .c ({signal_2124, signal_1385}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1222 ( .a ({signal_2013, signal_1274}), .b ({signal_2057, signal_1318}), .c ({signal_2125, signal_1386}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1223 ( .a ({signal_1977, signal_1238}), .b ({signal_2073, signal_1334}), .c ({signal_2126, signal_1387}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1224 ( .a ({signal_1914, signal_1201}), .b ({signal_2057, signal_1318}), .c ({signal_2127, signal_1388}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1225 ( .a ({signal_2016, signal_1277}), .b ({signal_2058, signal_1319}), .c ({signal_2128, signal_1389}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1226 ( .a ({signal_1978, signal_1239}), .b ({signal_2074, signal_1335}), .c ({signal_2129, signal_1390}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1227 ( .a ({signal_1918, signal_1203}), .b ({signal_2058, signal_1319}), .c ({signal_2130, signal_1391}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1228 ( .a ({signal_2019, signal_1280}), .b ({signal_2059, signal_1320}), .c ({signal_2131, signal_1392}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1229 ( .a ({signal_1979, signal_1240}), .b ({signal_2075, signal_1336}), .c ({signal_2132, signal_1393}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1230 ( .a ({signal_1922, signal_1205}), .b ({signal_2059, signal_1320}), .c ({signal_2133, signal_1394}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1231 ( .a ({signal_2022, signal_1283}), .b ({signal_2060, signal_1321}), .c ({signal_2134, signal_1395}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1232 ( .a ({signal_1980, signal_1241}), .b ({signal_2076, signal_1337}), .c ({signal_2135, signal_1396}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1233 ( .a ({signal_1926, signal_1207}), .b ({signal_2060, signal_1321}), .c ({signal_2136, signal_1397}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1234 ( .a ({signal_2025, signal_1286}), .b ({signal_2061, signal_1322}), .c ({signal_2137, signal_1398}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1235 ( .a ({signal_1981, signal_1242}), .b ({signal_2077, signal_1338}), .c ({signal_2138, signal_1399}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1236 ( .a ({signal_1930, signal_1209}), .b ({signal_2061, signal_1322}), .c ({signal_2139, signal_1400}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1237 ( .a ({signal_2028, signal_1289}), .b ({signal_2062, signal_1323}), .c ({signal_2140, signal_1401}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1238 ( .a ({signal_1982, signal_1243}), .b ({signal_2078, signal_1339}), .c ({signal_2141, signal_1402}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1239 ( .a ({signal_1934, signal_1211}), .b ({signal_2062, signal_1323}), .c ({signal_2142, signal_1403}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1240 ( .a ({1'b0, 1'b0}), .b ({signal_2094, signal_1355}), .c ({signal_2143, signal_1404}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1241 ( .a ({1'b0, 1'b0}), .b ({signal_2090, signal_1351}), .c ({signal_2144, signal_1405}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1242 ( .a ({1'b0, 1'b0}), .b ({signal_2087, signal_1348}), .c ({signal_2145, signal_1406}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1243 ( .a ({1'b0, 1'b0}), .b ({signal_2088, signal_1349}), .c ({signal_2146, signal_1407}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1244 ( .a ({1'b0, 1'b0}), .b ({signal_2089, signal_1350}), .c ({signal_2147, signal_1408}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1245 ( .a ({1'b0, 1'b0}), .b ({signal_2091, signal_1352}), .c ({signal_2148, signal_1409}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1246 ( .a ({1'b0, 1'b0}), .b ({signal_2092, signal_1353}), .c ({signal_2149, signal_1410}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1247 ( .a ({1'b0, 1'b0}), .b ({signal_2093, signal_1354}), .c ({signal_2150, signal_1411}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1248 ( .a ({signal_2082, signal_1343}), .b ({signal_2085, signal_1346}), .c ({signal_2151, signal_1412}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1249 ( .a ({signal_2079, signal_1340}), .b ({signal_2086, signal_1347}), .c ({signal_2152, signal_1413}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1250 ( .a ({signal_2080, signal_1341}), .b ({signal_2083, signal_1344}), .c ({signal_2153, signal_1414}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1251 ( .a ({signal_2081, signal_1342}), .b ({signal_2084, signal_1345}), .c ({signal_2154, signal_1415}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1284 ( .a ({signal_1967, signal_1228}), .b ({signal_2097, signal_1358}), .c ({signal_2187, signal_1448}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1285 ( .a ({signal_1968, signal_1229}), .b ({signal_2100, signal_1361}), .c ({signal_2188, signal_1449}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1286 ( .a ({signal_1969, signal_1230}), .b ({signal_2103, signal_1364}), .c ({signal_2189, signal_1450}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1287 ( .a ({signal_1970, signal_1231}), .b ({signal_2106, signal_1367}), .c ({signal_2190, signal_1451}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1288 ( .a ({signal_1971, signal_1232}), .b ({signal_2109, signal_1370}), .c ({signal_2191, signal_1452}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1289 ( .a ({signal_1972, signal_1233}), .b ({signal_2112, signal_1373}), .c ({signal_2192, signal_1453}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1290 ( .a ({signal_1973, signal_1234}), .b ({signal_2115, signal_1376}), .c ({signal_2193, signal_1454}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1291 ( .a ({signal_1974, signal_1235}), .b ({signal_2118, signal_1379}), .c ({signal_2194, signal_1455}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1292 ( .a ({signal_1975, signal_1236}), .b ({signal_2121, signal_1382}), .c ({signal_2195, signal_1456}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1293 ( .a ({signal_1976, signal_1237}), .b ({signal_2124, signal_1385}), .c ({signal_2196, signal_1457}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1294 ( .a ({signal_1977, signal_1238}), .b ({signal_2127, signal_1388}), .c ({signal_2197, signal_1458}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1295 ( .a ({signal_1978, signal_1239}), .b ({signal_2130, signal_1391}), .c ({signal_2198, signal_1459}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1296 ( .a ({signal_1979, signal_1240}), .b ({signal_2133, signal_1394}), .c ({signal_2199, signal_1460}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1297 ( .a ({signal_1980, signal_1241}), .b ({signal_2136, signal_1397}), .c ({signal_2200, signal_1461}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1298 ( .a ({signal_1981, signal_1242}), .b ({signal_2139, signal_1400}), .c ({signal_2201, signal_1462}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1299 ( .a ({signal_1982, signal_1243}), .b ({signal_2142, signal_1403}), .c ({signal_2202, signal_1463}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1300 ( .a ({1'b0, signal_1026}), .b ({signal_2143, signal_1404}), .c ({signal_2203, signal_1464}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1301 ( .a ({1'b0, 1'b0}), .b ({signal_2144, signal_1405}), .c ({signal_2204, signal_1465}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1302 ( .a ({signal_1653, signal_1161}), .b ({signal_2145, signal_1406}), .c ({signal_2205, signal_1466}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1303 ( .a ({signal_1665, signal_1157}), .b ({signal_2146, signal_1407}), .c ({signal_2206, signal_1467}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1304 ( .a ({signal_1677, signal_1153}), .b ({signal_2147, signal_1408}), .c ({signal_2207, signal_1468}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1305 ( .a ({signal_1701, signal_1145}), .b ({signal_2148, signal_1409}), .c ({signal_2208, signal_1469}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1306 ( .a ({signal_1713, signal_1141}), .b ({signal_2149, signal_1410}), .c ({signal_2209, signal_1470}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1307 ( .a ({signal_1725, signal_1137}), .b ({signal_2150, signal_1411}), .c ({signal_2210, signal_1471}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1308 ( .a ({signal_2208, signal_1469}), .b ({signal_2211, signal_805}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1309 ( .a ({signal_2209, signal_1470}), .b ({signal_2212, signal_801}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1310 ( .a ({signal_2210, signal_1471}), .b ({signal_2213, signal_797}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1327 ( .a ({1'b0, 1'b0}), .b ({signal_2202, signal_1463}), .c ({signal_2230, signal_1488}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1328 ( .a ({1'b0, 1'b0}), .b ({signal_2198, signal_1459}), .c ({signal_2231, signal_1489}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1329 ( .a ({1'b0, 1'b0}), .b ({signal_2195, signal_1456}), .c ({signal_2232, signal_1490}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1330 ( .a ({1'b0, 1'b0}), .b ({signal_2196, signal_1457}), .c ({signal_2233, signal_1491}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1331 ( .a ({1'b0, 1'b0}), .b ({signal_2197, signal_1458}), .c ({signal_2234, signal_1492}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1332 ( .a ({1'b0, 1'b0}), .b ({signal_2199, signal_1460}), .c ({signal_2235, signal_1493}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1333 ( .a ({1'b0, 1'b0}), .b ({signal_2200, signal_1461}), .c ({signal_2236, signal_1494}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1334 ( .a ({1'b0, 1'b0}), .b ({signal_2201, signal_1462}), .c ({signal_2237, signal_1495}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1335 ( .a ({signal_2190, signal_1451}), .b ({signal_2193, signal_1454}), .c ({signal_2238, signal_1496}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1336 ( .a ({signal_2187, signal_1448}), .b ({signal_2194, signal_1455}), .c ({signal_2239, signal_1497}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1337 ( .a ({signal_2188, signal_1449}), .b ({signal_2191, signal_1452}), .c ({signal_2240, signal_1498}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1338 ( .a ({signal_2189, signal_1450}), .b ({signal_2192, signal_1453}), .c ({signal_2241, signal_1499}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1339 ( .a ({1'b0, 1'b0}), .b ({signal_2204, signal_1465}), .c ({signal_2242, signal_1500}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1340 ( .a ({1'b0, 1'b0}), .b ({signal_2203, signal_1464}), .c ({signal_2243, signal_1501}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1341 ( .a ({1'b0, 1'b0}), .b ({signal_2208, signal_1469}), .c ({signal_2244, signal_1502}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1342 ( .a ({1'b0, 1'b0}), .b ({signal_2209, signal_1470}), .c ({signal_2245, signal_1503}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1343 ( .a ({1'b0, 1'b0}), .b ({signal_2210, signal_1471}), .c ({signal_2246, signal_1504}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1344 ( .a ({1'b0, 1'b0}), .b ({signal_2206, signal_1467}), .c ({signal_2247, signal_1505}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1345 ( .a ({1'b0, 1'b0}), .b ({signal_2207, signal_1468}), .c ({signal_2248, signal_1506}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1346 ( .a ({1'b0, 1'b0}), .b ({signal_2205, signal_1466}), .c ({signal_2249, signal_1507}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1379 ( .a ({1'b0, signal_1025}), .b ({signal_2230, signal_1488}), .c ({signal_2288, signal_1540}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1380 ( .a ({1'b0, 1'b0}), .b ({signal_2231, signal_1489}), .c ({signal_2289, signal_1541}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1381 ( .a ({signal_1656, signal_1160}), .b ({signal_2232, signal_1490}), .c ({signal_2290, signal_1542}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1382 ( .a ({signal_1668, signal_1156}), .b ({signal_2233, signal_1491}), .c ({signal_2291, signal_1543}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1383 ( .a ({signal_1680, signal_1152}), .b ({signal_2234, signal_1492}), .c ({signal_2292, signal_1544}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1384 ( .a ({signal_1704, signal_1144}), .b ({signal_2235, signal_1493}), .c ({signal_2293, signal_1545}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1385 ( .a ({signal_1716, signal_1140}), .b ({signal_2236, signal_1494}), .c ({signal_2294, signal_1546}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1386 ( .a ({signal_1728, signal_1136}), .b ({signal_2237, signal_1495}), .c ({signal_2295, signal_1547}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1387 ( .a ({signal_1689, signal_1149}), .b ({signal_2242, signal_1500}), .c ({signal_2296, signal_1548}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1388 ( .a ({signal_1737, signal_1133}), .b ({signal_2243, signal_1501}), .c ({signal_2297, signal_1549}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1389 ( .a ({signal_2151, signal_1412}), .b ({signal_2244, signal_1502}), .c ({signal_2298, signal_1550}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1390 ( .a ({signal_2152, signal_1413}), .b ({signal_2245, signal_1503}), .c ({signal_2299, signal_1551}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1391 ( .a ({signal_2153, signal_1414}), .b ({signal_2246, signal_1504}), .c ({signal_2300, signal_1552}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1392 ( .a ({signal_2085, signal_1346}), .b ({signal_2247, signal_1505}), .c ({signal_2301, signal_821}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1393 ( .a ({signal_2086, signal_1347}), .b ({signal_2248, signal_1506}), .c ({signal_2302, signal_817}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1394 ( .a ({signal_2084, signal_1345}), .b ({signal_2249, signal_1507}), .c ({signal_2303, signal_809}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1395 ( .a ({signal_2085, signal_1346}), .b ({signal_2244, signal_1502}), .c ({signal_2304, signal_837}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1396 ( .a ({signal_2086, signal_1347}), .b ({signal_2245, signal_1503}), .c ({signal_2305, signal_833}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1397 ( .a ({signal_2083, signal_1344}), .b ({signal_2246, signal_1504}), .c ({signal_2306, signal_829}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1398 ( .a ({signal_2293, signal_1545}), .b ({signal_2319, signal_804}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1399 ( .a ({signal_2294, signal_1546}), .b ({signal_2320, signal_800}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1400 ( .a ({signal_2295, signal_1547}), .b ({signal_2321, signal_796}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1401 ( .a ({signal_2297, signal_1549}), .b ({signal_2322, signal_793}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1402 ( .a ({signal_2298, signal_1550}), .b ({signal_2323, signal_789}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1403 ( .a ({signal_2299, signal_1551}), .b ({signal_2324, signal_785}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1404 ( .a ({signal_2300, signal_1552}), .b ({signal_2325, signal_781}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1433 ( .a ({1'b0, 1'b0}), .b ({signal_2289, signal_1541}), .c ({signal_2354, signal_1581}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1434 ( .a ({1'b0, 1'b0}), .b ({signal_2288, signal_1540}), .c ({signal_2355, signal_1582}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1435 ( .a ({1'b0, 1'b0}), .b ({signal_2293, signal_1545}), .c ({signal_2356, signal_1583}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1436 ( .a ({1'b0, 1'b0}), .b ({signal_2294, signal_1546}), .c ({signal_2357, signal_1584}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1437 ( .a ({1'b0, 1'b0}), .b ({signal_2295, signal_1547}), .c ({signal_2358, signal_1585}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1438 ( .a ({1'b0, 1'b0}), .b ({signal_2291, signal_1543}), .c ({signal_2359, signal_1586}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1439 ( .a ({1'b0, 1'b0}), .b ({signal_2292, signal_1544}), .c ({signal_2360, signal_1587}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1440 ( .a ({1'b0, 1'b0}), .b ({signal_2290, signal_1542}), .c ({signal_2361, signal_1588}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1441 ( .a ({1'b0, 1'b0}), .b ({signal_2297, signal_1549}), .c ({signal_2362, signal_1589}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1442 ( .a ({1'b0, 1'b0}), .b ({signal_2296, signal_1548}), .c ({signal_2363, signal_1590}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1462 ( .a ({signal_1692, signal_1148}), .b ({signal_2354, signal_1581}), .c ({signal_2397, signal_1607}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1463 ( .a ({signal_1740, signal_1132}), .b ({signal_2355, signal_1582}), .c ({signal_2398, signal_1608}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1464 ( .a ({signal_2238, signal_1496}), .b ({signal_2356, signal_1583}), .c ({signal_2399, signal_1609}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1466 ( .a ({signal_2239, signal_1497}), .b ({signal_2357, signal_1584}), .c ({signal_2401, signal_1611}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1467 ( .a ({signal_2240, signal_1498}), .b ({signal_2358, signal_1585}), .c ({signal_2402, signal_1612}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1468 ( .a ({signal_2193, signal_1454}), .b ({signal_2359, signal_1586}), .c ({signal_2403, signal_820}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1469 ( .a ({signal_2194, signal_1455}), .b ({signal_2360, signal_1587}), .c ({signal_2404, signal_816}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1470 ( .a ({signal_2192, signal_1453}), .b ({signal_2361, signal_1588}), .c ({signal_2405, signal_808}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1471 ( .a ({signal_2193, signal_1454}), .b ({signal_2356, signal_1583}), .c ({signal_2406, signal_836}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1472 ( .a ({signal_2194, signal_1455}), .b ({signal_2357, signal_1584}), .c ({signal_2407, signal_832}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1473 ( .a ({signal_2191, signal_1452}), .b ({signal_2358, signal_1585}), .c ({signal_2408, signal_828}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1474 ( .a ({signal_2154, signal_1415}), .b ({signal_2362, signal_1589}), .c ({signal_2409, signal_1613}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1475 ( .a ({signal_2083, signal_1344}), .b ({signal_2363, signal_1590}), .c ({signal_2410, signal_813}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1476 ( .a ({signal_2084, signal_1345}), .b ({signal_2362, signal_1589}), .c ({signal_2411, signal_825}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1477 ( .a ({signal_2398, signal_1608}), .b ({signal_2434, signal_792}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1478 ( .a ({signal_2399, signal_1609}), .b ({signal_2435, signal_788}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1479 ( .a ({signal_2401, signal_1611}), .b ({signal_2436, signal_784}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1480 ( .a ({signal_2402, signal_1612}), .b ({signal_2437, signal_780}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1481 ( .a ({signal_2409, signal_1613}), .b ({signal_2438, signal_777}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1498 ( .a ({1'b0, 1'b0}), .b ({signal_2398, signal_1608}), .c ({signal_2455, signal_1627}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1499 ( .a ({1'b0, 1'b0}), .b ({signal_2397, signal_1607}), .c ({signal_2456, signal_1628}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1519 ( .a ({signal_2241, signal_1499}), .b ({signal_2455, signal_1627}), .c ({signal_2492, signal_1638}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1520 ( .a ({signal_2191, signal_1452}), .b ({signal_2456, signal_1628}), .c ({signal_2493, signal_812}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1521 ( .a ({signal_2192, signal_1453}), .b ({signal_2455, signal_1627}), .c ({signal_2494, signal_824}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1522 ( .a ({signal_2492, signal_1638}), .b ({signal_2519, signal_776}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    mux2_masked #(.security_order(1), .pipeline(0)) cell_0 ( .s (rst), .b ({signal_2489, signal_839}), .a ({Plaintext_s1[0], Plaintext_s0[0]}), .c ({signal_2496, signal_903}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1 ( .s (rst), .b ({signal_2530, signal_838}), .a ({Plaintext_s1[1], Plaintext_s0[1]}), .c ({signal_2534, signal_902}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_4 ( .s (rst), .b ({signal_2490, signal_835}), .a ({Plaintext_s1[4], Plaintext_s0[4]}), .c ({signal_2498, signal_899}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_5 ( .s (rst), .b ({signal_2551, signal_834}), .a ({Plaintext_s1[5], Plaintext_s0[5]}), .c ({signal_2558, signal_898}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_8 ( .s (rst), .b ({signal_2491, signal_831}), .a ({Plaintext_s1[8], Plaintext_s0[8]}), .c ({signal_2500, signal_895}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_9 ( .s (rst), .b ({signal_2532, signal_830}), .a ({Plaintext_s1[9], Plaintext_s0[9]}), .c ({signal_2536, signal_894}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_12 ( .s (rst), .b ({signal_2556, signal_827}), .a ({Plaintext_s1[12], Plaintext_s0[12]}), .c ({signal_2560, signal_891}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_13 ( .s (rst), .b ({signal_2571, signal_826}), .a ({Plaintext_s1[13], Plaintext_s0[13]}), .c ({signal_2573, signal_890}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_16 ( .s (rst), .b ({signal_2483, signal_823}), .a ({Plaintext_s1[16], Plaintext_s0[16]}), .c ({signal_2504, signal_887}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_17 ( .s (rst), .b ({signal_2526, signal_822}), .a ({Plaintext_s1[17], Plaintext_s0[17]}), .c ({signal_2538, signal_886}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_20 ( .s (rst), .b ({signal_2485, signal_819}), .a ({Plaintext_s1[20], Plaintext_s0[20]}), .c ({signal_2506, signal_883}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_21 ( .s (rst), .b ({signal_2550, signal_818}), .a ({Plaintext_s1[21], Plaintext_s0[21]}), .c ({signal_2562, signal_882}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_24 ( .s (rst), .b ({signal_2554, signal_815}), .a ({Plaintext_s1[24], Plaintext_s0[24]}), .c ({signal_2564, signal_879}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_25 ( .s (rst), .b ({signal_2570, signal_814}), .a ({Plaintext_s1[25], Plaintext_s0[25]}), .c ({signal_2575, signal_878}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_28 ( .s (rst), .b ({signal_2487, signal_811}), .a ({Plaintext_s1[28], Plaintext_s0[28]}), .c ({signal_2510, signal_875}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_29 ( .s (rst), .b ({signal_2529, signal_810}), .a ({Plaintext_s1[29], Plaintext_s0[29]}), .c ({signal_2540, signal_874}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_32 ( .s (rst), .b ({signal_2388, signal_807}), .a ({Plaintext_s1[32], Plaintext_s0[32]}), .c ({signal_2429, signal_871}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_33 ( .s (rst), .b ({signal_2445, signal_806}), .a ({Plaintext_s1[33], Plaintext_s0[33]}), .c ({signal_2458, signal_870}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_36 ( .s (rst), .b ({signal_2390, signal_803}), .a ({Plaintext_s1[36], Plaintext_s0[36]}), .c ({signal_2431, signal_867}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_37 ( .s (rst), .b ({signal_2446, signal_802}), .a ({Plaintext_s1[37], Plaintext_s0[37]}), .c ({signal_2460, signal_866}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_40 ( .s (rst), .b ({signal_2392, signal_799}), .a ({Plaintext_s1[40], Plaintext_s0[40]}), .c ({signal_2433, signal_863}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_41 ( .s (rst), .b ({signal_2447, signal_798}), .a ({Plaintext_s1[41], Plaintext_s0[41]}), .c ({signal_2462, signal_862}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_44 ( .s (rst), .b ({signal_2475, signal_795}), .a ({Plaintext_s1[44], Plaintext_s0[44]}), .c ({signal_2512, signal_859}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_45 ( .s (rst), .b ({signal_2521, signal_794}), .a ({Plaintext_s1[45], Plaintext_s0[45]}), .c ({signal_2542, signal_858}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_48 ( .s (rst), .b ({signal_2477, signal_791}), .a ({Plaintext_s1[48], Plaintext_s0[48]}), .c ({signal_2514, signal_855}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_49 ( .s (rst), .b ({signal_2522, signal_790}), .a ({Plaintext_s1[49], Plaintext_s0[49]}), .c ({signal_2544, signal_854}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_52 ( .s (rst), .b ({signal_2479, signal_787}), .a ({Plaintext_s1[52], Plaintext_s0[52]}), .c ({signal_2516, signal_851}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_53 ( .s (rst), .b ({signal_2549, signal_786}), .a ({Plaintext_s1[53], Plaintext_s0[53]}), .c ({signal_2566, signal_850}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_56 ( .s (rst), .b ({signal_2481, signal_783}), .a ({Plaintext_s1[56], Plaintext_s0[56]}), .c ({signal_2518, signal_847}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_57 ( .s (rst), .b ({signal_2524, signal_782}), .a ({Plaintext_s1[57], Plaintext_s0[57]}), .c ({signal_2546, signal_846}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_60 ( .s (rst), .b ({signal_2552, signal_779}), .a ({Plaintext_s1[60], Plaintext_s0[60]}), .c ({signal_2568, signal_843}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_61 ( .s (rst), .b ({signal_2569, signal_778}), .a ({Plaintext_s1[61], Plaintext_s0[61]}), .c ({signal_2577, signal_842}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1252 ( .a ({Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({signal_2095, signal_1356}), .clk (clk), .r (Fresh[32]), .c ({signal_2155, signal_1416}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1253 ( .a ({signal_2031, signal_1292}), .b ({signal_2096, signal_1357}), .clk (clk), .r (Fresh[33]), .c ({signal_2156, signal_1417}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1254 ( .a ({Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({signal_2098, signal_1359}), .clk (clk), .r (Fresh[34]), .c ({signal_2157, signal_1418}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1255 ( .a ({signal_2032, signal_1293}), .b ({signal_2099, signal_1360}), .clk (clk), .r (Fresh[35]), .c ({signal_2158, signal_1419}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1256 ( .a ({Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({signal_2101, signal_1362}), .clk (clk), .r (Fresh[36]), .c ({signal_2159, signal_1420}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1257 ( .a ({signal_2033, signal_1294}), .b ({signal_2102, signal_1363}), .clk (clk), .r (Fresh[37]), .c ({signal_2160, signal_1421}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1258 ( .a ({Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({signal_2104, signal_1365}), .clk (clk), .r (Fresh[38]), .c ({signal_2161, signal_1422}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1259 ( .a ({signal_2034, signal_1295}), .b ({signal_2105, signal_1366}), .clk (clk), .r (Fresh[39]), .c ({signal_2162, signal_1423}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1260 ( .a ({Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({signal_2107, signal_1368}), .clk (clk), .r (Fresh[40]), .c ({signal_2163, signal_1424}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1261 ( .a ({signal_2035, signal_1296}), .b ({signal_2108, signal_1369}), .clk (clk), .r (Fresh[41]), .c ({signal_2164, signal_1425}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1262 ( .a ({Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({signal_2110, signal_1371}), .clk (clk), .r (Fresh[42]), .c ({signal_2165, signal_1426}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1263 ( .a ({signal_2036, signal_1297}), .b ({signal_2111, signal_1372}), .clk (clk), .r (Fresh[43]), .c ({signal_2166, signal_1427}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1264 ( .a ({Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({signal_2113, signal_1374}), .clk (clk), .r (Fresh[44]), .c ({signal_2167, signal_1428}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1265 ( .a ({signal_2037, signal_1298}), .b ({signal_2114, signal_1375}), .clk (clk), .r (Fresh[45]), .c ({signal_2168, signal_1429}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1266 ( .a ({Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({signal_2116, signal_1377}), .clk (clk), .r (Fresh[46]), .c ({signal_2169, signal_1430}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1267 ( .a ({signal_2038, signal_1299}), .b ({signal_2117, signal_1378}), .clk (clk), .r (Fresh[47]), .c ({signal_2170, signal_1431}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1268 ( .a ({Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({signal_2119, signal_1380}), .clk (clk), .r (Fresh[48]), .c ({signal_2171, signal_1432}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1269 ( .a ({signal_2039, signal_1300}), .b ({signal_2120, signal_1381}), .clk (clk), .r (Fresh[49]), .c ({signal_2172, signal_1433}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1270 ( .a ({Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({signal_2122, signal_1383}), .clk (clk), .r (Fresh[50]), .c ({signal_2173, signal_1434}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1271 ( .a ({signal_2040, signal_1301}), .b ({signal_2123, signal_1384}), .clk (clk), .r (Fresh[51]), .c ({signal_2174, signal_1435}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1272 ( .a ({Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({signal_2125, signal_1386}), .clk (clk), .r (Fresh[52]), .c ({signal_2175, signal_1436}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1273 ( .a ({signal_2041, signal_1302}), .b ({signal_2126, signal_1387}), .clk (clk), .r (Fresh[53]), .c ({signal_2176, signal_1437}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1274 ( .a ({Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({signal_2128, signal_1389}), .clk (clk), .r (Fresh[54]), .c ({signal_2177, signal_1438}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1275 ( .a ({signal_2042, signal_1303}), .b ({signal_2129, signal_1390}), .clk (clk), .r (Fresh[55]), .c ({signal_2178, signal_1439}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1276 ( .a ({Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({signal_2131, signal_1392}), .clk (clk), .r (Fresh[56]), .c ({signal_2179, signal_1440}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1277 ( .a ({signal_2043, signal_1304}), .b ({signal_2132, signal_1393}), .clk (clk), .r (Fresh[57]), .c ({signal_2180, signal_1441}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1278 ( .a ({Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({signal_2134, signal_1395}), .clk (clk), .r (Fresh[58]), .c ({signal_2181, signal_1442}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1279 ( .a ({signal_2044, signal_1305}), .b ({signal_2135, signal_1396}), .clk (clk), .r (Fresh[59]), .c ({signal_2182, signal_1443}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1280 ( .a ({Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({signal_2137, signal_1398}), .clk (clk), .r (Fresh[60]), .c ({signal_2183, signal_1444}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1281 ( .a ({signal_2045, signal_1306}), .b ({signal_2138, signal_1399}), .clk (clk), .r (Fresh[61]), .c ({signal_2184, signal_1445}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1282 ( .a ({Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({signal_2140, signal_1401}), .clk (clk), .r (Fresh[62]), .c ({signal_2185, signal_1446}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1283 ( .a ({signal_2046, signal_1307}), .b ({signal_2141, signal_1402}), .clk (clk), .r (Fresh[63]), .c ({signal_2186, signal_1447}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1311 ( .a ({signal_1967, signal_1228}), .b ({signal_2155, signal_1416}), .c ({signal_2214, signal_1472}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1312 ( .a ({signal_1968, signal_1229}), .b ({signal_2157, signal_1418}), .c ({signal_2215, signal_1473}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1313 ( .a ({signal_1969, signal_1230}), .b ({signal_2159, signal_1420}), .c ({signal_2216, signal_1474}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1314 ( .a ({signal_1970, signal_1231}), .b ({signal_2161, signal_1422}), .c ({signal_2217, signal_1475}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1315 ( .a ({signal_1971, signal_1232}), .b ({signal_2163, signal_1424}), .c ({signal_2218, signal_1476}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1316 ( .a ({signal_1972, signal_1233}), .b ({signal_2165, signal_1426}), .c ({signal_2219, signal_1477}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1317 ( .a ({signal_1973, signal_1234}), .b ({signal_2167, signal_1428}), .c ({signal_2220, signal_1478}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1318 ( .a ({signal_1974, signal_1235}), .b ({signal_2169, signal_1430}), .c ({signal_2221, signal_1479}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1319 ( .a ({signal_1975, signal_1236}), .b ({signal_2171, signal_1432}), .c ({signal_2222, signal_1480}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1320 ( .a ({signal_1976, signal_1237}), .b ({signal_2173, signal_1434}), .c ({signal_2223, signal_1481}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1321 ( .a ({signal_1977, signal_1238}), .b ({signal_2175, signal_1436}), .c ({signal_2224, signal_1482}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1322 ( .a ({signal_1978, signal_1239}), .b ({signal_2177, signal_1438}), .c ({signal_2225, signal_1483}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1323 ( .a ({signal_1979, signal_1240}), .b ({signal_2179, signal_1440}), .c ({signal_2226, signal_1484}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1324 ( .a ({signal_1980, signal_1241}), .b ({signal_2181, signal_1442}), .c ({signal_2227, signal_1485}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1325 ( .a ({signal_1981, signal_1242}), .b ({signal_2183, signal_1444}), .c ({signal_2228, signal_1486}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1326 ( .a ({signal_1982, signal_1243}), .b ({signal_2185, signal_1446}), .c ({signal_2229, signal_1487}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1347 ( .a ({signal_1936, signal_1212}), .b ({signal_2214, signal_1472}), .c ({signal_2256, signal_1508}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1348 ( .a ({signal_2156, signal_1417}), .b ({signal_2214, signal_1472}), .c ({signal_2257, signal_1509}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1349 ( .a ({signal_1938, signal_1213}), .b ({signal_2215, signal_1473}), .c ({signal_2258, signal_1510}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1350 ( .a ({signal_2158, signal_1419}), .b ({signal_2215, signal_1473}), .c ({signal_2259, signal_1511}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1351 ( .a ({signal_1940, signal_1214}), .b ({signal_2216, signal_1474}), .c ({signal_2260, signal_1512}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1352 ( .a ({signal_2160, signal_1421}), .b ({signal_2216, signal_1474}), .c ({signal_2261, signal_1513}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1353 ( .a ({signal_1942, signal_1215}), .b ({signal_2217, signal_1475}), .c ({signal_2262, signal_1514}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1354 ( .a ({signal_2162, signal_1423}), .b ({signal_2217, signal_1475}), .c ({signal_2263, signal_1515}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1355 ( .a ({signal_1944, signal_1216}), .b ({signal_2218, signal_1476}), .c ({signal_2264, signal_1516}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1356 ( .a ({signal_2164, signal_1425}), .b ({signal_2218, signal_1476}), .c ({signal_2265, signal_1517}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1357 ( .a ({signal_1946, signal_1217}), .b ({signal_2219, signal_1477}), .c ({signal_2266, signal_1518}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1358 ( .a ({signal_2166, signal_1427}), .b ({signal_2219, signal_1477}), .c ({signal_2267, signal_1519}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1359 ( .a ({signal_1948, signal_1218}), .b ({signal_2220, signal_1478}), .c ({signal_2268, signal_1520}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1360 ( .a ({signal_2168, signal_1429}), .b ({signal_2220, signal_1478}), .c ({signal_2269, signal_1521}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1361 ( .a ({signal_1950, signal_1219}), .b ({signal_2221, signal_1479}), .c ({signal_2270, signal_1522}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1362 ( .a ({signal_2170, signal_1431}), .b ({signal_2221, signal_1479}), .c ({signal_2271, signal_1523}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1363 ( .a ({signal_1952, signal_1220}), .b ({signal_2222, signal_1480}), .c ({signal_2272, signal_1524}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1364 ( .a ({signal_2172, signal_1433}), .b ({signal_2222, signal_1480}), .c ({signal_2273, signal_1525}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1365 ( .a ({signal_1954, signal_1221}), .b ({signal_2223, signal_1481}), .c ({signal_2274, signal_1526}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1366 ( .a ({signal_2174, signal_1435}), .b ({signal_2223, signal_1481}), .c ({signal_2275, signal_1527}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1367 ( .a ({signal_1956, signal_1222}), .b ({signal_2224, signal_1482}), .c ({signal_2276, signal_1528}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1368 ( .a ({signal_2176, signal_1437}), .b ({signal_2224, signal_1482}), .c ({signal_2277, signal_1529}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1369 ( .a ({signal_1958, signal_1223}), .b ({signal_2225, signal_1483}), .c ({signal_2278, signal_1530}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1370 ( .a ({signal_2178, signal_1439}), .b ({signal_2225, signal_1483}), .c ({signal_2279, signal_1531}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1371 ( .a ({signal_1960, signal_1224}), .b ({signal_2226, signal_1484}), .c ({signal_2280, signal_1532}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1372 ( .a ({signal_2180, signal_1441}), .b ({signal_2226, signal_1484}), .c ({signal_2281, signal_1533}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1373 ( .a ({signal_1962, signal_1225}), .b ({signal_2227, signal_1485}), .c ({signal_2282, signal_1534}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1374 ( .a ({signal_2182, signal_1443}), .b ({signal_2227, signal_1485}), .c ({signal_2283, signal_1535}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1375 ( .a ({signal_1964, signal_1226}), .b ({signal_2228, signal_1486}), .c ({signal_2284, signal_1536}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1376 ( .a ({signal_2184, signal_1445}), .b ({signal_2228, signal_1486}), .c ({signal_2285, signal_1537}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1377 ( .a ({signal_1966, signal_1227}), .b ({signal_2229, signal_1487}), .c ({signal_2286, signal_1538}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1378 ( .a ({signal_2186, signal_1447}), .b ({signal_2229, signal_1487}), .c ({signal_2287, signal_1539}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1405 ( .a ({signal_2187, signal_1448}), .b ({signal_2256, signal_1508}), .c ({signal_2326, signal_1553}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1406 ( .a ({signal_2188, signal_1449}), .b ({signal_2258, signal_1510}), .c ({signal_2327, signal_1554}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1407 ( .a ({signal_2189, signal_1450}), .b ({signal_2260, signal_1512}), .c ({signal_2328, signal_1555}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1408 ( .a ({signal_2190, signal_1451}), .b ({signal_2262, signal_1514}), .c ({signal_2329, signal_1556}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1409 ( .a ({signal_2191, signal_1452}), .b ({signal_2264, signal_1516}), .c ({signal_2330, signal_1557}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1410 ( .a ({signal_2192, signal_1453}), .b ({signal_2266, signal_1518}), .c ({signal_2331, signal_1558}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1411 ( .a ({signal_2193, signal_1454}), .b ({signal_2268, signal_1520}), .c ({signal_2332, signal_1559}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1412 ( .a ({signal_2194, signal_1455}), .b ({signal_2270, signal_1522}), .c ({signal_2333, signal_1560}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1413 ( .a ({signal_2195, signal_1456}), .b ({signal_2272, signal_1524}), .c ({signal_2334, signal_1561}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1414 ( .a ({signal_2196, signal_1457}), .b ({signal_2274, signal_1526}), .c ({signal_2335, signal_1562}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1415 ( .a ({signal_2197, signal_1458}), .b ({signal_2276, signal_1528}), .c ({signal_2336, signal_1563}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1416 ( .a ({signal_2198, signal_1459}), .b ({signal_2278, signal_1530}), .c ({signal_2337, signal_1564}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1417 ( .a ({signal_2199, signal_1460}), .b ({signal_2280, signal_1532}), .c ({signal_2338, signal_1565}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1418 ( .a ({signal_2200, signal_1461}), .b ({signal_2282, signal_1534}), .c ({signal_2339, signal_1566}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1419 ( .a ({signal_2201, signal_1462}), .b ({signal_2284, signal_1536}), .c ({signal_2340, signal_1567}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1420 ( .a ({signal_2202, signal_1463}), .b ({signal_2286, signal_1538}), .c ({signal_2341, signal_1568}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1421 ( .a ({1'b0, 1'b0}), .b ({signal_2287, signal_1539}), .c ({signal_2342, signal_1569}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1422 ( .a ({1'b0, 1'b0}), .b ({signal_2279, signal_1531}), .c ({signal_2343, signal_1570}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1423 ( .a ({1'b0, 1'b0}), .b ({signal_2273, signal_1525}), .c ({signal_2344, signal_1571}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1424 ( .a ({1'b0, 1'b0}), .b ({signal_2275, signal_1527}), .c ({signal_2345, signal_1572}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1425 ( .a ({1'b0, 1'b0}), .b ({signal_2277, signal_1529}), .c ({signal_2346, signal_1573}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1426 ( .a ({1'b0, 1'b0}), .b ({signal_2281, signal_1533}), .c ({signal_2347, signal_1574}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1427 ( .a ({1'b0, 1'b0}), .b ({signal_2283, signal_1535}), .c ({signal_2348, signal_1575}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1428 ( .a ({1'b0, 1'b0}), .b ({signal_2285, signal_1537}), .c ({signal_2349, signal_1576}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1429 ( .a ({signal_2263, signal_1515}), .b ({signal_2269, signal_1521}), .c ({signal_2350, signal_1577}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1430 ( .a ({signal_2257, signal_1509}), .b ({signal_2271, signal_1523}), .c ({signal_2351, signal_1578}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1431 ( .a ({signal_2259, signal_1511}), .b ({signal_2265, signal_1517}), .c ({signal_2352, signal_1579}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1432 ( .a ({signal_2261, signal_1513}), .b ({signal_2267, signal_1519}), .c ({signal_2353, signal_1580}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1443 ( .a ({1'b0, signal_1028}), .b ({signal_2342, signal_1569}), .c ({signal_2378, signal_1591}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1444 ( .a ({1'b0, 1'b0}), .b ({signal_2341, signal_1568}), .c ({signal_2379, signal_1592}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1445 ( .a ({1'b0, signal_940}), .b ({signal_2343, signal_1570}), .c ({signal_2380, signal_1593}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1446 ( .a ({1'b0, 1'b0}), .b ({signal_2337, signal_1564}), .c ({signal_2381, signal_1594}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1447 ( .a ({signal_1647, signal_1163}), .b ({signal_2344, signal_1571}), .c ({signal_2382, signal_1595}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1448 ( .a ({1'b0, 1'b0}), .b ({signal_2334, signal_1561}), .c ({signal_2383, signal_1596}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1449 ( .a ({signal_1659, signal_1159}), .b ({signal_2345, signal_1572}), .c ({signal_2384, signal_1597}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1450 ( .a ({1'b0, 1'b0}), .b ({signal_2335, signal_1562}), .c ({signal_2385, signal_1598}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1451 ( .a ({signal_1671, signal_1155}), .b ({signal_2346, signal_1573}), .c ({signal_2386, signal_1599}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1452 ( .a ({1'b0, 1'b0}), .b ({signal_2336, signal_1563}), .c ({signal_2387, signal_1600}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1453 ( .a ({signal_1695, signal_1147}), .b ({signal_2347, signal_1574}), .c ({signal_2388, signal_807}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1454 ( .a ({1'b0, 1'b0}), .b ({signal_2338, signal_1565}), .c ({signal_2389, signal_1601}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1455 ( .a ({signal_1707, signal_1143}), .b ({signal_2348, signal_1575}), .c ({signal_2390, signal_803}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1456 ( .a ({1'b0, 1'b0}), .b ({signal_2339, signal_1566}), .c ({signal_2391, signal_1602}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1457 ( .a ({signal_1719, signal_1139}), .b ({signal_2349, signal_1576}), .c ({signal_2392, signal_799}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1458 ( .a ({1'b0, 1'b0}), .b ({signal_2340, signal_1567}), .c ({signal_2393, signal_1603}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1459 ( .a ({signal_2329, signal_1556}), .b ({signal_2332, signal_1559}), .c ({signal_2394, signal_1604}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1460 ( .a ({signal_2327, signal_1554}), .b ({signal_2330, signal_1557}), .c ({signal_2395, signal_1605}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1461 ( .a ({signal_2328, signal_1555}), .b ({signal_2331, signal_1558}), .c ({signal_2396, signal_1606}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1465 ( .a ({signal_2326, signal_1553}), .b ({signal_2333, signal_1560}), .c ({signal_2400, signal_1610}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1482 ( .a ({1'b0, signal_943}), .b ({signal_2379, signal_1592}), .c ({signal_2439, signal_1614}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1483 ( .a ({1'b0, signal_939}), .b ({signal_2381, signal_1594}), .c ({signal_2440, signal_1615}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1484 ( .a ({signal_1650, signal_1162}), .b ({signal_2383, signal_1596}), .c ({signal_2441, signal_1616}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1485 ( .a ({signal_1662, signal_1158}), .b ({signal_2385, signal_1598}), .c ({signal_2442, signal_1617}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1486 ( .a ({signal_1674, signal_1154}), .b ({signal_2387, signal_1600}), .c ({signal_2443, signal_1618}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1487 ( .a ({1'b0, 1'b0}), .b ({signal_2380, signal_1593}), .c ({signal_2444, signal_1619}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1488 ( .a ({signal_1698, signal_1146}), .b ({signal_2389, signal_1601}), .c ({signal_2445, signal_806}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1489 ( .a ({signal_1710, signal_1142}), .b ({signal_2391, signal_1602}), .c ({signal_2446, signal_802}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1490 ( .a ({signal_1722, signal_1138}), .b ({signal_2393, signal_1603}), .c ({signal_2447, signal_798}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1491 ( .a ({1'b0, 1'b0}), .b ({signal_2378, signal_1591}), .c ({signal_2448, signal_1620}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1492 ( .a ({1'b0, 1'b0}), .b ({signal_2388, signal_807}), .c ({signal_2449, signal_1621}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1493 ( .a ({1'b0, 1'b0}), .b ({signal_2390, signal_803}), .c ({signal_2450, signal_1622}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1494 ( .a ({1'b0, 1'b0}), .b ({signal_2392, signal_799}), .c ({signal_2451, signal_1623}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1495 ( .a ({1'b0, 1'b0}), .b ({signal_2384, signal_1597}), .c ({signal_2452, signal_1624}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1496 ( .a ({1'b0, 1'b0}), .b ({signal_2386, signal_1599}), .c ({signal_2453, signal_1625}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1497 ( .a ({1'b0, 1'b0}), .b ({signal_2382, signal_1595}), .c ({signal_2454, signal_1626}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1500 ( .a ({signal_1683, signal_1151}), .b ({signal_2444, signal_1619}), .c ({signal_2473, signal_1629}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1501 ( .a ({1'b0, 1'b0}), .b ({signal_2440, signal_1615}), .c ({signal_2474, signal_1630}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1502 ( .a ({signal_1731, signal_1135}), .b ({signal_2448, signal_1620}), .c ({signal_2475, signal_795}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1503 ( .a ({1'b0, 1'b0}), .b ({signal_2439, signal_1614}), .c ({signal_2476, signal_1631}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1504 ( .a ({signal_2350, signal_1577}), .b ({signal_2449, signal_1621}), .c ({signal_2477, signal_791}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1505 ( .a ({1'b0, 1'b0}), .b ({signal_2445, signal_806}), .c ({signal_2478, signal_1632}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1506 ( .a ({signal_2351, signal_1578}), .b ({signal_2450, signal_1622}), .c ({signal_2479, signal_787}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1507 ( .a ({1'b0, 1'b0}), .b ({signal_2446, signal_802}), .c ({signal_2480, signal_1633}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1508 ( .a ({signal_2352, signal_1579}), .b ({signal_2451, signal_1623}), .c ({signal_2481, signal_783}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1509 ( .a ({1'b0, 1'b0}), .b ({signal_2447, signal_798}), .c ({signal_2482, signal_1634}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1510 ( .a ({signal_2269, signal_1521}), .b ({signal_2452, signal_1624}), .c ({signal_2483, signal_823}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1511 ( .a ({1'b0, 1'b0}), .b ({signal_2442, signal_1617}), .c ({signal_2484, signal_1635}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1512 ( .a ({signal_2271, signal_1523}), .b ({signal_2453, signal_1625}), .c ({signal_2485, signal_819}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1513 ( .a ({1'b0, 1'b0}), .b ({signal_2443, signal_1618}), .c ({signal_2486, signal_1636}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1514 ( .a ({signal_2267, signal_1519}), .b ({signal_2454, signal_1626}), .c ({signal_2487, signal_811}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1515 ( .a ({1'b0, 1'b0}), .b ({signal_2441, signal_1616}), .c ({signal_2488, signal_1637}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1516 ( .a ({signal_2269, signal_1521}), .b ({signal_2449, signal_1621}), .c ({signal_2489, signal_839}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1517 ( .a ({signal_2271, signal_1523}), .b ({signal_2450, signal_1622}), .c ({signal_2490, signal_835}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1518 ( .a ({signal_2265, signal_1517}), .b ({signal_2451, signal_1623}), .c ({signal_2491, signal_831}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1523 ( .a ({signal_1686, signal_1150}), .b ({signal_2474, signal_1630}), .c ({signal_2520, signal_1639}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1524 ( .a ({signal_1734, signal_1134}), .b ({signal_2476, signal_1631}), .c ({signal_2521, signal_794}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1525 ( .a ({signal_2394, signal_1604}), .b ({signal_2478, signal_1632}), .c ({signal_2522, signal_790}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1526 ( .a ({signal_2400, signal_1610}), .b ({signal_2480, signal_1633}), .c ({signal_2523, signal_1640}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1527 ( .a ({signal_2395, signal_1605}), .b ({signal_2482, signal_1634}), .c ({signal_2524, signal_782}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1528 ( .a ({1'b0, 1'b0}), .b ({signal_2475, signal_795}), .c ({signal_2525, signal_1641}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1529 ( .a ({signal_2332, signal_1559}), .b ({signal_2484, signal_1635}), .c ({signal_2526, signal_822}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1530 ( .a ({signal_2333, signal_1560}), .b ({signal_2486, signal_1636}), .c ({signal_2527, signal_1642}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1531 ( .a ({1'b0, 1'b0}), .b ({signal_2473, signal_1629}), .c ({signal_2528, signal_1643}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1532 ( .a ({signal_2331, signal_1558}), .b ({signal_2488, signal_1637}), .c ({signal_2529, signal_810}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1533 ( .a ({signal_2332, signal_1559}), .b ({signal_2478, signal_1632}), .c ({signal_2530, signal_838}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1534 ( .a ({signal_2333, signal_1560}), .b ({signal_2480, signal_1633}), .c ({signal_2531, signal_1644}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1535 ( .a ({signal_2330, signal_1557}), .b ({signal_2482, signal_1634}), .c ({signal_2532, signal_830}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1536 ( .a ({signal_2523, signal_1640}), .b ({signal_2549, signal_786}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1537 ( .a ({signal_2527, signal_1642}), .b ({signal_2550, signal_818}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1538 ( .a ({signal_2531, signal_1644}), .b ({signal_2551, signal_834}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1539 ( .a ({signal_2353, signal_1580}), .b ({signal_2525, signal_1641}), .c ({signal_2552, signal_779}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1540 ( .a ({1'b0, 1'b0}), .b ({signal_2521, signal_794}), .c ({signal_2553, signal_1645}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1541 ( .a ({signal_2265, signal_1517}), .b ({signal_2528, signal_1643}), .c ({signal_2554, signal_815}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1542 ( .a ({1'b0, 1'b0}), .b ({signal_2520, signal_1639}), .c ({signal_2555, signal_1646}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1543 ( .a ({signal_2267, signal_1519}), .b ({signal_2525, signal_1641}), .c ({signal_2556, signal_827}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1544 ( .a ({signal_2396, signal_1606}), .b ({signal_2553, signal_1645}), .c ({signal_2569, signal_778}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1545 ( .a ({signal_2330, signal_1557}), .b ({signal_2555, signal_1646}), .c ({signal_2570, signal_814}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1546 ( .a ({signal_2331, signal_1558}), .b ({signal_2553, signal_1645}), .c ({signal_2571, signal_826}) ) ;

    /* register cells */
    reg_masked #(.security_order(1), .pipeline(0)) cell_65 ( .clk (signal_2642), .D ({signal_2548, signal_840}), .Q ({Ciphertext_s1[63], Ciphertext_s0[63]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_67 ( .clk (signal_2642), .D ({signal_2472, signal_841}), .Q ({Ciphertext_s1[62], Ciphertext_s0[62]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_69 ( .clk (signal_2642), .D ({signal_2577, signal_842}), .Q ({Ciphertext_s1[61], Ciphertext_s0[61]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_71 ( .clk (signal_2642), .D ({signal_2568, signal_843}), .Q ({Ciphertext_s1[60], Ciphertext_s0[60]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_73 ( .clk (signal_2642), .D ({signal_2470, signal_844}), .Q ({Ciphertext_s1[59], Ciphertext_s0[59]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_75 ( .clk (signal_2642), .D ({signal_2377, signal_845}), .Q ({Ciphertext_s1[58], Ciphertext_s0[58]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_77 ( .clk (signal_2642), .D ({signal_2546, signal_846}), .Q ({Ciphertext_s1[57], Ciphertext_s0[57]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_79 ( .clk (signal_2642), .D ({signal_2518, signal_847}), .Q ({Ciphertext_s1[56], Ciphertext_s0[56]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_81 ( .clk (signal_2642), .D ({signal_2468, signal_848}), .Q ({Ciphertext_s1[55], Ciphertext_s0[55]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_83 ( .clk (signal_2642), .D ({signal_2375, signal_849}), .Q ({Ciphertext_s1[54], Ciphertext_s0[54]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_85 ( .clk (signal_2642), .D ({signal_2566, signal_850}), .Q ({Ciphertext_s1[53], Ciphertext_s0[53]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_87 ( .clk (signal_2642), .D ({signal_2516, signal_851}), .Q ({Ciphertext_s1[52], Ciphertext_s0[52]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_89 ( .clk (signal_2642), .D ({signal_2466, signal_852}), .Q ({Ciphertext_s1[51], Ciphertext_s0[51]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_91 ( .clk (signal_2642), .D ({signal_2373, signal_853}), .Q ({Ciphertext_s1[50], Ciphertext_s0[50]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_93 ( .clk (signal_2642), .D ({signal_2544, signal_854}), .Q ({Ciphertext_s1[49], Ciphertext_s0[49]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_95 ( .clk (signal_2642), .D ({signal_2514, signal_855}), .Q ({Ciphertext_s1[48], Ciphertext_s0[48]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_97 ( .clk (signal_2642), .D ({signal_2464, signal_856}), .Q ({Ciphertext_s1[47], Ciphertext_s0[47]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_99 ( .clk (signal_2642), .D ({signal_2371, signal_857}), .Q ({Ciphertext_s1[46], Ciphertext_s0[46]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_101 ( .clk (signal_2642), .D ({signal_2542, signal_858}), .Q ({Ciphertext_s1[45], Ciphertext_s0[45]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_103 ( .clk (signal_2642), .D ({signal_2512, signal_859}), .Q ({Ciphertext_s1[44], Ciphertext_s0[44]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_105 ( .clk (signal_2642), .D ({signal_2369, signal_860}), .Q ({Ciphertext_s1[43], Ciphertext_s0[43]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_107 ( .clk (signal_2642), .D ({signal_2255, signal_861}), .Q ({Ciphertext_s1[42], Ciphertext_s0[42]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_109 ( .clk (signal_2642), .D ({signal_2462, signal_862}), .Q ({Ciphertext_s1[41], Ciphertext_s0[41]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_111 ( .clk (signal_2642), .D ({signal_2433, signal_863}), .Q ({Ciphertext_s1[40], Ciphertext_s0[40]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_113 ( .clk (signal_2642), .D ({signal_2367, signal_864}), .Q ({Ciphertext_s1[39], Ciphertext_s0[39]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_115 ( .clk (signal_2642), .D ({signal_2253, signal_865}), .Q ({Ciphertext_s1[38], Ciphertext_s0[38]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_117 ( .clk (signal_2642), .D ({signal_2460, signal_866}), .Q ({Ciphertext_s1[37], Ciphertext_s0[37]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_119 ( .clk (signal_2642), .D ({signal_2431, signal_867}), .Q ({Ciphertext_s1[36], Ciphertext_s0[36]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_121 ( .clk (signal_2642), .D ({signal_2365, signal_868}), .Q ({Ciphertext_s1[35], Ciphertext_s0[35]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_123 ( .clk (signal_2642), .D ({signal_2251, signal_869}), .Q ({Ciphertext_s1[34], Ciphertext_s0[34]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_125 ( .clk (signal_2642), .D ({signal_2458, signal_870}), .Q ({Ciphertext_s1[33], Ciphertext_s0[33]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_127 ( .clk (signal_2642), .D ({signal_2429, signal_871}), .Q ({Ciphertext_s1[32], Ciphertext_s0[32]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_129 ( .clk (signal_2642), .D ({signal_2427, signal_872}), .Q ({Ciphertext_s1[31], Ciphertext_s0[31]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_131 ( .clk (signal_2642), .D ({signal_2318, signal_873}), .Q ({Ciphertext_s1[30], Ciphertext_s0[30]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_133 ( .clk (signal_2642), .D ({signal_2540, signal_874}), .Q ({Ciphertext_s1[29], Ciphertext_s0[29]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_135 ( .clk (signal_2642), .D ({signal_2510, signal_875}), .Q ({Ciphertext_s1[28], Ciphertext_s0[28]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_137 ( .clk (signal_2642), .D ({signal_2508, signal_876}), .Q ({Ciphertext_s1[27], Ciphertext_s0[27]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_139 ( .clk (signal_2642), .D ({signal_2425, signal_877}), .Q ({Ciphertext_s1[26], Ciphertext_s0[26]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_141 ( .clk (signal_2642), .D ({signal_2575, signal_878}), .Q ({Ciphertext_s1[25], Ciphertext_s0[25]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_143 ( .clk (signal_2642), .D ({signal_2564, signal_879}), .Q ({Ciphertext_s1[24], Ciphertext_s0[24]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_145 ( .clk (signal_2642), .D ({signal_2423, signal_880}), .Q ({Ciphertext_s1[23], Ciphertext_s0[23]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_147 ( .clk (signal_2642), .D ({signal_2316, signal_881}), .Q ({Ciphertext_s1[22], Ciphertext_s0[22]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_149 ( .clk (signal_2642), .D ({signal_2562, signal_882}), .Q ({Ciphertext_s1[21], Ciphertext_s0[21]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_151 ( .clk (signal_2642), .D ({signal_2506, signal_883}), .Q ({Ciphertext_s1[20], Ciphertext_s0[20]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_153 ( .clk (signal_2642), .D ({signal_2421, signal_884}), .Q ({Ciphertext_s1[19], Ciphertext_s0[19]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_155 ( .clk (signal_2642), .D ({signal_2314, signal_885}), .Q ({Ciphertext_s1[18], Ciphertext_s0[18]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_157 ( .clk (signal_2642), .D ({signal_2538, signal_886}), .Q ({Ciphertext_s1[17], Ciphertext_s0[17]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_159 ( .clk (signal_2642), .D ({signal_2504, signal_887}), .Q ({Ciphertext_s1[16], Ciphertext_s0[16]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_161 ( .clk (signal_2642), .D ({signal_2502, signal_888}), .Q ({Ciphertext_s1[15], Ciphertext_s0[15]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_163 ( .clk (signal_2642), .D ({signal_2419, signal_889}), .Q ({Ciphertext_s1[14], Ciphertext_s0[14]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_165 ( .clk (signal_2642), .D ({signal_2573, signal_890}), .Q ({Ciphertext_s1[13], Ciphertext_s0[13]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_167 ( .clk (signal_2642), .D ({signal_2560, signal_891}), .Q ({Ciphertext_s1[12], Ciphertext_s0[12]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_169 ( .clk (signal_2642), .D ({signal_2417, signal_892}), .Q ({Ciphertext_s1[11], Ciphertext_s0[11]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_171 ( .clk (signal_2642), .D ({signal_2312, signal_893}), .Q ({Ciphertext_s1[10], Ciphertext_s0[10]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_173 ( .clk (signal_2642), .D ({signal_2536, signal_894}), .Q ({Ciphertext_s1[9], Ciphertext_s0[9]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_175 ( .clk (signal_2642), .D ({signal_2500, signal_895}), .Q ({Ciphertext_s1[8], Ciphertext_s0[8]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_177 ( .clk (signal_2642), .D ({signal_2415, signal_896}), .Q ({Ciphertext_s1[7], Ciphertext_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_179 ( .clk (signal_2642), .D ({signal_2310, signal_897}), .Q ({Ciphertext_s1[6], Ciphertext_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_181 ( .clk (signal_2642), .D ({signal_2558, signal_898}), .Q ({Ciphertext_s1[5], Ciphertext_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_183 ( .clk (signal_2642), .D ({signal_2498, signal_899}), .Q ({Ciphertext_s1[4], Ciphertext_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_185 ( .clk (signal_2642), .D ({signal_2413, signal_900}), .Q ({Ciphertext_s1[3], Ciphertext_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_187 ( .clk (signal_2642), .D ({signal_2308, signal_901}), .Q ({Ciphertext_s1[2], Ciphertext_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_189 ( .clk (signal_2642), .D ({signal_2534, signal_902}), .Q ({Ciphertext_s1[1], Ciphertext_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_191 ( .clk (signal_2642), .D ({signal_2496, signal_903}), .Q ({Ciphertext_s1[0], Ciphertext_s0[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_834 ( .clk (signal_2642), .D ({signal_1838, signal_1036}), .Q ({signal_1740, signal_1132}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_836 ( .clk (signal_2642), .D ({signal_1835, signal_1037}), .Q ({signal_1737, signal_1133}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_838 ( .clk (signal_2642), .D ({signal_1832, signal_1038}), .Q ({signal_1734, signal_1134}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_840 ( .clk (signal_2642), .D ({signal_1829, signal_1039}), .Q ({signal_1731, signal_1135}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_842 ( .clk (signal_2642), .D ({signal_1826, signal_1040}), .Q ({signal_1728, signal_1136}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_844 ( .clk (signal_2642), .D ({signal_1823, signal_1041}), .Q ({signal_1725, signal_1137}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_846 ( .clk (signal_2642), .D ({signal_1820, signal_1042}), .Q ({signal_1722, signal_1138}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_848 ( .clk (signal_2642), .D ({signal_1817, signal_1043}), .Q ({signal_1719, signal_1139}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_850 ( .clk (signal_2642), .D ({signal_1814, signal_1044}), .Q ({signal_1716, signal_1140}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_852 ( .clk (signal_2642), .D ({signal_1811, signal_1045}), .Q ({signal_1713, signal_1141}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_854 ( .clk (signal_2642), .D ({signal_1808, signal_1046}), .Q ({signal_1710, signal_1142}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_856 ( .clk (signal_2642), .D ({signal_1805, signal_1047}), .Q ({signal_1707, signal_1143}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_858 ( .clk (signal_2642), .D ({signal_1802, signal_1048}), .Q ({signal_1704, signal_1144}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_860 ( .clk (signal_2642), .D ({signal_1799, signal_1049}), .Q ({signal_1701, signal_1145}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_862 ( .clk (signal_2642), .D ({signal_1796, signal_1050}), .Q ({signal_1698, signal_1146}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_864 ( .clk (signal_2642), .D ({signal_1793, signal_1051}), .Q ({signal_1695, signal_1147}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_866 ( .clk (signal_2642), .D ({signal_1790, signal_1052}), .Q ({signal_1692, signal_1148}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_868 ( .clk (signal_2642), .D ({signal_1787, signal_1053}), .Q ({signal_1689, signal_1149}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_870 ( .clk (signal_2642), .D ({signal_1784, signal_1054}), .Q ({signal_1686, signal_1150}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_872 ( .clk (signal_2642), .D ({signal_1781, signal_1055}), .Q ({signal_1683, signal_1151}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_874 ( .clk (signal_2642), .D ({signal_1778, signal_1056}), .Q ({signal_1680, signal_1152}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_876 ( .clk (signal_2642), .D ({signal_1775, signal_1057}), .Q ({signal_1677, signal_1153}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_878 ( .clk (signal_2642), .D ({signal_1772, signal_1058}), .Q ({signal_1674, signal_1154}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_880 ( .clk (signal_2642), .D ({signal_1769, signal_1059}), .Q ({signal_1671, signal_1155}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_882 ( .clk (signal_2642), .D ({signal_1766, signal_1060}), .Q ({signal_1668, signal_1156}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_884 ( .clk (signal_2642), .D ({signal_1763, signal_1061}), .Q ({signal_1665, signal_1157}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_886 ( .clk (signal_2642), .D ({signal_1760, signal_1062}), .Q ({signal_1662, signal_1158}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_888 ( .clk (signal_2642), .D ({signal_1757, signal_1063}), .Q ({signal_1659, signal_1159}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_890 ( .clk (signal_2642), .D ({signal_1754, signal_1064}), .Q ({signal_1656, signal_1160}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_892 ( .clk (signal_2642), .D ({signal_1751, signal_1065}), .Q ({signal_1653, signal_1161}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_894 ( .clk (signal_2642), .D ({signal_1748, signal_1066}), .Q ({signal_1650, signal_1162}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_896 ( .clk (signal_2642), .D ({signal_1745, signal_1067}), .Q ({signal_1647, signal_1163}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_898 ( .clk (signal_2642), .D ({signal_1742, signal_1068}), .Q ({signal_1812, signal_1108}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_900 ( .clk (signal_2642), .D ({signal_1739, signal_1069}), .Q ({signal_1809, signal_1109}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_902 ( .clk (signal_2642), .D ({signal_1736, signal_1070}), .Q ({signal_1806, signal_1110}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_904 ( .clk (signal_2642), .D ({signal_1733, signal_1071}), .Q ({signal_1803, signal_1111}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_906 ( .clk (signal_2642), .D ({signal_1730, signal_1072}), .Q ({signal_1836, signal_1100}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_908 ( .clk (signal_2642), .D ({signal_1727, signal_1073}), .Q ({signal_1833, signal_1101}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_910 ( .clk (signal_2642), .D ({signal_1724, signal_1074}), .Q ({signal_1830, signal_1102}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_912 ( .clk (signal_2642), .D ({signal_1721, signal_1075}), .Q ({signal_1827, signal_1103}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_914 ( .clk (signal_2642), .D ({signal_1718, signal_1076}), .Q ({signal_1788, signal_1116}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_916 ( .clk (signal_2642), .D ({signal_1715, signal_1077}), .Q ({signal_1785, signal_1117}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_918 ( .clk (signal_2642), .D ({signal_1712, signal_1078}), .Q ({signal_1782, signal_1118}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_920 ( .clk (signal_2642), .D ({signal_1709, signal_1079}), .Q ({signal_1779, signal_1119}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_922 ( .clk (signal_2642), .D ({signal_1706, signal_1080}), .Q ({signal_1752, signal_1128}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_924 ( .clk (signal_2642), .D ({signal_1703, signal_1081}), .Q ({signal_1749, signal_1129}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_926 ( .clk (signal_2642), .D ({signal_1700, signal_1082}), .Q ({signal_1746, signal_1130}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_928 ( .clk (signal_2642), .D ({signal_1697, signal_1083}), .Q ({signal_1743, signal_1131}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_930 ( .clk (signal_2642), .D ({signal_1694, signal_1084}), .Q ({signal_1764, signal_1124}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_932 ( .clk (signal_2642), .D ({signal_1691, signal_1085}), .Q ({signal_1761, signal_1125}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_934 ( .clk (signal_2642), .D ({signal_1688, signal_1086}), .Q ({signal_1758, signal_1126}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_936 ( .clk (signal_2642), .D ({signal_1685, signal_1087}), .Q ({signal_1755, signal_1127}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_938 ( .clk (signal_2642), .D ({signal_1682, signal_1088}), .Q ({signal_1800, signal_1112}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_940 ( .clk (signal_2642), .D ({signal_1679, signal_1089}), .Q ({signal_1797, signal_1113}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_942 ( .clk (signal_2642), .D ({signal_1676, signal_1090}), .Q ({signal_1794, signal_1114}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_944 ( .clk (signal_2642), .D ({signal_1673, signal_1091}), .Q ({signal_1791, signal_1115}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_946 ( .clk (signal_2642), .D ({signal_1670, signal_1092}), .Q ({signal_1776, signal_1120}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_948 ( .clk (signal_2642), .D ({signal_1667, signal_1093}), .Q ({signal_1773, signal_1121}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_950 ( .clk (signal_2642), .D ({signal_1664, signal_1094}), .Q ({signal_1770, signal_1122}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_952 ( .clk (signal_2642), .D ({signal_1661, signal_1095}), .Q ({signal_1767, signal_1123}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_954 ( .clk (signal_2642), .D ({signal_1658, signal_1096}), .Q ({signal_1824, signal_1104}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_956 ( .clk (signal_2642), .D ({signal_1655, signal_1097}), .Q ({signal_1821, signal_1105}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_958 ( .clk (signal_2642), .D ({signal_1652, signal_1098}), .Q ({signal_1818, signal_1106}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_960 ( .clk (signal_2642), .D ({signal_1649, signal_1099}), .Q ({signal_1815, signal_1107}) ) ;
    DFF_X1 cell_968 ( .CK (signal_2642), .D (signal_1030), .Q (signal_939), .QN () ) ;
    DFF_X1 cell_970 ( .CK (signal_2642), .D (signal_1031), .Q (signal_940), .QN () ) ;
    DFF_X1 cell_972 ( .CK (signal_2642), .D (signal_1032), .Q (signal_1025), .QN () ) ;
    DFF_X1 cell_974 ( .CK (signal_2642), .D (signal_1033), .Q (signal_1026), .QN () ) ;
    DFF_X1 cell_976 ( .CK (signal_2642), .D (signal_1034), .Q (signal_943), .QN () ) ;
    DFF_X1 cell_978 ( .CK (signal_2642), .D (signal_1035), .Q (signal_1028), .QN () ) ;
endmodule
