/* modified netlist. Source: module CRAFT in file Designs/CRAFT_round-based/AGEMA/CRAFT.v */
/* 2 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 3 register stage(s) in total */

module CRAFT_GHPC_ANF_Pipeline_d1 (plaintext_s0, key_s0, clk, rst, key_s1, plaintext_s1, Fresh, ciphertext_s0, done, ciphertext_s1);
    input [63:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input rst ;
    input [127:0] key_s1 ;
    input [63:0] plaintext_s1 ;
    input [63:0] Fresh ;
    output [63:0] ciphertext_s0 ;
    output done ;
    output [63:0] ciphertext_s1 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_285 ;
    wire signal_286 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_295 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_352 ;
    wire signal_353 ;
    wire signal_354 ;
    wire signal_355 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_359 ;
    wire signal_360 ;
    wire signal_361 ;
    wire signal_362 ;
    wire signal_363 ;
    wire signal_364 ;
    wire signal_365 ;
    wire signal_366 ;
    wire signal_367 ;
    wire signal_368 ;
    wire signal_369 ;
    wire signal_370 ;
    wire signal_371 ;
    wire signal_372 ;
    wire signal_373 ;
    wire signal_374 ;
    wire signal_375 ;
    wire signal_376 ;
    wire signal_377 ;
    wire signal_378 ;
    wire signal_379 ;
    wire signal_380 ;
    wire signal_381 ;
    wire signal_382 ;
    wire signal_383 ;
    wire signal_384 ;
    wire signal_385 ;
    wire signal_386 ;
    wire signal_387 ;
    wire signal_692 ;
    wire signal_693 ;
    wire signal_694 ;
    wire signal_702 ;
    wire signal_703 ;
    wire signal_704 ;
    wire signal_705 ;
    wire signal_706 ;
    wire signal_707 ;
    wire signal_711 ;
    wire signal_712 ;
    wire signal_713 ;
    wire signal_714 ;
    wire signal_715 ;
    wire signal_716 ;
    wire signal_717 ;
    wire signal_718 ;
    wire signal_719 ;
    wire signal_720 ;
    wire signal_721 ;
    wire signal_722 ;
    wire signal_723 ;
    wire signal_724 ;
    wire signal_725 ;
    wire signal_726 ;
    wire signal_727 ;
    wire signal_728 ;
    wire signal_729 ;
    wire signal_730 ;
    wire signal_731 ;
    wire signal_732 ;
    wire signal_733 ;
    wire signal_734 ;
    wire signal_735 ;
    wire signal_736 ;
    wire signal_737 ;
    wire signal_738 ;
    wire signal_739 ;
    wire signal_740 ;
    wire signal_741 ;
    wire signal_742 ;
    wire signal_743 ;
    wire signal_744 ;
    wire signal_745 ;
    wire signal_746 ;
    wire signal_747 ;
    wire signal_748 ;
    wire signal_749 ;
    wire signal_750 ;
    wire signal_751 ;
    wire signal_752 ;
    wire signal_753 ;
    wire signal_754 ;
    wire signal_755 ;
    wire signal_756 ;
    wire signal_757 ;
    wire signal_758 ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_768 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_771 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_774 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_777 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_780 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_783 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_786 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_789 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_792 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_809 ;
    wire signal_810 ;
    wire signal_811 ;
    wire signal_812 ;
    wire signal_813 ;
    wire signal_814 ;
    wire signal_815 ;
    wire signal_816 ;
    wire signal_817 ;
    wire signal_818 ;
    wire signal_819 ;
    wire signal_820 ;
    wire signal_821 ;
    wire signal_822 ;
    wire signal_823 ;
    wire signal_824 ;
    wire signal_825 ;
    wire signal_826 ;
    wire signal_827 ;
    wire signal_828 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_831 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_834 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_837 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_840 ;
    wire signal_841 ;
    wire signal_842 ;
    wire signal_843 ;
    wire signal_844 ;
    wire signal_845 ;
    wire signal_846 ;
    wire signal_847 ;
    wire signal_848 ;
    wire signal_849 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_852 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_855 ;
    wire signal_856 ;
    wire signal_857 ;
    wire signal_858 ;
    wire signal_859 ;
    wire signal_860 ;
    wire signal_861 ;
    wire signal_862 ;
    wire signal_863 ;
    wire signal_864 ;
    wire signal_865 ;
    wire signal_866 ;
    wire signal_867 ;
    wire signal_868 ;
    wire signal_869 ;
    wire signal_870 ;
    wire signal_871 ;
    wire signal_872 ;
    wire signal_873 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_879 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_885 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_888 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_891 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_894 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_897 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_900 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_903 ;
    wire signal_904 ;
    wire signal_905 ;
    wire signal_906 ;
    wire signal_907 ;
    wire signal_908 ;
    wire signal_909 ;
    wire signal_910 ;
    wire signal_911 ;
    wire signal_912 ;
    wire signal_913 ;
    wire signal_914 ;
    wire signal_915 ;
    wire signal_916 ;
    wire signal_917 ;
    wire signal_918 ;
    wire signal_919 ;
    wire signal_920 ;
    wire signal_921 ;
    wire signal_922 ;
    wire signal_923 ;
    wire signal_924 ;
    wire signal_925 ;
    wire signal_926 ;
    wire signal_927 ;
    wire signal_928 ;
    wire signal_929 ;
    wire signal_930 ;
    wire signal_931 ;
    wire signal_932 ;
    wire signal_933 ;
    wire signal_934 ;
    wire signal_935 ;
    wire signal_936 ;
    wire signal_937 ;
    wire signal_938 ;
    wire signal_939 ;
    wire signal_940 ;
    wire signal_941 ;
    wire signal_942 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1021 ;
    wire signal_1024 ;
    wire signal_1027 ;
    wire signal_1030 ;
    wire signal_1033 ;
    wire signal_1036 ;
    wire signal_1039 ;
    wire signal_1042 ;
    wire signal_1045 ;
    wire signal_1048 ;
    wire signal_1051 ;
    wire signal_1054 ;
    wire signal_1057 ;
    wire signal_1060 ;
    wire signal_1063 ;
    wire signal_1066 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1196 ;
    wire signal_1198 ;
    wire signal_1200 ;
    wire signal_1202 ;
    wire signal_1204 ;
    wire signal_1206 ;
    wire signal_1208 ;
    wire signal_1210 ;
    wire signal_1212 ;
    wire signal_1214 ;
    wire signal_1216 ;
    wire signal_1218 ;
    wire signal_1220 ;
    wire signal_1222 ;
    wire signal_1224 ;
    wire signal_1226 ;
    wire signal_1228 ;
    wire signal_1230 ;
    wire signal_1232 ;
    wire signal_1234 ;
    wire signal_1236 ;
    wire signal_1238 ;
    wire signal_1240 ;
    wire signal_1242 ;
    wire signal_1244 ;
    wire signal_1246 ;
    wire signal_1248 ;
    wire signal_1250 ;
    wire signal_1252 ;
    wire signal_1254 ;
    wire signal_1256 ;
    wire signal_1258 ;
    wire signal_1260 ;
    wire signal_1262 ;
    wire signal_1264 ;
    wire signal_1266 ;
    wire signal_1268 ;
    wire signal_1270 ;
    wire signal_1272 ;
    wire signal_1274 ;
    wire signal_1276 ;
    wire signal_1278 ;
    wire signal_1280 ;
    wire signal_1282 ;
    wire signal_1284 ;
    wire signal_1286 ;
    wire signal_1288 ;
    wire signal_1290 ;
    wire signal_1292 ;
    wire signal_1294 ;
    wire signal_1296 ;
    wire signal_1298 ;
    wire signal_1300 ;
    wire signal_1302 ;
    wire signal_1304 ;
    wire signal_1306 ;
    wire signal_1308 ;
    wire signal_1310 ;
    wire signal_1312 ;
    wire signal_1314 ;
    wire signal_1316 ;
    wire signal_1318 ;
    wire signal_1320 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1405 ;
    wire signal_1408 ;
    wire signal_1411 ;
    wire signal_1414 ;
    wire signal_1417 ;
    wire signal_1420 ;
    wire signal_1423 ;
    wire signal_1426 ;
    wire signal_1429 ;
    wire signal_1432 ;
    wire signal_1435 ;
    wire signal_1438 ;
    wire signal_1441 ;
    wire signal_1444 ;
    wire signal_1447 ;
    wire signal_1450 ;
    wire signal_1453 ;
    wire signal_1456 ;
    wire signal_1459 ;
    wire signal_1462 ;
    wire signal_1465 ;
    wire signal_1468 ;
    wire signal_1471 ;
    wire signal_1474 ;
    wire signal_1477 ;
    wire signal_1480 ;
    wire signal_1483 ;
    wire signal_1486 ;
    wire signal_1489 ;
    wire signal_1492 ;
    wire signal_1495 ;
    wire signal_1498 ;
    wire signal_1501 ;
    wire signal_1504 ;
    wire signal_1507 ;
    wire signal_1510 ;
    wire signal_1513 ;
    wire signal_1516 ;
    wire signal_1519 ;
    wire signal_1522 ;
    wire signal_1525 ;
    wire signal_1528 ;
    wire signal_1531 ;
    wire signal_1534 ;
    wire signal_1537 ;
    wire signal_1540 ;
    wire signal_1543 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1564 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1623 ;
    wire signal_1624 ;
    wire signal_1625 ;
    wire signal_1626 ;
    wire signal_1627 ;
    wire signal_1628 ;
    wire signal_1629 ;
    wire signal_1630 ;
    wire signal_1631 ;
    wire signal_1632 ;
    wire signal_1633 ;
    wire signal_1634 ;
    wire signal_1635 ;
    wire signal_1636 ;
    wire signal_1637 ;
    wire signal_1638 ;
    wire signal_1639 ;
    wire signal_1640 ;
    wire signal_1641 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1657 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1660 ;
    wire signal_1661 ;
    wire signal_1662 ;
    wire signal_1663 ;
    wire signal_1664 ;
    wire signal_1665 ;
    wire signal_1666 ;
    wire signal_1667 ;
    wire signal_1668 ;
    wire signal_1669 ;
    wire signal_1670 ;
    wire signal_1671 ;
    wire signal_1672 ;
    wire signal_1673 ;
    wire signal_1674 ;
    wire signal_1675 ;
    wire signal_1676 ;
    wire signal_1677 ;
    wire signal_1678 ;
    wire signal_1679 ;
    wire signal_1680 ;
    wire signal_1681 ;
    wire signal_1682 ;
    wire signal_1747 ;
    wire signal_1748 ;
    wire signal_1749 ;
    wire signal_1750 ;
    wire signal_1751 ;
    wire signal_1752 ;
    wire signal_1753 ;
    wire signal_1754 ;
    wire signal_1755 ;
    wire signal_1756 ;
    wire signal_1757 ;
    wire signal_1758 ;
    wire signal_1759 ;
    wire signal_1760 ;
    wire signal_1761 ;
    wire signal_1762 ;
    wire signal_1763 ;
    wire signal_1764 ;
    wire signal_1765 ;
    wire signal_1766 ;
    wire signal_1767 ;
    wire signal_1768 ;
    wire signal_1769 ;
    wire signal_1770 ;
    wire signal_1771 ;
    wire signal_1772 ;
    wire signal_1773 ;
    wire signal_1774 ;
    wire signal_1775 ;
    wire signal_1776 ;
    wire signal_1777 ;
    wire signal_1778 ;
    wire signal_1779 ;
    wire signal_1780 ;
    wire signal_1781 ;
    wire signal_1782 ;
    wire signal_1783 ;
    wire signal_1784 ;
    wire signal_1785 ;
    wire signal_1786 ;
    wire signal_1787 ;
    wire signal_1788 ;
    wire signal_1789 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1792 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1795 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1813 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1844 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1854 ;
    wire signal_1855 ;
    wire signal_1856 ;
    wire signal_1857 ;
    wire signal_1858 ;
    wire signal_1859 ;
    wire signal_1860 ;
    wire signal_1861 ;
    wire signal_1862 ;
    wire signal_1863 ;
    wire signal_1864 ;
    wire signal_1865 ;
    wire signal_1866 ;
    wire signal_1867 ;
    wire signal_1868 ;
    wire signal_1869 ;
    wire signal_1870 ;
    wire signal_1871 ;
    wire signal_1872 ;
    wire signal_1873 ;
    wire signal_1874 ;
    wire signal_1875 ;
    wire signal_1876 ;
    wire signal_1877 ;
    wire signal_1878 ;
    wire signal_1879 ;
    wire signal_1880 ;
    wire signal_1881 ;
    wire signal_1882 ;
    wire signal_1883 ;
    wire signal_1884 ;
    wire signal_1885 ;
    wire signal_1886 ;
    wire signal_1887 ;
    wire signal_1888 ;
    wire signal_1889 ;
    wire signal_1890 ;
    wire signal_1891 ;
    wire signal_1892 ;
    wire signal_1893 ;
    wire signal_1894 ;
    wire signal_1895 ;
    wire signal_1896 ;
    wire signal_1897 ;
    wire signal_1898 ;
    wire signal_1899 ;
    wire signal_1900 ;
    wire signal_1901 ;
    wire signal_1902 ;
    wire signal_1903 ;
    wire signal_1904 ;
    wire signal_1905 ;
    wire signal_1906 ;
    wire signal_1907 ;
    wire signal_1908 ;
    wire signal_1909 ;
    wire signal_1910 ;
    wire signal_1911 ;
    wire signal_1912 ;
    wire signal_1913 ;
    wire signal_1914 ;
    wire signal_1915 ;
    wire signal_1916 ;
    wire signal_1917 ;
    wire signal_1918 ;
    wire signal_1919 ;
    wire signal_1920 ;
    wire signal_1921 ;
    wire signal_1922 ;
    wire signal_1923 ;
    wire signal_1924 ;
    wire signal_1925 ;
    wire signal_1926 ;
    wire signal_1927 ;
    wire signal_1928 ;
    wire signal_1929 ;
    wire signal_1930 ;
    wire signal_1931 ;
    wire signal_1932 ;
    wire signal_1933 ;
    wire signal_1934 ;
    wire signal_1935 ;
    wire signal_1936 ;
    wire signal_1937 ;
    wire signal_1938 ;
    wire signal_1939 ;
    wire signal_1940 ;
    wire signal_1941 ;
    wire signal_1942 ;
    wire signal_1943 ;
    wire signal_1944 ;
    wire signal_1945 ;
    wire signal_1946 ;
    wire signal_1947 ;
    wire signal_1948 ;
    wire signal_1949 ;
    wire signal_1950 ;
    wire signal_1951 ;
    wire signal_1952 ;
    wire signal_1953 ;
    wire signal_1954 ;
    wire signal_1955 ;
    wire signal_1956 ;
    wire signal_1957 ;
    wire signal_1958 ;
    wire signal_1959 ;
    wire signal_1960 ;
    wire signal_1961 ;
    wire signal_1962 ;
    wire signal_1963 ;
    wire signal_1964 ;
    wire signal_1965 ;
    wire signal_1966 ;
    wire signal_1967 ;
    wire signal_1968 ;
    wire signal_1969 ;
    wire signal_1970 ;
    wire signal_1971 ;
    wire signal_1972 ;
    wire signal_1973 ;
    wire signal_1974 ;
    wire signal_1975 ;
    wire signal_1976 ;
    wire signal_1977 ;
    wire signal_1978 ;
    wire signal_1979 ;
    wire signal_1980 ;
    wire signal_1981 ;
    wire signal_1982 ;
    wire signal_1983 ;
    wire signal_1984 ;
    wire signal_1985 ;
    wire signal_1986 ;
    wire signal_1987 ;
    wire signal_1988 ;
    wire signal_1989 ;
    wire signal_1990 ;
    wire signal_1991 ;
    wire signal_1992 ;
    wire signal_1993 ;
    wire signal_1994 ;
    wire signal_1995 ;
    wire signal_1996 ;
    wire signal_1997 ;
    wire signal_1998 ;
    wire signal_1999 ;
    wire signal_2000 ;
    wire signal_2001 ;
    wire signal_2002 ;
    wire signal_2003 ;
    wire signal_2004 ;
    wire signal_2005 ;
    wire signal_2006 ;
    wire signal_2007 ;
    wire signal_2008 ;
    wire signal_2009 ;
    wire signal_2010 ;
    wire signal_2011 ;
    wire signal_2012 ;
    wire signal_2013 ;
    wire signal_2014 ;
    wire signal_2015 ;
    wire signal_2016 ;
    wire signal_2017 ;
    wire signal_2018 ;
    wire signal_2019 ;
    wire signal_2020 ;
    wire signal_2021 ;
    wire signal_2022 ;
    wire signal_2023 ;
    wire signal_2024 ;
    wire signal_2025 ;
    wire signal_2026 ;
    wire signal_2027 ;
    wire signal_2028 ;
    wire signal_2029 ;
    wire signal_2030 ;
    wire signal_2031 ;
    wire signal_2032 ;
    wire signal_2033 ;
    wire signal_2034 ;
    wire signal_2035 ;
    wire signal_2036 ;
    wire signal_2037 ;
    wire signal_2038 ;
    wire signal_2039 ;
    wire signal_2040 ;
    wire signal_2041 ;
    wire signal_2042 ;
    wire signal_2043 ;
    wire signal_2044 ;
    wire signal_2045 ;
    wire signal_2046 ;
    wire signal_2047 ;
    wire signal_2048 ;
    wire signal_2049 ;
    wire signal_2050 ;
    wire signal_2051 ;
    wire signal_2052 ;
    wire signal_2053 ;
    wire signal_2054 ;
    wire signal_2055 ;
    wire signal_2056 ;
    wire signal_2057 ;
    wire signal_2058 ;
    wire signal_2059 ;
    wire signal_2060 ;
    wire signal_2061 ;
    wire signal_2062 ;
    wire signal_2063 ;
    wire signal_2064 ;
    wire signal_2065 ;
    wire signal_2066 ;
    wire signal_2067 ;
    wire signal_2068 ;
    wire signal_2069 ;
    wire signal_2070 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2079 ;
    wire signal_2080 ;
    wire signal_2081 ;
    wire signal_2082 ;
    wire signal_2083 ;
    wire signal_2084 ;
    wire signal_2085 ;
    wire signal_2086 ;
    wire signal_2087 ;
    wire signal_2088 ;
    wire signal_2089 ;
    wire signal_2090 ;
    wire signal_2091 ;
    wire signal_2092 ;
    wire signal_2093 ;
    wire signal_2094 ;
    wire signal_2095 ;
    wire signal_2096 ;
    wire signal_2097 ;
    wire signal_2098 ;
    wire signal_2099 ;
    wire signal_2100 ;
    wire signal_2101 ;
    wire signal_2102 ;
    wire signal_2103 ;
    wire signal_2104 ;
    wire signal_2105 ;
    wire signal_2106 ;
    wire signal_2107 ;
    wire signal_2108 ;
    wire signal_2109 ;
    wire signal_2110 ;
    wire signal_2111 ;
    wire signal_2112 ;
    wire signal_2113 ;
    wire signal_2114 ;
    wire signal_2115 ;
    wire signal_2116 ;
    wire signal_2117 ;
    wire signal_2118 ;
    wire signal_2119 ;
    wire signal_2120 ;
    wire signal_2121 ;
    wire signal_2122 ;
    wire signal_2123 ;
    wire signal_2124 ;
    wire signal_2125 ;
    wire signal_2126 ;
    wire signal_2127 ;
    wire signal_2128 ;
    wire signal_2129 ;
    wire signal_2130 ;
    wire signal_2131 ;
    wire signal_2132 ;
    wire signal_2133 ;
    wire signal_2134 ;
    wire signal_2135 ;
    wire signal_2136 ;
    wire signal_2137 ;
    wire signal_2138 ;
    wire signal_2139 ;
    wire signal_2140 ;
    wire signal_2141 ;
    wire signal_2142 ;
    wire signal_2143 ;
    wire signal_2144 ;
    wire signal_2145 ;
    wire signal_2146 ;
    wire signal_2147 ;
    wire signal_2148 ;
    wire signal_2149 ;
    wire signal_2150 ;
    wire signal_2151 ;
    wire signal_2152 ;
    wire signal_2153 ;
    wire signal_2154 ;
    wire signal_2155 ;
    wire signal_2156 ;
    wire signal_2157 ;
    wire signal_2158 ;
    wire signal_2159 ;
    wire signal_2160 ;
    wire signal_2161 ;
    wire signal_2162 ;
    wire signal_2163 ;
    wire signal_2164 ;
    wire signal_2165 ;
    wire signal_2166 ;
    wire signal_2167 ;
    wire signal_2168 ;
    wire signal_2169 ;
    wire signal_2170 ;
    wire signal_2171 ;
    wire signal_2172 ;
    wire signal_2173 ;
    wire signal_2174 ;
    wire signal_2175 ;
    wire signal_2176 ;
    wire signal_2177 ;
    wire signal_2178 ;
    wire signal_2179 ;
    wire signal_2180 ;
    wire signal_2181 ;
    wire signal_2182 ;
    wire signal_2183 ;
    wire signal_2184 ;
    wire signal_2185 ;
    wire signal_2186 ;
    wire signal_2187 ;
    wire signal_2188 ;
    wire signal_2189 ;
    wire signal_2190 ;
    wire signal_2191 ;
    wire signal_2192 ;
    wire signal_2193 ;
    wire signal_2194 ;
    wire signal_2195 ;
    wire signal_2196 ;
    wire signal_2197 ;
    wire signal_2198 ;
    wire signal_2199 ;
    wire signal_2200 ;
    wire signal_2201 ;
    wire signal_2202 ;
    wire signal_2203 ;
    wire signal_2204 ;
    wire signal_2205 ;
    wire signal_2206 ;
    wire signal_2207 ;
    wire signal_2208 ;
    wire signal_2209 ;
    wire signal_2210 ;
    wire signal_2211 ;
    wire signal_2212 ;
    wire signal_2213 ;
    wire signal_2214 ;
    wire signal_2215 ;
    wire signal_2216 ;
    wire signal_2217 ;
    wire signal_2218 ;
    wire signal_2219 ;
    wire signal_2220 ;
    wire signal_2221 ;
    wire signal_2222 ;
    wire signal_2223 ;
    wire signal_2224 ;
    wire signal_2225 ;
    wire signal_2226 ;
    wire signal_2227 ;
    wire signal_2228 ;
    wire signal_2229 ;
    wire signal_2230 ;
    wire signal_2231 ;
    wire signal_2232 ;
    wire signal_2233 ;
    wire signal_2234 ;
    wire signal_2235 ;
    wire signal_2236 ;
    wire signal_2237 ;
    wire signal_2238 ;
    wire signal_2239 ;
    wire signal_2240 ;
    wire signal_2241 ;
    wire signal_2242 ;
    wire signal_2243 ;
    wire signal_2244 ;
    wire signal_2245 ;
    wire signal_2246 ;
    wire signal_2247 ;
    wire signal_2248 ;
    wire signal_2249 ;
    wire signal_2250 ;
    wire signal_2251 ;
    wire signal_2252 ;
    wire signal_2253 ;
    wire signal_2254 ;
    wire signal_2255 ;
    wire signal_2256 ;
    wire signal_2257 ;
    wire signal_2258 ;
    wire signal_2259 ;
    wire signal_2260 ;
    wire signal_2261 ;
    wire signal_2262 ;
    wire signal_2263 ;
    wire signal_2264 ;
    wire signal_2265 ;
    wire signal_2266 ;
    wire signal_2267 ;
    wire signal_2268 ;
    wire signal_2269 ;
    wire signal_2270 ;
    wire signal_2271 ;
    wire signal_2272 ;
    wire signal_2273 ;
    wire signal_2274 ;
    wire signal_2275 ;
    wire signal_2276 ;
    wire signal_2277 ;
    wire signal_2278 ;
    wire signal_2279 ;
    wire signal_2280 ;

    /* cells in depth 0 */
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_177 ( .a ({signal_1492, signal_894}), .b ({1'b0, signal_266}), .c ({signal_1579, signal_333}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_180 ( .a ({signal_1495, signal_893}), .b ({1'b0, signal_1014}), .c ({signal_1580, signal_335}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_183 ( .a ({signal_1498, signal_892}), .b ({1'b0, signal_1013}), .c ({signal_1581, signal_337}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_186 ( .a ({signal_1501, signal_891}), .b ({1'b0, 1'b0}), .c ({signal_1582, signal_339}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_189 ( .a ({signal_1504, signal_890}), .b ({1'b0, signal_265}), .c ({signal_1583, signal_341}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_192 ( .a ({signal_1507, signal_889}), .b ({1'b0, signal_1011}), .c ({signal_1584, signal_343}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_195 ( .a ({signal_1510, signal_888}), .b ({1'b0, signal_1010}), .c ({signal_1585, signal_345}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_198 ( .a ({signal_1513, signal_887}), .b ({1'b0, signal_1009}), .c ({signal_1586, signal_347}) ) ;
    INV_X1 cell_712 ( .A (signal_1000), .ZN (signal_692) ) ;
    INV_X1 cell_713 ( .A (signal_692), .ZN (signal_693) ) ;
    INV_X1 cell_714 ( .A (signal_692), .ZN (signal_694) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_715 ( .s (signal_1000), .b ({key_s1[64], key_s0[64]}), .a ({key_s1[0], key_s0[0]}), .c ({signal_1021, signal_934}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_716 ( .s (signal_693), .b ({key_s1[65], key_s0[65]}), .a ({key_s1[1], key_s0[1]}), .c ({signal_1405, signal_933}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_717 ( .s (signal_1000), .b ({key_s1[66], key_s0[66]}), .a ({key_s1[2], key_s0[2]}), .c ({signal_1024, signal_932}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_718 ( .s (signal_693), .b ({key_s1[67], key_s0[67]}), .a ({key_s1[3], key_s0[3]}), .c ({signal_1408, signal_931}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_719 ( .s (signal_693), .b ({key_s1[68], key_s0[68]}), .a ({key_s1[4], key_s0[4]}), .c ({signal_1411, signal_930}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_720 ( .s (signal_693), .b ({key_s1[69], key_s0[69]}), .a ({key_s1[5], key_s0[5]}), .c ({signal_1414, signal_929}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_721 ( .s (signal_693), .b ({key_s1[70], key_s0[70]}), .a ({key_s1[6], key_s0[6]}), .c ({signal_1417, signal_928}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_722 ( .s (signal_693), .b ({key_s1[71], key_s0[71]}), .a ({key_s1[7], key_s0[7]}), .c ({signal_1420, signal_927}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_723 ( .s (signal_693), .b ({key_s1[72], key_s0[72]}), .a ({key_s1[8], key_s0[8]}), .c ({signal_1423, signal_926}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_724 ( .s (signal_693), .b ({key_s1[73], key_s0[73]}), .a ({key_s1[9], key_s0[9]}), .c ({signal_1426, signal_925}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_725 ( .s (signal_693), .b ({key_s1[74], key_s0[74]}), .a ({key_s1[10], key_s0[10]}), .c ({signal_1429, signal_924}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_726 ( .s (signal_693), .b ({key_s1[75], key_s0[75]}), .a ({key_s1[11], key_s0[11]}), .c ({signal_1432, signal_923}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_727 ( .s (signal_693), .b ({key_s1[76], key_s0[76]}), .a ({key_s1[12], key_s0[12]}), .c ({signal_1435, signal_922}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_728 ( .s (signal_693), .b ({key_s1[77], key_s0[77]}), .a ({key_s1[13], key_s0[13]}), .c ({signal_1438, signal_921}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_729 ( .s (signal_693), .b ({key_s1[78], key_s0[78]}), .a ({key_s1[14], key_s0[14]}), .c ({signal_1441, signal_920}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_730 ( .s (signal_693), .b ({key_s1[79], key_s0[79]}), .a ({key_s1[15], key_s0[15]}), .c ({signal_1444, signal_919}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_731 ( .s (signal_693), .b ({key_s1[80], key_s0[80]}), .a ({key_s1[16], key_s0[16]}), .c ({signal_1447, signal_918}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_732 ( .s (signal_693), .b ({key_s1[81], key_s0[81]}), .a ({key_s1[17], key_s0[17]}), .c ({signal_1450, signal_917}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_733 ( .s (signal_693), .b ({key_s1[82], key_s0[82]}), .a ({key_s1[18], key_s0[18]}), .c ({signal_1453, signal_916}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_734 ( .s (signal_693), .b ({key_s1[83], key_s0[83]}), .a ({key_s1[19], key_s0[19]}), .c ({signal_1456, signal_915}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_735 ( .s (signal_693), .b ({key_s1[84], key_s0[84]}), .a ({key_s1[20], key_s0[20]}), .c ({signal_1459, signal_914}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_736 ( .s (signal_693), .b ({key_s1[85], key_s0[85]}), .a ({key_s1[21], key_s0[21]}), .c ({signal_1462, signal_913}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_737 ( .s (signal_1000), .b ({key_s1[86], key_s0[86]}), .a ({key_s1[22], key_s0[22]}), .c ({signal_1027, signal_912}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_738 ( .s (signal_1000), .b ({key_s1[87], key_s0[87]}), .a ({key_s1[23], key_s0[23]}), .c ({signal_1030, signal_911}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_739 ( .s (signal_1000), .b ({key_s1[88], key_s0[88]}), .a ({key_s1[24], key_s0[24]}), .c ({signal_1033, signal_910}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_740 ( .s (signal_1000), .b ({key_s1[89], key_s0[89]}), .a ({key_s1[25], key_s0[25]}), .c ({signal_1036, signal_909}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_741 ( .s (signal_1000), .b ({key_s1[90], key_s0[90]}), .a ({key_s1[26], key_s0[26]}), .c ({signal_1039, signal_908}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_742 ( .s (signal_1000), .b ({key_s1[91], key_s0[91]}), .a ({key_s1[27], key_s0[27]}), .c ({signal_1042, signal_907}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_743 ( .s (signal_694), .b ({key_s1[92], key_s0[92]}), .a ({key_s1[28], key_s0[28]}), .c ({signal_1465, signal_906}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_744 ( .s (signal_694), .b ({key_s1[93], key_s0[93]}), .a ({key_s1[29], key_s0[29]}), .c ({signal_1468, signal_905}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_745 ( .s (signal_694), .b ({key_s1[94], key_s0[94]}), .a ({key_s1[30], key_s0[30]}), .c ({signal_1471, signal_904}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_746 ( .s (signal_694), .b ({key_s1[95], key_s0[95]}), .a ({key_s1[31], key_s0[31]}), .c ({signal_1474, signal_903}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_747 ( .s (signal_694), .b ({key_s1[96], key_s0[96]}), .a ({key_s1[32], key_s0[32]}), .c ({signal_1477, signal_902}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_748 ( .s (signal_1000), .b ({key_s1[97], key_s0[97]}), .a ({key_s1[33], key_s0[33]}), .c ({signal_1045, signal_901}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_749 ( .s (signal_694), .b ({key_s1[98], key_s0[98]}), .a ({key_s1[34], key_s0[34]}), .c ({signal_1480, signal_900}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_750 ( .s (signal_694), .b ({key_s1[99], key_s0[99]}), .a ({key_s1[35], key_s0[35]}), .c ({signal_1483, signal_899}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_751 ( .s (signal_1000), .b ({key_s1[100], key_s0[100]}), .a ({key_s1[36], key_s0[36]}), .c ({signal_1048, signal_898}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_752 ( .s (signal_694), .b ({key_s1[101], key_s0[101]}), .a ({key_s1[37], key_s0[37]}), .c ({signal_1486, signal_897}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_753 ( .s (signal_694), .b ({key_s1[102], key_s0[102]}), .a ({key_s1[38], key_s0[38]}), .c ({signal_1489, signal_896}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_754 ( .s (signal_1000), .b ({key_s1[103], key_s0[103]}), .a ({key_s1[39], key_s0[39]}), .c ({signal_1051, signal_895}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_755 ( .s (signal_694), .b ({key_s1[104], key_s0[104]}), .a ({key_s1[40], key_s0[40]}), .c ({signal_1492, signal_894}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_756 ( .s (signal_694), .b ({key_s1[105], key_s0[105]}), .a ({key_s1[41], key_s0[41]}), .c ({signal_1495, signal_893}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_757 ( .s (signal_694), .b ({key_s1[106], key_s0[106]}), .a ({key_s1[42], key_s0[42]}), .c ({signal_1498, signal_892}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_758 ( .s (signal_694), .b ({key_s1[107], key_s0[107]}), .a ({key_s1[43], key_s0[43]}), .c ({signal_1501, signal_891}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_759 ( .s (signal_694), .b ({key_s1[108], key_s0[108]}), .a ({key_s1[44], key_s0[44]}), .c ({signal_1504, signal_890}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_760 ( .s (signal_694), .b ({key_s1[109], key_s0[109]}), .a ({key_s1[45], key_s0[45]}), .c ({signal_1507, signal_889}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_761 ( .s (signal_694), .b ({key_s1[110], key_s0[110]}), .a ({key_s1[46], key_s0[46]}), .c ({signal_1510, signal_888}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_762 ( .s (signal_694), .b ({key_s1[111], key_s0[111]}), .a ({key_s1[47], key_s0[47]}), .c ({signal_1513, signal_887}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_763 ( .s (signal_694), .b ({key_s1[112], key_s0[112]}), .a ({key_s1[48], key_s0[48]}), .c ({signal_1516, signal_886}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_764 ( .s (signal_694), .b ({key_s1[113], key_s0[113]}), .a ({key_s1[49], key_s0[49]}), .c ({signal_1519, signal_885}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_765 ( .s (signal_694), .b ({key_s1[114], key_s0[114]}), .a ({key_s1[50], key_s0[50]}), .c ({signal_1522, signal_884}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_766 ( .s (signal_694), .b ({key_s1[115], key_s0[115]}), .a ({key_s1[51], key_s0[51]}), .c ({signal_1525, signal_883}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_767 ( .s (signal_694), .b ({key_s1[116], key_s0[116]}), .a ({key_s1[52], key_s0[52]}), .c ({signal_1528, signal_882}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_768 ( .s (signal_1000), .b ({key_s1[117], key_s0[117]}), .a ({key_s1[53], key_s0[53]}), .c ({signal_1054, signal_881}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_769 ( .s (signal_1000), .b ({key_s1[118], key_s0[118]}), .a ({key_s1[54], key_s0[54]}), .c ({signal_1057, signal_880}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_770 ( .s (signal_694), .b ({key_s1[119], key_s0[119]}), .a ({key_s1[55], key_s0[55]}), .c ({signal_1531, signal_879}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_771 ( .s (signal_1000), .b ({key_s1[120], key_s0[120]}), .a ({key_s1[56], key_s0[56]}), .c ({signal_1060, signal_878}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_772 ( .s (signal_694), .b ({key_s1[121], key_s0[121]}), .a ({key_s1[57], key_s0[57]}), .c ({signal_1534, signal_877}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_773 ( .s (signal_694), .b ({key_s1[122], key_s0[122]}), .a ({key_s1[58], key_s0[58]}), .c ({signal_1537, signal_876}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_774 ( .s (signal_1000), .b ({key_s1[123], key_s0[123]}), .a ({key_s1[59], key_s0[59]}), .c ({signal_1063, signal_875}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_775 ( .s (signal_694), .b ({key_s1[124], key_s0[124]}), .a ({key_s1[60], key_s0[60]}), .c ({signal_1540, signal_874}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_776 ( .s (signal_694), .b ({key_s1[125], key_s0[125]}), .a ({key_s1[61], key_s0[61]}), .c ({signal_1543, signal_873}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_777 ( .s (signal_1000), .b ({key_s1[126], key_s0[126]}), .a ({key_s1[62], key_s0[62]}), .c ({signal_1066, signal_872}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_778 ( .s (signal_694), .b ({key_s1[127], key_s0[127]}), .a ({key_s1[63], key_s0[63]}), .c ({signal_1546, signal_871}) ) ;
    MUX2_X1 cell_779 ( .S (rst), .A (signal_1007), .B (1'b1), .Z (signal_266) ) ;
    MUX2_X1 cell_780 ( .S (rst), .A (signal_1006), .B (1'b0), .Z (signal_1014) ) ;
    MUX2_X1 cell_781 ( .S (rst), .A (signal_1005), .B (1'b0), .Z (signal_1013) ) ;
    MUX2_X1 cell_782 ( .S (rst), .A (signal_1004), .B (1'b1), .Z (signal_265) ) ;
    MUX2_X1 cell_783 ( .S (rst), .A (signal_1003), .B (1'b0), .Z (signal_1011) ) ;
    MUX2_X1 cell_784 ( .S (rst), .A (signal_1002), .B (1'b0), .Z (signal_1010) ) ;
    MUX2_X1 cell_785 ( .S (rst), .A (signal_1001), .B (1'b0), .Z (signal_1009) ) ;
    XOR2_X1 cell_786 ( .A (signal_265), .B (signal_1011), .Z (signal_1008) ) ;
    XOR2_X1 cell_787 ( .A (signal_1014), .B (signal_266), .Z (signal_1012) ) ;
    AND2_X1 cell_802 ( .A1 (signal_1009), .A2 (signal_702), .ZN (signal_267) ) ;
    NOR2_X1 cell_803 ( .A1 (signal_703), .A2 (signal_704), .ZN (signal_702) ) ;
    NAND2_X1 cell_804 ( .A1 (signal_705), .A2 (signal_706), .ZN (signal_704) ) ;
    NOR2_X1 cell_805 ( .A1 (signal_1011), .A2 (signal_1010), .ZN (signal_706) ) ;
    NOR2_X1 cell_806 ( .A1 (signal_1014), .A2 (signal_265), .ZN (signal_705) ) ;
    NAND2_X1 cell_807 ( .A1 (signal_266), .A2 (signal_1013), .ZN (signal_703) ) ;
    MUX2_X1 cell_808 ( .S (rst), .A (signal_1016), .B (1'b0), .Z (signal_1000) ) ;
    MUX2_X1 cell_809 ( .S (rst), .A (signal_1015), .B (1'b0), .Z (signal_999) ) ;
    XNOR2_X1 cell_810 ( .A (signal_707), .B (signal_999), .ZN (signal_1017) ) ;
    XNOR2_X1 cell_811 ( .A (signal_1000), .B (1'b0), .ZN (signal_707) ) ;
    INV_X1 cell_812 ( .A (signal_1000), .ZN (signal_1018) ) ;

    /* cells in depth 1 */
    buf_clk cell_820 ( .C (clk), .D (rst), .Q (signal_1747) ) ;
    buf_clk cell_822 ( .C (clk), .D (plaintext_s0[0]), .Q (signal_1749) ) ;
    buf_clk cell_824 ( .C (clk), .D (plaintext_s1[0]), .Q (signal_1751) ) ;
    buf_clk cell_826 ( .C (clk), .D (plaintext_s0[1]), .Q (signal_1753) ) ;
    buf_clk cell_828 ( .C (clk), .D (plaintext_s1[1]), .Q (signal_1755) ) ;
    buf_clk cell_830 ( .C (clk), .D (plaintext_s0[2]), .Q (signal_1757) ) ;
    buf_clk cell_832 ( .C (clk), .D (plaintext_s1[2]), .Q (signal_1759) ) ;
    buf_clk cell_834 ( .C (clk), .D (plaintext_s0[3]), .Q (signal_1761) ) ;
    buf_clk cell_836 ( .C (clk), .D (plaintext_s1[3]), .Q (signal_1763) ) ;
    buf_clk cell_838 ( .C (clk), .D (plaintext_s0[4]), .Q (signal_1765) ) ;
    buf_clk cell_840 ( .C (clk), .D (plaintext_s1[4]), .Q (signal_1767) ) ;
    buf_clk cell_842 ( .C (clk), .D (plaintext_s0[5]), .Q (signal_1769) ) ;
    buf_clk cell_844 ( .C (clk), .D (plaintext_s1[5]), .Q (signal_1771) ) ;
    buf_clk cell_846 ( .C (clk), .D (plaintext_s0[6]), .Q (signal_1773) ) ;
    buf_clk cell_848 ( .C (clk), .D (plaintext_s1[6]), .Q (signal_1775) ) ;
    buf_clk cell_850 ( .C (clk), .D (plaintext_s0[7]), .Q (signal_1777) ) ;
    buf_clk cell_852 ( .C (clk), .D (plaintext_s1[7]), .Q (signal_1779) ) ;
    buf_clk cell_854 ( .C (clk), .D (plaintext_s0[8]), .Q (signal_1781) ) ;
    buf_clk cell_856 ( .C (clk), .D (plaintext_s1[8]), .Q (signal_1783) ) ;
    buf_clk cell_858 ( .C (clk), .D (plaintext_s0[9]), .Q (signal_1785) ) ;
    buf_clk cell_860 ( .C (clk), .D (plaintext_s1[9]), .Q (signal_1787) ) ;
    buf_clk cell_862 ( .C (clk), .D (plaintext_s0[10]), .Q (signal_1789) ) ;
    buf_clk cell_864 ( .C (clk), .D (plaintext_s1[10]), .Q (signal_1791) ) ;
    buf_clk cell_866 ( .C (clk), .D (plaintext_s0[11]), .Q (signal_1793) ) ;
    buf_clk cell_868 ( .C (clk), .D (plaintext_s1[11]), .Q (signal_1795) ) ;
    buf_clk cell_870 ( .C (clk), .D (plaintext_s0[12]), .Q (signal_1797) ) ;
    buf_clk cell_872 ( .C (clk), .D (plaintext_s1[12]), .Q (signal_1799) ) ;
    buf_clk cell_874 ( .C (clk), .D (plaintext_s0[13]), .Q (signal_1801) ) ;
    buf_clk cell_876 ( .C (clk), .D (plaintext_s1[13]), .Q (signal_1803) ) ;
    buf_clk cell_878 ( .C (clk), .D (plaintext_s0[14]), .Q (signal_1805) ) ;
    buf_clk cell_880 ( .C (clk), .D (plaintext_s1[14]), .Q (signal_1807) ) ;
    buf_clk cell_882 ( .C (clk), .D (plaintext_s0[15]), .Q (signal_1809) ) ;
    buf_clk cell_884 ( .C (clk), .D (plaintext_s1[15]), .Q (signal_1811) ) ;
    buf_clk cell_886 ( .C (clk), .D (plaintext_s0[16]), .Q (signal_1813) ) ;
    buf_clk cell_888 ( .C (clk), .D (plaintext_s1[16]), .Q (signal_1815) ) ;
    buf_clk cell_890 ( .C (clk), .D (plaintext_s0[17]), .Q (signal_1817) ) ;
    buf_clk cell_892 ( .C (clk), .D (plaintext_s1[17]), .Q (signal_1819) ) ;
    buf_clk cell_894 ( .C (clk), .D (plaintext_s0[18]), .Q (signal_1821) ) ;
    buf_clk cell_896 ( .C (clk), .D (plaintext_s1[18]), .Q (signal_1823) ) ;
    buf_clk cell_898 ( .C (clk), .D (plaintext_s0[19]), .Q (signal_1825) ) ;
    buf_clk cell_900 ( .C (clk), .D (plaintext_s1[19]), .Q (signal_1827) ) ;
    buf_clk cell_902 ( .C (clk), .D (plaintext_s0[20]), .Q (signal_1829) ) ;
    buf_clk cell_904 ( .C (clk), .D (plaintext_s1[20]), .Q (signal_1831) ) ;
    buf_clk cell_906 ( .C (clk), .D (plaintext_s0[21]), .Q (signal_1833) ) ;
    buf_clk cell_908 ( .C (clk), .D (plaintext_s1[21]), .Q (signal_1835) ) ;
    buf_clk cell_910 ( .C (clk), .D (plaintext_s0[22]), .Q (signal_1837) ) ;
    buf_clk cell_912 ( .C (clk), .D (plaintext_s1[22]), .Q (signal_1839) ) ;
    buf_clk cell_914 ( .C (clk), .D (plaintext_s0[23]), .Q (signal_1841) ) ;
    buf_clk cell_916 ( .C (clk), .D (plaintext_s1[23]), .Q (signal_1843) ) ;
    buf_clk cell_918 ( .C (clk), .D (plaintext_s0[24]), .Q (signal_1845) ) ;
    buf_clk cell_920 ( .C (clk), .D (plaintext_s1[24]), .Q (signal_1847) ) ;
    buf_clk cell_922 ( .C (clk), .D (plaintext_s0[25]), .Q (signal_1849) ) ;
    buf_clk cell_924 ( .C (clk), .D (plaintext_s1[25]), .Q (signal_1851) ) ;
    buf_clk cell_926 ( .C (clk), .D (plaintext_s0[26]), .Q (signal_1853) ) ;
    buf_clk cell_928 ( .C (clk), .D (plaintext_s1[26]), .Q (signal_1855) ) ;
    buf_clk cell_930 ( .C (clk), .D (plaintext_s0[27]), .Q (signal_1857) ) ;
    buf_clk cell_932 ( .C (clk), .D (plaintext_s1[27]), .Q (signal_1859) ) ;
    buf_clk cell_934 ( .C (clk), .D (plaintext_s0[28]), .Q (signal_1861) ) ;
    buf_clk cell_936 ( .C (clk), .D (plaintext_s1[28]), .Q (signal_1863) ) ;
    buf_clk cell_938 ( .C (clk), .D (plaintext_s0[29]), .Q (signal_1865) ) ;
    buf_clk cell_940 ( .C (clk), .D (plaintext_s1[29]), .Q (signal_1867) ) ;
    buf_clk cell_942 ( .C (clk), .D (plaintext_s0[30]), .Q (signal_1869) ) ;
    buf_clk cell_944 ( .C (clk), .D (plaintext_s1[30]), .Q (signal_1871) ) ;
    buf_clk cell_946 ( .C (clk), .D (plaintext_s0[31]), .Q (signal_1873) ) ;
    buf_clk cell_948 ( .C (clk), .D (plaintext_s1[31]), .Q (signal_1875) ) ;
    buf_clk cell_950 ( .C (clk), .D (plaintext_s0[32]), .Q (signal_1877) ) ;
    buf_clk cell_952 ( .C (clk), .D (plaintext_s1[32]), .Q (signal_1879) ) ;
    buf_clk cell_954 ( .C (clk), .D (plaintext_s0[33]), .Q (signal_1881) ) ;
    buf_clk cell_956 ( .C (clk), .D (plaintext_s1[33]), .Q (signal_1883) ) ;
    buf_clk cell_958 ( .C (clk), .D (plaintext_s0[34]), .Q (signal_1885) ) ;
    buf_clk cell_960 ( .C (clk), .D (plaintext_s1[34]), .Q (signal_1887) ) ;
    buf_clk cell_962 ( .C (clk), .D (plaintext_s0[35]), .Q (signal_1889) ) ;
    buf_clk cell_964 ( .C (clk), .D (plaintext_s1[35]), .Q (signal_1891) ) ;
    buf_clk cell_966 ( .C (clk), .D (plaintext_s0[36]), .Q (signal_1893) ) ;
    buf_clk cell_968 ( .C (clk), .D (plaintext_s1[36]), .Q (signal_1895) ) ;
    buf_clk cell_970 ( .C (clk), .D (plaintext_s0[37]), .Q (signal_1897) ) ;
    buf_clk cell_972 ( .C (clk), .D (plaintext_s1[37]), .Q (signal_1899) ) ;
    buf_clk cell_974 ( .C (clk), .D (plaintext_s0[38]), .Q (signal_1901) ) ;
    buf_clk cell_976 ( .C (clk), .D (plaintext_s1[38]), .Q (signal_1903) ) ;
    buf_clk cell_978 ( .C (clk), .D (plaintext_s0[39]), .Q (signal_1905) ) ;
    buf_clk cell_980 ( .C (clk), .D (plaintext_s1[39]), .Q (signal_1907) ) ;
    buf_clk cell_982 ( .C (clk), .D (plaintext_s0[40]), .Q (signal_1909) ) ;
    buf_clk cell_984 ( .C (clk), .D (plaintext_s1[40]), .Q (signal_1911) ) ;
    buf_clk cell_986 ( .C (clk), .D (plaintext_s0[41]), .Q (signal_1913) ) ;
    buf_clk cell_988 ( .C (clk), .D (plaintext_s1[41]), .Q (signal_1915) ) ;
    buf_clk cell_990 ( .C (clk), .D (plaintext_s0[42]), .Q (signal_1917) ) ;
    buf_clk cell_992 ( .C (clk), .D (plaintext_s1[42]), .Q (signal_1919) ) ;
    buf_clk cell_994 ( .C (clk), .D (plaintext_s0[43]), .Q (signal_1921) ) ;
    buf_clk cell_996 ( .C (clk), .D (plaintext_s1[43]), .Q (signal_1923) ) ;
    buf_clk cell_998 ( .C (clk), .D (plaintext_s0[44]), .Q (signal_1925) ) ;
    buf_clk cell_1000 ( .C (clk), .D (plaintext_s1[44]), .Q (signal_1927) ) ;
    buf_clk cell_1002 ( .C (clk), .D (plaintext_s0[45]), .Q (signal_1929) ) ;
    buf_clk cell_1004 ( .C (clk), .D (plaintext_s1[45]), .Q (signal_1931) ) ;
    buf_clk cell_1006 ( .C (clk), .D (plaintext_s0[46]), .Q (signal_1933) ) ;
    buf_clk cell_1008 ( .C (clk), .D (plaintext_s1[46]), .Q (signal_1935) ) ;
    buf_clk cell_1010 ( .C (clk), .D (plaintext_s0[47]), .Q (signal_1937) ) ;
    buf_clk cell_1012 ( .C (clk), .D (plaintext_s1[47]), .Q (signal_1939) ) ;
    buf_clk cell_1014 ( .C (clk), .D (plaintext_s0[48]), .Q (signal_1941) ) ;
    buf_clk cell_1016 ( .C (clk), .D (plaintext_s1[48]), .Q (signal_1943) ) ;
    buf_clk cell_1018 ( .C (clk), .D (plaintext_s0[49]), .Q (signal_1945) ) ;
    buf_clk cell_1020 ( .C (clk), .D (plaintext_s1[49]), .Q (signal_1947) ) ;
    buf_clk cell_1022 ( .C (clk), .D (plaintext_s0[50]), .Q (signal_1949) ) ;
    buf_clk cell_1024 ( .C (clk), .D (plaintext_s1[50]), .Q (signal_1951) ) ;
    buf_clk cell_1026 ( .C (clk), .D (plaintext_s0[51]), .Q (signal_1953) ) ;
    buf_clk cell_1028 ( .C (clk), .D (plaintext_s1[51]), .Q (signal_1955) ) ;
    buf_clk cell_1030 ( .C (clk), .D (plaintext_s0[52]), .Q (signal_1957) ) ;
    buf_clk cell_1032 ( .C (clk), .D (plaintext_s1[52]), .Q (signal_1959) ) ;
    buf_clk cell_1034 ( .C (clk), .D (plaintext_s0[53]), .Q (signal_1961) ) ;
    buf_clk cell_1036 ( .C (clk), .D (plaintext_s1[53]), .Q (signal_1963) ) ;
    buf_clk cell_1038 ( .C (clk), .D (plaintext_s0[54]), .Q (signal_1965) ) ;
    buf_clk cell_1040 ( .C (clk), .D (plaintext_s1[54]), .Q (signal_1967) ) ;
    buf_clk cell_1042 ( .C (clk), .D (plaintext_s0[55]), .Q (signal_1969) ) ;
    buf_clk cell_1044 ( .C (clk), .D (plaintext_s1[55]), .Q (signal_1971) ) ;
    buf_clk cell_1046 ( .C (clk), .D (plaintext_s0[56]), .Q (signal_1973) ) ;
    buf_clk cell_1048 ( .C (clk), .D (plaintext_s1[56]), .Q (signal_1975) ) ;
    buf_clk cell_1050 ( .C (clk), .D (plaintext_s0[57]), .Q (signal_1977) ) ;
    buf_clk cell_1052 ( .C (clk), .D (plaintext_s1[57]), .Q (signal_1979) ) ;
    buf_clk cell_1054 ( .C (clk), .D (plaintext_s0[58]), .Q (signal_1981) ) ;
    buf_clk cell_1056 ( .C (clk), .D (plaintext_s1[58]), .Q (signal_1983) ) ;
    buf_clk cell_1058 ( .C (clk), .D (plaintext_s0[59]), .Q (signal_1985) ) ;
    buf_clk cell_1060 ( .C (clk), .D (plaintext_s1[59]), .Q (signal_1987) ) ;
    buf_clk cell_1062 ( .C (clk), .D (plaintext_s0[60]), .Q (signal_1989) ) ;
    buf_clk cell_1064 ( .C (clk), .D (plaintext_s1[60]), .Q (signal_1991) ) ;
    buf_clk cell_1066 ( .C (clk), .D (plaintext_s0[61]), .Q (signal_1993) ) ;
    buf_clk cell_1068 ( .C (clk), .D (plaintext_s1[61]), .Q (signal_1995) ) ;
    buf_clk cell_1070 ( .C (clk), .D (plaintext_s0[62]), .Q (signal_1997) ) ;
    buf_clk cell_1072 ( .C (clk), .D (plaintext_s1[62]), .Q (signal_1999) ) ;
    buf_clk cell_1074 ( .C (clk), .D (plaintext_s0[63]), .Q (signal_2001) ) ;
    buf_clk cell_1076 ( .C (clk), .D (plaintext_s1[63]), .Q (signal_2003) ) ;
    buf_clk cell_1078 ( .C (clk), .D (signal_886), .Q (signal_2005) ) ;
    buf_clk cell_1080 ( .C (clk), .D (signal_1516), .Q (signal_2007) ) ;
    buf_clk cell_1082 ( .C (clk), .D (signal_885), .Q (signal_2009) ) ;
    buf_clk cell_1084 ( .C (clk), .D (signal_1519), .Q (signal_2011) ) ;
    buf_clk cell_1086 ( .C (clk), .D (signal_884), .Q (signal_2013) ) ;
    buf_clk cell_1088 ( .C (clk), .D (signal_1522), .Q (signal_2015) ) ;
    buf_clk cell_1090 ( .C (clk), .D (signal_883), .Q (signal_2017) ) ;
    buf_clk cell_1092 ( .C (clk), .D (signal_1525), .Q (signal_2019) ) ;
    buf_clk cell_1094 ( .C (clk), .D (signal_882), .Q (signal_2021) ) ;
    buf_clk cell_1096 ( .C (clk), .D (signal_1528), .Q (signal_2023) ) ;
    buf_clk cell_1098 ( .C (clk), .D (signal_881), .Q (signal_2025) ) ;
    buf_clk cell_1100 ( .C (clk), .D (signal_1054), .Q (signal_2027) ) ;
    buf_clk cell_1102 ( .C (clk), .D (signal_880), .Q (signal_2029) ) ;
    buf_clk cell_1104 ( .C (clk), .D (signal_1057), .Q (signal_2031) ) ;
    buf_clk cell_1106 ( .C (clk), .D (signal_879), .Q (signal_2033) ) ;
    buf_clk cell_1108 ( .C (clk), .D (signal_1531), .Q (signal_2035) ) ;
    buf_clk cell_1110 ( .C (clk), .D (signal_878), .Q (signal_2037) ) ;
    buf_clk cell_1112 ( .C (clk), .D (signal_1060), .Q (signal_2039) ) ;
    buf_clk cell_1114 ( .C (clk), .D (signal_877), .Q (signal_2041) ) ;
    buf_clk cell_1116 ( .C (clk), .D (signal_1534), .Q (signal_2043) ) ;
    buf_clk cell_1118 ( .C (clk), .D (signal_876), .Q (signal_2045) ) ;
    buf_clk cell_1120 ( .C (clk), .D (signal_1537), .Q (signal_2047) ) ;
    buf_clk cell_1122 ( .C (clk), .D (signal_875), .Q (signal_2049) ) ;
    buf_clk cell_1124 ( .C (clk), .D (signal_1063), .Q (signal_2051) ) ;
    buf_clk cell_1126 ( .C (clk), .D (signal_874), .Q (signal_2053) ) ;
    buf_clk cell_1128 ( .C (clk), .D (signal_1540), .Q (signal_2055) ) ;
    buf_clk cell_1130 ( .C (clk), .D (signal_873), .Q (signal_2057) ) ;
    buf_clk cell_1132 ( .C (clk), .D (signal_1543), .Q (signal_2059) ) ;
    buf_clk cell_1134 ( .C (clk), .D (signal_872), .Q (signal_2061) ) ;
    buf_clk cell_1136 ( .C (clk), .D (signal_1066), .Q (signal_2063) ) ;
    buf_clk cell_1138 ( .C (clk), .D (signal_871), .Q (signal_2065) ) ;
    buf_clk cell_1140 ( .C (clk), .D (signal_1546), .Q (signal_2067) ) ;
    buf_clk cell_1142 ( .C (clk), .D (signal_333), .Q (signal_2069) ) ;
    buf_clk cell_1144 ( .C (clk), .D (signal_1579), .Q (signal_2071) ) ;
    buf_clk cell_1146 ( .C (clk), .D (signal_335), .Q (signal_2073) ) ;
    buf_clk cell_1148 ( .C (clk), .D (signal_1580), .Q (signal_2075) ) ;
    buf_clk cell_1150 ( .C (clk), .D (signal_337), .Q (signal_2077) ) ;
    buf_clk cell_1152 ( .C (clk), .D (signal_1581), .Q (signal_2079) ) ;
    buf_clk cell_1154 ( .C (clk), .D (signal_339), .Q (signal_2081) ) ;
    buf_clk cell_1156 ( .C (clk), .D (signal_1582), .Q (signal_2083) ) ;
    buf_clk cell_1158 ( .C (clk), .D (signal_341), .Q (signal_2085) ) ;
    buf_clk cell_1160 ( .C (clk), .D (signal_1583), .Q (signal_2087) ) ;
    buf_clk cell_1162 ( .C (clk), .D (signal_343), .Q (signal_2089) ) ;
    buf_clk cell_1164 ( .C (clk), .D (signal_1584), .Q (signal_2091) ) ;
    buf_clk cell_1166 ( .C (clk), .D (signal_345), .Q (signal_2093) ) ;
    buf_clk cell_1168 ( .C (clk), .D (signal_1585), .Q (signal_2095) ) ;
    buf_clk cell_1170 ( .C (clk), .D (signal_347), .Q (signal_2097) ) ;
    buf_clk cell_1172 ( .C (clk), .D (signal_1586), .Q (signal_2099) ) ;
    buf_clk cell_1174 ( .C (clk), .D (signal_934), .Q (signal_2101) ) ;
    buf_clk cell_1176 ( .C (clk), .D (signal_1021), .Q (signal_2103) ) ;
    buf_clk cell_1178 ( .C (clk), .D (signal_933), .Q (signal_2105) ) ;
    buf_clk cell_1180 ( .C (clk), .D (signal_1405), .Q (signal_2107) ) ;
    buf_clk cell_1182 ( .C (clk), .D (signal_932), .Q (signal_2109) ) ;
    buf_clk cell_1184 ( .C (clk), .D (signal_1024), .Q (signal_2111) ) ;
    buf_clk cell_1186 ( .C (clk), .D (signal_931), .Q (signal_2113) ) ;
    buf_clk cell_1188 ( .C (clk), .D (signal_1408), .Q (signal_2115) ) ;
    buf_clk cell_1190 ( .C (clk), .D (signal_930), .Q (signal_2117) ) ;
    buf_clk cell_1192 ( .C (clk), .D (signal_1411), .Q (signal_2119) ) ;
    buf_clk cell_1194 ( .C (clk), .D (signal_929), .Q (signal_2121) ) ;
    buf_clk cell_1196 ( .C (clk), .D (signal_1414), .Q (signal_2123) ) ;
    buf_clk cell_1198 ( .C (clk), .D (signal_928), .Q (signal_2125) ) ;
    buf_clk cell_1200 ( .C (clk), .D (signal_1417), .Q (signal_2127) ) ;
    buf_clk cell_1202 ( .C (clk), .D (signal_927), .Q (signal_2129) ) ;
    buf_clk cell_1204 ( .C (clk), .D (signal_1420), .Q (signal_2131) ) ;
    buf_clk cell_1206 ( .C (clk), .D (signal_926), .Q (signal_2133) ) ;
    buf_clk cell_1208 ( .C (clk), .D (signal_1423), .Q (signal_2135) ) ;
    buf_clk cell_1210 ( .C (clk), .D (signal_925), .Q (signal_2137) ) ;
    buf_clk cell_1212 ( .C (clk), .D (signal_1426), .Q (signal_2139) ) ;
    buf_clk cell_1214 ( .C (clk), .D (signal_924), .Q (signal_2141) ) ;
    buf_clk cell_1216 ( .C (clk), .D (signal_1429), .Q (signal_2143) ) ;
    buf_clk cell_1218 ( .C (clk), .D (signal_923), .Q (signal_2145) ) ;
    buf_clk cell_1220 ( .C (clk), .D (signal_1432), .Q (signal_2147) ) ;
    buf_clk cell_1222 ( .C (clk), .D (signal_922), .Q (signal_2149) ) ;
    buf_clk cell_1224 ( .C (clk), .D (signal_1435), .Q (signal_2151) ) ;
    buf_clk cell_1226 ( .C (clk), .D (signal_921), .Q (signal_2153) ) ;
    buf_clk cell_1228 ( .C (clk), .D (signal_1438), .Q (signal_2155) ) ;
    buf_clk cell_1230 ( .C (clk), .D (signal_920), .Q (signal_2157) ) ;
    buf_clk cell_1232 ( .C (clk), .D (signal_1441), .Q (signal_2159) ) ;
    buf_clk cell_1234 ( .C (clk), .D (signal_919), .Q (signal_2161) ) ;
    buf_clk cell_1236 ( .C (clk), .D (signal_1444), .Q (signal_2163) ) ;
    buf_clk cell_1238 ( .C (clk), .D (signal_918), .Q (signal_2165) ) ;
    buf_clk cell_1240 ( .C (clk), .D (signal_1447), .Q (signal_2167) ) ;
    buf_clk cell_1242 ( .C (clk), .D (signal_917), .Q (signal_2169) ) ;
    buf_clk cell_1244 ( .C (clk), .D (signal_1450), .Q (signal_2171) ) ;
    buf_clk cell_1246 ( .C (clk), .D (signal_916), .Q (signal_2173) ) ;
    buf_clk cell_1248 ( .C (clk), .D (signal_1453), .Q (signal_2175) ) ;
    buf_clk cell_1250 ( .C (clk), .D (signal_915), .Q (signal_2177) ) ;
    buf_clk cell_1252 ( .C (clk), .D (signal_1456), .Q (signal_2179) ) ;
    buf_clk cell_1254 ( .C (clk), .D (signal_914), .Q (signal_2181) ) ;
    buf_clk cell_1256 ( .C (clk), .D (signal_1459), .Q (signal_2183) ) ;
    buf_clk cell_1258 ( .C (clk), .D (signal_913), .Q (signal_2185) ) ;
    buf_clk cell_1260 ( .C (clk), .D (signal_1462), .Q (signal_2187) ) ;
    buf_clk cell_1262 ( .C (clk), .D (signal_912), .Q (signal_2189) ) ;
    buf_clk cell_1264 ( .C (clk), .D (signal_1027), .Q (signal_2191) ) ;
    buf_clk cell_1266 ( .C (clk), .D (signal_911), .Q (signal_2193) ) ;
    buf_clk cell_1268 ( .C (clk), .D (signal_1030), .Q (signal_2195) ) ;
    buf_clk cell_1270 ( .C (clk), .D (signal_910), .Q (signal_2197) ) ;
    buf_clk cell_1272 ( .C (clk), .D (signal_1033), .Q (signal_2199) ) ;
    buf_clk cell_1274 ( .C (clk), .D (signal_909), .Q (signal_2201) ) ;
    buf_clk cell_1276 ( .C (clk), .D (signal_1036), .Q (signal_2203) ) ;
    buf_clk cell_1278 ( .C (clk), .D (signal_908), .Q (signal_2205) ) ;
    buf_clk cell_1280 ( .C (clk), .D (signal_1039), .Q (signal_2207) ) ;
    buf_clk cell_1282 ( .C (clk), .D (signal_907), .Q (signal_2209) ) ;
    buf_clk cell_1284 ( .C (clk), .D (signal_1042), .Q (signal_2211) ) ;
    buf_clk cell_1286 ( .C (clk), .D (signal_906), .Q (signal_2213) ) ;
    buf_clk cell_1288 ( .C (clk), .D (signal_1465), .Q (signal_2215) ) ;
    buf_clk cell_1290 ( .C (clk), .D (signal_905), .Q (signal_2217) ) ;
    buf_clk cell_1292 ( .C (clk), .D (signal_1468), .Q (signal_2219) ) ;
    buf_clk cell_1294 ( .C (clk), .D (signal_904), .Q (signal_2221) ) ;
    buf_clk cell_1296 ( .C (clk), .D (signal_1471), .Q (signal_2223) ) ;
    buf_clk cell_1298 ( .C (clk), .D (signal_903), .Q (signal_2225) ) ;
    buf_clk cell_1300 ( .C (clk), .D (signal_1474), .Q (signal_2227) ) ;
    buf_clk cell_1302 ( .C (clk), .D (signal_902), .Q (signal_2229) ) ;
    buf_clk cell_1304 ( .C (clk), .D (signal_1477), .Q (signal_2231) ) ;
    buf_clk cell_1306 ( .C (clk), .D (signal_901), .Q (signal_2233) ) ;
    buf_clk cell_1308 ( .C (clk), .D (signal_1045), .Q (signal_2235) ) ;
    buf_clk cell_1310 ( .C (clk), .D (signal_900), .Q (signal_2237) ) ;
    buf_clk cell_1312 ( .C (clk), .D (signal_1480), .Q (signal_2239) ) ;
    buf_clk cell_1314 ( .C (clk), .D (signal_899), .Q (signal_2241) ) ;
    buf_clk cell_1316 ( .C (clk), .D (signal_1483), .Q (signal_2243) ) ;
    buf_clk cell_1318 ( .C (clk), .D (signal_898), .Q (signal_2245) ) ;
    buf_clk cell_1320 ( .C (clk), .D (signal_1048), .Q (signal_2247) ) ;
    buf_clk cell_1322 ( .C (clk), .D (signal_897), .Q (signal_2249) ) ;
    buf_clk cell_1324 ( .C (clk), .D (signal_1486), .Q (signal_2251) ) ;
    buf_clk cell_1326 ( .C (clk), .D (signal_896), .Q (signal_2253) ) ;
    buf_clk cell_1328 ( .C (clk), .D (signal_1489), .Q (signal_2255) ) ;
    buf_clk cell_1330 ( .C (clk), .D (signal_895), .Q (signal_2257) ) ;
    buf_clk cell_1332 ( .C (clk), .D (signal_1051), .Q (signal_2259) ) ;
    buf_clk cell_1334 ( .C (clk), .D (signal_1008), .Q (signal_2261) ) ;
    buf_clk cell_1336 ( .C (clk), .D (signal_1009), .Q (signal_2263) ) ;
    buf_clk cell_1338 ( .C (clk), .D (signal_1010), .Q (signal_2265) ) ;
    buf_clk cell_1340 ( .C (clk), .D (signal_1011), .Q (signal_2267) ) ;
    buf_clk cell_1342 ( .C (clk), .D (signal_1012), .Q (signal_2269) ) ;
    buf_clk cell_1344 ( .C (clk), .D (signal_1013), .Q (signal_2271) ) ;
    buf_clk cell_1346 ( .C (clk), .D (signal_1014), .Q (signal_2273) ) ;
    buf_clk cell_1348 ( .C (clk), .D (signal_1017), .Q (signal_2275) ) ;
    buf_clk cell_1350 ( .C (clk), .D (signal_1018), .Q (signal_2277) ) ;
    buf_clk cell_1352 ( .C (clk), .D (signal_267), .Q (signal_2279) ) ;

    /* cells in depth 2 */
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_0 ( .s (signal_1748), .b ({signal_1194, signal_774}), .a ({signal_1752, signal_1750}), .c ({signal_1196, signal_870}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1 ( .s (signal_1748), .b ({signal_1193, signal_773}), .a ({signal_1756, signal_1754}), .c ({signal_1198, signal_869}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_2 ( .s (signal_1748), .b ({signal_1192, signal_772}), .a ({signal_1760, signal_1758}), .c ({signal_1200, signal_868}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3 ( .s (signal_1748), .b ({signal_1191, signal_771}), .a ({signal_1764, signal_1762}), .c ({signal_1202, signal_867}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_4 ( .s (signal_1748), .b ({signal_1190, signal_770}), .a ({signal_1768, signal_1766}), .c ({signal_1204, signal_866}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_5 ( .s (signal_1748), .b ({signal_1189, signal_769}), .a ({signal_1772, signal_1770}), .c ({signal_1206, signal_865}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_6 ( .s (signal_1748), .b ({signal_1188, signal_768}), .a ({signal_1776, signal_1774}), .c ({signal_1208, signal_864}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_7 ( .s (signal_1748), .b ({signal_1187, signal_767}), .a ({signal_1780, signal_1778}), .c ({signal_1210, signal_863}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_8 ( .s (signal_1748), .b ({signal_1186, signal_766}), .a ({signal_1784, signal_1782}), .c ({signal_1212, signal_862}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_9 ( .s (signal_1748), .b ({signal_1185, signal_765}), .a ({signal_1788, signal_1786}), .c ({signal_1214, signal_861}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_10 ( .s (signal_1748), .b ({signal_1184, signal_764}), .a ({signal_1792, signal_1790}), .c ({signal_1216, signal_860}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_11 ( .s (signal_1748), .b ({signal_1183, signal_763}), .a ({signal_1796, signal_1794}), .c ({signal_1218, signal_859}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_12 ( .s (signal_1748), .b ({signal_1182, signal_762}), .a ({signal_1800, signal_1798}), .c ({signal_1220, signal_858}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_13 ( .s (signal_1748), .b ({signal_1181, signal_761}), .a ({signal_1804, signal_1802}), .c ({signal_1222, signal_857}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_14 ( .s (signal_1748), .b ({signal_1180, signal_760}), .a ({signal_1808, signal_1806}), .c ({signal_1224, signal_856}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_15 ( .s (signal_1748), .b ({signal_1179, signal_759}), .a ({signal_1812, signal_1810}), .c ({signal_1226, signal_855}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_16 ( .s (signal_1748), .b ({signal_1178, signal_758}), .a ({signal_1816, signal_1814}), .c ({signal_1228, signal_854}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_17 ( .s (signal_1748), .b ({signal_1177, signal_757}), .a ({signal_1820, signal_1818}), .c ({signal_1230, signal_853}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_18 ( .s (signal_1748), .b ({signal_1176, signal_756}), .a ({signal_1824, signal_1822}), .c ({signal_1232, signal_852}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_19 ( .s (signal_1748), .b ({signal_1175, signal_755}), .a ({signal_1828, signal_1826}), .c ({signal_1234, signal_851}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_20 ( .s (signal_1748), .b ({signal_1174, signal_754}), .a ({signal_1832, signal_1830}), .c ({signal_1236, signal_850}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_21 ( .s (signal_1748), .b ({signal_1173, signal_753}), .a ({signal_1836, signal_1834}), .c ({signal_1238, signal_849}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_22 ( .s (signal_1748), .b ({signal_1172, signal_752}), .a ({signal_1840, signal_1838}), .c ({signal_1240, signal_848}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_23 ( .s (signal_1748), .b ({signal_1171, signal_751}), .a ({signal_1844, signal_1842}), .c ({signal_1242, signal_847}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_24 ( .s (signal_1748), .b ({signal_1170, signal_750}), .a ({signal_1848, signal_1846}), .c ({signal_1244, signal_846}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_25 ( .s (signal_1748), .b ({signal_1169, signal_749}), .a ({signal_1852, signal_1850}), .c ({signal_1246, signal_845}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_26 ( .s (signal_1748), .b ({signal_1168, signal_748}), .a ({signal_1856, signal_1854}), .c ({signal_1248, signal_844}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_27 ( .s (signal_1748), .b ({signal_1167, signal_747}), .a ({signal_1860, signal_1858}), .c ({signal_1250, signal_843}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_28 ( .s (signal_1748), .b ({signal_1166, signal_746}), .a ({signal_1864, signal_1862}), .c ({signal_1252, signal_842}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_29 ( .s (signal_1748), .b ({signal_1165, signal_745}), .a ({signal_1868, signal_1866}), .c ({signal_1254, signal_841}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_30 ( .s (signal_1748), .b ({signal_1164, signal_744}), .a ({signal_1872, signal_1870}), .c ({signal_1256, signal_840}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_31 ( .s (signal_1748), .b ({signal_1163, signal_743}), .a ({signal_1876, signal_1874}), .c ({signal_1258, signal_839}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_32 ( .s (signal_1748), .b ({signal_1162, signal_742}), .a ({signal_1880, signal_1878}), .c ({signal_1260, signal_806}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_33 ( .s (signal_1748), .b ({signal_1161, signal_741}), .a ({signal_1884, signal_1882}), .c ({signal_1262, signal_805}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_34 ( .s (signal_1748), .b ({signal_1160, signal_740}), .a ({signal_1888, signal_1886}), .c ({signal_1264, signal_804}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_35 ( .s (signal_1748), .b ({signal_1159, signal_739}), .a ({signal_1892, signal_1890}), .c ({signal_1266, signal_803}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_36 ( .s (signal_1748), .b ({signal_1158, signal_738}), .a ({signal_1896, signal_1894}), .c ({signal_1268, signal_802}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_37 ( .s (signal_1748), .b ({signal_1157, signal_737}), .a ({signal_1900, signal_1898}), .c ({signal_1270, signal_801}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_38 ( .s (signal_1748), .b ({signal_1156, signal_736}), .a ({signal_1904, signal_1902}), .c ({signal_1272, signal_800}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_39 ( .s (signal_1748), .b ({signal_1155, signal_735}), .a ({signal_1908, signal_1906}), .c ({signal_1274, signal_799}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_40 ( .s (signal_1748), .b ({signal_1154, signal_734}), .a ({signal_1912, signal_1910}), .c ({signal_1276, signal_798}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_41 ( .s (signal_1748), .b ({signal_1153, signal_733}), .a ({signal_1916, signal_1914}), .c ({signal_1278, signal_797}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_42 ( .s (signal_1748), .b ({signal_1152, signal_732}), .a ({signal_1920, signal_1918}), .c ({signal_1280, signal_796}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_43 ( .s (signal_1748), .b ({signal_1151, signal_731}), .a ({signal_1924, signal_1922}), .c ({signal_1282, signal_795}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_44 ( .s (signal_1748), .b ({signal_1150, signal_730}), .a ({signal_1928, signal_1926}), .c ({signal_1284, signal_794}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_45 ( .s (signal_1748), .b ({signal_1149, signal_729}), .a ({signal_1932, signal_1930}), .c ({signal_1286, signal_793}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_46 ( .s (signal_1748), .b ({signal_1148, signal_728}), .a ({signal_1936, signal_1934}), .c ({signal_1288, signal_792}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_47 ( .s (signal_1748), .b ({signal_1147, signal_727}), .a ({signal_1940, signal_1938}), .c ({signal_1290, signal_791}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_48 ( .s (signal_1748), .b ({signal_1146, signal_726}), .a ({signal_1944, signal_1942}), .c ({signal_1292, signal_790}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_49 ( .s (signal_1748), .b ({signal_1145, signal_725}), .a ({signal_1948, signal_1946}), .c ({signal_1294, signal_789}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_50 ( .s (signal_1748), .b ({signal_1144, signal_724}), .a ({signal_1952, signal_1950}), .c ({signal_1296, signal_788}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_51 ( .s (signal_1748), .b ({signal_1143, signal_723}), .a ({signal_1956, signal_1954}), .c ({signal_1298, signal_787}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_52 ( .s (signal_1748), .b ({signal_1142, signal_722}), .a ({signal_1960, signal_1958}), .c ({signal_1300, signal_786}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_53 ( .s (signal_1748), .b ({signal_1141, signal_721}), .a ({signal_1964, signal_1962}), .c ({signal_1302, signal_785}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_54 ( .s (signal_1748), .b ({signal_1140, signal_720}), .a ({signal_1968, signal_1966}), .c ({signal_1304, signal_784}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_55 ( .s (signal_1748), .b ({signal_1139, signal_719}), .a ({signal_1972, signal_1970}), .c ({signal_1306, signal_783}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_56 ( .s (signal_1748), .b ({signal_1138, signal_718}), .a ({signal_1976, signal_1974}), .c ({signal_1308, signal_782}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_57 ( .s (signal_1748), .b ({signal_1137, signal_717}), .a ({signal_1980, signal_1978}), .c ({signal_1310, signal_781}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_58 ( .s (signal_1748), .b ({signal_1136, signal_716}), .a ({signal_1984, signal_1982}), .c ({signal_1312, signal_780}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_59 ( .s (signal_1748), .b ({signal_1135, signal_715}), .a ({signal_1988, signal_1986}), .c ({signal_1314, signal_779}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_60 ( .s (signal_1748), .b ({signal_1134, signal_714}), .a ({signal_1992, signal_1990}), .c ({signal_1316, signal_778}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_61 ( .s (signal_1748), .b ({signal_1133, signal_713}), .a ({signal_1996, signal_1994}), .c ({signal_1318, signal_777}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_62 ( .s (signal_1748), .b ({signal_1132, signal_712}), .a ({signal_2000, signal_1998}), .c ({signal_1320, signal_776}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_63 ( .s (signal_1748), .b ({signal_1131, signal_711}), .a ({signal_2004, signal_2002}), .c ({signal_1322, signal_775}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_64 ( .a ({signal_1324, signal_268}), .b ({signal_1323, signal_269}), .c ({signal_1547, signal_822}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_65 ( .a ({signal_1228, signal_854}), .b ({signal_1196, signal_870}), .c ({signal_1323, signal_269}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_66 ( .a ({1'b0, 1'b0}), .b ({signal_1292, signal_790}), .c ({signal_1324, signal_268}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_67 ( .a ({signal_1325, signal_270}), .b ({signal_1196, signal_870}), .c ({signal_1548, signal_838}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_68 ( .a ({1'b0, 1'b0}), .b ({signal_1260, signal_806}), .c ({signal_1325, signal_270}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_69 ( .a ({signal_1327, signal_271}), .b ({signal_1326, signal_272}), .c ({signal_1549, signal_821}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_70 ( .a ({signal_1230, signal_853}), .b ({signal_1198, signal_869}), .c ({signal_1326, signal_272}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_71 ( .a ({1'b0, 1'b0}), .b ({signal_1294, signal_789}), .c ({signal_1327, signal_271}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_72 ( .a ({signal_1328, signal_273}), .b ({signal_1198, signal_869}), .c ({signal_1550, signal_837}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_73 ( .a ({1'b0, 1'b0}), .b ({signal_1262, signal_805}), .c ({signal_1328, signal_273}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_74 ( .a ({signal_1330, signal_274}), .b ({signal_1329, signal_275}), .c ({signal_1551, signal_820}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_75 ( .a ({signal_1232, signal_852}), .b ({signal_1200, signal_868}), .c ({signal_1329, signal_275}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_76 ( .a ({1'b0, 1'b0}), .b ({signal_1296, signal_788}), .c ({signal_1330, signal_274}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_77 ( .a ({signal_1331, signal_276}), .b ({signal_1200, signal_868}), .c ({signal_1552, signal_836}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_78 ( .a ({1'b0, 1'b0}), .b ({signal_1264, signal_804}), .c ({signal_1331, signal_276}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_79 ( .a ({signal_1333, signal_277}), .b ({signal_1332, signal_278}), .c ({signal_1553, signal_819}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_80 ( .a ({signal_1234, signal_851}), .b ({signal_1202, signal_867}), .c ({signal_1332, signal_278}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_81 ( .a ({1'b0, 1'b0}), .b ({signal_1298, signal_787}), .c ({signal_1333, signal_277}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_82 ( .a ({signal_1334, signal_279}), .b ({signal_1202, signal_867}), .c ({signal_1554, signal_835}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_83 ( .a ({1'b0, 1'b0}), .b ({signal_1266, signal_803}), .c ({signal_1334, signal_279}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_84 ( .a ({signal_1336, signal_280}), .b ({signal_1335, signal_281}), .c ({signal_1555, signal_818}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_85 ( .a ({signal_1236, signal_850}), .b ({signal_1204, signal_866}), .c ({signal_1335, signal_281}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_86 ( .a ({1'b0, 1'b0}), .b ({signal_1300, signal_786}), .c ({signal_1336, signal_280}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_87 ( .a ({signal_1337, signal_282}), .b ({signal_1204, signal_866}), .c ({signal_1556, signal_834}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_88 ( .a ({1'b0, 1'b0}), .b ({signal_1268, signal_802}), .c ({signal_1337, signal_282}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_89 ( .a ({signal_1339, signal_283}), .b ({signal_1338, signal_284}), .c ({signal_1557, signal_817}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_90 ( .a ({signal_1238, signal_849}), .b ({signal_1206, signal_865}), .c ({signal_1338, signal_284}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_91 ( .a ({1'b0, 1'b0}), .b ({signal_1302, signal_785}), .c ({signal_1339, signal_283}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_92 ( .a ({signal_1340, signal_285}), .b ({signal_1206, signal_865}), .c ({signal_1558, signal_833}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_93 ( .a ({1'b0, 1'b0}), .b ({signal_1270, signal_801}), .c ({signal_1340, signal_285}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_94 ( .a ({signal_1342, signal_286}), .b ({signal_1341, signal_287}), .c ({signal_1559, signal_816}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_95 ( .a ({signal_1240, signal_848}), .b ({signal_1208, signal_864}), .c ({signal_1341, signal_287}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_96 ( .a ({1'b0, 1'b0}), .b ({signal_1304, signal_784}), .c ({signal_1342, signal_286}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_97 ( .a ({signal_1343, signal_288}), .b ({signal_1208, signal_864}), .c ({signal_1560, signal_832}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_98 ( .a ({1'b0, 1'b0}), .b ({signal_1272, signal_800}), .c ({signal_1343, signal_288}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_99 ( .a ({signal_1345, signal_289}), .b ({signal_1344, signal_290}), .c ({signal_1561, signal_815}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_100 ( .a ({signal_1242, signal_847}), .b ({signal_1210, signal_863}), .c ({signal_1344, signal_290}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_101 ( .a ({1'b0, 1'b0}), .b ({signal_1306, signal_783}), .c ({signal_1345, signal_289}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_102 ( .a ({signal_1346, signal_291}), .b ({signal_1210, signal_863}), .c ({signal_1562, signal_831}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_103 ( .a ({1'b0, 1'b0}), .b ({signal_1274, signal_799}), .c ({signal_1346, signal_291}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_104 ( .a ({signal_1348, signal_292}), .b ({signal_1347, signal_293}), .c ({signal_1563, signal_814}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_105 ( .a ({signal_1244, signal_846}), .b ({signal_1212, signal_862}), .c ({signal_1347, signal_293}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_106 ( .a ({1'b0, 1'b0}), .b ({signal_1308, signal_782}), .c ({signal_1348, signal_292}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_107 ( .a ({signal_1349, signal_294}), .b ({signal_1212, signal_862}), .c ({signal_1564, signal_830}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_108 ( .a ({1'b0, 1'b0}), .b ({signal_1276, signal_798}), .c ({signal_1349, signal_294}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_109 ( .a ({signal_1351, signal_295}), .b ({signal_1350, signal_296}), .c ({signal_1565, signal_813}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_110 ( .a ({signal_1246, signal_845}), .b ({signal_1214, signal_861}), .c ({signal_1350, signal_296}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_111 ( .a ({1'b0, 1'b0}), .b ({signal_1310, signal_781}), .c ({signal_1351, signal_295}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_112 ( .a ({signal_1352, signal_297}), .b ({signal_1214, signal_861}), .c ({signal_1566, signal_829}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_113 ( .a ({1'b0, 1'b0}), .b ({signal_1278, signal_797}), .c ({signal_1352, signal_297}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_114 ( .a ({signal_1354, signal_298}), .b ({signal_1353, signal_299}), .c ({signal_1567, signal_812}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_115 ( .a ({signal_1248, signal_844}), .b ({signal_1216, signal_860}), .c ({signal_1353, signal_299}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_116 ( .a ({1'b0, 1'b0}), .b ({signal_1312, signal_780}), .c ({signal_1354, signal_298}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_117 ( .a ({signal_1355, signal_300}), .b ({signal_1216, signal_860}), .c ({signal_1568, signal_828}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_118 ( .a ({1'b0, 1'b0}), .b ({signal_1280, signal_796}), .c ({signal_1355, signal_300}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_119 ( .a ({signal_1357, signal_301}), .b ({signal_1356, signal_302}), .c ({signal_1569, signal_811}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_120 ( .a ({signal_1250, signal_843}), .b ({signal_1218, signal_859}), .c ({signal_1356, signal_302}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_121 ( .a ({1'b0, 1'b0}), .b ({signal_1314, signal_779}), .c ({signal_1357, signal_301}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_122 ( .a ({signal_1358, signal_303}), .b ({signal_1218, signal_859}), .c ({signal_1570, signal_827}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_123 ( .a ({1'b0, 1'b0}), .b ({signal_1282, signal_795}), .c ({signal_1358, signal_303}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_124 ( .a ({signal_1360, signal_304}), .b ({signal_1359, signal_305}), .c ({signal_1571, signal_810}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_125 ( .a ({signal_1252, signal_842}), .b ({signal_1220, signal_858}), .c ({signal_1359, signal_305}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_126 ( .a ({1'b0, 1'b0}), .b ({signal_1316, signal_778}), .c ({signal_1360, signal_304}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_127 ( .a ({signal_1361, signal_306}), .b ({signal_1220, signal_858}), .c ({signal_1572, signal_826}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_128 ( .a ({1'b0, 1'b0}), .b ({signal_1284, signal_794}), .c ({signal_1361, signal_306}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_129 ( .a ({signal_1363, signal_307}), .b ({signal_1362, signal_308}), .c ({signal_1573, signal_809}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_130 ( .a ({signal_1254, signal_841}), .b ({signal_1222, signal_857}), .c ({signal_1362, signal_308}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_131 ( .a ({1'b0, 1'b0}), .b ({signal_1318, signal_777}), .c ({signal_1363, signal_307}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_132 ( .a ({signal_1364, signal_309}), .b ({signal_1222, signal_857}), .c ({signal_1574, signal_825}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_133 ( .a ({1'b0, 1'b0}), .b ({signal_1286, signal_793}), .c ({signal_1364, signal_309}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_134 ( .a ({signal_1366, signal_310}), .b ({signal_1365, signal_311}), .c ({signal_1575, signal_808}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_135 ( .a ({signal_1256, signal_840}), .b ({signal_1224, signal_856}), .c ({signal_1365, signal_311}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_136 ( .a ({1'b0, 1'b0}), .b ({signal_1320, signal_776}), .c ({signal_1366, signal_310}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_137 ( .a ({signal_1367, signal_312}), .b ({signal_1224, signal_856}), .c ({signal_1576, signal_824}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_138 ( .a ({1'b0, 1'b0}), .b ({signal_1288, signal_792}), .c ({signal_1367, signal_312}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_139 ( .a ({signal_1369, signal_313}), .b ({signal_1368, signal_314}), .c ({signal_1577, signal_807}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_140 ( .a ({signal_1258, signal_839}), .b ({signal_1226, signal_855}), .c ({signal_1368, signal_314}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_141 ( .a ({1'b0, 1'b0}), .b ({signal_1322, signal_775}), .c ({signal_1369, signal_313}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_142 ( .a ({signal_1370, signal_315}), .b ({signal_1226, signal_855}), .c ({signal_1578, signal_823}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_143 ( .a ({1'b0, 1'b0}), .b ({signal_1290, signal_791}), .c ({signal_1370, signal_315}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_144 ( .a ({signal_1619, signal_316}), .b ({signal_2008, signal_2006}), .c ({signal_1651, signal_950}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_145 ( .a ({1'b0, 1'b0}), .b ({signal_1547, signal_822}), .c ({signal_1619, signal_316}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_146 ( .a ({signal_1620, signal_317}), .b ({signal_2012, signal_2010}), .c ({signal_1652, signal_949}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_147 ( .a ({1'b0, 1'b0}), .b ({signal_1549, signal_821}), .c ({signal_1620, signal_317}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_148 ( .a ({signal_1621, signal_318}), .b ({signal_2016, signal_2014}), .c ({signal_1653, signal_948}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_149 ( .a ({1'b0, 1'b0}), .b ({signal_1551, signal_820}), .c ({signal_1621, signal_318}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_150 ( .a ({signal_1622, signal_319}), .b ({signal_2020, signal_2018}), .c ({signal_1654, signal_947}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_151 ( .a ({1'b0, 1'b0}), .b ({signal_1553, signal_819}), .c ({signal_1622, signal_319}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_152 ( .a ({signal_1623, signal_320}), .b ({signal_2024, signal_2022}), .c ({signal_1655, signal_946}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_153 ( .a ({1'b0, 1'b0}), .b ({signal_1555, signal_818}), .c ({signal_1623, signal_320}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_154 ( .a ({signal_1624, signal_321}), .b ({signal_2028, signal_2026}), .c ({signal_1656, signal_945}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_155 ( .a ({1'b0, 1'b0}), .b ({signal_1557, signal_817}), .c ({signal_1624, signal_321}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_156 ( .a ({signal_1625, signal_322}), .b ({signal_2032, signal_2030}), .c ({signal_1657, signal_944}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_157 ( .a ({1'b0, 1'b0}), .b ({signal_1559, signal_816}), .c ({signal_1625, signal_322}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_158 ( .a ({signal_1626, signal_323}), .b ({signal_2036, signal_2034}), .c ({signal_1658, signal_943}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_159 ( .a ({1'b0, 1'b0}), .b ({signal_1561, signal_815}), .c ({signal_1626, signal_323}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_160 ( .a ({signal_1627, signal_324}), .b ({signal_2040, signal_2038}), .c ({signal_1659, signal_942}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_161 ( .a ({1'b0, 1'b0}), .b ({signal_1563, signal_814}), .c ({signal_1627, signal_324}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_162 ( .a ({signal_1628, signal_325}), .b ({signal_2044, signal_2042}), .c ({signal_1660, signal_941}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_163 ( .a ({1'b0, 1'b0}), .b ({signal_1565, signal_813}), .c ({signal_1628, signal_325}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_164 ( .a ({signal_1629, signal_326}), .b ({signal_2048, signal_2046}), .c ({signal_1661, signal_940}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_165 ( .a ({1'b0, 1'b0}), .b ({signal_1567, signal_812}), .c ({signal_1629, signal_326}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_166 ( .a ({signal_1630, signal_327}), .b ({signal_2052, signal_2050}), .c ({signal_1662, signal_939}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_167 ( .a ({1'b0, 1'b0}), .b ({signal_1569, signal_811}), .c ({signal_1630, signal_327}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_168 ( .a ({signal_1631, signal_328}), .b ({signal_2056, signal_2054}), .c ({signal_1663, signal_938}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_169 ( .a ({1'b0, 1'b0}), .b ({signal_1571, signal_810}), .c ({signal_1631, signal_328}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_170 ( .a ({signal_1632, signal_329}), .b ({signal_2060, signal_2058}), .c ({signal_1664, signal_937}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_171 ( .a ({1'b0, 1'b0}), .b ({signal_1573, signal_809}), .c ({signal_1632, signal_329}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_172 ( .a ({signal_1633, signal_330}), .b ({signal_2064, signal_2062}), .c ({signal_1665, signal_936}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_173 ( .a ({1'b0, 1'b0}), .b ({signal_1575, signal_808}), .c ({signal_1633, signal_330}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_174 ( .a ({signal_1634, signal_331}), .b ({signal_2068, signal_2066}), .c ({signal_1666, signal_935}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_175 ( .a ({1'b0, 1'b0}), .b ({signal_1577, signal_807}), .c ({signal_1634, signal_331}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_176 ( .a ({signal_1635, signal_332}), .b ({signal_2072, signal_2070}), .c ({signal_1667, signal_958}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_178 ( .a ({1'b0, 1'b0}), .b ({signal_1564, signal_830}), .c ({signal_1635, signal_332}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_179 ( .a ({signal_1636, signal_334}), .b ({signal_2076, signal_2074}), .c ({signal_1668, signal_957}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_181 ( .a ({1'b0, 1'b0}), .b ({signal_1566, signal_829}), .c ({signal_1636, signal_334}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_182 ( .a ({signal_1637, signal_336}), .b ({signal_2080, signal_2078}), .c ({signal_1669, signal_956}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_184 ( .a ({1'b0, 1'b0}), .b ({signal_1568, signal_828}), .c ({signal_1637, signal_336}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_185 ( .a ({signal_1638, signal_338}), .b ({signal_2084, signal_2082}), .c ({signal_1670, signal_955}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_187 ( .a ({1'b0, 1'b0}), .b ({signal_1570, signal_827}), .c ({signal_1638, signal_338}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_188 ( .a ({signal_1639, signal_340}), .b ({signal_2088, signal_2086}), .c ({signal_1671, signal_954}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_190 ( .a ({1'b0, 1'b0}), .b ({signal_1572, signal_826}), .c ({signal_1639, signal_340}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_191 ( .a ({signal_1640, signal_342}), .b ({signal_2092, signal_2090}), .c ({signal_1672, signal_953}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_193 ( .a ({1'b0, 1'b0}), .b ({signal_1574, signal_825}), .c ({signal_1640, signal_342}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_194 ( .a ({signal_1641, signal_344}), .b ({signal_2096, signal_2094}), .c ({signal_1673, signal_952}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_196 ( .a ({1'b0, 1'b0}), .b ({signal_1576, signal_824}), .c ({signal_1641, signal_344}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_197 ( .a ({signal_1642, signal_346}), .b ({signal_2100, signal_2098}), .c ({signal_1674, signal_951}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_199 ( .a ({1'b0, 1'b0}), .b ({signal_1578, signal_823}), .c ({signal_1642, signal_346}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_200 ( .a ({signal_1371, signal_348}), .b ({signal_2104, signal_2102}), .c ({signal_1587, signal_998}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_201 ( .a ({1'b0, 1'b0}), .b ({signal_1196, signal_870}), .c ({signal_1371, signal_348}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_202 ( .a ({signal_1372, signal_349}), .b ({signal_2108, signal_2106}), .c ({signal_1588, signal_997}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_203 ( .a ({1'b0, 1'b0}), .b ({signal_1198, signal_869}), .c ({signal_1372, signal_349}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_204 ( .a ({signal_1373, signal_350}), .b ({signal_2112, signal_2110}), .c ({signal_1589, signal_996}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_205 ( .a ({1'b0, 1'b0}), .b ({signal_1200, signal_868}), .c ({signal_1373, signal_350}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_206 ( .a ({signal_1374, signal_351}), .b ({signal_2116, signal_2114}), .c ({signal_1590, signal_995}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_207 ( .a ({1'b0, 1'b0}), .b ({signal_1202, signal_867}), .c ({signal_1374, signal_351}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_208 ( .a ({signal_1375, signal_352}), .b ({signal_2120, signal_2118}), .c ({signal_1591, signal_994}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_209 ( .a ({1'b0, 1'b0}), .b ({signal_1204, signal_866}), .c ({signal_1375, signal_352}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_210 ( .a ({signal_1376, signal_353}), .b ({signal_2124, signal_2122}), .c ({signal_1592, signal_993}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_211 ( .a ({1'b0, 1'b0}), .b ({signal_1206, signal_865}), .c ({signal_1376, signal_353}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_212 ( .a ({signal_1377, signal_354}), .b ({signal_2128, signal_2126}), .c ({signal_1593, signal_992}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_213 ( .a ({1'b0, 1'b0}), .b ({signal_1208, signal_864}), .c ({signal_1377, signal_354}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_214 ( .a ({signal_1378, signal_355}), .b ({signal_2132, signal_2130}), .c ({signal_1594, signal_991}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_215 ( .a ({1'b0, 1'b0}), .b ({signal_1210, signal_863}), .c ({signal_1378, signal_355}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_216 ( .a ({signal_1379, signal_356}), .b ({signal_2136, signal_2134}), .c ({signal_1595, signal_990}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_217 ( .a ({1'b0, 1'b0}), .b ({signal_1212, signal_862}), .c ({signal_1379, signal_356}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_218 ( .a ({signal_1380, signal_357}), .b ({signal_2140, signal_2138}), .c ({signal_1596, signal_989}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_219 ( .a ({1'b0, 1'b0}), .b ({signal_1214, signal_861}), .c ({signal_1380, signal_357}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_220 ( .a ({signal_1381, signal_358}), .b ({signal_2144, signal_2142}), .c ({signal_1597, signal_988}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_221 ( .a ({1'b0, 1'b0}), .b ({signal_1216, signal_860}), .c ({signal_1381, signal_358}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_222 ( .a ({signal_1382, signal_359}), .b ({signal_2148, signal_2146}), .c ({signal_1598, signal_987}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_223 ( .a ({1'b0, 1'b0}), .b ({signal_1218, signal_859}), .c ({signal_1382, signal_359}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_224 ( .a ({signal_1383, signal_360}), .b ({signal_2152, signal_2150}), .c ({signal_1599, signal_986}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_225 ( .a ({1'b0, 1'b0}), .b ({signal_1220, signal_858}), .c ({signal_1383, signal_360}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_226 ( .a ({signal_1384, signal_361}), .b ({signal_2156, signal_2154}), .c ({signal_1600, signal_985}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_227 ( .a ({1'b0, 1'b0}), .b ({signal_1222, signal_857}), .c ({signal_1384, signal_361}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_228 ( .a ({signal_1385, signal_362}), .b ({signal_2160, signal_2158}), .c ({signal_1601, signal_984}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_229 ( .a ({1'b0, 1'b0}), .b ({signal_1224, signal_856}), .c ({signal_1385, signal_362}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_230 ( .a ({signal_1386, signal_363}), .b ({signal_2164, signal_2162}), .c ({signal_1602, signal_983}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_231 ( .a ({1'b0, 1'b0}), .b ({signal_1226, signal_855}), .c ({signal_1386, signal_363}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_232 ( .a ({signal_1387, signal_364}), .b ({signal_2168, signal_2166}), .c ({signal_1603, signal_982}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_233 ( .a ({1'b0, 1'b0}), .b ({signal_1228, signal_854}), .c ({signal_1387, signal_364}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_234 ( .a ({signal_1388, signal_365}), .b ({signal_2172, signal_2170}), .c ({signal_1604, signal_981}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_235 ( .a ({1'b0, 1'b0}), .b ({signal_1230, signal_853}), .c ({signal_1388, signal_365}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_236 ( .a ({signal_1389, signal_366}), .b ({signal_2176, signal_2174}), .c ({signal_1605, signal_980}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_237 ( .a ({1'b0, 1'b0}), .b ({signal_1232, signal_852}), .c ({signal_1389, signal_366}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_238 ( .a ({signal_1390, signal_367}), .b ({signal_2180, signal_2178}), .c ({signal_1606, signal_979}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_239 ( .a ({1'b0, 1'b0}), .b ({signal_1234, signal_851}), .c ({signal_1390, signal_367}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_240 ( .a ({signal_1391, signal_368}), .b ({signal_2184, signal_2182}), .c ({signal_1607, signal_978}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_241 ( .a ({1'b0, 1'b0}), .b ({signal_1236, signal_850}), .c ({signal_1391, signal_368}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_242 ( .a ({signal_1392, signal_369}), .b ({signal_2188, signal_2186}), .c ({signal_1608, signal_977}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_243 ( .a ({1'b0, 1'b0}), .b ({signal_1238, signal_849}), .c ({signal_1392, signal_369}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_244 ( .a ({signal_1393, signal_370}), .b ({signal_2192, signal_2190}), .c ({signal_1609, signal_976}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_245 ( .a ({1'b0, 1'b0}), .b ({signal_1240, signal_848}), .c ({signal_1393, signal_370}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_246 ( .a ({signal_1394, signal_371}), .b ({signal_2196, signal_2194}), .c ({signal_1610, signal_975}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_247 ( .a ({1'b0, 1'b0}), .b ({signal_1242, signal_847}), .c ({signal_1394, signal_371}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_248 ( .a ({signal_1395, signal_372}), .b ({signal_2200, signal_2198}), .c ({signal_1611, signal_974}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_249 ( .a ({1'b0, 1'b0}), .b ({signal_1244, signal_846}), .c ({signal_1395, signal_372}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_250 ( .a ({signal_1396, signal_373}), .b ({signal_2204, signal_2202}), .c ({signal_1612, signal_973}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_251 ( .a ({1'b0, 1'b0}), .b ({signal_1246, signal_845}), .c ({signal_1396, signal_373}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_252 ( .a ({signal_1397, signal_374}), .b ({signal_2208, signal_2206}), .c ({signal_1613, signal_972}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_253 ( .a ({1'b0, 1'b0}), .b ({signal_1248, signal_844}), .c ({signal_1397, signal_374}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_254 ( .a ({signal_1398, signal_375}), .b ({signal_2212, signal_2210}), .c ({signal_1614, signal_971}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_255 ( .a ({1'b0, 1'b0}), .b ({signal_1250, signal_843}), .c ({signal_1398, signal_375}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_256 ( .a ({signal_1399, signal_376}), .b ({signal_2216, signal_2214}), .c ({signal_1615, signal_970}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_257 ( .a ({1'b0, 1'b0}), .b ({signal_1252, signal_842}), .c ({signal_1399, signal_376}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_258 ( .a ({signal_1400, signal_377}), .b ({signal_2220, signal_2218}), .c ({signal_1616, signal_969}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_259 ( .a ({1'b0, 1'b0}), .b ({signal_1254, signal_841}), .c ({signal_1400, signal_377}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_260 ( .a ({signal_1401, signal_378}), .b ({signal_2224, signal_2222}), .c ({signal_1617, signal_968}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_261 ( .a ({1'b0, 1'b0}), .b ({signal_1256, signal_840}), .c ({signal_1401, signal_378}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_262 ( .a ({signal_1402, signal_379}), .b ({signal_2228, signal_2226}), .c ({signal_1618, signal_967}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_263 ( .a ({1'b0, 1'b0}), .b ({signal_1258, signal_839}), .c ({signal_1402, signal_379}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_264 ( .a ({signal_1643, signal_380}), .b ({signal_2232, signal_2230}), .c ({signal_1675, signal_966}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_265 ( .a ({1'b0, 1'b0}), .b ({signal_1548, signal_838}), .c ({signal_1643, signal_380}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_266 ( .a ({signal_1644, signal_381}), .b ({signal_2236, signal_2234}), .c ({signal_1676, signal_965}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_267 ( .a ({1'b0, 1'b0}), .b ({signal_1550, signal_837}), .c ({signal_1644, signal_381}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_268 ( .a ({signal_1645, signal_382}), .b ({signal_2240, signal_2238}), .c ({signal_1677, signal_964}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_269 ( .a ({1'b0, 1'b0}), .b ({signal_1552, signal_836}), .c ({signal_1645, signal_382}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_270 ( .a ({signal_1646, signal_383}), .b ({signal_2244, signal_2242}), .c ({signal_1678, signal_963}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_271 ( .a ({1'b0, 1'b0}), .b ({signal_1554, signal_835}), .c ({signal_1646, signal_383}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_272 ( .a ({signal_1647, signal_384}), .b ({signal_2248, signal_2246}), .c ({signal_1679, signal_962}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_273 ( .a ({1'b0, 1'b0}), .b ({signal_1556, signal_834}), .c ({signal_1647, signal_384}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_274 ( .a ({signal_1648, signal_385}), .b ({signal_2252, signal_2250}), .c ({signal_1680, signal_961}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_275 ( .a ({1'b0, 1'b0}), .b ({signal_1558, signal_833}), .c ({signal_1648, signal_385}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_276 ( .a ({signal_1649, signal_386}), .b ({signal_2256, signal_2254}), .c ({signal_1681, signal_960}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_277 ( .a ({1'b0, 1'b0}), .b ({signal_1560, signal_832}), .c ({signal_1649, signal_386}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_278 ( .a ({signal_1650, signal_387}), .b ({signal_2260, signal_2258}), .c ({signal_1682, signal_959}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_279 ( .a ({1'b0, 1'b0}), .b ({signal_1562, signal_831}), .c ({signal_1650, signal_387}) ) ;
    CRAFT_step2_ANF #(.low_latency(0), .pipeline(1)) cell_819 ( .in0 ({ciphertext_s0[0], ciphertext_s0[1], ciphertext_s0[2], ciphertext_s0[3], ciphertext_s0[4], ciphertext_s0[5], ciphertext_s0[6], ciphertext_s0[7], ciphertext_s0[8], ciphertext_s0[9], ciphertext_s0[10], ciphertext_s0[11], ciphertext_s0[12], ciphertext_s0[13], ciphertext_s0[14], ciphertext_s0[15], ciphertext_s0[16], ciphertext_s0[17], ciphertext_s0[18], ciphertext_s0[19], ciphertext_s0[20], ciphertext_s0[21], ciphertext_s0[22], ciphertext_s0[23], ciphertext_s0[24], ciphertext_s0[25], ciphertext_s0[26], ciphertext_s0[27], ciphertext_s0[28], ciphertext_s0[29], ciphertext_s0[30], ciphertext_s0[31], ciphertext_s0[32], ciphertext_s0[33], ciphertext_s0[34], ciphertext_s0[35], ciphertext_s0[36], ciphertext_s0[37], ciphertext_s0[38], ciphertext_s0[39], ciphertext_s0[40], ciphertext_s0[41], ciphertext_s0[42], ciphertext_s0[43], ciphertext_s0[44], ciphertext_s0[45], ciphertext_s0[46], ciphertext_s0[47], ciphertext_s0[48], ciphertext_s0[49], ciphertext_s0[50], ciphertext_s0[51], ciphertext_s0[52], ciphertext_s0[53], ciphertext_s0[54], ciphertext_s0[55], ciphertext_s0[56], ciphertext_s0[57], ciphertext_s0[58], ciphertext_s0[59], ciphertext_s0[60], ciphertext_s0[61], ciphertext_s0[62], ciphertext_s0[63]}), .in1 ({ciphertext_s1[0], ciphertext_s1[1], ciphertext_s1[2], ciphertext_s1[3], ciphertext_s1[4], ciphertext_s1[5], ciphertext_s1[6], ciphertext_s1[7], ciphertext_s1[8], ciphertext_s1[9], ciphertext_s1[10], ciphertext_s1[11], ciphertext_s1[12], ciphertext_s1[13], ciphertext_s1[14], ciphertext_s1[15], ciphertext_s1[16], ciphertext_s1[17], ciphertext_s1[18], ciphertext_s1[19], ciphertext_s1[20], ciphertext_s1[21], ciphertext_s1[22], ciphertext_s1[23], ciphertext_s1[24], ciphertext_s1[25], ciphertext_s1[26], ciphertext_s1[27], ciphertext_s1[28], ciphertext_s1[29], ciphertext_s1[30], ciphertext_s1[31], ciphertext_s1[32], ciphertext_s1[33], ciphertext_s1[34], ciphertext_s1[35], ciphertext_s1[36], ciphertext_s1[37], ciphertext_s1[38], ciphertext_s1[39], ciphertext_s1[40], ciphertext_s1[41], ciphertext_s1[42], ciphertext_s1[43], ciphertext_s1[44], ciphertext_s1[45], ciphertext_s1[46], ciphertext_s1[47], ciphertext_s1[48], ciphertext_s1[49], ciphertext_s1[50], ciphertext_s1[51], ciphertext_s1[52], ciphertext_s1[53], ciphertext_s1[54], ciphertext_s1[55], ciphertext_s1[56], ciphertext_s1[57], ciphertext_s1[58], ciphertext_s1[59], ciphertext_s1[60], ciphertext_s1[61], ciphertext_s1[62], ciphertext_s1[63]}), .clk (clk), .r ({Fresh[63], Fresh[62], Fresh[61], Fresh[60], Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48], Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30], Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .out0 ({signal_774, signal_773, signal_772, signal_771, signal_770, signal_769, signal_768, signal_767, signal_766, signal_765, signal_764, signal_763, signal_762, signal_761, signal_760, signal_759, signal_758, signal_757, signal_756, signal_755, signal_754, signal_753, signal_752, signal_751, signal_750, signal_749, signal_748, signal_747, signal_746, signal_745, signal_744, signal_743, signal_742, signal_741, signal_740, signal_739, signal_738, signal_737, signal_736, signal_735, signal_734, signal_733, signal_732, signal_731, signal_730, signal_729, signal_728, signal_727, signal_726, signal_725, signal_724, signal_723, signal_722, signal_721, signal_720, signal_719, signal_718, signal_717, signal_716, signal_715, signal_714, signal_713, signal_712, signal_711}), .out1 ({signal_1194, signal_1193, signal_1192, signal_1191, signal_1190, signal_1189, signal_1188, signal_1187, signal_1186, signal_1185, signal_1184, signal_1183, signal_1182, signal_1181, signal_1180, signal_1179, signal_1178, signal_1177, signal_1176, signal_1175, signal_1174, signal_1173, signal_1172, signal_1171, signal_1170, signal_1169, signal_1168, signal_1167, signal_1166, signal_1165, signal_1164, signal_1163, signal_1162, signal_1161, signal_1160, signal_1159, signal_1158, signal_1157, signal_1156, signal_1155, signal_1154, signal_1153, signal_1152, signal_1151, signal_1150, signal_1149, signal_1148, signal_1147, signal_1146, signal_1145, signal_1144, signal_1143, signal_1142, signal_1141, signal_1140, signal_1139, signal_1138, signal_1137, signal_1136, signal_1135, signal_1134, signal_1133, signal_1132, signal_1131}) ) ;
    buf_clk cell_821 ( .C (clk), .D (signal_1747), .Q (signal_1748) ) ;
    buf_clk cell_823 ( .C (clk), .D (signal_1749), .Q (signal_1750) ) ;
    buf_clk cell_825 ( .C (clk), .D (signal_1751), .Q (signal_1752) ) ;
    buf_clk cell_827 ( .C (clk), .D (signal_1753), .Q (signal_1754) ) ;
    buf_clk cell_829 ( .C (clk), .D (signal_1755), .Q (signal_1756) ) ;
    buf_clk cell_831 ( .C (clk), .D (signal_1757), .Q (signal_1758) ) ;
    buf_clk cell_833 ( .C (clk), .D (signal_1759), .Q (signal_1760) ) ;
    buf_clk cell_835 ( .C (clk), .D (signal_1761), .Q (signal_1762) ) ;
    buf_clk cell_837 ( .C (clk), .D (signal_1763), .Q (signal_1764) ) ;
    buf_clk cell_839 ( .C (clk), .D (signal_1765), .Q (signal_1766) ) ;
    buf_clk cell_841 ( .C (clk), .D (signal_1767), .Q (signal_1768) ) ;
    buf_clk cell_843 ( .C (clk), .D (signal_1769), .Q (signal_1770) ) ;
    buf_clk cell_845 ( .C (clk), .D (signal_1771), .Q (signal_1772) ) ;
    buf_clk cell_847 ( .C (clk), .D (signal_1773), .Q (signal_1774) ) ;
    buf_clk cell_849 ( .C (clk), .D (signal_1775), .Q (signal_1776) ) ;
    buf_clk cell_851 ( .C (clk), .D (signal_1777), .Q (signal_1778) ) ;
    buf_clk cell_853 ( .C (clk), .D (signal_1779), .Q (signal_1780) ) ;
    buf_clk cell_855 ( .C (clk), .D (signal_1781), .Q (signal_1782) ) ;
    buf_clk cell_857 ( .C (clk), .D (signal_1783), .Q (signal_1784) ) ;
    buf_clk cell_859 ( .C (clk), .D (signal_1785), .Q (signal_1786) ) ;
    buf_clk cell_861 ( .C (clk), .D (signal_1787), .Q (signal_1788) ) ;
    buf_clk cell_863 ( .C (clk), .D (signal_1789), .Q (signal_1790) ) ;
    buf_clk cell_865 ( .C (clk), .D (signal_1791), .Q (signal_1792) ) ;
    buf_clk cell_867 ( .C (clk), .D (signal_1793), .Q (signal_1794) ) ;
    buf_clk cell_869 ( .C (clk), .D (signal_1795), .Q (signal_1796) ) ;
    buf_clk cell_871 ( .C (clk), .D (signal_1797), .Q (signal_1798) ) ;
    buf_clk cell_873 ( .C (clk), .D (signal_1799), .Q (signal_1800) ) ;
    buf_clk cell_875 ( .C (clk), .D (signal_1801), .Q (signal_1802) ) ;
    buf_clk cell_877 ( .C (clk), .D (signal_1803), .Q (signal_1804) ) ;
    buf_clk cell_879 ( .C (clk), .D (signal_1805), .Q (signal_1806) ) ;
    buf_clk cell_881 ( .C (clk), .D (signal_1807), .Q (signal_1808) ) ;
    buf_clk cell_883 ( .C (clk), .D (signal_1809), .Q (signal_1810) ) ;
    buf_clk cell_885 ( .C (clk), .D (signal_1811), .Q (signal_1812) ) ;
    buf_clk cell_887 ( .C (clk), .D (signal_1813), .Q (signal_1814) ) ;
    buf_clk cell_889 ( .C (clk), .D (signal_1815), .Q (signal_1816) ) ;
    buf_clk cell_891 ( .C (clk), .D (signal_1817), .Q (signal_1818) ) ;
    buf_clk cell_893 ( .C (clk), .D (signal_1819), .Q (signal_1820) ) ;
    buf_clk cell_895 ( .C (clk), .D (signal_1821), .Q (signal_1822) ) ;
    buf_clk cell_897 ( .C (clk), .D (signal_1823), .Q (signal_1824) ) ;
    buf_clk cell_899 ( .C (clk), .D (signal_1825), .Q (signal_1826) ) ;
    buf_clk cell_901 ( .C (clk), .D (signal_1827), .Q (signal_1828) ) ;
    buf_clk cell_903 ( .C (clk), .D (signal_1829), .Q (signal_1830) ) ;
    buf_clk cell_905 ( .C (clk), .D (signal_1831), .Q (signal_1832) ) ;
    buf_clk cell_907 ( .C (clk), .D (signal_1833), .Q (signal_1834) ) ;
    buf_clk cell_909 ( .C (clk), .D (signal_1835), .Q (signal_1836) ) ;
    buf_clk cell_911 ( .C (clk), .D (signal_1837), .Q (signal_1838) ) ;
    buf_clk cell_913 ( .C (clk), .D (signal_1839), .Q (signal_1840) ) ;
    buf_clk cell_915 ( .C (clk), .D (signal_1841), .Q (signal_1842) ) ;
    buf_clk cell_917 ( .C (clk), .D (signal_1843), .Q (signal_1844) ) ;
    buf_clk cell_919 ( .C (clk), .D (signal_1845), .Q (signal_1846) ) ;
    buf_clk cell_921 ( .C (clk), .D (signal_1847), .Q (signal_1848) ) ;
    buf_clk cell_923 ( .C (clk), .D (signal_1849), .Q (signal_1850) ) ;
    buf_clk cell_925 ( .C (clk), .D (signal_1851), .Q (signal_1852) ) ;
    buf_clk cell_927 ( .C (clk), .D (signal_1853), .Q (signal_1854) ) ;
    buf_clk cell_929 ( .C (clk), .D (signal_1855), .Q (signal_1856) ) ;
    buf_clk cell_931 ( .C (clk), .D (signal_1857), .Q (signal_1858) ) ;
    buf_clk cell_933 ( .C (clk), .D (signal_1859), .Q (signal_1860) ) ;
    buf_clk cell_935 ( .C (clk), .D (signal_1861), .Q (signal_1862) ) ;
    buf_clk cell_937 ( .C (clk), .D (signal_1863), .Q (signal_1864) ) ;
    buf_clk cell_939 ( .C (clk), .D (signal_1865), .Q (signal_1866) ) ;
    buf_clk cell_941 ( .C (clk), .D (signal_1867), .Q (signal_1868) ) ;
    buf_clk cell_943 ( .C (clk), .D (signal_1869), .Q (signal_1870) ) ;
    buf_clk cell_945 ( .C (clk), .D (signal_1871), .Q (signal_1872) ) ;
    buf_clk cell_947 ( .C (clk), .D (signal_1873), .Q (signal_1874) ) ;
    buf_clk cell_949 ( .C (clk), .D (signal_1875), .Q (signal_1876) ) ;
    buf_clk cell_951 ( .C (clk), .D (signal_1877), .Q (signal_1878) ) ;
    buf_clk cell_953 ( .C (clk), .D (signal_1879), .Q (signal_1880) ) ;
    buf_clk cell_955 ( .C (clk), .D (signal_1881), .Q (signal_1882) ) ;
    buf_clk cell_957 ( .C (clk), .D (signal_1883), .Q (signal_1884) ) ;
    buf_clk cell_959 ( .C (clk), .D (signal_1885), .Q (signal_1886) ) ;
    buf_clk cell_961 ( .C (clk), .D (signal_1887), .Q (signal_1888) ) ;
    buf_clk cell_963 ( .C (clk), .D (signal_1889), .Q (signal_1890) ) ;
    buf_clk cell_965 ( .C (clk), .D (signal_1891), .Q (signal_1892) ) ;
    buf_clk cell_967 ( .C (clk), .D (signal_1893), .Q (signal_1894) ) ;
    buf_clk cell_969 ( .C (clk), .D (signal_1895), .Q (signal_1896) ) ;
    buf_clk cell_971 ( .C (clk), .D (signal_1897), .Q (signal_1898) ) ;
    buf_clk cell_973 ( .C (clk), .D (signal_1899), .Q (signal_1900) ) ;
    buf_clk cell_975 ( .C (clk), .D (signal_1901), .Q (signal_1902) ) ;
    buf_clk cell_977 ( .C (clk), .D (signal_1903), .Q (signal_1904) ) ;
    buf_clk cell_979 ( .C (clk), .D (signal_1905), .Q (signal_1906) ) ;
    buf_clk cell_981 ( .C (clk), .D (signal_1907), .Q (signal_1908) ) ;
    buf_clk cell_983 ( .C (clk), .D (signal_1909), .Q (signal_1910) ) ;
    buf_clk cell_985 ( .C (clk), .D (signal_1911), .Q (signal_1912) ) ;
    buf_clk cell_987 ( .C (clk), .D (signal_1913), .Q (signal_1914) ) ;
    buf_clk cell_989 ( .C (clk), .D (signal_1915), .Q (signal_1916) ) ;
    buf_clk cell_991 ( .C (clk), .D (signal_1917), .Q (signal_1918) ) ;
    buf_clk cell_993 ( .C (clk), .D (signal_1919), .Q (signal_1920) ) ;
    buf_clk cell_995 ( .C (clk), .D (signal_1921), .Q (signal_1922) ) ;
    buf_clk cell_997 ( .C (clk), .D (signal_1923), .Q (signal_1924) ) ;
    buf_clk cell_999 ( .C (clk), .D (signal_1925), .Q (signal_1926) ) ;
    buf_clk cell_1001 ( .C (clk), .D (signal_1927), .Q (signal_1928) ) ;
    buf_clk cell_1003 ( .C (clk), .D (signal_1929), .Q (signal_1930) ) ;
    buf_clk cell_1005 ( .C (clk), .D (signal_1931), .Q (signal_1932) ) ;
    buf_clk cell_1007 ( .C (clk), .D (signal_1933), .Q (signal_1934) ) ;
    buf_clk cell_1009 ( .C (clk), .D (signal_1935), .Q (signal_1936) ) ;
    buf_clk cell_1011 ( .C (clk), .D (signal_1937), .Q (signal_1938) ) ;
    buf_clk cell_1013 ( .C (clk), .D (signal_1939), .Q (signal_1940) ) ;
    buf_clk cell_1015 ( .C (clk), .D (signal_1941), .Q (signal_1942) ) ;
    buf_clk cell_1017 ( .C (clk), .D (signal_1943), .Q (signal_1944) ) ;
    buf_clk cell_1019 ( .C (clk), .D (signal_1945), .Q (signal_1946) ) ;
    buf_clk cell_1021 ( .C (clk), .D (signal_1947), .Q (signal_1948) ) ;
    buf_clk cell_1023 ( .C (clk), .D (signal_1949), .Q (signal_1950) ) ;
    buf_clk cell_1025 ( .C (clk), .D (signal_1951), .Q (signal_1952) ) ;
    buf_clk cell_1027 ( .C (clk), .D (signal_1953), .Q (signal_1954) ) ;
    buf_clk cell_1029 ( .C (clk), .D (signal_1955), .Q (signal_1956) ) ;
    buf_clk cell_1031 ( .C (clk), .D (signal_1957), .Q (signal_1958) ) ;
    buf_clk cell_1033 ( .C (clk), .D (signal_1959), .Q (signal_1960) ) ;
    buf_clk cell_1035 ( .C (clk), .D (signal_1961), .Q (signal_1962) ) ;
    buf_clk cell_1037 ( .C (clk), .D (signal_1963), .Q (signal_1964) ) ;
    buf_clk cell_1039 ( .C (clk), .D (signal_1965), .Q (signal_1966) ) ;
    buf_clk cell_1041 ( .C (clk), .D (signal_1967), .Q (signal_1968) ) ;
    buf_clk cell_1043 ( .C (clk), .D (signal_1969), .Q (signal_1970) ) ;
    buf_clk cell_1045 ( .C (clk), .D (signal_1971), .Q (signal_1972) ) ;
    buf_clk cell_1047 ( .C (clk), .D (signal_1973), .Q (signal_1974) ) ;
    buf_clk cell_1049 ( .C (clk), .D (signal_1975), .Q (signal_1976) ) ;
    buf_clk cell_1051 ( .C (clk), .D (signal_1977), .Q (signal_1978) ) ;
    buf_clk cell_1053 ( .C (clk), .D (signal_1979), .Q (signal_1980) ) ;
    buf_clk cell_1055 ( .C (clk), .D (signal_1981), .Q (signal_1982) ) ;
    buf_clk cell_1057 ( .C (clk), .D (signal_1983), .Q (signal_1984) ) ;
    buf_clk cell_1059 ( .C (clk), .D (signal_1985), .Q (signal_1986) ) ;
    buf_clk cell_1061 ( .C (clk), .D (signal_1987), .Q (signal_1988) ) ;
    buf_clk cell_1063 ( .C (clk), .D (signal_1989), .Q (signal_1990) ) ;
    buf_clk cell_1065 ( .C (clk), .D (signal_1991), .Q (signal_1992) ) ;
    buf_clk cell_1067 ( .C (clk), .D (signal_1993), .Q (signal_1994) ) ;
    buf_clk cell_1069 ( .C (clk), .D (signal_1995), .Q (signal_1996) ) ;
    buf_clk cell_1071 ( .C (clk), .D (signal_1997), .Q (signal_1998) ) ;
    buf_clk cell_1073 ( .C (clk), .D (signal_1999), .Q (signal_2000) ) ;
    buf_clk cell_1075 ( .C (clk), .D (signal_2001), .Q (signal_2002) ) ;
    buf_clk cell_1077 ( .C (clk), .D (signal_2003), .Q (signal_2004) ) ;
    buf_clk cell_1079 ( .C (clk), .D (signal_2005), .Q (signal_2006) ) ;
    buf_clk cell_1081 ( .C (clk), .D (signal_2007), .Q (signal_2008) ) ;
    buf_clk cell_1083 ( .C (clk), .D (signal_2009), .Q (signal_2010) ) ;
    buf_clk cell_1085 ( .C (clk), .D (signal_2011), .Q (signal_2012) ) ;
    buf_clk cell_1087 ( .C (clk), .D (signal_2013), .Q (signal_2014) ) ;
    buf_clk cell_1089 ( .C (clk), .D (signal_2015), .Q (signal_2016) ) ;
    buf_clk cell_1091 ( .C (clk), .D (signal_2017), .Q (signal_2018) ) ;
    buf_clk cell_1093 ( .C (clk), .D (signal_2019), .Q (signal_2020) ) ;
    buf_clk cell_1095 ( .C (clk), .D (signal_2021), .Q (signal_2022) ) ;
    buf_clk cell_1097 ( .C (clk), .D (signal_2023), .Q (signal_2024) ) ;
    buf_clk cell_1099 ( .C (clk), .D (signal_2025), .Q (signal_2026) ) ;
    buf_clk cell_1101 ( .C (clk), .D (signal_2027), .Q (signal_2028) ) ;
    buf_clk cell_1103 ( .C (clk), .D (signal_2029), .Q (signal_2030) ) ;
    buf_clk cell_1105 ( .C (clk), .D (signal_2031), .Q (signal_2032) ) ;
    buf_clk cell_1107 ( .C (clk), .D (signal_2033), .Q (signal_2034) ) ;
    buf_clk cell_1109 ( .C (clk), .D (signal_2035), .Q (signal_2036) ) ;
    buf_clk cell_1111 ( .C (clk), .D (signal_2037), .Q (signal_2038) ) ;
    buf_clk cell_1113 ( .C (clk), .D (signal_2039), .Q (signal_2040) ) ;
    buf_clk cell_1115 ( .C (clk), .D (signal_2041), .Q (signal_2042) ) ;
    buf_clk cell_1117 ( .C (clk), .D (signal_2043), .Q (signal_2044) ) ;
    buf_clk cell_1119 ( .C (clk), .D (signal_2045), .Q (signal_2046) ) ;
    buf_clk cell_1121 ( .C (clk), .D (signal_2047), .Q (signal_2048) ) ;
    buf_clk cell_1123 ( .C (clk), .D (signal_2049), .Q (signal_2050) ) ;
    buf_clk cell_1125 ( .C (clk), .D (signal_2051), .Q (signal_2052) ) ;
    buf_clk cell_1127 ( .C (clk), .D (signal_2053), .Q (signal_2054) ) ;
    buf_clk cell_1129 ( .C (clk), .D (signal_2055), .Q (signal_2056) ) ;
    buf_clk cell_1131 ( .C (clk), .D (signal_2057), .Q (signal_2058) ) ;
    buf_clk cell_1133 ( .C (clk), .D (signal_2059), .Q (signal_2060) ) ;
    buf_clk cell_1135 ( .C (clk), .D (signal_2061), .Q (signal_2062) ) ;
    buf_clk cell_1137 ( .C (clk), .D (signal_2063), .Q (signal_2064) ) ;
    buf_clk cell_1139 ( .C (clk), .D (signal_2065), .Q (signal_2066) ) ;
    buf_clk cell_1141 ( .C (clk), .D (signal_2067), .Q (signal_2068) ) ;
    buf_clk cell_1143 ( .C (clk), .D (signal_2069), .Q (signal_2070) ) ;
    buf_clk cell_1145 ( .C (clk), .D (signal_2071), .Q (signal_2072) ) ;
    buf_clk cell_1147 ( .C (clk), .D (signal_2073), .Q (signal_2074) ) ;
    buf_clk cell_1149 ( .C (clk), .D (signal_2075), .Q (signal_2076) ) ;
    buf_clk cell_1151 ( .C (clk), .D (signal_2077), .Q (signal_2078) ) ;
    buf_clk cell_1153 ( .C (clk), .D (signal_2079), .Q (signal_2080) ) ;
    buf_clk cell_1155 ( .C (clk), .D (signal_2081), .Q (signal_2082) ) ;
    buf_clk cell_1157 ( .C (clk), .D (signal_2083), .Q (signal_2084) ) ;
    buf_clk cell_1159 ( .C (clk), .D (signal_2085), .Q (signal_2086) ) ;
    buf_clk cell_1161 ( .C (clk), .D (signal_2087), .Q (signal_2088) ) ;
    buf_clk cell_1163 ( .C (clk), .D (signal_2089), .Q (signal_2090) ) ;
    buf_clk cell_1165 ( .C (clk), .D (signal_2091), .Q (signal_2092) ) ;
    buf_clk cell_1167 ( .C (clk), .D (signal_2093), .Q (signal_2094) ) ;
    buf_clk cell_1169 ( .C (clk), .D (signal_2095), .Q (signal_2096) ) ;
    buf_clk cell_1171 ( .C (clk), .D (signal_2097), .Q (signal_2098) ) ;
    buf_clk cell_1173 ( .C (clk), .D (signal_2099), .Q (signal_2100) ) ;
    buf_clk cell_1175 ( .C (clk), .D (signal_2101), .Q (signal_2102) ) ;
    buf_clk cell_1177 ( .C (clk), .D (signal_2103), .Q (signal_2104) ) ;
    buf_clk cell_1179 ( .C (clk), .D (signal_2105), .Q (signal_2106) ) ;
    buf_clk cell_1181 ( .C (clk), .D (signal_2107), .Q (signal_2108) ) ;
    buf_clk cell_1183 ( .C (clk), .D (signal_2109), .Q (signal_2110) ) ;
    buf_clk cell_1185 ( .C (clk), .D (signal_2111), .Q (signal_2112) ) ;
    buf_clk cell_1187 ( .C (clk), .D (signal_2113), .Q (signal_2114) ) ;
    buf_clk cell_1189 ( .C (clk), .D (signal_2115), .Q (signal_2116) ) ;
    buf_clk cell_1191 ( .C (clk), .D (signal_2117), .Q (signal_2118) ) ;
    buf_clk cell_1193 ( .C (clk), .D (signal_2119), .Q (signal_2120) ) ;
    buf_clk cell_1195 ( .C (clk), .D (signal_2121), .Q (signal_2122) ) ;
    buf_clk cell_1197 ( .C (clk), .D (signal_2123), .Q (signal_2124) ) ;
    buf_clk cell_1199 ( .C (clk), .D (signal_2125), .Q (signal_2126) ) ;
    buf_clk cell_1201 ( .C (clk), .D (signal_2127), .Q (signal_2128) ) ;
    buf_clk cell_1203 ( .C (clk), .D (signal_2129), .Q (signal_2130) ) ;
    buf_clk cell_1205 ( .C (clk), .D (signal_2131), .Q (signal_2132) ) ;
    buf_clk cell_1207 ( .C (clk), .D (signal_2133), .Q (signal_2134) ) ;
    buf_clk cell_1209 ( .C (clk), .D (signal_2135), .Q (signal_2136) ) ;
    buf_clk cell_1211 ( .C (clk), .D (signal_2137), .Q (signal_2138) ) ;
    buf_clk cell_1213 ( .C (clk), .D (signal_2139), .Q (signal_2140) ) ;
    buf_clk cell_1215 ( .C (clk), .D (signal_2141), .Q (signal_2142) ) ;
    buf_clk cell_1217 ( .C (clk), .D (signal_2143), .Q (signal_2144) ) ;
    buf_clk cell_1219 ( .C (clk), .D (signal_2145), .Q (signal_2146) ) ;
    buf_clk cell_1221 ( .C (clk), .D (signal_2147), .Q (signal_2148) ) ;
    buf_clk cell_1223 ( .C (clk), .D (signal_2149), .Q (signal_2150) ) ;
    buf_clk cell_1225 ( .C (clk), .D (signal_2151), .Q (signal_2152) ) ;
    buf_clk cell_1227 ( .C (clk), .D (signal_2153), .Q (signal_2154) ) ;
    buf_clk cell_1229 ( .C (clk), .D (signal_2155), .Q (signal_2156) ) ;
    buf_clk cell_1231 ( .C (clk), .D (signal_2157), .Q (signal_2158) ) ;
    buf_clk cell_1233 ( .C (clk), .D (signal_2159), .Q (signal_2160) ) ;
    buf_clk cell_1235 ( .C (clk), .D (signal_2161), .Q (signal_2162) ) ;
    buf_clk cell_1237 ( .C (clk), .D (signal_2163), .Q (signal_2164) ) ;
    buf_clk cell_1239 ( .C (clk), .D (signal_2165), .Q (signal_2166) ) ;
    buf_clk cell_1241 ( .C (clk), .D (signal_2167), .Q (signal_2168) ) ;
    buf_clk cell_1243 ( .C (clk), .D (signal_2169), .Q (signal_2170) ) ;
    buf_clk cell_1245 ( .C (clk), .D (signal_2171), .Q (signal_2172) ) ;
    buf_clk cell_1247 ( .C (clk), .D (signal_2173), .Q (signal_2174) ) ;
    buf_clk cell_1249 ( .C (clk), .D (signal_2175), .Q (signal_2176) ) ;
    buf_clk cell_1251 ( .C (clk), .D (signal_2177), .Q (signal_2178) ) ;
    buf_clk cell_1253 ( .C (clk), .D (signal_2179), .Q (signal_2180) ) ;
    buf_clk cell_1255 ( .C (clk), .D (signal_2181), .Q (signal_2182) ) ;
    buf_clk cell_1257 ( .C (clk), .D (signal_2183), .Q (signal_2184) ) ;
    buf_clk cell_1259 ( .C (clk), .D (signal_2185), .Q (signal_2186) ) ;
    buf_clk cell_1261 ( .C (clk), .D (signal_2187), .Q (signal_2188) ) ;
    buf_clk cell_1263 ( .C (clk), .D (signal_2189), .Q (signal_2190) ) ;
    buf_clk cell_1265 ( .C (clk), .D (signal_2191), .Q (signal_2192) ) ;
    buf_clk cell_1267 ( .C (clk), .D (signal_2193), .Q (signal_2194) ) ;
    buf_clk cell_1269 ( .C (clk), .D (signal_2195), .Q (signal_2196) ) ;
    buf_clk cell_1271 ( .C (clk), .D (signal_2197), .Q (signal_2198) ) ;
    buf_clk cell_1273 ( .C (clk), .D (signal_2199), .Q (signal_2200) ) ;
    buf_clk cell_1275 ( .C (clk), .D (signal_2201), .Q (signal_2202) ) ;
    buf_clk cell_1277 ( .C (clk), .D (signal_2203), .Q (signal_2204) ) ;
    buf_clk cell_1279 ( .C (clk), .D (signal_2205), .Q (signal_2206) ) ;
    buf_clk cell_1281 ( .C (clk), .D (signal_2207), .Q (signal_2208) ) ;
    buf_clk cell_1283 ( .C (clk), .D (signal_2209), .Q (signal_2210) ) ;
    buf_clk cell_1285 ( .C (clk), .D (signal_2211), .Q (signal_2212) ) ;
    buf_clk cell_1287 ( .C (clk), .D (signal_2213), .Q (signal_2214) ) ;
    buf_clk cell_1289 ( .C (clk), .D (signal_2215), .Q (signal_2216) ) ;
    buf_clk cell_1291 ( .C (clk), .D (signal_2217), .Q (signal_2218) ) ;
    buf_clk cell_1293 ( .C (clk), .D (signal_2219), .Q (signal_2220) ) ;
    buf_clk cell_1295 ( .C (clk), .D (signal_2221), .Q (signal_2222) ) ;
    buf_clk cell_1297 ( .C (clk), .D (signal_2223), .Q (signal_2224) ) ;
    buf_clk cell_1299 ( .C (clk), .D (signal_2225), .Q (signal_2226) ) ;
    buf_clk cell_1301 ( .C (clk), .D (signal_2227), .Q (signal_2228) ) ;
    buf_clk cell_1303 ( .C (clk), .D (signal_2229), .Q (signal_2230) ) ;
    buf_clk cell_1305 ( .C (clk), .D (signal_2231), .Q (signal_2232) ) ;
    buf_clk cell_1307 ( .C (clk), .D (signal_2233), .Q (signal_2234) ) ;
    buf_clk cell_1309 ( .C (clk), .D (signal_2235), .Q (signal_2236) ) ;
    buf_clk cell_1311 ( .C (clk), .D (signal_2237), .Q (signal_2238) ) ;
    buf_clk cell_1313 ( .C (clk), .D (signal_2239), .Q (signal_2240) ) ;
    buf_clk cell_1315 ( .C (clk), .D (signal_2241), .Q (signal_2242) ) ;
    buf_clk cell_1317 ( .C (clk), .D (signal_2243), .Q (signal_2244) ) ;
    buf_clk cell_1319 ( .C (clk), .D (signal_2245), .Q (signal_2246) ) ;
    buf_clk cell_1321 ( .C (clk), .D (signal_2247), .Q (signal_2248) ) ;
    buf_clk cell_1323 ( .C (clk), .D (signal_2249), .Q (signal_2250) ) ;
    buf_clk cell_1325 ( .C (clk), .D (signal_2251), .Q (signal_2252) ) ;
    buf_clk cell_1327 ( .C (clk), .D (signal_2253), .Q (signal_2254) ) ;
    buf_clk cell_1329 ( .C (clk), .D (signal_2255), .Q (signal_2256) ) ;
    buf_clk cell_1331 ( .C (clk), .D (signal_2257), .Q (signal_2258) ) ;
    buf_clk cell_1333 ( .C (clk), .D (signal_2259), .Q (signal_2260) ) ;
    buf_clk cell_1335 ( .C (clk), .D (signal_2261), .Q (signal_2262) ) ;
    buf_clk cell_1337 ( .C (clk), .D (signal_2263), .Q (signal_2264) ) ;
    buf_clk cell_1339 ( .C (clk), .D (signal_2265), .Q (signal_2266) ) ;
    buf_clk cell_1341 ( .C (clk), .D (signal_2267), .Q (signal_2268) ) ;
    buf_clk cell_1343 ( .C (clk), .D (signal_2269), .Q (signal_2270) ) ;
    buf_clk cell_1345 ( .C (clk), .D (signal_2271), .Q (signal_2272) ) ;
    buf_clk cell_1347 ( .C (clk), .D (signal_2273), .Q (signal_2274) ) ;
    buf_clk cell_1349 ( .C (clk), .D (signal_2275), .Q (signal_2276) ) ;
    buf_clk cell_1351 ( .C (clk), .D (signal_2277), .Q (signal_2278) ) ;
    buf_clk cell_1353 ( .C (clk), .D (signal_2279), .Q (signal_2280) ) ;

    /* register cells */
    reg_masked #(.low_latency(0), .pipeline(1)) cell_281 ( .clk (clk), .D ({signal_1666, signal_935}), .Q ({ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_283 ( .clk (clk), .D ({signal_1665, signal_936}), .Q ({ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_285 ( .clk (clk), .D ({signal_1664, signal_937}), .Q ({ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_287 ( .clk (clk), .D ({signal_1663, signal_938}), .Q ({ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_289 ( .clk (clk), .D ({signal_1662, signal_939}), .Q ({ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_291 ( .clk (clk), .D ({signal_1661, signal_940}), .Q ({ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_293 ( .clk (clk), .D ({signal_1660, signal_941}), .Q ({ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_295 ( .clk (clk), .D ({signal_1659, signal_942}), .Q ({ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_297 ( .clk (clk), .D ({signal_1658, signal_943}), .Q ({ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_299 ( .clk (clk), .D ({signal_1657, signal_944}), .Q ({ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_301 ( .clk (clk), .D ({signal_1656, signal_945}), .Q ({ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_303 ( .clk (clk), .D ({signal_1655, signal_946}), .Q ({ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_305 ( .clk (clk), .D ({signal_1654, signal_947}), .Q ({ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_307 ( .clk (clk), .D ({signal_1653, signal_948}), .Q ({ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_309 ( .clk (clk), .D ({signal_1652, signal_949}), .Q ({ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_311 ( .clk (clk), .D ({signal_1651, signal_950}), .Q ({ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_313 ( .clk (clk), .D ({signal_1674, signal_951}), .Q ({ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_315 ( .clk (clk), .D ({signal_1673, signal_952}), .Q ({ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_317 ( .clk (clk), .D ({signal_1672, signal_953}), .Q ({ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_319 ( .clk (clk), .D ({signal_1671, signal_954}), .Q ({ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_321 ( .clk (clk), .D ({signal_1670, signal_955}), .Q ({ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_323 ( .clk (clk), .D ({signal_1669, signal_956}), .Q ({ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_325 ( .clk (clk), .D ({signal_1668, signal_957}), .Q ({ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_327 ( .clk (clk), .D ({signal_1667, signal_958}), .Q ({ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_329 ( .clk (clk), .D ({signal_1682, signal_959}), .Q ({ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_331 ( .clk (clk), .D ({signal_1681, signal_960}), .Q ({ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_333 ( .clk (clk), .D ({signal_1680, signal_961}), .Q ({ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_335 ( .clk (clk), .D ({signal_1679, signal_962}), .Q ({ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_337 ( .clk (clk), .D ({signal_1678, signal_963}), .Q ({ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_339 ( .clk (clk), .D ({signal_1677, signal_964}), .Q ({ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_341 ( .clk (clk), .D ({signal_1676, signal_965}), .Q ({ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_343 ( .clk (clk), .D ({signal_1675, signal_966}), .Q ({ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_345 ( .clk (clk), .D ({signal_1618, signal_967}), .Q ({ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_347 ( .clk (clk), .D ({signal_1617, signal_968}), .Q ({ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_349 ( .clk (clk), .D ({signal_1616, signal_969}), .Q ({ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_351 ( .clk (clk), .D ({signal_1615, signal_970}), .Q ({ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_353 ( .clk (clk), .D ({signal_1614, signal_971}), .Q ({ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_355 ( .clk (clk), .D ({signal_1613, signal_972}), .Q ({ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_357 ( .clk (clk), .D ({signal_1612, signal_973}), .Q ({ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_359 ( .clk (clk), .D ({signal_1611, signal_974}), .Q ({ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_361 ( .clk (clk), .D ({signal_1610, signal_975}), .Q ({ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_363 ( .clk (clk), .D ({signal_1609, signal_976}), .Q ({ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_365 ( .clk (clk), .D ({signal_1608, signal_977}), .Q ({ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_367 ( .clk (clk), .D ({signal_1607, signal_978}), .Q ({ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_369 ( .clk (clk), .D ({signal_1606, signal_979}), .Q ({ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_371 ( .clk (clk), .D ({signal_1605, signal_980}), .Q ({ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_373 ( .clk (clk), .D ({signal_1604, signal_981}), .Q ({ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_375 ( .clk (clk), .D ({signal_1603, signal_982}), .Q ({ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_377 ( .clk (clk), .D ({signal_1602, signal_983}), .Q ({ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_379 ( .clk (clk), .D ({signal_1601, signal_984}), .Q ({ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_381 ( .clk (clk), .D ({signal_1600, signal_985}), .Q ({ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_383 ( .clk (clk), .D ({signal_1599, signal_986}), .Q ({ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_385 ( .clk (clk), .D ({signal_1598, signal_987}), .Q ({ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_387 ( .clk (clk), .D ({signal_1597, signal_988}), .Q ({ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_389 ( .clk (clk), .D ({signal_1596, signal_989}), .Q ({ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_391 ( .clk (clk), .D ({signal_1595, signal_990}), .Q ({ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_393 ( .clk (clk), .D ({signal_1594, signal_991}), .Q ({ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_395 ( .clk (clk), .D ({signal_1593, signal_992}), .Q ({ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_397 ( .clk (clk), .D ({signal_1592, signal_993}), .Q ({ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_399 ( .clk (clk), .D ({signal_1591, signal_994}), .Q ({ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_401 ( .clk (clk), .D ({signal_1590, signal_995}), .Q ({ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_403 ( .clk (clk), .D ({signal_1589, signal_996}), .Q ({ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_405 ( .clk (clk), .D ({signal_1588, signal_997}), .Q ({ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_407 ( .clk (clk), .D ({signal_1587, signal_998}), .Q ({ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    DFF_X1 cell_789 ( .CK (clk), .D (signal_2262), .Q (signal_1001), .QN () ) ;
    DFF_X1 cell_791 ( .CK (clk), .D (signal_2264), .Q (signal_1002), .QN () ) ;
    DFF_X1 cell_793 ( .CK (clk), .D (signal_2266), .Q (signal_1003), .QN () ) ;
    DFF_X1 cell_795 ( .CK (clk), .D (signal_2268), .Q (signal_1004), .QN () ) ;
    DFF_X1 cell_797 ( .CK (clk), .D (signal_2270), .Q (signal_1005), .QN () ) ;
    DFF_X1 cell_799 ( .CK (clk), .D (signal_2272), .Q (signal_1006), .QN () ) ;
    DFF_X1 cell_801 ( .CK (clk), .D (signal_2274), .Q (signal_1007), .QN () ) ;
    DFF_X1 cell_814 ( .CK (clk), .D (signal_2276), .Q (signal_1015), .QN () ) ;
    DFF_X1 cell_816 ( .CK (clk), .D (signal_2278), .Q (signal_1016), .QN () ) ;
    DFF_X1 cell_818 ( .CK (clk), .D (signal_2280), .Q (done), .QN () ) ;
endmodule
