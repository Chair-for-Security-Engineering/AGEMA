/* modified netlist. Source: module AES in file /mnt/c/Users/Amir/Desktop/Papers_in_progress/AGEMA/Designs/AES_serial/AGEMA/sbox_opt3/AES.v */
/* 4 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 5 register stage(s) in total */

module AES_GHPCLL_Pipeline_d1 (plaintext_s0, key_s0, clk, start, plaintext_s1, key_s1, Fresh, ciphertext_s0, done, ciphertext_s1);
    input [127:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input start ;
    input [127:0] plaintext_s1 ;
    input [127:0] key_s1 ;
    input [135:0] Fresh ;
    output [127:0] ciphertext_s0 ;
    output done ;
    output [127:0] ciphertext_s1 ;
    wire nReset ;
    wire selMC ;
    wire selSR ;
    wire selXOR ;
    wire enRCon ;
    wire finalStep ;
    wire intFinal ;
    wire intselXOR ;
    wire notFirst ;
    wire n10 ;
    wire n9 ;
    wire n12 ;
    wire n13 ;
    wire ctrl_n16 ;
    wire ctrl_n15 ;
    wire ctrl_n14 ;
    wire ctrl_n11 ;
    wire ctrl_n10 ;
    wire ctrl_n9 ;
    wire ctrl_n8 ;
    wire ctrl_n7 ;
    wire ctrl_n5 ;
    wire ctrl_n4 ;
    wire ctrl_n2 ;
    wire ctrl_n12 ;
    wire ctrl_n6 ;
    wire ctrl_N14 ;
    wire ctrl_seq4Out_1_ ;
    wire ctrl_seq4In_1_ ;
    wire ctrl_nRstSeq4 ;
    wire ctrl_n13 ;
    wire ctrl_seq6Out_4_ ;
    wire ctrl_seq6In_1_ ;
    wire ctrl_seq6In_2_ ;
    wire ctrl_seq6In_3_ ;
    wire ctrl_seq6In_4_ ;
    wire ctrl_seq6_SFF_0_QD ;
    wire ctrl_seq6_SFF_1_QD ;
    wire ctrl_seq6_SFF_2_QD ;
    wire ctrl_seq6_SFF_3_QD ;
    wire ctrl_seq6_SFF_4_QD ;
    wire ctrl_seq4_SFF_0_QD ;
    wire ctrl_seq4_SFF_1_QD ;
    wire stateArray_n33 ;
    wire stateArray_n32 ;
    wire stateArray_n31 ;
    wire stateArray_n30 ;
    wire stateArray_n29 ;
    wire stateArray_n28 ;
    wire stateArray_n27 ;
    wire stateArray_n26 ;
    wire stateArray_n25 ;
    wire stateArray_n24 ;
    wire stateArray_n23 ;
    wire stateArray_n22 ;
    wire stateArray_n21 ;
    wire stateArray_n20 ;
    wire stateArray_n19 ;
    wire stateArray_n18 ;
    wire stateArray_n17 ;
    wire stateArray_n16 ;
    wire stateArray_n15 ;
    wire stateArray_n14 ;
    wire stateArray_n13 ;
    wire stateArray_S00reg_gff_1_SFF_0_QD ;
    wire stateArray_S00reg_gff_1_SFF_1_QD ;
    wire stateArray_S00reg_gff_1_SFF_2_QD ;
    wire stateArray_S00reg_gff_1_SFF_3_QD ;
    wire stateArray_S00reg_gff_1_SFF_4_QD ;
    wire stateArray_S00reg_gff_1_SFF_5_QD ;
    wire stateArray_S00reg_gff_1_SFF_6_QD ;
    wire stateArray_S00reg_gff_1_SFF_7_QD ;
    wire stateArray_S01reg_gff_1_SFF_0_QD ;
    wire stateArray_S01reg_gff_1_SFF_1_QD ;
    wire stateArray_S01reg_gff_1_SFF_2_QD ;
    wire stateArray_S01reg_gff_1_SFF_3_QD ;
    wire stateArray_S01reg_gff_1_SFF_4_QD ;
    wire stateArray_S01reg_gff_1_SFF_5_QD ;
    wire stateArray_S01reg_gff_1_SFF_6_QD ;
    wire stateArray_S01reg_gff_1_SFF_7_QD ;
    wire stateArray_S02reg_gff_1_SFF_0_QD ;
    wire stateArray_S02reg_gff_1_SFF_1_QD ;
    wire stateArray_S02reg_gff_1_SFF_2_QD ;
    wire stateArray_S02reg_gff_1_SFF_3_QD ;
    wire stateArray_S02reg_gff_1_SFF_4_QD ;
    wire stateArray_S02reg_gff_1_SFF_5_QD ;
    wire stateArray_S02reg_gff_1_SFF_6_QD ;
    wire stateArray_S02reg_gff_1_SFF_7_QD ;
    wire stateArray_S03reg_gff_1_SFF_0_QD ;
    wire stateArray_S03reg_gff_1_SFF_1_QD ;
    wire stateArray_S03reg_gff_1_SFF_2_QD ;
    wire stateArray_S03reg_gff_1_SFF_3_QD ;
    wire stateArray_S03reg_gff_1_SFF_4_QD ;
    wire stateArray_S03reg_gff_1_SFF_5_QD ;
    wire stateArray_S03reg_gff_1_SFF_6_QD ;
    wire stateArray_S03reg_gff_1_SFF_7_QD ;
    wire stateArray_S10reg_gff_1_SFF_0_QD ;
    wire stateArray_S10reg_gff_1_SFF_1_QD ;
    wire stateArray_S10reg_gff_1_SFF_2_QD ;
    wire stateArray_S10reg_gff_1_SFF_3_QD ;
    wire stateArray_S10reg_gff_1_SFF_4_QD ;
    wire stateArray_S10reg_gff_1_SFF_5_QD ;
    wire stateArray_S10reg_gff_1_SFF_6_QD ;
    wire stateArray_S10reg_gff_1_SFF_7_QD ;
    wire stateArray_S11reg_gff_1_SFF_0_QD ;
    wire stateArray_S11reg_gff_1_SFF_1_QD ;
    wire stateArray_S11reg_gff_1_SFF_2_QD ;
    wire stateArray_S11reg_gff_1_SFF_3_QD ;
    wire stateArray_S11reg_gff_1_SFF_4_QD ;
    wire stateArray_S11reg_gff_1_SFF_5_QD ;
    wire stateArray_S11reg_gff_1_SFF_6_QD ;
    wire stateArray_S11reg_gff_1_SFF_7_QD ;
    wire stateArray_S12reg_gff_1_SFF_0_QD ;
    wire stateArray_S12reg_gff_1_SFF_1_QD ;
    wire stateArray_S12reg_gff_1_SFF_2_QD ;
    wire stateArray_S12reg_gff_1_SFF_3_QD ;
    wire stateArray_S12reg_gff_1_SFF_4_QD ;
    wire stateArray_S12reg_gff_1_SFF_5_QD ;
    wire stateArray_S12reg_gff_1_SFF_6_QD ;
    wire stateArray_S12reg_gff_1_SFF_7_QD ;
    wire stateArray_S13reg_gff_1_SFF_0_QD ;
    wire stateArray_S13reg_gff_1_SFF_1_QD ;
    wire stateArray_S13reg_gff_1_SFF_2_QD ;
    wire stateArray_S13reg_gff_1_SFF_3_QD ;
    wire stateArray_S13reg_gff_1_SFF_4_QD ;
    wire stateArray_S13reg_gff_1_SFF_5_QD ;
    wire stateArray_S13reg_gff_1_SFF_6_QD ;
    wire stateArray_S13reg_gff_1_SFF_7_QD ;
    wire stateArray_S20reg_gff_1_SFF_0_QD ;
    wire stateArray_S20reg_gff_1_SFF_1_QD ;
    wire stateArray_S20reg_gff_1_SFF_2_QD ;
    wire stateArray_S20reg_gff_1_SFF_3_QD ;
    wire stateArray_S20reg_gff_1_SFF_4_QD ;
    wire stateArray_S20reg_gff_1_SFF_5_QD ;
    wire stateArray_S20reg_gff_1_SFF_6_QD ;
    wire stateArray_S20reg_gff_1_SFF_7_QD ;
    wire stateArray_S21reg_gff_1_SFF_0_QD ;
    wire stateArray_S21reg_gff_1_SFF_1_QD ;
    wire stateArray_S21reg_gff_1_SFF_2_QD ;
    wire stateArray_S21reg_gff_1_SFF_3_QD ;
    wire stateArray_S21reg_gff_1_SFF_4_QD ;
    wire stateArray_S21reg_gff_1_SFF_5_QD ;
    wire stateArray_S21reg_gff_1_SFF_6_QD ;
    wire stateArray_S21reg_gff_1_SFF_7_QD ;
    wire stateArray_S22reg_gff_1_SFF_0_QD ;
    wire stateArray_S22reg_gff_1_SFF_1_QD ;
    wire stateArray_S22reg_gff_1_SFF_2_QD ;
    wire stateArray_S22reg_gff_1_SFF_3_QD ;
    wire stateArray_S22reg_gff_1_SFF_4_QD ;
    wire stateArray_S22reg_gff_1_SFF_5_QD ;
    wire stateArray_S22reg_gff_1_SFF_6_QD ;
    wire stateArray_S22reg_gff_1_SFF_7_QD ;
    wire stateArray_S23reg_gff_1_SFF_0_QD ;
    wire stateArray_S23reg_gff_1_SFF_1_QD ;
    wire stateArray_S23reg_gff_1_SFF_2_QD ;
    wire stateArray_S23reg_gff_1_SFF_3_QD ;
    wire stateArray_S23reg_gff_1_SFF_4_QD ;
    wire stateArray_S23reg_gff_1_SFF_5_QD ;
    wire stateArray_S23reg_gff_1_SFF_6_QD ;
    wire stateArray_S23reg_gff_1_SFF_7_QD ;
    wire stateArray_S30reg_gff_1_SFF_0_QD ;
    wire stateArray_S30reg_gff_1_SFF_1_QD ;
    wire stateArray_S30reg_gff_1_SFF_2_QD ;
    wire stateArray_S30reg_gff_1_SFF_3_QD ;
    wire stateArray_S30reg_gff_1_SFF_4_QD ;
    wire stateArray_S30reg_gff_1_SFF_5_QD ;
    wire stateArray_S30reg_gff_1_SFF_6_QD ;
    wire stateArray_S30reg_gff_1_SFF_7_QD ;
    wire stateArray_S31reg_gff_1_SFF_0_QD ;
    wire stateArray_S31reg_gff_1_SFF_1_QD ;
    wire stateArray_S31reg_gff_1_SFF_2_QD ;
    wire stateArray_S31reg_gff_1_SFF_3_QD ;
    wire stateArray_S31reg_gff_1_SFF_4_QD ;
    wire stateArray_S31reg_gff_1_SFF_5_QD ;
    wire stateArray_S31reg_gff_1_SFF_6_QD ;
    wire stateArray_S31reg_gff_1_SFF_7_QD ;
    wire stateArray_S32reg_gff_1_SFF_0_QD ;
    wire stateArray_S32reg_gff_1_SFF_1_QD ;
    wire stateArray_S32reg_gff_1_SFF_2_QD ;
    wire stateArray_S32reg_gff_1_SFF_3_QD ;
    wire stateArray_S32reg_gff_1_SFF_4_QD ;
    wire stateArray_S32reg_gff_1_SFF_5_QD ;
    wire stateArray_S32reg_gff_1_SFF_6_QD ;
    wire stateArray_S32reg_gff_1_SFF_7_QD ;
    wire stateArray_S33reg_gff_1_SFF_0_QD ;
    wire stateArray_S33reg_gff_1_SFF_1_QD ;
    wire stateArray_S33reg_gff_1_SFF_2_QD ;
    wire stateArray_S33reg_gff_1_SFF_3_QD ;
    wire stateArray_S33reg_gff_1_SFF_4_QD ;
    wire stateArray_S33reg_gff_1_SFF_5_QD ;
    wire stateArray_S33reg_gff_1_SFF_6_QD ;
    wire stateArray_S33reg_gff_1_SFF_7_QD ;
    wire MUX_StateInMC_n7 ;
    wire MUX_StateInMC_n6 ;
    wire MUX_StateInMC_n5 ;
    wire KeyArray_n55 ;
    wire KeyArray_n54 ;
    wire KeyArray_n53 ;
    wire KeyArray_n52 ;
    wire KeyArray_n51 ;
    wire KeyArray_n50 ;
    wire KeyArray_n49 ;
    wire KeyArray_n48 ;
    wire KeyArray_n47 ;
    wire KeyArray_n46 ;
    wire KeyArray_n45 ;
    wire KeyArray_n44 ;
    wire KeyArray_n43 ;
    wire KeyArray_n42 ;
    wire KeyArray_n41 ;
    wire KeyArray_n40 ;
    wire KeyArray_n39 ;
    wire KeyArray_n38 ;
    wire KeyArray_n37 ;
    wire KeyArray_n36 ;
    wire KeyArray_n35 ;
    wire KeyArray_n34 ;
    wire KeyArray_n33 ;
    wire KeyArray_n32 ;
    wire KeyArray_n31 ;
    wire KeyArray_n30 ;
    wire KeyArray_n29 ;
    wire KeyArray_n28 ;
    wire KeyArray_n27 ;
    wire KeyArray_n26 ;
    wire KeyArray_n25 ;
    wire KeyArray_n24 ;
    wire KeyArray_n23 ;
    wire KeyArray_n22 ;
    wire KeyArray_outS01ser_0_ ;
    wire KeyArray_outS01ser_1_ ;
    wire KeyArray_outS01ser_2_ ;
    wire KeyArray_outS01ser_3_ ;
    wire KeyArray_outS01ser_4_ ;
    wire KeyArray_outS01ser_5_ ;
    wire KeyArray_outS01ser_6_ ;
    wire KeyArray_outS01ser_7_ ;
    wire KeyArray_S00reg_gff_1_SFF_0_n5 ;
    wire KeyArray_S00reg_gff_1_SFF_0_QD ;
    wire KeyArray_S00reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S00reg_gff_1_SFF_1_QD ;
    wire KeyArray_S00reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S00reg_gff_1_SFF_2_QD ;
    wire KeyArray_S00reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S00reg_gff_1_SFF_3_QD ;
    wire KeyArray_S00reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S00reg_gff_1_SFF_4_QD ;
    wire KeyArray_S00reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S00reg_gff_1_SFF_5_QD ;
    wire KeyArray_S00reg_gff_1_SFF_6_n6 ;
    wire KeyArray_S00reg_gff_1_SFF_6_QD ;
    wire KeyArray_S00reg_gff_1_SFF_7_n6 ;
    wire KeyArray_S00reg_gff_1_SFF_7_QD ;
    wire KeyArray_S01reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S01reg_gff_1_SFF_0_QD ;
    wire KeyArray_S01reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S01reg_gff_1_SFF_1_QD ;
    wire KeyArray_S01reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S01reg_gff_1_SFF_2_QD ;
    wire KeyArray_S01reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S01reg_gff_1_SFF_3_QD ;
    wire KeyArray_S01reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S01reg_gff_1_SFF_4_QD ;
    wire KeyArray_S01reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S01reg_gff_1_SFF_5_QD ;
    wire KeyArray_S01reg_gff_1_SFF_6_n6 ;
    wire KeyArray_S01reg_gff_1_SFF_6_QD ;
    wire KeyArray_S01reg_gff_1_SFF_7_n6 ;
    wire KeyArray_S01reg_gff_1_SFF_7_QD ;
    wire KeyArray_S02reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S02reg_gff_1_SFF_0_QD ;
    wire KeyArray_S02reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S02reg_gff_1_SFF_1_QD ;
    wire KeyArray_S02reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S02reg_gff_1_SFF_2_QD ;
    wire KeyArray_S02reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S02reg_gff_1_SFF_3_QD ;
    wire KeyArray_S02reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S02reg_gff_1_SFF_4_QD ;
    wire KeyArray_S02reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S02reg_gff_1_SFF_5_QD ;
    wire KeyArray_S02reg_gff_1_SFF_6_n6 ;
    wire KeyArray_S02reg_gff_1_SFF_6_QD ;
    wire KeyArray_S02reg_gff_1_SFF_7_n6 ;
    wire KeyArray_S02reg_gff_1_SFF_7_QD ;
    wire KeyArray_S03reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S03reg_gff_1_SFF_0_QD ;
    wire KeyArray_S03reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S03reg_gff_1_SFF_1_QD ;
    wire KeyArray_S03reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S03reg_gff_1_SFF_2_QD ;
    wire KeyArray_S03reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S03reg_gff_1_SFF_3_QD ;
    wire KeyArray_S03reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S03reg_gff_1_SFF_4_QD ;
    wire KeyArray_S03reg_gff_1_SFF_5_n5 ;
    wire KeyArray_S03reg_gff_1_SFF_5_QD ;
    wire KeyArray_S03reg_gff_1_SFF_6_n5 ;
    wire KeyArray_S03reg_gff_1_SFF_6_QD ;
    wire KeyArray_S03reg_gff_1_SFF_7_n5 ;
    wire KeyArray_S03reg_gff_1_SFF_7_QD ;
    wire KeyArray_S10reg_gff_1_SFF_0_n5 ;
    wire KeyArray_S10reg_gff_1_SFF_0_QD ;
    wire KeyArray_S10reg_gff_1_SFF_1_n5 ;
    wire KeyArray_S10reg_gff_1_SFF_1_QD ;
    wire KeyArray_S10reg_gff_1_SFF_2_n5 ;
    wire KeyArray_S10reg_gff_1_SFF_2_QD ;
    wire KeyArray_S10reg_gff_1_SFF_3_n5 ;
    wire KeyArray_S10reg_gff_1_SFF_3_QD ;
    wire KeyArray_S10reg_gff_1_SFF_4_n5 ;
    wire KeyArray_S10reg_gff_1_SFF_4_QD ;
    wire KeyArray_S10reg_gff_1_SFF_5_n5 ;
    wire KeyArray_S10reg_gff_1_SFF_5_QD ;
    wire KeyArray_S10reg_gff_1_SFF_6_n5 ;
    wire KeyArray_S10reg_gff_1_SFF_6_QD ;
    wire KeyArray_S10reg_gff_1_SFF_7_n5 ;
    wire KeyArray_S10reg_gff_1_SFF_7_QD ;
    wire KeyArray_S11reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S11reg_gff_1_SFF_0_QD ;
    wire KeyArray_S11reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S11reg_gff_1_SFF_1_QD ;
    wire KeyArray_S11reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S11reg_gff_1_SFF_2_QD ;
    wire KeyArray_S11reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S11reg_gff_1_SFF_3_QD ;
    wire KeyArray_S11reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S11reg_gff_1_SFF_4_QD ;
    wire KeyArray_S11reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S11reg_gff_1_SFF_5_QD ;
    wire KeyArray_S11reg_gff_1_SFF_6_n6 ;
    wire KeyArray_S11reg_gff_1_SFF_6_QD ;
    wire KeyArray_S11reg_gff_1_SFF_7_n6 ;
    wire KeyArray_S11reg_gff_1_SFF_7_QD ;
    wire KeyArray_S12reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S12reg_gff_1_SFF_0_QD ;
    wire KeyArray_S12reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S12reg_gff_1_SFF_1_QD ;
    wire KeyArray_S12reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S12reg_gff_1_SFF_2_QD ;
    wire KeyArray_S12reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S12reg_gff_1_SFF_3_QD ;
    wire KeyArray_S12reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S12reg_gff_1_SFF_4_QD ;
    wire KeyArray_S12reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S12reg_gff_1_SFF_5_QD ;
    wire KeyArray_S12reg_gff_1_SFF_6_n6 ;
    wire KeyArray_S12reg_gff_1_SFF_6_QD ;
    wire KeyArray_S12reg_gff_1_SFF_7_n6 ;
    wire KeyArray_S12reg_gff_1_SFF_7_QD ;
    wire KeyArray_S13reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S13reg_gff_1_SFF_0_QD ;
    wire KeyArray_S13reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S13reg_gff_1_SFF_1_QD ;
    wire KeyArray_S13reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S13reg_gff_1_SFF_2_QD ;
    wire KeyArray_S13reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S13reg_gff_1_SFF_3_QD ;
    wire KeyArray_S13reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S13reg_gff_1_SFF_4_QD ;
    wire KeyArray_S13reg_gff_1_SFF_5_n5 ;
    wire KeyArray_S13reg_gff_1_SFF_5_QD ;
    wire KeyArray_S13reg_gff_1_SFF_6_n5 ;
    wire KeyArray_S13reg_gff_1_SFF_6_QD ;
    wire KeyArray_S13reg_gff_1_SFF_7_n5 ;
    wire KeyArray_S13reg_gff_1_SFF_7_QD ;
    wire KeyArray_S20reg_gff_1_SFF_0_n5 ;
    wire KeyArray_S20reg_gff_1_SFF_0_QD ;
    wire KeyArray_S20reg_gff_1_SFF_1_n5 ;
    wire KeyArray_S20reg_gff_1_SFF_1_QD ;
    wire KeyArray_S20reg_gff_1_SFF_2_n5 ;
    wire KeyArray_S20reg_gff_1_SFF_2_QD ;
    wire KeyArray_S20reg_gff_1_SFF_3_n5 ;
    wire KeyArray_S20reg_gff_1_SFF_3_QD ;
    wire KeyArray_S20reg_gff_1_SFF_4_n5 ;
    wire KeyArray_S20reg_gff_1_SFF_4_QD ;
    wire KeyArray_S20reg_gff_1_SFF_5_n5 ;
    wire KeyArray_S20reg_gff_1_SFF_5_QD ;
    wire KeyArray_S20reg_gff_1_SFF_6_n5 ;
    wire KeyArray_S20reg_gff_1_SFF_6_QD ;
    wire KeyArray_S20reg_gff_1_SFF_7_n5 ;
    wire KeyArray_S20reg_gff_1_SFF_7_QD ;
    wire KeyArray_S21reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S21reg_gff_1_SFF_0_QD ;
    wire KeyArray_S21reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S21reg_gff_1_SFF_1_QD ;
    wire KeyArray_S21reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S21reg_gff_1_SFF_2_QD ;
    wire KeyArray_S21reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S21reg_gff_1_SFF_3_QD ;
    wire KeyArray_S21reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S21reg_gff_1_SFF_4_QD ;
    wire KeyArray_S21reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S21reg_gff_1_SFF_5_QD ;
    wire KeyArray_S21reg_gff_1_SFF_6_n6 ;
    wire KeyArray_S21reg_gff_1_SFF_6_QD ;
    wire KeyArray_S21reg_gff_1_SFF_7_n6 ;
    wire KeyArray_S21reg_gff_1_SFF_7_QD ;
    wire KeyArray_S22reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S22reg_gff_1_SFF_0_QD ;
    wire KeyArray_S22reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S22reg_gff_1_SFF_1_QD ;
    wire KeyArray_S22reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S22reg_gff_1_SFF_2_QD ;
    wire KeyArray_S22reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S22reg_gff_1_SFF_3_QD ;
    wire KeyArray_S22reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S22reg_gff_1_SFF_4_QD ;
    wire KeyArray_S22reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S22reg_gff_1_SFF_5_QD ;
    wire KeyArray_S22reg_gff_1_SFF_6_n6 ;
    wire KeyArray_S22reg_gff_1_SFF_6_QD ;
    wire KeyArray_S22reg_gff_1_SFF_7_n6 ;
    wire KeyArray_S22reg_gff_1_SFF_7_QD ;
    wire KeyArray_S23reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S23reg_gff_1_SFF_0_QD ;
    wire KeyArray_S23reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S23reg_gff_1_SFF_1_QD ;
    wire KeyArray_S23reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S23reg_gff_1_SFF_2_QD ;
    wire KeyArray_S23reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S23reg_gff_1_SFF_3_QD ;
    wire KeyArray_S23reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S23reg_gff_1_SFF_4_QD ;
    wire KeyArray_S23reg_gff_1_SFF_5_n5 ;
    wire KeyArray_S23reg_gff_1_SFF_5_QD ;
    wire KeyArray_S23reg_gff_1_SFF_6_n5 ;
    wire KeyArray_S23reg_gff_1_SFF_6_QD ;
    wire KeyArray_S23reg_gff_1_SFF_7_n5 ;
    wire KeyArray_S23reg_gff_1_SFF_7_QD ;
    wire KeyArray_S30reg_gff_1_SFF_0_n5 ;
    wire KeyArray_S30reg_gff_1_SFF_0_QD ;
    wire KeyArray_S30reg_gff_1_SFF_1_n5 ;
    wire KeyArray_S30reg_gff_1_SFF_1_QD ;
    wire KeyArray_S30reg_gff_1_SFF_2_n5 ;
    wire KeyArray_S30reg_gff_1_SFF_2_QD ;
    wire KeyArray_S30reg_gff_1_SFF_3_n5 ;
    wire KeyArray_S30reg_gff_1_SFF_3_QD ;
    wire KeyArray_S30reg_gff_1_SFF_4_n5 ;
    wire KeyArray_S30reg_gff_1_SFF_4_QD ;
    wire KeyArray_S30reg_gff_1_SFF_5_n5 ;
    wire KeyArray_S30reg_gff_1_SFF_5_QD ;
    wire KeyArray_S30reg_gff_1_SFF_6_n5 ;
    wire KeyArray_S30reg_gff_1_SFF_6_QD ;
    wire KeyArray_S30reg_gff_1_SFF_7_n5 ;
    wire KeyArray_S30reg_gff_1_SFF_7_QD ;
    wire KeyArray_S31reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S31reg_gff_1_SFF_0_QD ;
    wire KeyArray_S31reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S31reg_gff_1_SFF_1_QD ;
    wire KeyArray_S31reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S31reg_gff_1_SFF_2_QD ;
    wire KeyArray_S31reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S31reg_gff_1_SFF_3_QD ;
    wire KeyArray_S31reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S31reg_gff_1_SFF_4_QD ;
    wire KeyArray_S31reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S31reg_gff_1_SFF_5_QD ;
    wire KeyArray_S31reg_gff_1_SFF_6_n6 ;
    wire KeyArray_S31reg_gff_1_SFF_6_QD ;
    wire KeyArray_S31reg_gff_1_SFF_7_n6 ;
    wire KeyArray_S31reg_gff_1_SFF_7_QD ;
    wire KeyArray_S32reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S32reg_gff_1_SFF_0_QD ;
    wire KeyArray_S32reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S32reg_gff_1_SFF_1_QD ;
    wire KeyArray_S32reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S32reg_gff_1_SFF_2_QD ;
    wire KeyArray_S32reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S32reg_gff_1_SFF_3_QD ;
    wire KeyArray_S32reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S32reg_gff_1_SFF_4_QD ;
    wire KeyArray_S32reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S32reg_gff_1_SFF_5_QD ;
    wire KeyArray_S32reg_gff_1_SFF_6_n5 ;
    wire KeyArray_S32reg_gff_1_SFF_6_QD ;
    wire KeyArray_S32reg_gff_1_SFF_7_n5 ;
    wire KeyArray_S32reg_gff_1_SFF_7_QD ;
    wire KeyArray_S33reg_gff_1_SFF_0_n5 ;
    wire KeyArray_S33reg_gff_1_SFF_0_QD ;
    wire KeyArray_S33reg_gff_1_SFF_1_n5 ;
    wire KeyArray_S33reg_gff_1_SFF_1_QD ;
    wire KeyArray_S33reg_gff_1_SFF_2_n5 ;
    wire KeyArray_S33reg_gff_1_SFF_2_QD ;
    wire KeyArray_S33reg_gff_1_SFF_3_n5 ;
    wire KeyArray_S33reg_gff_1_SFF_3_QD ;
    wire KeyArray_S33reg_gff_1_SFF_4_n5 ;
    wire KeyArray_S33reg_gff_1_SFF_4_QD ;
    wire KeyArray_S33reg_gff_1_SFF_5_n5 ;
    wire KeyArray_S33reg_gff_1_SFF_5_QD ;
    wire KeyArray_S33reg_gff_1_SFF_6_n5 ;
    wire KeyArray_S33reg_gff_1_SFF_6_QD ;
    wire KeyArray_S33reg_gff_1_SFF_7_n5 ;
    wire KeyArray_S33reg_gff_1_SFF_7_QD ;
    wire MixColumns_line0_n16 ;
    wire MixColumns_line0_n15 ;
    wire MixColumns_line0_n14 ;
    wire MixColumns_line0_n13 ;
    wire MixColumns_line0_n12 ;
    wire MixColumns_line0_n11 ;
    wire MixColumns_line0_n10 ;
    wire MixColumns_line0_n9 ;
    wire MixColumns_line0_n8 ;
    wire MixColumns_line0_n7 ;
    wire MixColumns_line0_n6 ;
    wire MixColumns_line0_n5 ;
    wire MixColumns_line0_n4 ;
    wire MixColumns_line0_n3 ;
    wire MixColumns_line0_n2 ;
    wire MixColumns_line0_n1 ;
    wire MixColumns_line1_n16 ;
    wire MixColumns_line1_n15 ;
    wire MixColumns_line1_n14 ;
    wire MixColumns_line1_n13 ;
    wire MixColumns_line1_n12 ;
    wire MixColumns_line1_n11 ;
    wire MixColumns_line1_n10 ;
    wire MixColumns_line1_n9 ;
    wire MixColumns_line1_n8 ;
    wire MixColumns_line1_n7 ;
    wire MixColumns_line1_n6 ;
    wire MixColumns_line1_n5 ;
    wire MixColumns_line1_n4 ;
    wire MixColumns_line1_n3 ;
    wire MixColumns_line1_n2 ;
    wire MixColumns_line1_n1 ;
    wire MixColumns_line1_S02_1_ ;
    wire MixColumns_line1_S02_3_ ;
    wire MixColumns_line1_S02_4_ ;
    wire MixColumns_line2_n16 ;
    wire MixColumns_line2_n15 ;
    wire MixColumns_line2_n14 ;
    wire MixColumns_line2_n13 ;
    wire MixColumns_line2_n12 ;
    wire MixColumns_line2_n11 ;
    wire MixColumns_line2_n10 ;
    wire MixColumns_line2_n9 ;
    wire MixColumns_line2_n8 ;
    wire MixColumns_line2_n7 ;
    wire MixColumns_line2_n6 ;
    wire MixColumns_line2_n5 ;
    wire MixColumns_line2_n4 ;
    wire MixColumns_line2_n3 ;
    wire MixColumns_line2_n2 ;
    wire MixColumns_line2_n1 ;
    wire MixColumns_line2_S02_1_ ;
    wire MixColumns_line2_S02_3_ ;
    wire MixColumns_line2_S02_4_ ;
    wire MixColumns_line3_n16 ;
    wire MixColumns_line3_n15 ;
    wire MixColumns_line3_n14 ;
    wire MixColumns_line3_n13 ;
    wire MixColumns_line3_n12 ;
    wire MixColumns_line3_n11 ;
    wire MixColumns_line3_n10 ;
    wire MixColumns_line3_n9 ;
    wire MixColumns_line3_n8 ;
    wire MixColumns_line3_n7 ;
    wire MixColumns_line3_n6 ;
    wire MixColumns_line3_n5 ;
    wire MixColumns_line3_n4 ;
    wire MixColumns_line3_n3 ;
    wire MixColumns_line3_n2 ;
    wire MixColumns_line3_n1 ;
    wire MixColumns_line3_S02_1_ ;
    wire MixColumns_line3_S02_3_ ;
    wire MixColumns_line3_S02_4_ ;
    wire MixColumns_line3_timesTHREE_input2_1_ ;
    wire MixColumns_line3_timesTHREE_input2_3_ ;
    wire MixColumns_line3_timesTHREE_input2_4_ ;
    wire calcRCon_n38 ;
    wire calcRCon_n37 ;
    wire calcRCon_n36 ;
    wire calcRCon_n35 ;
    wire calcRCon_n34 ;
    wire calcRCon_n33 ;
    wire calcRCon_n32 ;
    wire calcRCon_n31 ;
    wire calcRCon_n30 ;
    wire calcRCon_n29 ;
    wire calcRCon_n28 ;
    wire calcRCon_n27 ;
    wire calcRCon_n26 ;
    wire calcRCon_n25 ;
    wire calcRCon_n24 ;
    wire calcRCon_n23 ;
    wire calcRCon_n22 ;
    wire calcRCon_n21 ;
    wire calcRCon_n20 ;
    wire calcRCon_n19 ;
    wire calcRCon_n18 ;
    wire calcRCon_n17 ;
    wire calcRCon_n10 ;
    wire calcRCon_n9 ;
    wire calcRCon_n8 ;
    wire calcRCon_n7 ;
    wire calcRCon_n6 ;
    wire calcRCon_n5 ;
    wire calcRCon_n3 ;
    wire calcRCon_n11 ;
    wire calcRCon_n44 ;
    wire calcRCon_n16 ;
    wire calcRCon_n45 ;
    wire calcRCon_n46 ;
    wire calcRCon_n47 ;
    wire calcRCon_n15 ;
    wire calcRCon_n48 ;
    wire calcRCon_n12 ;
    wire calcRCon_n49 ;
    wire calcRCon_n14 ;
    wire calcRCon_n50 ;
    wire calcRCon_n13 ;
    wire calcRCon_s_current_state_0_ ;
    wire calcRCon_s_current_state_1_ ;
    wire calcRCon_s_current_state_2_ ;
    wire calcRCon_s_current_state_3_ ;
    wire calcRCon_s_current_state_4_ ;
    wire calcRCon_s_current_state_5_ ;
    wire calcRCon_s_current_state_6_ ;
    wire calcRCon_n51 ;
    wire Inst_bSbox_L29 ;
    wire Inst_bSbox_L28 ;
    wire Inst_bSbox_L27 ;
    wire Inst_bSbox_L26 ;
    wire Inst_bSbox_L25 ;
    wire Inst_bSbox_L24 ;
    wire Inst_bSbox_L23 ;
    wire Inst_bSbox_L22 ;
    wire Inst_bSbox_L21 ;
    wire Inst_bSbox_L20 ;
    wire Inst_bSbox_L19 ;
    wire Inst_bSbox_L18 ;
    wire Inst_bSbox_L17 ;
    wire Inst_bSbox_L16 ;
    wire Inst_bSbox_L15 ;
    wire Inst_bSbox_L14 ;
    wire Inst_bSbox_L13 ;
    wire Inst_bSbox_L12 ;
    wire Inst_bSbox_L11 ;
    wire Inst_bSbox_L10 ;
    wire Inst_bSbox_L9 ;
    wire Inst_bSbox_L8 ;
    wire Inst_bSbox_L7 ;
    wire Inst_bSbox_L6 ;
    wire Inst_bSbox_L5 ;
    wire Inst_bSbox_L4 ;
    wire Inst_bSbox_L3 ;
    wire Inst_bSbox_L2 ;
    wire Inst_bSbox_L1 ;
    wire Inst_bSbox_L0 ;
    wire Inst_bSbox_M63 ;
    wire Inst_bSbox_M62 ;
    wire Inst_bSbox_M61 ;
    wire Inst_bSbox_M60 ;
    wire Inst_bSbox_M59 ;
    wire Inst_bSbox_M58 ;
    wire Inst_bSbox_M57 ;
    wire Inst_bSbox_M56 ;
    wire Inst_bSbox_M55 ;
    wire Inst_bSbox_M54 ;
    wire Inst_bSbox_M53 ;
    wire Inst_bSbox_M52 ;
    wire Inst_bSbox_M51 ;
    wire Inst_bSbox_M50 ;
    wire Inst_bSbox_M49 ;
    wire Inst_bSbox_M48 ;
    wire Inst_bSbox_M47 ;
    wire Inst_bSbox_M46 ;
    wire Inst_bSbox_M45 ;
    wire Inst_bSbox_M44 ;
    wire Inst_bSbox_M43 ;
    wire Inst_bSbox_M42 ;
    wire Inst_bSbox_M41 ;
    wire Inst_bSbox_M40 ;
    wire Inst_bSbox_M39 ;
    wire Inst_bSbox_M38 ;
    wire Inst_bSbox_M37 ;
    wire Inst_bSbox_M36 ;
    wire Inst_bSbox_M35 ;
    wire Inst_bSbox_M34 ;
    wire Inst_bSbox_M33 ;
    wire Inst_bSbox_M32 ;
    wire Inst_bSbox_M31 ;
    wire Inst_bSbox_M30 ;
    wire Inst_bSbox_M29 ;
    wire Inst_bSbox_M28 ;
    wire Inst_bSbox_M27 ;
    wire Inst_bSbox_M26 ;
    wire Inst_bSbox_M25 ;
    wire Inst_bSbox_M24 ;
    wire Inst_bSbox_M23 ;
    wire Inst_bSbox_M22 ;
    wire Inst_bSbox_M21 ;
    wire Inst_bSbox_M20 ;
    wire Inst_bSbox_M19 ;
    wire Inst_bSbox_M18 ;
    wire Inst_bSbox_M17 ;
    wire Inst_bSbox_M16 ;
    wire Inst_bSbox_M15 ;
    wire Inst_bSbox_M14 ;
    wire Inst_bSbox_M13 ;
    wire Inst_bSbox_M12 ;
    wire Inst_bSbox_M11 ;
    wire Inst_bSbox_M10 ;
    wire Inst_bSbox_M9 ;
    wire Inst_bSbox_M8 ;
    wire Inst_bSbox_M7 ;
    wire Inst_bSbox_M6 ;
    wire Inst_bSbox_M5 ;
    wire Inst_bSbox_M4 ;
    wire Inst_bSbox_M3 ;
    wire Inst_bSbox_M2 ;
    wire Inst_bSbox_M1 ;
    wire Inst_bSbox_T27 ;
    wire Inst_bSbox_T26 ;
    wire Inst_bSbox_T25 ;
    wire Inst_bSbox_T24 ;
    wire Inst_bSbox_T23 ;
    wire Inst_bSbox_T22 ;
    wire Inst_bSbox_T21 ;
    wire Inst_bSbox_T20 ;
    wire Inst_bSbox_T19 ;
    wire Inst_bSbox_T18 ;
    wire Inst_bSbox_T17 ;
    wire Inst_bSbox_T16 ;
    wire Inst_bSbox_T15 ;
    wire Inst_bSbox_T14 ;
    wire Inst_bSbox_T13 ;
    wire Inst_bSbox_T12 ;
    wire Inst_bSbox_T11 ;
    wire Inst_bSbox_T10 ;
    wire Inst_bSbox_T9 ;
    wire Inst_bSbox_T8 ;
    wire Inst_bSbox_T7 ;
    wire Inst_bSbox_T6 ;
    wire Inst_bSbox_T5 ;
    wire Inst_bSbox_T4 ;
    wire Inst_bSbox_T3 ;
    wire Inst_bSbox_T2 ;
    wire Inst_bSbox_T1 ;
    wire [7:0] SboxOut ;
    wire [7:0] StateOutXORroundKey ;
    wire [7:0] StateIn ;
    wire [31:0] StateInMC ;
    wire [31:0] MCout ;
    wire [7:0] keyStateIn ;
    wire [7:0] roundConstant ;
    wire [7:0] keySBIn ;
    wire [7:0] SboxIn ;
    wire [7:0] stateArray_input_MC ;
    wire [7:0] stateArray_outS30ser_MC ;
    wire [7:0] stateArray_outS20ser_MC ;
    wire [7:0] stateArray_outS10ser_MC ;
    wire [7:0] stateArray_inS33ser ;
    wire [7:0] stateArray_inS32ser ;
    wire [7:0] stateArray_inS31ser ;
    wire [7:0] stateArray_inS30ser ;
    wire [7:0] stateArray_inS23ser ;
    wire [7:0] stateArray_inS22ser ;
    wire [7:0] stateArray_inS21ser ;
    wire [7:0] stateArray_inS20ser ;
    wire [7:0] stateArray_inS13ser ;
    wire [7:0] stateArray_inS12ser ;
    wire [7:0] stateArray_inS11ser ;
    wire [7:0] stateArray_inS10ser ;
    wire [7:0] stateArray_inS03ser ;
    wire [7:0] stateArray_inS02ser ;
    wire [7:0] stateArray_inS01ser ;
    wire [7:0] stateArray_inS00ser ;
    wire [7:0] KeyArray_outS01ser_p ;
    wire [7:0] KeyArray_outS01ser_XOR_00 ;
    wire [7:0] KeyArray_outS33ser ;
    wire [7:0] KeyArray_inS33ser ;
    wire [7:0] KeyArray_outS32ser ;
    wire [7:0] KeyArray_inS32ser ;
    wire [7:0] KeyArray_outS31ser ;
    wire [7:0] KeyArray_inS31ser ;
    wire [7:0] KeyArray_outS30ser ;
    wire [7:0] KeyArray_inS30par ;
    wire [7:0] KeyArray_inS30ser ;
    wire [7:0] KeyArray_outS23ser ;
    wire [7:0] KeyArray_inS23ser ;
    wire [7:0] KeyArray_outS22ser ;
    wire [7:0] KeyArray_inS22ser ;
    wire [7:0] KeyArray_outS21ser ;
    wire [7:0] KeyArray_inS21ser ;
    wire [7:0] KeyArray_outS20ser ;
    wire [7:0] KeyArray_inS20ser ;
    wire [7:0] KeyArray_inS13ser ;
    wire [7:0] KeyArray_outS12ser ;
    wire [7:0] KeyArray_inS12ser ;
    wire [7:0] KeyArray_outS11ser ;
    wire [7:0] KeyArray_inS11ser ;
    wire [7:0] KeyArray_outS10ser ;
    wire [7:0] KeyArray_inS10ser ;
    wire [7:0] KeyArray_outS03ser ;
    wire [7:0] KeyArray_inS03ser ;
    wire [7:0] KeyArray_outS02ser ;
    wire [7:0] KeyArray_inS02ser ;
    wire [7:0] KeyArray_inS01ser ;
    wire [7:0] KeyArray_inS00ser ;
    wire [7:0] MixColumns_line0_S13 ;
    wire [4:1] MixColumns_line0_S02 ;
    wire [4:1] MixColumns_line0_timesTHREE_input2 ;
    wire [7:0] MixColumns_line1_S13 ;
    wire [4:1] MixColumns_line1_timesTHREE_input2 ;
    wire [7:0] MixColumns_line2_S13 ;
    wire [4:1] MixColumns_line2_timesTHREE_input2 ;
    wire [7:0] MixColumns_line3_S13 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1986 ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1989 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1995 ;
    wire new_AGEMA_signal_1996 ;
    wire new_AGEMA_signal_1998 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2004 ;
    wire new_AGEMA_signal_2005 ;
    wire new_AGEMA_signal_2006 ;
    wire new_AGEMA_signal_2007 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2014 ;
    wire new_AGEMA_signal_2015 ;
    wire new_AGEMA_signal_2016 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2051 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2086 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2097 ;
    wire new_AGEMA_signal_2098 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2102 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2104 ;
    wire new_AGEMA_signal_2105 ;
    wire new_AGEMA_signal_2106 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2114 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2116 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2120 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2122 ;
    wire new_AGEMA_signal_2123 ;
    wire new_AGEMA_signal_2124 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2127 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2130 ;
    wire new_AGEMA_signal_2131 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2133 ;
    wire new_AGEMA_signal_2134 ;
    wire new_AGEMA_signal_2135 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2139 ;
    wire new_AGEMA_signal_2140 ;
    wire new_AGEMA_signal_2141 ;
    wire new_AGEMA_signal_2142 ;
    wire new_AGEMA_signal_2143 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2147 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2150 ;
    wire new_AGEMA_signal_2151 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2156 ;
    wire new_AGEMA_signal_2159 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2168 ;
    wire new_AGEMA_signal_2171 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2183 ;
    wire new_AGEMA_signal_2186 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2195 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2222 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2228 ;
    wire new_AGEMA_signal_2231 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2240 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2264 ;
    wire new_AGEMA_signal_2267 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2276 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2282 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2294 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2300 ;
    wire new_AGEMA_signal_2303 ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2312 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2324 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2330 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2375 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2826 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2914 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2926 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2934 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2942 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2950 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2962 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2966 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2970 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2976 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2988 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2992 ;
    wire new_AGEMA_signal_2993 ;
    wire new_AGEMA_signal_2994 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2996 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3000 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3004 ;
    wire new_AGEMA_signal_3005 ;
    wire new_AGEMA_signal_3006 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3012 ;
    wire new_AGEMA_signal_3013 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3016 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3020 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3022 ;
    wire new_AGEMA_signal_3023 ;
    wire new_AGEMA_signal_3024 ;
    wire new_AGEMA_signal_3025 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3028 ;
    wire new_AGEMA_signal_3029 ;
    wire new_AGEMA_signal_3030 ;
    wire new_AGEMA_signal_3031 ;
    wire new_AGEMA_signal_3032 ;
    wire new_AGEMA_signal_3033 ;
    wire new_AGEMA_signal_3034 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3036 ;
    wire new_AGEMA_signal_3037 ;
    wire new_AGEMA_signal_3038 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3040 ;
    wire new_AGEMA_signal_3041 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3043 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3056 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3060 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3074 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3078 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3086 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3132 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3139 ;
    wire new_AGEMA_signal_3140 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3374 ;
    wire new_AGEMA_signal_3375 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3391 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3411 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3418 ;
    wire new_AGEMA_signal_3419 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3423 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3427 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3447 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3483 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_3723 ;
    wire new_AGEMA_signal_3724 ;
    wire new_AGEMA_signal_3725 ;
    wire new_AGEMA_signal_3726 ;
    wire new_AGEMA_signal_3727 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3730 ;
    wire new_AGEMA_signal_3731 ;
    wire new_AGEMA_signal_3732 ;
    wire new_AGEMA_signal_3733 ;
    wire new_AGEMA_signal_3734 ;
    wire new_AGEMA_signal_3735 ;
    wire new_AGEMA_signal_3736 ;
    wire new_AGEMA_signal_3737 ;
    wire new_AGEMA_signal_3738 ;
    wire new_AGEMA_signal_3739 ;
    wire new_AGEMA_signal_3740 ;
    wire new_AGEMA_signal_3741 ;
    wire new_AGEMA_signal_3742 ;
    wire new_AGEMA_signal_3743 ;
    wire new_AGEMA_signal_3744 ;
    wire new_AGEMA_signal_3745 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3747 ;
    wire new_AGEMA_signal_3748 ;
    wire new_AGEMA_signal_3749 ;
    wire new_AGEMA_signal_3750 ;
    wire new_AGEMA_signal_3751 ;
    wire new_AGEMA_signal_3752 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3754 ;
    wire new_AGEMA_signal_3755 ;
    wire new_AGEMA_signal_3756 ;
    wire new_AGEMA_signal_3757 ;
    wire new_AGEMA_signal_3758 ;
    wire new_AGEMA_signal_3759 ;
    wire new_AGEMA_signal_3760 ;
    wire new_AGEMA_signal_3761 ;
    wire new_AGEMA_signal_3762 ;
    wire new_AGEMA_signal_3763 ;
    wire new_AGEMA_signal_3764 ;
    wire new_AGEMA_signal_3765 ;
    wire new_AGEMA_signal_3766 ;
    wire new_AGEMA_signal_3767 ;
    wire new_AGEMA_signal_3768 ;
    wire new_AGEMA_signal_3769 ;
    wire new_AGEMA_signal_3770 ;
    wire new_AGEMA_signal_3771 ;
    wire new_AGEMA_signal_3772 ;
    wire new_AGEMA_signal_3773 ;
    wire new_AGEMA_signal_3774 ;
    wire new_AGEMA_signal_3775 ;
    wire new_AGEMA_signal_3776 ;
    wire new_AGEMA_signal_3777 ;
    wire new_AGEMA_signal_3778 ;
    wire new_AGEMA_signal_3779 ;
    wire new_AGEMA_signal_3780 ;
    wire new_AGEMA_signal_3781 ;
    wire new_AGEMA_signal_3782 ;
    wire new_AGEMA_signal_3783 ;
    wire new_AGEMA_signal_3784 ;
    wire new_AGEMA_signal_3785 ;
    wire new_AGEMA_signal_3786 ;
    wire new_AGEMA_signal_3787 ;
    wire new_AGEMA_signal_3788 ;
    wire new_AGEMA_signal_3789 ;
    wire new_AGEMA_signal_3790 ;
    wire new_AGEMA_signal_3791 ;
    wire new_AGEMA_signal_3792 ;
    wire new_AGEMA_signal_3793 ;
    wire new_AGEMA_signal_3794 ;
    wire new_AGEMA_signal_3795 ;
    wire new_AGEMA_signal_3796 ;
    wire new_AGEMA_signal_3797 ;
    wire new_AGEMA_signal_3798 ;
    wire new_AGEMA_signal_3799 ;
    wire new_AGEMA_signal_3800 ;
    wire new_AGEMA_signal_3801 ;
    wire new_AGEMA_signal_3802 ;
    wire new_AGEMA_signal_3803 ;
    wire new_AGEMA_signal_3804 ;
    wire new_AGEMA_signal_3805 ;
    wire new_AGEMA_signal_3806 ;
    wire new_AGEMA_signal_3807 ;
    wire new_AGEMA_signal_3808 ;
    wire new_AGEMA_signal_3809 ;
    wire new_AGEMA_signal_3810 ;
    wire new_AGEMA_signal_3811 ;
    wire new_AGEMA_signal_3812 ;
    wire new_AGEMA_signal_3813 ;
    wire new_AGEMA_signal_3814 ;
    wire new_AGEMA_signal_3815 ;
    wire new_AGEMA_signal_3816 ;
    wire new_AGEMA_signal_3817 ;
    wire new_AGEMA_signal_3818 ;
    wire new_AGEMA_signal_3819 ;
    wire new_AGEMA_signal_3820 ;
    wire new_AGEMA_signal_3821 ;
    wire new_AGEMA_signal_3822 ;
    wire new_AGEMA_signal_3823 ;
    wire new_AGEMA_signal_3824 ;
    wire new_AGEMA_signal_3825 ;
    wire new_AGEMA_signal_3826 ;
    wire new_AGEMA_signal_3827 ;
    wire new_AGEMA_signal_3828 ;
    wire new_AGEMA_signal_3829 ;
    wire new_AGEMA_signal_3830 ;
    wire new_AGEMA_signal_3831 ;
    wire new_AGEMA_signal_3832 ;
    wire new_AGEMA_signal_3833 ;
    wire new_AGEMA_signal_3834 ;
    wire new_AGEMA_signal_3835 ;
    wire new_AGEMA_signal_3836 ;
    wire new_AGEMA_signal_3837 ;
    wire new_AGEMA_signal_3838 ;
    wire new_AGEMA_signal_3839 ;
    wire new_AGEMA_signal_3840 ;
    wire new_AGEMA_signal_3841 ;
    wire new_AGEMA_signal_3842 ;
    wire new_AGEMA_signal_3843 ;
    wire new_AGEMA_signal_3844 ;
    wire new_AGEMA_signal_3845 ;
    wire new_AGEMA_signal_3846 ;
    wire new_AGEMA_signal_3847 ;
    wire new_AGEMA_signal_3848 ;
    wire new_AGEMA_signal_3849 ;
    wire new_AGEMA_signal_3850 ;
    wire new_AGEMA_signal_3851 ;
    wire new_AGEMA_signal_3852 ;
    wire new_AGEMA_signal_3853 ;
    wire new_AGEMA_signal_3854 ;
    wire new_AGEMA_signal_3855 ;
    wire new_AGEMA_signal_3856 ;
    wire new_AGEMA_signal_3857 ;
    wire new_AGEMA_signal_3858 ;
    wire new_AGEMA_signal_3859 ;
    wire new_AGEMA_signal_3860 ;
    wire new_AGEMA_signal_3861 ;
    wire new_AGEMA_signal_3862 ;
    wire new_AGEMA_signal_3863 ;
    wire new_AGEMA_signal_3864 ;
    wire new_AGEMA_signal_3865 ;
    wire new_AGEMA_signal_3866 ;
    wire new_AGEMA_signal_3867 ;
    wire new_AGEMA_signal_3868 ;
    wire new_AGEMA_signal_3869 ;
    wire new_AGEMA_signal_3870 ;
    wire new_AGEMA_signal_3871 ;
    wire new_AGEMA_signal_3872 ;
    wire new_AGEMA_signal_3873 ;
    wire new_AGEMA_signal_3874 ;
    wire new_AGEMA_signal_3875 ;
    wire new_AGEMA_signal_3876 ;
    wire new_AGEMA_signal_3877 ;
    wire new_AGEMA_signal_3878 ;
    wire new_AGEMA_signal_3879 ;
    wire new_AGEMA_signal_3880 ;
    wire new_AGEMA_signal_3881 ;
    wire new_AGEMA_signal_3882 ;
    wire new_AGEMA_signal_3883 ;
    wire new_AGEMA_signal_3884 ;
    wire new_AGEMA_signal_3885 ;
    wire new_AGEMA_signal_3886 ;
    wire new_AGEMA_signal_3887 ;
    wire new_AGEMA_signal_3888 ;
    wire new_AGEMA_signal_3889 ;
    wire new_AGEMA_signal_3890 ;
    wire new_AGEMA_signal_3891 ;
    wire new_AGEMA_signal_3892 ;
    wire new_AGEMA_signal_3893 ;
    wire new_AGEMA_signal_3894 ;
    wire new_AGEMA_signal_3895 ;
    wire new_AGEMA_signal_3896 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3898 ;
    wire new_AGEMA_signal_3899 ;
    wire new_AGEMA_signal_3900 ;
    wire new_AGEMA_signal_3901 ;
    wire new_AGEMA_signal_3902 ;
    wire new_AGEMA_signal_3903 ;
    wire new_AGEMA_signal_3904 ;
    wire new_AGEMA_signal_3905 ;
    wire new_AGEMA_signal_3906 ;
    wire new_AGEMA_signal_3907 ;
    wire new_AGEMA_signal_3908 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3910 ;
    wire new_AGEMA_signal_3911 ;
    wire new_AGEMA_signal_3912 ;
    wire new_AGEMA_signal_3913 ;
    wire new_AGEMA_signal_3914 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3916 ;
    wire new_AGEMA_signal_3917 ;
    wire new_AGEMA_signal_3918 ;
    wire new_AGEMA_signal_3919 ;
    wire new_AGEMA_signal_3920 ;
    wire new_AGEMA_signal_3921 ;
    wire new_AGEMA_signal_3922 ;
    wire new_AGEMA_signal_3923 ;
    wire new_AGEMA_signal_3924 ;
    wire new_AGEMA_signal_3925 ;
    wire new_AGEMA_signal_3926 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3928 ;
    wire new_AGEMA_signal_3929 ;
    wire new_AGEMA_signal_3930 ;
    wire new_AGEMA_signal_3931 ;
    wire new_AGEMA_signal_3932 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3934 ;
    wire new_AGEMA_signal_3935 ;
    wire new_AGEMA_signal_3936 ;
    wire new_AGEMA_signal_3937 ;
    wire new_AGEMA_signal_3938 ;
    wire new_AGEMA_signal_3939 ;
    wire new_AGEMA_signal_3940 ;
    wire new_AGEMA_signal_3941 ;
    wire new_AGEMA_signal_3942 ;
    wire new_AGEMA_signal_3943 ;
    wire new_AGEMA_signal_3944 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3946 ;
    wire new_AGEMA_signal_3947 ;
    wire new_AGEMA_signal_3948 ;
    wire new_AGEMA_signal_3949 ;
    wire new_AGEMA_signal_3950 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_3952 ;
    wire new_AGEMA_signal_3953 ;
    wire new_AGEMA_signal_3954 ;
    wire new_AGEMA_signal_3955 ;
    wire new_AGEMA_signal_3956 ;
    wire new_AGEMA_signal_3957 ;
    wire new_AGEMA_signal_3958 ;
    wire new_AGEMA_signal_3959 ;
    wire new_AGEMA_signal_3960 ;
    wire new_AGEMA_signal_3961 ;
    wire new_AGEMA_signal_3962 ;
    wire new_AGEMA_signal_3963 ;
    wire new_AGEMA_signal_3964 ;
    wire new_AGEMA_signal_3965 ;
    wire new_AGEMA_signal_3966 ;
    wire new_AGEMA_signal_3967 ;
    wire new_AGEMA_signal_3968 ;
    wire new_AGEMA_signal_3969 ;
    wire new_AGEMA_signal_3970 ;
    wire new_AGEMA_signal_3971 ;
    wire new_AGEMA_signal_3972 ;
    wire new_AGEMA_signal_3973 ;
    wire new_AGEMA_signal_3974 ;
    wire new_AGEMA_signal_3975 ;
    wire new_AGEMA_signal_3976 ;
    wire new_AGEMA_signal_3977 ;
    wire new_AGEMA_signal_3978 ;
    wire new_AGEMA_signal_3979 ;
    wire new_AGEMA_signal_3980 ;
    wire new_AGEMA_signal_3981 ;
    wire new_AGEMA_signal_3982 ;
    wire new_AGEMA_signal_3983 ;
    wire new_AGEMA_signal_3984 ;
    wire new_AGEMA_signal_3985 ;
    wire new_AGEMA_signal_3986 ;
    wire new_AGEMA_signal_3987 ;
    wire new_AGEMA_signal_3988 ;
    wire new_AGEMA_signal_3989 ;
    wire new_AGEMA_signal_3990 ;
    wire new_AGEMA_signal_3991 ;
    wire new_AGEMA_signal_3992 ;
    wire new_AGEMA_signal_3993 ;
    wire new_AGEMA_signal_3994 ;
    wire new_AGEMA_signal_3995 ;
    wire new_AGEMA_signal_3996 ;
    wire new_AGEMA_signal_3997 ;
    wire new_AGEMA_signal_3998 ;
    wire new_AGEMA_signal_3999 ;
    wire new_AGEMA_signal_4000 ;
    wire new_AGEMA_signal_4001 ;
    wire new_AGEMA_signal_4002 ;
    wire new_AGEMA_signal_4003 ;
    wire new_AGEMA_signal_4004 ;
    wire new_AGEMA_signal_4005 ;
    wire new_AGEMA_signal_4006 ;
    wire new_AGEMA_signal_4007 ;
    wire new_AGEMA_signal_4008 ;
    wire new_AGEMA_signal_4009 ;
    wire new_AGEMA_signal_4010 ;
    wire new_AGEMA_signal_4011 ;
    wire new_AGEMA_signal_4012 ;
    wire new_AGEMA_signal_4013 ;
    wire new_AGEMA_signal_4014 ;
    wire new_AGEMA_signal_4015 ;
    wire new_AGEMA_signal_4016 ;
    wire new_AGEMA_signal_4017 ;
    wire new_AGEMA_signal_4018 ;
    wire new_AGEMA_signal_4019 ;
    wire new_AGEMA_signal_4020 ;
    wire new_AGEMA_signal_4021 ;
    wire new_AGEMA_signal_4022 ;
    wire new_AGEMA_signal_4023 ;
    wire new_AGEMA_signal_4024 ;
    wire new_AGEMA_signal_4025 ;
    wire new_AGEMA_signal_4026 ;
    wire new_AGEMA_signal_4027 ;
    wire new_AGEMA_signal_4028 ;
    wire new_AGEMA_signal_4029 ;
    wire new_AGEMA_signal_4030 ;
    wire new_AGEMA_signal_4031 ;
    wire new_AGEMA_signal_4032 ;
    wire new_AGEMA_signal_4033 ;
    wire new_AGEMA_signal_4034 ;
    wire new_AGEMA_signal_4035 ;
    wire new_AGEMA_signal_4036 ;
    wire new_AGEMA_signal_4037 ;
    wire new_AGEMA_signal_4038 ;
    wire new_AGEMA_signal_4039 ;
    wire new_AGEMA_signal_4040 ;
    wire new_AGEMA_signal_4041 ;
    wire new_AGEMA_signal_4042 ;
    wire new_AGEMA_signal_4043 ;
    wire new_AGEMA_signal_4044 ;
    wire new_AGEMA_signal_4045 ;
    wire new_AGEMA_signal_4046 ;
    wire new_AGEMA_signal_4047 ;
    wire new_AGEMA_signal_4048 ;
    wire new_AGEMA_signal_4049 ;
    wire new_AGEMA_signal_4050 ;
    wire new_AGEMA_signal_4051 ;
    wire new_AGEMA_signal_4052 ;
    wire new_AGEMA_signal_4053 ;
    wire new_AGEMA_signal_4054 ;
    wire new_AGEMA_signal_4055 ;
    wire new_AGEMA_signal_4056 ;
    wire new_AGEMA_signal_4057 ;
    wire new_AGEMA_signal_4058 ;
    wire new_AGEMA_signal_4059 ;
    wire new_AGEMA_signal_4060 ;
    wire new_AGEMA_signal_4061 ;
    wire new_AGEMA_signal_4062 ;
    wire new_AGEMA_signal_4063 ;
    wire new_AGEMA_signal_4064 ;
    wire new_AGEMA_signal_4065 ;
    wire new_AGEMA_signal_4066 ;
    wire new_AGEMA_signal_4067 ;
    wire new_AGEMA_signal_4068 ;
    wire new_AGEMA_signal_4069 ;
    wire new_AGEMA_signal_4070 ;
    wire new_AGEMA_signal_4071 ;
    wire new_AGEMA_signal_4072 ;
    wire new_AGEMA_signal_4073 ;
    wire new_AGEMA_signal_4074 ;
    wire new_AGEMA_signal_4075 ;
    wire new_AGEMA_signal_4076 ;
    wire new_AGEMA_signal_4077 ;
    wire new_AGEMA_signal_4078 ;
    wire new_AGEMA_signal_4079 ;
    wire new_AGEMA_signal_4080 ;
    wire new_AGEMA_signal_4081 ;
    wire new_AGEMA_signal_4082 ;
    wire new_AGEMA_signal_4083 ;
    wire new_AGEMA_signal_4084 ;
    wire new_AGEMA_signal_4085 ;
    wire new_AGEMA_signal_4086 ;
    wire new_AGEMA_signal_4087 ;
    wire new_AGEMA_signal_4088 ;
    wire new_AGEMA_signal_4089 ;
    wire new_AGEMA_signal_4090 ;
    wire new_AGEMA_signal_4091 ;
    wire new_AGEMA_signal_4092 ;
    wire new_AGEMA_signal_4093 ;
    wire new_AGEMA_signal_4094 ;
    wire new_AGEMA_signal_4095 ;
    wire new_AGEMA_signal_4096 ;
    wire new_AGEMA_signal_4097 ;
    wire new_AGEMA_signal_4098 ;
    wire new_AGEMA_signal_4099 ;
    wire new_AGEMA_signal_4100 ;
    wire new_AGEMA_signal_4101 ;
    wire new_AGEMA_signal_4102 ;
    wire new_AGEMA_signal_4103 ;
    wire new_AGEMA_signal_4104 ;
    wire new_AGEMA_signal_4105 ;
    wire new_AGEMA_signal_4106 ;
    wire new_AGEMA_signal_4107 ;
    wire new_AGEMA_signal_4108 ;
    wire new_AGEMA_signal_4109 ;
    wire new_AGEMA_signal_4110 ;
    wire new_AGEMA_signal_4111 ;
    wire new_AGEMA_signal_4112 ;
    wire new_AGEMA_signal_4113 ;
    wire new_AGEMA_signal_4114 ;
    wire new_AGEMA_signal_4115 ;
    wire new_AGEMA_signal_4116 ;
    wire new_AGEMA_signal_4117 ;
    wire new_AGEMA_signal_4118 ;
    wire new_AGEMA_signal_4119 ;
    wire new_AGEMA_signal_4120 ;
    wire new_AGEMA_signal_4121 ;
    wire new_AGEMA_signal_4122 ;
    wire new_AGEMA_signal_4123 ;
    wire new_AGEMA_signal_4124 ;
    wire new_AGEMA_signal_4125 ;
    wire new_AGEMA_signal_4126 ;
    wire new_AGEMA_signal_4127 ;
    wire new_AGEMA_signal_4128 ;
    wire new_AGEMA_signal_4129 ;
    wire new_AGEMA_signal_4130 ;
    wire new_AGEMA_signal_4131 ;
    wire new_AGEMA_signal_4132 ;
    wire new_AGEMA_signal_4133 ;
    wire new_AGEMA_signal_4134 ;
    wire new_AGEMA_signal_4135 ;
    wire new_AGEMA_signal_4136 ;
    wire new_AGEMA_signal_4137 ;
    wire new_AGEMA_signal_4138 ;
    wire new_AGEMA_signal_4139 ;
    wire new_AGEMA_signal_4140 ;
    wire new_AGEMA_signal_4141 ;
    wire new_AGEMA_signal_4142 ;
    wire new_AGEMA_signal_4143 ;
    wire new_AGEMA_signal_4144 ;
    wire new_AGEMA_signal_4145 ;
    wire new_AGEMA_signal_4146 ;
    wire new_AGEMA_signal_4147 ;
    wire new_AGEMA_signal_4148 ;
    wire new_AGEMA_signal_4149 ;
    wire new_AGEMA_signal_4150 ;
    wire new_AGEMA_signal_4151 ;
    wire new_AGEMA_signal_4152 ;
    wire new_AGEMA_signal_4153 ;
    wire new_AGEMA_signal_4154 ;
    wire new_AGEMA_signal_4155 ;
    wire new_AGEMA_signal_4156 ;
    wire new_AGEMA_signal_4157 ;
    wire new_AGEMA_signal_4158 ;
    wire new_AGEMA_signal_4159 ;
    wire new_AGEMA_signal_4160 ;
    wire new_AGEMA_signal_4161 ;
    wire new_AGEMA_signal_4162 ;
    wire new_AGEMA_signal_4163 ;
    wire new_AGEMA_signal_4164 ;
    wire new_AGEMA_signal_4165 ;
    wire new_AGEMA_signal_4166 ;
    wire new_AGEMA_signal_4167 ;
    wire new_AGEMA_signal_4168 ;
    wire new_AGEMA_signal_4169 ;
    wire new_AGEMA_signal_4170 ;
    wire new_AGEMA_signal_4171 ;
    wire new_AGEMA_signal_4172 ;
    wire new_AGEMA_signal_4173 ;
    wire new_AGEMA_signal_4174 ;
    wire new_AGEMA_signal_4175 ;
    wire new_AGEMA_signal_4176 ;
    wire new_AGEMA_signal_4177 ;
    wire new_AGEMA_signal_4178 ;
    wire new_AGEMA_signal_4179 ;
    wire new_AGEMA_signal_4180 ;
    wire new_AGEMA_signal_4181 ;
    wire new_AGEMA_signal_4182 ;
    wire new_AGEMA_signal_4183 ;
    wire new_AGEMA_signal_4184 ;
    wire new_AGEMA_signal_4185 ;
    wire new_AGEMA_signal_4186 ;
    wire new_AGEMA_signal_4187 ;
    wire new_AGEMA_signal_4188 ;
    wire new_AGEMA_signal_4189 ;
    wire new_AGEMA_signal_4190 ;
    wire new_AGEMA_signal_4191 ;
    wire new_AGEMA_signal_4192 ;
    wire new_AGEMA_signal_4193 ;
    wire new_AGEMA_signal_4194 ;
    wire new_AGEMA_signal_4195 ;
    wire new_AGEMA_signal_4196 ;
    wire new_AGEMA_signal_4197 ;
    wire new_AGEMA_signal_4198 ;
    wire new_AGEMA_signal_4199 ;
    wire new_AGEMA_signal_4200 ;
    wire new_AGEMA_signal_4201 ;
    wire new_AGEMA_signal_4202 ;
    wire new_AGEMA_signal_4203 ;
    wire new_AGEMA_signal_4204 ;
    wire new_AGEMA_signal_4205 ;
    wire new_AGEMA_signal_4206 ;
    wire new_AGEMA_signal_4207 ;
    wire new_AGEMA_signal_4208 ;
    wire new_AGEMA_signal_4209 ;
    wire new_AGEMA_signal_4210 ;
    wire new_AGEMA_signal_4211 ;
    wire new_AGEMA_signal_4212 ;
    wire new_AGEMA_signal_4213 ;
    wire new_AGEMA_signal_4214 ;
    wire new_AGEMA_signal_4215 ;
    wire new_AGEMA_signal_4216 ;
    wire new_AGEMA_signal_4217 ;
    wire new_AGEMA_signal_4218 ;
    wire new_AGEMA_signal_4219 ;
    wire new_AGEMA_signal_4220 ;
    wire new_AGEMA_signal_4221 ;
    wire new_AGEMA_signal_4222 ;
    wire new_AGEMA_signal_4223 ;
    wire new_AGEMA_signal_4224 ;
    wire new_AGEMA_signal_4225 ;
    wire new_AGEMA_signal_4226 ;
    wire new_AGEMA_signal_4227 ;
    wire new_AGEMA_signal_4228 ;
    wire new_AGEMA_signal_4229 ;
    wire new_AGEMA_signal_4230 ;
    wire new_AGEMA_signal_4231 ;
    wire new_AGEMA_signal_4232 ;
    wire new_AGEMA_signal_4233 ;
    wire new_AGEMA_signal_4234 ;
    wire new_AGEMA_signal_4235 ;
    wire new_AGEMA_signal_4236 ;
    wire new_AGEMA_signal_4237 ;
    wire new_AGEMA_signal_4238 ;
    wire new_AGEMA_signal_4239 ;
    wire new_AGEMA_signal_4240 ;
    wire new_AGEMA_signal_4241 ;
    wire new_AGEMA_signal_4242 ;
    wire new_AGEMA_signal_4243 ;
    wire new_AGEMA_signal_4244 ;
    wire new_AGEMA_signal_4245 ;
    wire new_AGEMA_signal_4246 ;
    wire new_AGEMA_signal_4247 ;
    wire new_AGEMA_signal_4248 ;
    wire new_AGEMA_signal_4249 ;
    wire new_AGEMA_signal_4250 ;
    wire new_AGEMA_signal_4251 ;
    wire new_AGEMA_signal_4252 ;
    wire new_AGEMA_signal_4253 ;
    wire new_AGEMA_signal_4254 ;
    wire new_AGEMA_signal_4255 ;
    wire new_AGEMA_signal_4256 ;
    wire new_AGEMA_signal_4257 ;
    wire new_AGEMA_signal_4258 ;
    wire new_AGEMA_signal_4259 ;
    wire new_AGEMA_signal_4260 ;
    wire new_AGEMA_signal_4261 ;
    wire new_AGEMA_signal_4262 ;
    wire new_AGEMA_signal_4263 ;
    wire new_AGEMA_signal_4264 ;
    wire new_AGEMA_signal_4265 ;
    wire new_AGEMA_signal_4266 ;
    wire new_AGEMA_signal_4267 ;
    wire new_AGEMA_signal_4268 ;
    wire new_AGEMA_signal_4269 ;
    wire new_AGEMA_signal_4270 ;
    wire new_AGEMA_signal_4271 ;
    wire new_AGEMA_signal_4272 ;
    wire new_AGEMA_signal_4273 ;
    wire new_AGEMA_signal_4274 ;
    wire new_AGEMA_signal_4275 ;
    wire new_AGEMA_signal_4276 ;
    wire new_AGEMA_signal_4277 ;
    wire new_AGEMA_signal_4278 ;
    wire new_AGEMA_signal_4279 ;
    wire new_AGEMA_signal_4280 ;
    wire new_AGEMA_signal_4281 ;
    wire new_AGEMA_signal_4282 ;
    wire new_AGEMA_signal_4283 ;
    wire new_AGEMA_signal_4284 ;
    wire new_AGEMA_signal_4285 ;
    wire new_AGEMA_signal_4286 ;
    wire new_AGEMA_signal_4287 ;
    wire new_AGEMA_signal_4288 ;
    wire new_AGEMA_signal_4289 ;
    wire new_AGEMA_signal_4290 ;
    wire new_AGEMA_signal_4291 ;
    wire new_AGEMA_signal_4292 ;
    wire new_AGEMA_signal_4293 ;
    wire new_AGEMA_signal_4294 ;
    wire new_AGEMA_signal_4295 ;
    wire new_AGEMA_signal_4296 ;
    wire new_AGEMA_signal_4297 ;
    wire new_AGEMA_signal_4298 ;
    wire new_AGEMA_signal_4299 ;
    wire new_AGEMA_signal_4300 ;
    wire new_AGEMA_signal_4301 ;
    wire new_AGEMA_signal_4302 ;
    wire new_AGEMA_signal_4303 ;
    wire new_AGEMA_signal_4304 ;
    wire new_AGEMA_signal_4305 ;
    wire new_AGEMA_signal_4306 ;
    wire new_AGEMA_signal_4307 ;
    wire new_AGEMA_signal_4308 ;
    wire new_AGEMA_signal_4309 ;
    wire new_AGEMA_signal_4310 ;
    wire new_AGEMA_signal_4311 ;
    wire new_AGEMA_signal_4312 ;
    wire new_AGEMA_signal_4313 ;
    wire new_AGEMA_signal_4314 ;
    wire new_AGEMA_signal_4315 ;
    wire new_AGEMA_signal_4316 ;
    wire new_AGEMA_signal_4317 ;
    wire new_AGEMA_signal_4318 ;
    wire new_AGEMA_signal_4319 ;
    wire new_AGEMA_signal_4320 ;
    wire new_AGEMA_signal_4321 ;
    wire new_AGEMA_signal_4322 ;
    wire new_AGEMA_signal_4323 ;
    wire new_AGEMA_signal_4324 ;
    wire new_AGEMA_signal_4325 ;
    wire new_AGEMA_signal_4326 ;
    wire new_AGEMA_signal_4327 ;
    wire new_AGEMA_signal_4328 ;
    wire new_AGEMA_signal_4329 ;
    wire new_AGEMA_signal_4330 ;
    wire new_AGEMA_signal_4331 ;
    wire new_AGEMA_signal_4332 ;
    wire new_AGEMA_signal_4333 ;
    wire new_AGEMA_signal_4334 ;
    wire new_AGEMA_signal_4335 ;
    wire new_AGEMA_signal_4336 ;
    wire new_AGEMA_signal_4337 ;
    wire new_AGEMA_signal_4338 ;
    wire new_AGEMA_signal_4339 ;
    wire new_AGEMA_signal_4340 ;
    wire new_AGEMA_signal_4341 ;
    wire new_AGEMA_signal_4342 ;
    wire new_AGEMA_signal_4343 ;
    wire new_AGEMA_signal_4344 ;
    wire new_AGEMA_signal_4345 ;
    wire new_AGEMA_signal_4346 ;
    wire new_AGEMA_signal_4347 ;
    wire new_AGEMA_signal_4348 ;
    wire new_AGEMA_signal_4349 ;
    wire new_AGEMA_signal_4350 ;
    wire new_AGEMA_signal_4351 ;
    wire new_AGEMA_signal_4352 ;
    wire new_AGEMA_signal_4353 ;
    wire new_AGEMA_signal_4354 ;
    wire new_AGEMA_signal_4355 ;
    wire new_AGEMA_signal_4356 ;
    wire new_AGEMA_signal_4357 ;
    wire new_AGEMA_signal_4358 ;
    wire new_AGEMA_signal_4359 ;
    wire new_AGEMA_signal_4360 ;
    wire new_AGEMA_signal_4361 ;
    wire new_AGEMA_signal_4362 ;
    wire new_AGEMA_signal_4363 ;
    wire new_AGEMA_signal_4364 ;
    wire new_AGEMA_signal_4365 ;
    wire new_AGEMA_signal_4366 ;
    wire new_AGEMA_signal_4367 ;
    wire new_AGEMA_signal_4368 ;
    wire new_AGEMA_signal_4369 ;
    wire new_AGEMA_signal_4370 ;
    wire new_AGEMA_signal_4371 ;
    wire new_AGEMA_signal_4372 ;
    wire new_AGEMA_signal_4373 ;
    wire new_AGEMA_signal_4374 ;
    wire new_AGEMA_signal_4375 ;
    wire new_AGEMA_signal_4376 ;
    wire new_AGEMA_signal_4377 ;
    wire new_AGEMA_signal_4378 ;
    wire new_AGEMA_signal_4379 ;
    wire new_AGEMA_signal_4380 ;
    wire new_AGEMA_signal_4381 ;
    wire new_AGEMA_signal_4382 ;
    wire new_AGEMA_signal_4383 ;
    wire new_AGEMA_signal_4384 ;
    wire new_AGEMA_signal_4385 ;
    wire new_AGEMA_signal_4386 ;
    wire new_AGEMA_signal_4387 ;
    wire new_AGEMA_signal_4388 ;
    wire new_AGEMA_signal_4389 ;
    wire new_AGEMA_signal_4390 ;
    wire new_AGEMA_signal_4391 ;
    wire new_AGEMA_signal_4392 ;
    wire new_AGEMA_signal_4393 ;
    wire new_AGEMA_signal_4394 ;
    wire new_AGEMA_signal_4395 ;
    wire new_AGEMA_signal_4396 ;
    wire new_AGEMA_signal_4397 ;
    wire new_AGEMA_signal_4398 ;
    wire new_AGEMA_signal_4399 ;
    wire new_AGEMA_signal_4400 ;
    wire new_AGEMA_signal_4401 ;
    wire new_AGEMA_signal_4402 ;
    wire new_AGEMA_signal_4403 ;
    wire new_AGEMA_signal_4404 ;
    wire new_AGEMA_signal_4405 ;
    wire new_AGEMA_signal_4406 ;
    wire new_AGEMA_signal_4407 ;
    wire new_AGEMA_signal_4408 ;
    wire new_AGEMA_signal_4409 ;
    wire new_AGEMA_signal_4410 ;
    wire new_AGEMA_signal_4411 ;
    wire new_AGEMA_signal_4412 ;
    wire new_AGEMA_signal_4413 ;
    wire new_AGEMA_signal_4414 ;
    wire new_AGEMA_signal_4415 ;
    wire new_AGEMA_signal_4416 ;
    wire new_AGEMA_signal_4417 ;
    wire new_AGEMA_signal_4418 ;
    wire new_AGEMA_signal_4419 ;
    wire new_AGEMA_signal_4420 ;
    wire new_AGEMA_signal_4421 ;
    wire new_AGEMA_signal_4422 ;
    wire new_AGEMA_signal_4423 ;
    wire new_AGEMA_signal_4424 ;
    wire new_AGEMA_signal_4425 ;
    wire new_AGEMA_signal_4426 ;
    wire new_AGEMA_signal_4427 ;
    wire new_AGEMA_signal_4428 ;
    wire new_AGEMA_signal_4429 ;
    wire new_AGEMA_signal_4430 ;
    wire new_AGEMA_signal_4431 ;
    wire new_AGEMA_signal_4432 ;
    wire new_AGEMA_signal_4433 ;
    wire new_AGEMA_signal_4434 ;
    wire new_AGEMA_signal_4435 ;
    wire new_AGEMA_signal_4436 ;
    wire new_AGEMA_signal_4437 ;
    wire new_AGEMA_signal_4438 ;
    wire new_AGEMA_signal_4439 ;
    wire new_AGEMA_signal_4440 ;
    wire new_AGEMA_signal_4441 ;
    wire new_AGEMA_signal_4442 ;
    wire new_AGEMA_signal_4443 ;
    wire new_AGEMA_signal_4444 ;
    wire new_AGEMA_signal_4445 ;
    wire new_AGEMA_signal_4446 ;
    wire new_AGEMA_signal_4447 ;
    wire new_AGEMA_signal_4448 ;
    wire new_AGEMA_signal_4449 ;
    wire new_AGEMA_signal_4450 ;
    wire new_AGEMA_signal_4451 ;
    wire new_AGEMA_signal_4452 ;
    wire new_AGEMA_signal_4453 ;
    wire new_AGEMA_signal_4454 ;
    wire new_AGEMA_signal_4455 ;
    wire new_AGEMA_signal_4456 ;
    wire new_AGEMA_signal_4457 ;
    wire new_AGEMA_signal_4458 ;
    wire new_AGEMA_signal_4459 ;
    wire new_AGEMA_signal_4460 ;
    wire new_AGEMA_signal_4461 ;
    wire new_AGEMA_signal_4462 ;
    wire new_AGEMA_signal_4463 ;
    wire new_AGEMA_signal_4464 ;
    wire new_AGEMA_signal_4465 ;
    wire new_AGEMA_signal_4466 ;
    wire new_AGEMA_signal_4467 ;
    wire new_AGEMA_signal_4468 ;
    wire new_AGEMA_signal_4469 ;
    wire new_AGEMA_signal_4470 ;
    wire new_AGEMA_signal_4471 ;
    wire new_AGEMA_signal_4472 ;
    wire new_AGEMA_signal_4473 ;
    wire new_AGEMA_signal_4474 ;
    wire new_AGEMA_signal_4475 ;
    wire new_AGEMA_signal_4476 ;
    wire new_AGEMA_signal_4477 ;
    wire new_AGEMA_signal_4478 ;
    wire new_AGEMA_signal_4479 ;
    wire new_AGEMA_signal_4480 ;
    wire new_AGEMA_signal_4481 ;
    wire new_AGEMA_signal_4482 ;
    wire new_AGEMA_signal_4483 ;
    wire new_AGEMA_signal_4484 ;
    wire new_AGEMA_signal_4485 ;
    wire new_AGEMA_signal_4486 ;
    wire new_AGEMA_signal_4487 ;
    wire new_AGEMA_signal_4488 ;
    wire new_AGEMA_signal_4489 ;
    wire new_AGEMA_signal_4490 ;
    wire new_AGEMA_signal_4491 ;
    wire new_AGEMA_signal_4492 ;
    wire new_AGEMA_signal_4493 ;
    wire new_AGEMA_signal_4494 ;
    wire new_AGEMA_signal_4495 ;
    wire new_AGEMA_signal_4496 ;
    wire new_AGEMA_signal_4497 ;
    wire new_AGEMA_signal_4498 ;
    wire new_AGEMA_signal_4499 ;
    wire new_AGEMA_signal_4500 ;
    wire new_AGEMA_signal_4501 ;
    wire new_AGEMA_signal_4502 ;
    wire new_AGEMA_signal_4503 ;
    wire new_AGEMA_signal_4504 ;
    wire new_AGEMA_signal_4505 ;
    wire new_AGEMA_signal_4506 ;
    wire new_AGEMA_signal_4507 ;
    wire new_AGEMA_signal_4508 ;
    wire new_AGEMA_signal_4509 ;
    wire new_AGEMA_signal_4510 ;
    wire new_AGEMA_signal_4511 ;
    wire new_AGEMA_signal_4512 ;
    wire new_AGEMA_signal_4513 ;
    wire new_AGEMA_signal_4514 ;
    wire new_AGEMA_signal_4515 ;
    wire new_AGEMA_signal_4516 ;
    wire new_AGEMA_signal_4517 ;
    wire new_AGEMA_signal_4518 ;
    wire new_AGEMA_signal_4519 ;
    wire new_AGEMA_signal_4520 ;
    wire new_AGEMA_signal_4521 ;
    wire new_AGEMA_signal_4522 ;
    wire new_AGEMA_signal_4523 ;
    wire new_AGEMA_signal_4524 ;
    wire new_AGEMA_signal_4525 ;
    wire new_AGEMA_signal_4526 ;
    wire new_AGEMA_signal_4527 ;
    wire new_AGEMA_signal_4528 ;
    wire new_AGEMA_signal_4529 ;
    wire new_AGEMA_signal_4530 ;
    wire new_AGEMA_signal_4531 ;
    wire new_AGEMA_signal_4532 ;
    wire new_AGEMA_signal_4533 ;
    wire new_AGEMA_signal_4534 ;
    wire new_AGEMA_signal_4535 ;
    wire new_AGEMA_signal_4536 ;
    wire new_AGEMA_signal_4537 ;
    wire new_AGEMA_signal_4538 ;
    wire new_AGEMA_signal_4539 ;
    wire new_AGEMA_signal_4540 ;
    wire new_AGEMA_signal_4541 ;
    wire new_AGEMA_signal_4542 ;
    wire new_AGEMA_signal_4543 ;
    wire new_AGEMA_signal_4544 ;
    wire new_AGEMA_signal_4545 ;
    wire new_AGEMA_signal_4546 ;
    wire new_AGEMA_signal_4547 ;
    wire new_AGEMA_signal_4548 ;
    wire new_AGEMA_signal_4549 ;
    wire new_AGEMA_signal_4550 ;
    wire new_AGEMA_signal_4551 ;
    wire new_AGEMA_signal_4552 ;
    wire new_AGEMA_signal_4553 ;
    wire new_AGEMA_signal_4554 ;
    wire new_AGEMA_signal_4555 ;
    wire new_AGEMA_signal_4556 ;
    wire new_AGEMA_signal_4557 ;
    wire new_AGEMA_signal_4558 ;
    wire new_AGEMA_signal_4559 ;
    wire new_AGEMA_signal_4560 ;
    wire new_AGEMA_signal_4561 ;
    wire new_AGEMA_signal_4562 ;
    wire new_AGEMA_signal_4563 ;
    wire new_AGEMA_signal_4564 ;
    wire new_AGEMA_signal_4565 ;
    wire new_AGEMA_signal_4566 ;
    wire new_AGEMA_signal_4567 ;
    wire new_AGEMA_signal_4568 ;
    wire new_AGEMA_signal_4569 ;
    wire new_AGEMA_signal_4570 ;
    wire new_AGEMA_signal_4571 ;
    wire new_AGEMA_signal_4572 ;
    wire new_AGEMA_signal_4573 ;
    wire new_AGEMA_signal_4574 ;
    wire new_AGEMA_signal_4575 ;
    wire new_AGEMA_signal_4576 ;
    wire new_AGEMA_signal_4577 ;
    wire new_AGEMA_signal_4578 ;
    wire new_AGEMA_signal_4579 ;
    wire new_AGEMA_signal_4580 ;
    wire new_AGEMA_signal_4581 ;
    wire new_AGEMA_signal_4582 ;
    wire new_AGEMA_signal_4583 ;
    wire new_AGEMA_signal_4584 ;
    wire new_AGEMA_signal_4585 ;
    wire new_AGEMA_signal_4586 ;
    wire new_AGEMA_signal_4587 ;
    wire new_AGEMA_signal_4588 ;
    wire new_AGEMA_signal_4589 ;
    wire new_AGEMA_signal_4590 ;
    wire new_AGEMA_signal_4591 ;
    wire new_AGEMA_signal_4592 ;
    wire new_AGEMA_signal_4593 ;
    wire new_AGEMA_signal_4594 ;
    wire new_AGEMA_signal_4595 ;
    wire new_AGEMA_signal_4596 ;
    wire new_AGEMA_signal_4597 ;
    wire new_AGEMA_signal_4598 ;
    wire new_AGEMA_signal_4599 ;
    wire new_AGEMA_signal_4600 ;
    wire new_AGEMA_signal_4601 ;
    wire new_AGEMA_signal_4602 ;
    wire new_AGEMA_signal_4603 ;
    wire new_AGEMA_signal_4604 ;
    wire new_AGEMA_signal_4605 ;
    wire new_AGEMA_signal_4606 ;
    wire new_AGEMA_signal_4607 ;
    wire new_AGEMA_signal_4608 ;
    wire new_AGEMA_signal_4609 ;
    wire new_AGEMA_signal_4610 ;
    wire new_AGEMA_signal_4611 ;
    wire new_AGEMA_signal_4612 ;
    wire new_AGEMA_signal_4613 ;
    wire new_AGEMA_signal_4614 ;
    wire new_AGEMA_signal_4615 ;
    wire new_AGEMA_signal_4616 ;
    wire new_AGEMA_signal_4617 ;
    wire new_AGEMA_signal_4618 ;
    wire new_AGEMA_signal_4619 ;
    wire new_AGEMA_signal_4620 ;
    wire new_AGEMA_signal_4621 ;
    wire new_AGEMA_signal_4622 ;
    wire new_AGEMA_signal_4623 ;
    wire new_AGEMA_signal_4624 ;
    wire new_AGEMA_signal_4625 ;
    wire new_AGEMA_signal_4626 ;
    wire new_AGEMA_signal_4627 ;
    wire new_AGEMA_signal_4628 ;
    wire new_AGEMA_signal_4629 ;
    wire new_AGEMA_signal_4630 ;
    wire new_AGEMA_signal_4631 ;
    wire new_AGEMA_signal_4632 ;
    wire new_AGEMA_signal_4633 ;
    wire new_AGEMA_signal_4634 ;
    wire new_AGEMA_signal_4635 ;
    wire new_AGEMA_signal_4636 ;
    wire new_AGEMA_signal_4637 ;
    wire new_AGEMA_signal_4638 ;
    wire new_AGEMA_signal_4639 ;
    wire new_AGEMA_signal_4640 ;
    wire new_AGEMA_signal_4641 ;
    wire new_AGEMA_signal_4642 ;
    wire new_AGEMA_signal_4643 ;
    wire new_AGEMA_signal_4644 ;
    wire new_AGEMA_signal_4645 ;
    wire new_AGEMA_signal_4646 ;
    wire new_AGEMA_signal_4647 ;
    wire new_AGEMA_signal_4648 ;
    wire new_AGEMA_signal_4649 ;
    wire new_AGEMA_signal_4650 ;
    wire new_AGEMA_signal_4651 ;
    wire new_AGEMA_signal_4652 ;
    wire new_AGEMA_signal_4653 ;
    wire new_AGEMA_signal_4654 ;
    wire new_AGEMA_signal_4655 ;
    wire new_AGEMA_signal_4656 ;
    wire new_AGEMA_signal_4657 ;
    wire new_AGEMA_signal_4658 ;
    wire new_AGEMA_signal_4659 ;
    wire new_AGEMA_signal_4660 ;
    wire new_AGEMA_signal_4661 ;
    wire new_AGEMA_signal_4662 ;
    wire new_AGEMA_signal_4663 ;
    wire new_AGEMA_signal_4664 ;
    wire new_AGEMA_signal_4665 ;
    wire new_AGEMA_signal_4666 ;
    wire new_AGEMA_signal_4667 ;
    wire new_AGEMA_signal_4668 ;
    wire new_AGEMA_signal_4669 ;
    wire new_AGEMA_signal_4670 ;
    wire new_AGEMA_signal_4671 ;
    wire new_AGEMA_signal_4672 ;
    wire new_AGEMA_signal_4673 ;
    wire new_AGEMA_signal_4674 ;
    wire new_AGEMA_signal_4675 ;
    wire new_AGEMA_signal_4676 ;
    wire new_AGEMA_signal_4677 ;
    wire new_AGEMA_signal_4678 ;
    wire new_AGEMA_signal_4679 ;
    wire new_AGEMA_signal_4680 ;
    wire new_AGEMA_signal_4681 ;
    wire new_AGEMA_signal_4682 ;
    wire new_AGEMA_signal_4683 ;
    wire new_AGEMA_signal_4684 ;
    wire new_AGEMA_signal_4685 ;
    wire new_AGEMA_signal_4686 ;
    wire new_AGEMA_signal_4687 ;
    wire new_AGEMA_signal_4688 ;
    wire new_AGEMA_signal_4689 ;
    wire new_AGEMA_signal_4690 ;
    wire new_AGEMA_signal_4691 ;
    wire new_AGEMA_signal_4692 ;
    wire new_AGEMA_signal_4693 ;
    wire new_AGEMA_signal_4694 ;
    wire new_AGEMA_signal_4695 ;
    wire new_AGEMA_signal_4696 ;
    wire new_AGEMA_signal_4697 ;
    wire new_AGEMA_signal_4698 ;
    wire new_AGEMA_signal_4699 ;
    wire new_AGEMA_signal_4700 ;
    wire new_AGEMA_signal_4701 ;
    wire new_AGEMA_signal_4702 ;
    wire new_AGEMA_signal_4703 ;
    wire new_AGEMA_signal_4704 ;
    wire new_AGEMA_signal_4705 ;
    wire new_AGEMA_signal_4706 ;
    wire new_AGEMA_signal_4707 ;
    wire new_AGEMA_signal_4708 ;
    wire new_AGEMA_signal_4709 ;
    wire new_AGEMA_signal_4710 ;
    wire new_AGEMA_signal_4711 ;
    wire new_AGEMA_signal_4712 ;
    wire new_AGEMA_signal_4713 ;
    wire new_AGEMA_signal_4714 ;
    wire new_AGEMA_signal_4715 ;
    wire new_AGEMA_signal_4716 ;
    wire new_AGEMA_signal_4717 ;
    wire new_AGEMA_signal_4718 ;
    wire new_AGEMA_signal_4719 ;
    wire new_AGEMA_signal_4720 ;
    wire new_AGEMA_signal_4721 ;
    wire new_AGEMA_signal_4722 ;
    wire new_AGEMA_signal_4723 ;
    wire new_AGEMA_signal_4724 ;
    wire new_AGEMA_signal_4725 ;
    wire new_AGEMA_signal_4726 ;
    wire new_AGEMA_signal_4727 ;
    wire new_AGEMA_signal_4728 ;
    wire new_AGEMA_signal_4729 ;
    wire new_AGEMA_signal_4730 ;
    wire new_AGEMA_signal_4731 ;
    wire new_AGEMA_signal_4732 ;
    wire new_AGEMA_signal_4733 ;
    wire new_AGEMA_signal_4734 ;
    wire new_AGEMA_signal_4735 ;
    wire new_AGEMA_signal_4736 ;
    wire new_AGEMA_signal_4737 ;
    wire new_AGEMA_signal_4738 ;
    wire new_AGEMA_signal_4739 ;
    wire new_AGEMA_signal_4740 ;
    wire new_AGEMA_signal_4741 ;
    wire new_AGEMA_signal_4742 ;
    wire new_AGEMA_signal_4743 ;
    wire new_AGEMA_signal_4744 ;
    wire new_AGEMA_signal_4745 ;
    wire new_AGEMA_signal_4746 ;
    wire new_AGEMA_signal_4747 ;
    wire new_AGEMA_signal_4748 ;
    wire new_AGEMA_signal_4749 ;
    wire new_AGEMA_signal_4750 ;
    wire new_AGEMA_signal_4751 ;
    wire new_AGEMA_signal_4752 ;
    wire new_AGEMA_signal_4753 ;
    wire new_AGEMA_signal_4754 ;
    wire new_AGEMA_signal_4755 ;
    wire new_AGEMA_signal_4756 ;
    wire new_AGEMA_signal_4757 ;
    wire new_AGEMA_signal_4758 ;
    wire new_AGEMA_signal_4759 ;
    wire new_AGEMA_signal_4760 ;
    wire new_AGEMA_signal_4761 ;
    wire new_AGEMA_signal_4762 ;
    wire new_AGEMA_signal_4763 ;
    wire new_AGEMA_signal_4764 ;
    wire new_AGEMA_signal_4765 ;
    wire new_AGEMA_signal_4766 ;
    wire new_AGEMA_signal_4767 ;
    wire new_AGEMA_signal_4768 ;
    wire new_AGEMA_signal_4769 ;
    wire new_AGEMA_signal_4770 ;
    wire new_AGEMA_signal_4771 ;
    wire new_AGEMA_signal_4772 ;
    wire new_AGEMA_signal_4773 ;
    wire new_AGEMA_signal_4774 ;
    wire new_AGEMA_signal_4775 ;
    wire new_AGEMA_signal_4776 ;
    wire new_AGEMA_signal_4777 ;
    wire new_AGEMA_signal_4778 ;
    wire new_AGEMA_signal_4779 ;
    wire new_AGEMA_signal_4780 ;
    wire new_AGEMA_signal_4781 ;
    wire new_AGEMA_signal_4782 ;
    wire new_AGEMA_signal_4783 ;
    wire new_AGEMA_signal_4784 ;
    wire new_AGEMA_signal_4785 ;
    wire new_AGEMA_signal_4786 ;
    wire new_AGEMA_signal_4787 ;
    wire new_AGEMA_signal_4788 ;
    wire new_AGEMA_signal_4789 ;
    wire new_AGEMA_signal_4790 ;
    wire new_AGEMA_signal_4791 ;
    wire new_AGEMA_signal_4792 ;
    wire new_AGEMA_signal_4793 ;
    wire new_AGEMA_signal_4794 ;
    wire new_AGEMA_signal_4795 ;
    wire new_AGEMA_signal_4796 ;
    wire new_AGEMA_signal_4797 ;
    wire new_AGEMA_signal_4798 ;
    wire new_AGEMA_signal_4799 ;
    wire new_AGEMA_signal_4800 ;
    wire new_AGEMA_signal_4801 ;
    wire new_AGEMA_signal_4802 ;
    wire new_AGEMA_signal_4803 ;
    wire new_AGEMA_signal_4804 ;
    wire new_AGEMA_signal_4805 ;
    wire new_AGEMA_signal_4806 ;
    wire new_AGEMA_signal_4807 ;
    wire new_AGEMA_signal_4808 ;
    wire new_AGEMA_signal_4809 ;
    wire new_AGEMA_signal_4810 ;
    wire new_AGEMA_signal_4811 ;
    wire new_AGEMA_signal_4812 ;
    wire new_AGEMA_signal_4813 ;
    wire new_AGEMA_signal_4814 ;
    wire new_AGEMA_signal_4815 ;
    wire new_AGEMA_signal_4816 ;
    wire new_AGEMA_signal_4817 ;
    wire new_AGEMA_signal_4818 ;
    wire new_AGEMA_signal_4819 ;
    wire new_AGEMA_signal_4820 ;
    wire new_AGEMA_signal_4821 ;
    wire new_AGEMA_signal_4822 ;
    wire new_AGEMA_signal_4823 ;
    wire new_AGEMA_signal_4824 ;
    wire new_AGEMA_signal_4825 ;
    wire new_AGEMA_signal_4826 ;
    wire new_AGEMA_signal_4827 ;
    wire new_AGEMA_signal_4828 ;
    wire new_AGEMA_signal_4829 ;
    wire new_AGEMA_signal_4830 ;
    wire new_AGEMA_signal_4831 ;
    wire new_AGEMA_signal_4832 ;
    wire new_AGEMA_signal_4833 ;
    wire new_AGEMA_signal_4834 ;
    wire new_AGEMA_signal_4835 ;
    wire new_AGEMA_signal_4836 ;
    wire new_AGEMA_signal_4837 ;
    wire new_AGEMA_signal_4838 ;
    wire new_AGEMA_signal_4839 ;
    wire new_AGEMA_signal_4840 ;
    wire new_AGEMA_signal_4841 ;
    wire new_AGEMA_signal_4842 ;
    wire new_AGEMA_signal_4843 ;
    wire new_AGEMA_signal_4844 ;
    wire new_AGEMA_signal_4845 ;
    wire new_AGEMA_signal_4846 ;
    wire new_AGEMA_signal_4847 ;
    wire new_AGEMA_signal_4848 ;
    wire new_AGEMA_signal_4849 ;
    wire new_AGEMA_signal_4850 ;
    wire new_AGEMA_signal_4851 ;
    wire new_AGEMA_signal_4852 ;
    wire new_AGEMA_signal_4853 ;
    wire new_AGEMA_signal_4854 ;
    wire new_AGEMA_signal_4855 ;
    wire new_AGEMA_signal_4856 ;
    wire new_AGEMA_signal_4857 ;
    wire new_AGEMA_signal_4858 ;
    wire new_AGEMA_signal_4859 ;
    wire new_AGEMA_signal_4860 ;
    wire new_AGEMA_signal_4861 ;
    wire new_AGEMA_signal_4862 ;
    wire new_AGEMA_signal_4863 ;
    wire new_AGEMA_signal_4864 ;
    wire new_AGEMA_signal_4865 ;
    wire new_AGEMA_signal_4866 ;
    wire new_AGEMA_signal_4867 ;
    wire new_AGEMA_signal_4868 ;
    wire new_AGEMA_signal_4869 ;
    wire new_AGEMA_signal_4870 ;
    wire new_AGEMA_signal_4871 ;
    wire new_AGEMA_signal_4872 ;
    wire new_AGEMA_signal_4873 ;
    wire new_AGEMA_signal_4874 ;
    wire new_AGEMA_signal_4875 ;
    wire new_AGEMA_signal_4876 ;
    wire new_AGEMA_signal_4877 ;
    wire new_AGEMA_signal_4878 ;
    wire new_AGEMA_signal_4879 ;
    wire new_AGEMA_signal_4880 ;
    wire new_AGEMA_signal_4881 ;
    wire new_AGEMA_signal_4882 ;
    wire new_AGEMA_signal_4883 ;
    wire new_AGEMA_signal_4884 ;
    wire new_AGEMA_signal_4885 ;
    wire new_AGEMA_signal_4886 ;
    wire new_AGEMA_signal_4887 ;
    wire new_AGEMA_signal_4888 ;
    wire new_AGEMA_signal_4889 ;
    wire new_AGEMA_signal_4890 ;
    wire new_AGEMA_signal_4891 ;
    wire new_AGEMA_signal_4892 ;
    wire new_AGEMA_signal_4893 ;
    wire new_AGEMA_signal_4894 ;
    wire new_AGEMA_signal_4895 ;
    wire new_AGEMA_signal_4896 ;
    wire new_AGEMA_signal_4897 ;
    wire new_AGEMA_signal_4898 ;
    wire new_AGEMA_signal_4899 ;
    wire new_AGEMA_signal_4900 ;
    wire new_AGEMA_signal_4901 ;
    wire new_AGEMA_signal_4902 ;
    wire new_AGEMA_signal_4903 ;
    wire new_AGEMA_signal_4904 ;
    wire new_AGEMA_signal_4905 ;
    wire new_AGEMA_signal_4906 ;
    wire new_AGEMA_signal_4907 ;
    wire new_AGEMA_signal_4908 ;
    wire new_AGEMA_signal_4909 ;
    wire new_AGEMA_signal_4910 ;
    wire new_AGEMA_signal_4911 ;
    wire new_AGEMA_signal_4912 ;
    wire new_AGEMA_signal_4913 ;
    wire new_AGEMA_signal_4914 ;
    wire new_AGEMA_signal_4915 ;
    wire new_AGEMA_signal_4916 ;
    wire new_AGEMA_signal_4917 ;
    wire new_AGEMA_signal_4918 ;
    wire new_AGEMA_signal_4919 ;
    wire new_AGEMA_signal_4920 ;
    wire new_AGEMA_signal_4921 ;
    wire new_AGEMA_signal_4922 ;
    wire new_AGEMA_signal_4923 ;
    wire new_AGEMA_signal_4924 ;
    wire new_AGEMA_signal_4925 ;
    wire new_AGEMA_signal_4926 ;
    wire new_AGEMA_signal_4927 ;
    wire new_AGEMA_signal_4928 ;
    wire new_AGEMA_signal_4929 ;
    wire new_AGEMA_signal_4930 ;
    wire new_AGEMA_signal_4931 ;
    wire new_AGEMA_signal_4932 ;
    wire new_AGEMA_signal_4933 ;
    wire new_AGEMA_signal_4934 ;
    wire new_AGEMA_signal_4935 ;
    wire new_AGEMA_signal_4936 ;
    wire new_AGEMA_signal_4937 ;
    wire new_AGEMA_signal_4938 ;
    wire new_AGEMA_signal_4939 ;
    wire new_AGEMA_signal_4940 ;
    wire new_AGEMA_signal_4941 ;
    wire new_AGEMA_signal_4942 ;
    wire new_AGEMA_signal_4943 ;
    wire new_AGEMA_signal_4944 ;
    wire new_AGEMA_signal_4945 ;
    wire new_AGEMA_signal_4946 ;
    wire new_AGEMA_signal_4947 ;
    wire new_AGEMA_signal_4948 ;
    wire new_AGEMA_signal_4949 ;
    wire new_AGEMA_signal_4950 ;
    wire new_AGEMA_signal_4951 ;
    wire new_AGEMA_signal_4952 ;
    wire new_AGEMA_signal_4953 ;
    wire new_AGEMA_signal_4954 ;
    wire new_AGEMA_signal_4955 ;
    wire new_AGEMA_signal_4956 ;
    wire new_AGEMA_signal_4957 ;
    wire new_AGEMA_signal_4958 ;
    wire new_AGEMA_signal_4959 ;
    wire new_AGEMA_signal_4960 ;
    wire new_AGEMA_signal_4961 ;
    wire new_AGEMA_signal_4962 ;
    wire new_AGEMA_signal_4963 ;
    wire new_AGEMA_signal_4964 ;
    wire new_AGEMA_signal_4965 ;
    wire new_AGEMA_signal_4966 ;
    wire new_AGEMA_signal_4967 ;
    wire new_AGEMA_signal_4968 ;
    wire new_AGEMA_signal_4969 ;
    wire new_AGEMA_signal_4970 ;
    wire new_AGEMA_signal_4971 ;
    wire new_AGEMA_signal_4972 ;
    wire new_AGEMA_signal_4973 ;
    wire new_AGEMA_signal_4974 ;
    wire new_AGEMA_signal_4975 ;
    wire new_AGEMA_signal_4976 ;
    wire new_AGEMA_signal_4977 ;
    wire new_AGEMA_signal_4978 ;
    wire new_AGEMA_signal_4979 ;
    wire new_AGEMA_signal_4980 ;
    wire new_AGEMA_signal_4981 ;
    wire new_AGEMA_signal_4982 ;
    wire new_AGEMA_signal_4983 ;
    wire new_AGEMA_signal_4984 ;
    wire new_AGEMA_signal_4985 ;
    wire new_AGEMA_signal_4986 ;
    wire new_AGEMA_signal_4987 ;
    wire new_AGEMA_signal_4988 ;
    wire new_AGEMA_signal_4989 ;
    wire new_AGEMA_signal_4990 ;
    wire new_AGEMA_signal_4991 ;
    wire new_AGEMA_signal_4992 ;
    wire new_AGEMA_signal_4993 ;
    wire new_AGEMA_signal_4994 ;
    wire new_AGEMA_signal_4995 ;
    wire new_AGEMA_signal_4996 ;
    wire new_AGEMA_signal_4997 ;
    wire new_AGEMA_signal_4998 ;
    wire new_AGEMA_signal_4999 ;
    wire new_AGEMA_signal_5000 ;
    wire new_AGEMA_signal_5001 ;
    wire new_AGEMA_signal_5002 ;
    wire new_AGEMA_signal_5003 ;
    wire new_AGEMA_signal_5004 ;
    wire new_AGEMA_signal_5005 ;
    wire new_AGEMA_signal_5006 ;
    wire new_AGEMA_signal_5007 ;
    wire new_AGEMA_signal_5008 ;
    wire new_AGEMA_signal_5009 ;
    wire new_AGEMA_signal_5010 ;
    wire new_AGEMA_signal_5011 ;
    wire new_AGEMA_signal_5012 ;
    wire new_AGEMA_signal_5013 ;
    wire new_AGEMA_signal_5014 ;
    wire new_AGEMA_signal_5015 ;
    wire new_AGEMA_signal_5016 ;
    wire new_AGEMA_signal_5017 ;
    wire new_AGEMA_signal_5018 ;
    wire new_AGEMA_signal_5019 ;
    wire new_AGEMA_signal_5020 ;
    wire new_AGEMA_signal_5021 ;
    wire new_AGEMA_signal_5022 ;
    wire new_AGEMA_signal_5023 ;
    wire new_AGEMA_signal_5024 ;
    wire new_AGEMA_signal_5025 ;
    wire new_AGEMA_signal_5026 ;
    wire new_AGEMA_signal_5027 ;
    wire new_AGEMA_signal_5028 ;
    wire new_AGEMA_signal_5029 ;
    wire new_AGEMA_signal_5030 ;
    wire new_AGEMA_signal_5031 ;
    wire new_AGEMA_signal_5032 ;
    wire new_AGEMA_signal_5033 ;
    wire new_AGEMA_signal_5034 ;
    wire new_AGEMA_signal_5035 ;
    wire new_AGEMA_signal_5036 ;
    wire new_AGEMA_signal_5037 ;
    wire new_AGEMA_signal_5038 ;
    wire new_AGEMA_signal_5039 ;
    wire new_AGEMA_signal_5040 ;
    wire new_AGEMA_signal_5041 ;
    wire new_AGEMA_signal_5042 ;
    wire new_AGEMA_signal_5043 ;
    wire new_AGEMA_signal_5044 ;
    wire new_AGEMA_signal_5045 ;
    wire new_AGEMA_signal_5046 ;
    wire new_AGEMA_signal_5047 ;
    wire new_AGEMA_signal_5048 ;
    wire new_AGEMA_signal_5049 ;
    wire new_AGEMA_signal_5050 ;
    wire new_AGEMA_signal_5051 ;
    wire new_AGEMA_signal_5052 ;
    wire new_AGEMA_signal_5053 ;
    wire new_AGEMA_signal_5054 ;
    wire new_AGEMA_signal_5055 ;
    wire new_AGEMA_signal_5056 ;
    wire new_AGEMA_signal_5057 ;
    wire new_AGEMA_signal_5058 ;
    wire new_AGEMA_signal_5059 ;
    wire new_AGEMA_signal_5060 ;
    wire new_AGEMA_signal_5061 ;
    wire new_AGEMA_signal_5062 ;
    wire new_AGEMA_signal_5063 ;
    wire new_AGEMA_signal_5064 ;
    wire new_AGEMA_signal_5065 ;
    wire new_AGEMA_signal_5066 ;
    wire new_AGEMA_signal_5067 ;
    wire new_AGEMA_signal_5068 ;
    wire new_AGEMA_signal_5069 ;
    wire new_AGEMA_signal_5070 ;
    wire new_AGEMA_signal_5071 ;
    wire new_AGEMA_signal_5072 ;
    wire new_AGEMA_signal_5073 ;
    wire new_AGEMA_signal_5074 ;
    wire new_AGEMA_signal_5075 ;
    wire new_AGEMA_signal_5076 ;
    wire new_AGEMA_signal_5077 ;
    wire new_AGEMA_signal_5078 ;
    wire new_AGEMA_signal_5079 ;
    wire new_AGEMA_signal_5080 ;
    wire new_AGEMA_signal_5081 ;
    wire new_AGEMA_signal_5082 ;
    wire new_AGEMA_signal_5083 ;
    wire new_AGEMA_signal_5084 ;
    wire new_AGEMA_signal_5085 ;
    wire new_AGEMA_signal_5086 ;
    wire new_AGEMA_signal_5087 ;
    wire new_AGEMA_signal_5088 ;
    wire new_AGEMA_signal_5089 ;
    wire new_AGEMA_signal_5090 ;
    wire new_AGEMA_signal_5091 ;
    wire new_AGEMA_signal_5092 ;
    wire new_AGEMA_signal_5093 ;
    wire new_AGEMA_signal_5094 ;
    wire new_AGEMA_signal_5095 ;
    wire new_AGEMA_signal_5096 ;
    wire new_AGEMA_signal_5097 ;
    wire new_AGEMA_signal_5098 ;
    wire new_AGEMA_signal_5099 ;
    wire new_AGEMA_signal_5100 ;
    wire new_AGEMA_signal_5101 ;
    wire new_AGEMA_signal_5102 ;
    wire new_AGEMA_signal_5103 ;
    wire new_AGEMA_signal_5104 ;
    wire new_AGEMA_signal_5105 ;
    wire new_AGEMA_signal_5106 ;
    wire new_AGEMA_signal_5107 ;
    wire new_AGEMA_signal_5108 ;
    wire new_AGEMA_signal_5109 ;
    wire new_AGEMA_signal_5110 ;
    wire new_AGEMA_signal_5111 ;
    wire new_AGEMA_signal_5112 ;
    wire new_AGEMA_signal_5113 ;
    wire new_AGEMA_signal_5114 ;
    wire new_AGEMA_signal_5115 ;
    wire new_AGEMA_signal_5116 ;
    wire new_AGEMA_signal_5117 ;
    wire new_AGEMA_signal_5118 ;
    wire new_AGEMA_signal_5119 ;
    wire new_AGEMA_signal_5120 ;
    wire new_AGEMA_signal_5121 ;
    wire new_AGEMA_signal_5122 ;
    wire new_AGEMA_signal_5123 ;
    wire new_AGEMA_signal_5124 ;
    wire new_AGEMA_signal_5125 ;
    wire new_AGEMA_signal_5126 ;
    wire new_AGEMA_signal_5127 ;
    wire new_AGEMA_signal_5128 ;
    wire new_AGEMA_signal_5129 ;
    wire new_AGEMA_signal_5130 ;
    wire new_AGEMA_signal_5131 ;
    wire new_AGEMA_signal_5132 ;
    wire new_AGEMA_signal_5133 ;
    wire new_AGEMA_signal_5134 ;
    wire new_AGEMA_signal_5135 ;
    wire new_AGEMA_signal_5136 ;
    wire new_AGEMA_signal_5137 ;
    wire new_AGEMA_signal_5138 ;
    wire new_AGEMA_signal_5139 ;
    wire new_AGEMA_signal_5140 ;
    wire new_AGEMA_signal_5141 ;
    wire new_AGEMA_signal_5142 ;
    wire new_AGEMA_signal_5143 ;
    wire new_AGEMA_signal_5144 ;
    wire new_AGEMA_signal_5145 ;
    wire new_AGEMA_signal_5146 ;
    wire new_AGEMA_signal_5147 ;
    wire new_AGEMA_signal_5148 ;
    wire new_AGEMA_signal_5149 ;
    wire new_AGEMA_signal_5150 ;
    wire new_AGEMA_signal_5151 ;
    wire new_AGEMA_signal_5152 ;
    wire new_AGEMA_signal_5153 ;
    wire new_AGEMA_signal_5154 ;
    wire new_AGEMA_signal_5155 ;
    wire new_AGEMA_signal_5156 ;
    wire new_AGEMA_signal_5157 ;
    wire new_AGEMA_signal_5158 ;
    wire new_AGEMA_signal_5159 ;
    wire new_AGEMA_signal_5160 ;
    wire new_AGEMA_signal_5161 ;
    wire new_AGEMA_signal_5162 ;
    wire new_AGEMA_signal_5163 ;
    wire new_AGEMA_signal_5164 ;
    wire new_AGEMA_signal_5165 ;
    wire new_AGEMA_signal_5166 ;
    wire new_AGEMA_signal_5167 ;
    wire new_AGEMA_signal_5168 ;
    wire new_AGEMA_signal_5169 ;
    wire new_AGEMA_signal_5170 ;
    wire new_AGEMA_signal_5171 ;
    wire new_AGEMA_signal_5172 ;
    wire new_AGEMA_signal_5173 ;
    wire new_AGEMA_signal_5174 ;
    wire new_AGEMA_signal_5175 ;
    wire new_AGEMA_signal_5176 ;
    wire new_AGEMA_signal_5177 ;
    wire new_AGEMA_signal_5178 ;
    wire new_AGEMA_signal_5179 ;
    wire new_AGEMA_signal_5180 ;
    wire new_AGEMA_signal_5181 ;
    wire new_AGEMA_signal_5182 ;
    wire new_AGEMA_signal_5183 ;
    wire new_AGEMA_signal_5184 ;
    wire new_AGEMA_signal_5185 ;
    wire new_AGEMA_signal_5186 ;
    wire new_AGEMA_signal_5187 ;
    wire new_AGEMA_signal_5188 ;
    wire new_AGEMA_signal_5189 ;
    wire new_AGEMA_signal_5190 ;
    wire new_AGEMA_signal_5191 ;
    wire new_AGEMA_signal_5192 ;
    wire new_AGEMA_signal_5193 ;
    wire new_AGEMA_signal_5194 ;
    wire new_AGEMA_signal_5195 ;
    wire new_AGEMA_signal_5196 ;
    wire new_AGEMA_signal_5197 ;
    wire new_AGEMA_signal_5198 ;
    wire new_AGEMA_signal_5199 ;
    wire new_AGEMA_signal_5200 ;
    wire new_AGEMA_signal_5201 ;
    wire new_AGEMA_signal_5202 ;
    wire new_AGEMA_signal_5203 ;
    wire new_AGEMA_signal_5204 ;
    wire new_AGEMA_signal_5205 ;
    wire new_AGEMA_signal_5206 ;
    wire new_AGEMA_signal_5207 ;
    wire new_AGEMA_signal_5208 ;
    wire new_AGEMA_signal_5209 ;
    wire new_AGEMA_signal_5210 ;
    wire new_AGEMA_signal_5211 ;
    wire new_AGEMA_signal_5212 ;
    wire new_AGEMA_signal_5213 ;
    wire new_AGEMA_signal_5214 ;
    wire new_AGEMA_signal_5215 ;
    wire new_AGEMA_signal_5216 ;
    wire new_AGEMA_signal_5217 ;
    wire new_AGEMA_signal_5218 ;
    wire new_AGEMA_signal_5219 ;
    wire new_AGEMA_signal_5220 ;
    wire new_AGEMA_signal_5221 ;
    wire new_AGEMA_signal_5222 ;
    wire new_AGEMA_signal_5223 ;
    wire new_AGEMA_signal_5224 ;
    wire new_AGEMA_signal_5225 ;
    wire new_AGEMA_signal_5226 ;
    wire new_AGEMA_signal_5227 ;
    wire new_AGEMA_signal_5228 ;
    wire new_AGEMA_signal_5229 ;
    wire new_AGEMA_signal_5230 ;
    wire new_AGEMA_signal_5231 ;
    wire new_AGEMA_signal_5232 ;
    wire new_AGEMA_signal_5233 ;
    wire new_AGEMA_signal_5234 ;
    wire new_AGEMA_signal_5235 ;
    wire new_AGEMA_signal_5236 ;
    wire new_AGEMA_signal_5237 ;
    wire new_AGEMA_signal_5238 ;
    wire new_AGEMA_signal_5239 ;
    wire new_AGEMA_signal_5240 ;
    wire new_AGEMA_signal_5241 ;
    wire new_AGEMA_signal_5242 ;
    wire new_AGEMA_signal_5243 ;
    wire new_AGEMA_signal_5244 ;
    wire new_AGEMA_signal_5245 ;
    wire new_AGEMA_signal_5246 ;
    wire new_AGEMA_signal_5247 ;
    wire new_AGEMA_signal_5248 ;
    wire new_AGEMA_signal_5249 ;
    wire new_AGEMA_signal_5250 ;
    wire new_AGEMA_signal_5251 ;
    wire new_AGEMA_signal_5252 ;
    wire new_AGEMA_signal_5253 ;
    wire new_AGEMA_signal_5254 ;
    wire new_AGEMA_signal_5255 ;
    wire new_AGEMA_signal_5256 ;
    wire new_AGEMA_signal_5257 ;
    wire new_AGEMA_signal_5258 ;
    wire new_AGEMA_signal_5259 ;
    wire new_AGEMA_signal_5260 ;
    wire new_AGEMA_signal_5261 ;
    wire new_AGEMA_signal_5262 ;
    wire new_AGEMA_signal_5263 ;
    wire new_AGEMA_signal_5264 ;
    wire new_AGEMA_signal_5265 ;
    wire new_AGEMA_signal_5266 ;
    wire new_AGEMA_signal_5267 ;
    wire new_AGEMA_signal_5268 ;
    wire new_AGEMA_signal_5269 ;
    wire new_AGEMA_signal_5270 ;
    wire new_AGEMA_signal_5271 ;
    wire new_AGEMA_signal_5272 ;
    wire new_AGEMA_signal_5273 ;
    wire new_AGEMA_signal_5274 ;
    wire new_AGEMA_signal_5275 ;
    wire new_AGEMA_signal_5276 ;
    wire new_AGEMA_signal_5277 ;
    wire new_AGEMA_signal_5278 ;
    wire new_AGEMA_signal_5279 ;
    wire new_AGEMA_signal_5280 ;
    wire new_AGEMA_signal_5281 ;
    wire new_AGEMA_signal_5282 ;
    wire new_AGEMA_signal_5283 ;
    wire new_AGEMA_signal_5284 ;
    wire new_AGEMA_signal_5285 ;
    wire new_AGEMA_signal_5286 ;
    wire new_AGEMA_signal_5287 ;
    wire new_AGEMA_signal_5288 ;
    wire new_AGEMA_signal_5289 ;
    wire new_AGEMA_signal_5290 ;
    wire new_AGEMA_signal_5291 ;
    wire new_AGEMA_signal_5292 ;
    wire new_AGEMA_signal_5293 ;
    wire new_AGEMA_signal_5294 ;
    wire new_AGEMA_signal_5295 ;
    wire new_AGEMA_signal_5296 ;
    wire new_AGEMA_signal_5297 ;
    wire new_AGEMA_signal_5298 ;
    wire new_AGEMA_signal_5299 ;
    wire new_AGEMA_signal_5300 ;
    wire new_AGEMA_signal_5301 ;
    wire new_AGEMA_signal_5302 ;
    wire new_AGEMA_signal_5303 ;
    wire new_AGEMA_signal_5304 ;
    wire new_AGEMA_signal_5305 ;
    wire new_AGEMA_signal_5306 ;
    wire new_AGEMA_signal_5307 ;
    wire new_AGEMA_signal_5308 ;
    wire new_AGEMA_signal_5309 ;
    wire new_AGEMA_signal_5310 ;
    wire new_AGEMA_signal_5311 ;
    wire new_AGEMA_signal_5312 ;
    wire new_AGEMA_signal_5313 ;
    wire new_AGEMA_signal_5314 ;
    wire new_AGEMA_signal_5315 ;
    wire new_AGEMA_signal_5316 ;
    wire new_AGEMA_signal_5317 ;
    wire new_AGEMA_signal_5318 ;
    wire new_AGEMA_signal_5319 ;
    wire new_AGEMA_signal_5320 ;
    wire new_AGEMA_signal_5321 ;
    wire new_AGEMA_signal_5322 ;
    wire new_AGEMA_signal_5323 ;
    wire new_AGEMA_signal_5324 ;
    wire new_AGEMA_signal_5325 ;
    wire new_AGEMA_signal_5326 ;
    wire new_AGEMA_signal_5327 ;
    wire new_AGEMA_signal_5328 ;
    wire new_AGEMA_signal_5329 ;
    wire new_AGEMA_signal_5330 ;
    wire new_AGEMA_signal_5331 ;
    wire new_AGEMA_signal_5332 ;
    wire new_AGEMA_signal_5333 ;
    wire new_AGEMA_signal_5334 ;
    wire new_AGEMA_signal_5335 ;
    wire new_AGEMA_signal_5336 ;
    wire new_AGEMA_signal_5337 ;
    wire new_AGEMA_signal_5338 ;
    wire new_AGEMA_signal_5339 ;
    wire new_AGEMA_signal_5340 ;
    wire new_AGEMA_signal_5341 ;
    wire new_AGEMA_signal_5342 ;
    wire new_AGEMA_signal_5343 ;
    wire new_AGEMA_signal_5344 ;
    wire new_AGEMA_signal_5345 ;
    wire new_AGEMA_signal_5346 ;
    wire new_AGEMA_signal_5347 ;
    wire new_AGEMA_signal_5348 ;
    wire new_AGEMA_signal_5349 ;
    wire new_AGEMA_signal_5350 ;
    wire new_AGEMA_signal_5351 ;
    wire new_AGEMA_signal_5352 ;
    wire new_AGEMA_signal_5353 ;
    wire new_AGEMA_signal_5354 ;
    wire new_AGEMA_signal_5355 ;
    wire new_AGEMA_signal_5356 ;
    wire new_AGEMA_signal_5357 ;
    wire new_AGEMA_signal_5358 ;
    wire new_AGEMA_signal_5359 ;
    wire new_AGEMA_signal_5360 ;
    wire new_AGEMA_signal_5361 ;
    wire new_AGEMA_signal_5362 ;
    wire new_AGEMA_signal_5363 ;
    wire new_AGEMA_signal_5364 ;
    wire new_AGEMA_signal_5365 ;
    wire new_AGEMA_signal_5366 ;
    wire new_AGEMA_signal_5367 ;
    wire new_AGEMA_signal_5368 ;
    wire new_AGEMA_signal_5369 ;
    wire new_AGEMA_signal_5370 ;
    wire new_AGEMA_signal_5371 ;
    wire new_AGEMA_signal_5372 ;
    wire new_AGEMA_signal_5373 ;
    wire new_AGEMA_signal_5374 ;
    wire new_AGEMA_signal_5375 ;
    wire new_AGEMA_signal_5376 ;
    wire new_AGEMA_signal_5377 ;
    wire new_AGEMA_signal_5378 ;
    wire new_AGEMA_signal_5379 ;
    wire new_AGEMA_signal_5380 ;
    wire new_AGEMA_signal_5381 ;
    wire new_AGEMA_signal_5382 ;
    wire new_AGEMA_signal_5383 ;
    wire new_AGEMA_signal_5384 ;
    wire new_AGEMA_signal_5385 ;
    wire new_AGEMA_signal_5386 ;
    wire new_AGEMA_signal_5387 ;
    wire new_AGEMA_signal_5388 ;
    wire new_AGEMA_signal_5389 ;
    wire new_AGEMA_signal_5390 ;
    wire new_AGEMA_signal_5391 ;
    wire new_AGEMA_signal_5392 ;
    wire new_AGEMA_signal_5393 ;
    wire new_AGEMA_signal_5394 ;
    wire new_AGEMA_signal_5395 ;
    wire new_AGEMA_signal_5396 ;
    wire new_AGEMA_signal_5397 ;
    wire new_AGEMA_signal_5398 ;
    wire new_AGEMA_signal_5399 ;
    wire new_AGEMA_signal_5400 ;
    wire new_AGEMA_signal_5401 ;
    wire new_AGEMA_signal_5402 ;
    wire new_AGEMA_signal_5403 ;
    wire new_AGEMA_signal_5404 ;
    wire new_AGEMA_signal_5405 ;
    wire new_AGEMA_signal_5406 ;
    wire new_AGEMA_signal_5407 ;
    wire new_AGEMA_signal_5408 ;
    wire new_AGEMA_signal_5409 ;
    wire new_AGEMA_signal_5410 ;
    wire new_AGEMA_signal_5411 ;
    wire new_AGEMA_signal_5412 ;
    wire new_AGEMA_signal_5413 ;
    wire new_AGEMA_signal_5414 ;
    wire new_AGEMA_signal_5415 ;
    wire new_AGEMA_signal_5416 ;
    wire new_AGEMA_signal_5417 ;
    wire new_AGEMA_signal_5418 ;
    wire new_AGEMA_signal_5419 ;
    wire new_AGEMA_signal_5420 ;
    wire new_AGEMA_signal_5421 ;
    wire new_AGEMA_signal_5422 ;
    wire new_AGEMA_signal_5423 ;
    wire new_AGEMA_signal_5424 ;
    wire new_AGEMA_signal_5425 ;
    wire new_AGEMA_signal_5426 ;
    wire new_AGEMA_signal_5427 ;
    wire new_AGEMA_signal_5428 ;
    wire new_AGEMA_signal_5429 ;
    wire new_AGEMA_signal_5430 ;
    wire new_AGEMA_signal_5431 ;
    wire new_AGEMA_signal_5432 ;
    wire new_AGEMA_signal_5433 ;
    wire new_AGEMA_signal_5434 ;
    wire new_AGEMA_signal_5435 ;
    wire new_AGEMA_signal_5436 ;
    wire new_AGEMA_signal_5437 ;
    wire new_AGEMA_signal_5438 ;
    wire new_AGEMA_signal_5439 ;
    wire new_AGEMA_signal_5440 ;
    wire new_AGEMA_signal_5441 ;
    wire new_AGEMA_signal_5442 ;
    wire new_AGEMA_signal_5443 ;
    wire new_AGEMA_signal_5444 ;
    wire new_AGEMA_signal_5445 ;
    wire new_AGEMA_signal_5446 ;
    wire new_AGEMA_signal_5447 ;
    wire new_AGEMA_signal_5448 ;
    wire new_AGEMA_signal_5449 ;
    wire new_AGEMA_signal_5450 ;
    wire new_AGEMA_signal_5451 ;
    wire new_AGEMA_signal_5452 ;
    wire new_AGEMA_signal_5453 ;
    wire new_AGEMA_signal_5454 ;
    wire new_AGEMA_signal_5455 ;
    wire new_AGEMA_signal_5456 ;
    wire new_AGEMA_signal_5457 ;
    wire new_AGEMA_signal_5458 ;
    wire new_AGEMA_signal_5459 ;
    wire new_AGEMA_signal_5460 ;
    wire new_AGEMA_signal_5461 ;
    wire new_AGEMA_signal_5462 ;
    wire new_AGEMA_signal_5463 ;
    wire new_AGEMA_signal_5464 ;
    wire new_AGEMA_signal_5465 ;
    wire new_AGEMA_signal_5466 ;
    wire new_AGEMA_signal_5467 ;
    wire new_AGEMA_signal_5468 ;
    wire new_AGEMA_signal_5469 ;
    wire new_AGEMA_signal_5470 ;
    wire new_AGEMA_signal_5471 ;
    wire new_AGEMA_signal_5472 ;
    wire new_AGEMA_signal_5473 ;
    wire new_AGEMA_signal_5474 ;
    wire new_AGEMA_signal_5475 ;
    wire new_AGEMA_signal_5476 ;
    wire new_AGEMA_signal_5477 ;
    wire new_AGEMA_signal_5478 ;
    wire new_AGEMA_signal_5479 ;
    wire new_AGEMA_signal_5480 ;
    wire new_AGEMA_signal_5481 ;
    wire new_AGEMA_signal_5482 ;
    wire new_AGEMA_signal_5483 ;
    wire new_AGEMA_signal_5484 ;
    wire new_AGEMA_signal_5485 ;
    wire new_AGEMA_signal_5486 ;
    wire new_AGEMA_signal_5487 ;
    wire new_AGEMA_signal_5488 ;
    wire new_AGEMA_signal_5489 ;
    wire new_AGEMA_signal_5490 ;
    wire new_AGEMA_signal_5491 ;
    wire new_AGEMA_signal_5492 ;
    wire new_AGEMA_signal_5493 ;
    wire new_AGEMA_signal_5494 ;
    wire new_AGEMA_signal_5495 ;
    wire new_AGEMA_signal_5496 ;
    wire new_AGEMA_signal_5497 ;
    wire new_AGEMA_signal_5498 ;
    wire new_AGEMA_signal_5499 ;
    wire new_AGEMA_signal_5500 ;
    wire new_AGEMA_signal_5501 ;
    wire new_AGEMA_signal_5502 ;
    wire new_AGEMA_signal_5503 ;
    wire new_AGEMA_signal_5504 ;
    wire new_AGEMA_signal_5505 ;
    wire new_AGEMA_signal_5506 ;
    wire new_AGEMA_signal_5507 ;
    wire new_AGEMA_signal_5508 ;
    wire new_AGEMA_signal_5509 ;
    wire new_AGEMA_signal_5510 ;
    wire new_AGEMA_signal_5511 ;
    wire new_AGEMA_signal_5512 ;
    wire new_AGEMA_signal_5513 ;
    wire new_AGEMA_signal_5514 ;
    wire new_AGEMA_signal_5515 ;
    wire new_AGEMA_signal_5516 ;
    wire new_AGEMA_signal_5517 ;
    wire new_AGEMA_signal_5518 ;
    wire new_AGEMA_signal_5519 ;
    wire new_AGEMA_signal_5520 ;
    wire new_AGEMA_signal_5521 ;
    wire new_AGEMA_signal_5522 ;
    wire new_AGEMA_signal_5523 ;
    wire new_AGEMA_signal_5524 ;
    wire new_AGEMA_signal_5525 ;
    wire new_AGEMA_signal_5526 ;
    wire new_AGEMA_signal_5527 ;
    wire new_AGEMA_signal_5528 ;
    wire new_AGEMA_signal_5529 ;
    wire new_AGEMA_signal_5530 ;
    wire new_AGEMA_signal_5531 ;
    wire new_AGEMA_signal_5532 ;
    wire new_AGEMA_signal_5533 ;
    wire new_AGEMA_signal_5534 ;
    wire new_AGEMA_signal_5535 ;
    wire new_AGEMA_signal_5536 ;
    wire new_AGEMA_signal_5537 ;
    wire new_AGEMA_signal_5538 ;
    wire new_AGEMA_signal_5539 ;
    wire new_AGEMA_signal_5540 ;
    wire new_AGEMA_signal_5541 ;
    wire new_AGEMA_signal_5542 ;
    wire new_AGEMA_signal_5543 ;
    wire new_AGEMA_signal_5544 ;
    wire new_AGEMA_signal_5545 ;
    wire new_AGEMA_signal_5546 ;
    wire new_AGEMA_signal_5547 ;
    wire new_AGEMA_signal_5548 ;
    wire new_AGEMA_signal_5549 ;
    wire new_AGEMA_signal_5550 ;
    wire new_AGEMA_signal_5551 ;
    wire new_AGEMA_signal_5552 ;
    wire new_AGEMA_signal_5553 ;
    wire new_AGEMA_signal_5554 ;
    wire new_AGEMA_signal_5555 ;
    wire new_AGEMA_signal_5556 ;
    wire new_AGEMA_signal_5557 ;
    wire new_AGEMA_signal_5558 ;
    wire new_AGEMA_signal_5559 ;
    wire new_AGEMA_signal_5560 ;
    wire new_AGEMA_signal_5561 ;
    wire new_AGEMA_signal_5562 ;
    wire new_AGEMA_signal_5563 ;
    wire new_AGEMA_signal_5564 ;
    wire new_AGEMA_signal_5565 ;
    wire new_AGEMA_signal_5566 ;
    wire new_AGEMA_signal_5567 ;
    wire new_AGEMA_signal_5568 ;
    wire new_AGEMA_signal_5569 ;
    wire new_AGEMA_signal_5570 ;
    wire new_AGEMA_signal_5571 ;
    wire new_AGEMA_signal_5572 ;
    wire new_AGEMA_signal_5573 ;
    wire new_AGEMA_signal_5574 ;
    wire new_AGEMA_signal_5575 ;
    wire new_AGEMA_signal_5576 ;
    wire new_AGEMA_signal_5577 ;
    wire new_AGEMA_signal_5578 ;
    wire new_AGEMA_signal_5579 ;
    wire new_AGEMA_signal_5580 ;
    wire new_AGEMA_signal_5581 ;
    wire new_AGEMA_signal_5582 ;
    wire new_AGEMA_signal_5583 ;
    wire new_AGEMA_signal_5584 ;
    wire new_AGEMA_signal_5585 ;
    wire new_AGEMA_signal_5586 ;
    wire new_AGEMA_signal_5587 ;
    wire new_AGEMA_signal_5588 ;
    wire new_AGEMA_signal_5589 ;
    wire new_AGEMA_signal_5590 ;
    wire new_AGEMA_signal_5591 ;
    wire new_AGEMA_signal_5592 ;
    wire new_AGEMA_signal_5593 ;
    wire new_AGEMA_signal_5594 ;
    wire new_AGEMA_signal_5595 ;
    wire new_AGEMA_signal_5596 ;
    wire new_AGEMA_signal_5597 ;
    wire new_AGEMA_signal_5598 ;
    wire new_AGEMA_signal_5599 ;
    wire new_AGEMA_signal_5600 ;
    wire new_AGEMA_signal_5601 ;
    wire new_AGEMA_signal_5602 ;
    wire new_AGEMA_signal_5603 ;
    wire new_AGEMA_signal_5604 ;
    wire new_AGEMA_signal_5605 ;
    wire new_AGEMA_signal_5606 ;
    wire new_AGEMA_signal_5607 ;
    wire new_AGEMA_signal_5608 ;
    wire new_AGEMA_signal_5609 ;
    wire new_AGEMA_signal_5610 ;
    wire new_AGEMA_signal_5611 ;
    wire new_AGEMA_signal_5612 ;
    wire new_AGEMA_signal_5613 ;
    wire new_AGEMA_signal_5614 ;
    wire new_AGEMA_signal_5615 ;
    wire new_AGEMA_signal_5616 ;
    wire new_AGEMA_signal_5617 ;
    wire new_AGEMA_signal_5618 ;
    wire new_AGEMA_signal_5619 ;
    wire new_AGEMA_signal_5620 ;
    wire new_AGEMA_signal_5621 ;
    wire new_AGEMA_signal_5622 ;
    wire new_AGEMA_signal_5623 ;
    wire new_AGEMA_signal_5624 ;
    wire new_AGEMA_signal_5625 ;
    wire new_AGEMA_signal_5626 ;
    wire new_AGEMA_signal_5627 ;
    wire new_AGEMA_signal_5628 ;
    wire new_AGEMA_signal_5629 ;
    wire new_AGEMA_signal_5630 ;
    wire new_AGEMA_signal_5631 ;
    wire new_AGEMA_signal_5632 ;
    wire new_AGEMA_signal_5633 ;
    wire new_AGEMA_signal_5634 ;
    wire new_AGEMA_signal_5635 ;
    wire new_AGEMA_signal_5636 ;
    wire new_AGEMA_signal_5637 ;
    wire new_AGEMA_signal_5638 ;
    wire new_AGEMA_signal_5639 ;
    wire new_AGEMA_signal_5640 ;
    wire new_AGEMA_signal_5641 ;
    wire new_AGEMA_signal_5642 ;
    wire new_AGEMA_signal_5643 ;
    wire new_AGEMA_signal_5644 ;
    wire new_AGEMA_signal_5645 ;
    wire new_AGEMA_signal_5646 ;
    wire new_AGEMA_signal_5647 ;
    wire new_AGEMA_signal_5648 ;
    wire new_AGEMA_signal_5649 ;
    wire new_AGEMA_signal_5650 ;
    wire new_AGEMA_signal_5651 ;
    wire new_AGEMA_signal_5652 ;
    wire new_AGEMA_signal_5653 ;
    wire new_AGEMA_signal_5654 ;
    wire new_AGEMA_signal_5655 ;
    wire new_AGEMA_signal_5656 ;
    wire new_AGEMA_signal_5657 ;
    wire new_AGEMA_signal_5658 ;
    wire new_AGEMA_signal_5659 ;
    wire new_AGEMA_signal_5660 ;
    wire new_AGEMA_signal_5661 ;
    wire new_AGEMA_signal_5662 ;
    wire new_AGEMA_signal_5663 ;
    wire new_AGEMA_signal_5664 ;
    wire new_AGEMA_signal_5665 ;
    wire new_AGEMA_signal_5666 ;
    wire new_AGEMA_signal_5667 ;
    wire new_AGEMA_signal_5668 ;
    wire new_AGEMA_signal_5669 ;
    wire new_AGEMA_signal_5670 ;
    wire new_AGEMA_signal_5671 ;
    wire new_AGEMA_signal_5672 ;
    wire new_AGEMA_signal_5673 ;
    wire new_AGEMA_signal_5674 ;
    wire new_AGEMA_signal_5675 ;
    wire new_AGEMA_signal_5676 ;
    wire new_AGEMA_signal_5677 ;
    wire new_AGEMA_signal_5678 ;
    wire new_AGEMA_signal_5679 ;
    wire new_AGEMA_signal_5680 ;
    wire new_AGEMA_signal_5681 ;
    wire new_AGEMA_signal_5682 ;
    wire new_AGEMA_signal_5683 ;
    wire new_AGEMA_signal_5684 ;
    wire new_AGEMA_signal_5685 ;
    wire new_AGEMA_signal_5686 ;
    wire new_AGEMA_signal_5687 ;
    wire new_AGEMA_signal_5688 ;
    wire new_AGEMA_signal_5689 ;
    wire new_AGEMA_signal_5690 ;
    wire new_AGEMA_signal_5691 ;
    wire new_AGEMA_signal_5692 ;
    wire new_AGEMA_signal_5693 ;
    wire new_AGEMA_signal_5694 ;
    wire new_AGEMA_signal_5695 ;
    wire new_AGEMA_signal_5696 ;
    wire new_AGEMA_signal_5697 ;
    wire new_AGEMA_signal_5698 ;
    wire new_AGEMA_signal_5699 ;
    wire new_AGEMA_signal_5700 ;
    wire new_AGEMA_signal_5701 ;
    wire new_AGEMA_signal_5702 ;
    wire new_AGEMA_signal_5703 ;
    wire new_AGEMA_signal_5704 ;
    wire new_AGEMA_signal_5705 ;
    wire new_AGEMA_signal_5706 ;
    wire new_AGEMA_signal_5707 ;
    wire new_AGEMA_signal_5708 ;
    wire new_AGEMA_signal_5709 ;
    wire new_AGEMA_signal_5710 ;
    wire new_AGEMA_signal_5711 ;
    wire new_AGEMA_signal_5712 ;
    wire new_AGEMA_signal_5713 ;
    wire new_AGEMA_signal_5714 ;
    wire new_AGEMA_signal_5715 ;
    wire new_AGEMA_signal_5716 ;
    wire new_AGEMA_signal_5717 ;
    wire new_AGEMA_signal_5718 ;
    wire new_AGEMA_signal_5719 ;
    wire new_AGEMA_signal_5720 ;
    wire new_AGEMA_signal_5721 ;
    wire new_AGEMA_signal_5722 ;
    wire new_AGEMA_signal_5723 ;
    wire new_AGEMA_signal_5724 ;
    wire new_AGEMA_signal_5725 ;
    wire new_AGEMA_signal_5726 ;
    wire new_AGEMA_signal_5727 ;
    wire new_AGEMA_signal_5728 ;
    wire new_AGEMA_signal_5729 ;
    wire new_AGEMA_signal_5730 ;
    wire new_AGEMA_signal_5731 ;
    wire new_AGEMA_signal_5732 ;
    wire new_AGEMA_signal_5733 ;
    wire new_AGEMA_signal_5734 ;
    wire new_AGEMA_signal_5735 ;
    wire new_AGEMA_signal_5736 ;
    wire new_AGEMA_signal_5737 ;
    wire new_AGEMA_signal_5738 ;
    wire new_AGEMA_signal_5739 ;
    wire new_AGEMA_signal_5740 ;
    wire new_AGEMA_signal_5741 ;
    wire new_AGEMA_signal_5742 ;
    wire new_AGEMA_signal_5743 ;
    wire new_AGEMA_signal_5744 ;
    wire new_AGEMA_signal_5745 ;
    wire new_AGEMA_signal_5746 ;
    wire new_AGEMA_signal_5747 ;
    wire new_AGEMA_signal_5748 ;
    wire new_AGEMA_signal_5749 ;
    wire new_AGEMA_signal_5750 ;
    wire new_AGEMA_signal_5751 ;
    wire new_AGEMA_signal_5752 ;
    wire new_AGEMA_signal_5753 ;
    wire new_AGEMA_signal_5754 ;
    wire new_AGEMA_signal_5755 ;
    wire new_AGEMA_signal_5756 ;
    wire new_AGEMA_signal_5757 ;
    wire new_AGEMA_signal_5758 ;
    wire new_AGEMA_signal_5759 ;
    wire new_AGEMA_signal_5760 ;
    wire new_AGEMA_signal_5761 ;
    wire new_AGEMA_signal_5762 ;
    wire new_AGEMA_signal_5763 ;
    wire new_AGEMA_signal_5764 ;
    wire new_AGEMA_signal_5765 ;
    wire new_AGEMA_signal_5766 ;
    wire new_AGEMA_signal_5767 ;
    wire new_AGEMA_signal_5768 ;
    wire new_AGEMA_signal_5769 ;
    wire new_AGEMA_signal_5770 ;
    wire new_AGEMA_signal_5771 ;
    wire new_AGEMA_signal_5772 ;
    wire new_AGEMA_signal_5773 ;
    wire new_AGEMA_signal_5774 ;
    wire new_AGEMA_signal_5775 ;
    wire new_AGEMA_signal_5776 ;
    wire new_AGEMA_signal_5777 ;
    wire new_AGEMA_signal_5778 ;
    wire new_AGEMA_signal_5779 ;
    wire new_AGEMA_signal_5780 ;
    wire new_AGEMA_signal_5781 ;
    wire new_AGEMA_signal_5782 ;
    wire new_AGEMA_signal_5783 ;
    wire new_AGEMA_signal_5784 ;
    wire new_AGEMA_signal_5785 ;
    wire new_AGEMA_signal_5786 ;
    wire new_AGEMA_signal_5787 ;
    wire new_AGEMA_signal_5788 ;
    wire new_AGEMA_signal_5789 ;
    wire new_AGEMA_signal_5790 ;
    wire new_AGEMA_signal_5791 ;
    wire new_AGEMA_signal_5792 ;
    wire new_AGEMA_signal_5793 ;
    wire new_AGEMA_signal_5794 ;
    wire new_AGEMA_signal_5795 ;
    wire new_AGEMA_signal_5796 ;
    wire new_AGEMA_signal_5797 ;
    wire new_AGEMA_signal_5798 ;
    wire new_AGEMA_signal_5799 ;
    wire new_AGEMA_signal_5800 ;
    wire new_AGEMA_signal_5801 ;
    wire new_AGEMA_signal_5802 ;
    wire new_AGEMA_signal_5803 ;
    wire new_AGEMA_signal_5804 ;
    wire new_AGEMA_signal_5805 ;
    wire new_AGEMA_signal_5806 ;
    wire new_AGEMA_signal_5807 ;
    wire new_AGEMA_signal_5808 ;
    wire new_AGEMA_signal_5809 ;
    wire new_AGEMA_signal_5810 ;
    wire new_AGEMA_signal_5811 ;
    wire new_AGEMA_signal_5812 ;
    wire new_AGEMA_signal_5813 ;
    wire new_AGEMA_signal_5814 ;
    wire new_AGEMA_signal_5815 ;
    wire new_AGEMA_signal_5816 ;
    wire new_AGEMA_signal_5817 ;
    wire new_AGEMA_signal_5818 ;
    wire new_AGEMA_signal_5819 ;
    wire new_AGEMA_signal_5820 ;
    wire new_AGEMA_signal_5821 ;
    wire new_AGEMA_signal_5822 ;
    wire new_AGEMA_signal_5823 ;
    wire new_AGEMA_signal_5824 ;
    wire new_AGEMA_signal_5825 ;
    wire new_AGEMA_signal_5826 ;
    wire new_AGEMA_signal_5827 ;
    wire new_AGEMA_signal_5828 ;
    wire new_AGEMA_signal_5829 ;
    wire new_AGEMA_signal_5830 ;
    wire new_AGEMA_signal_5831 ;
    wire new_AGEMA_signal_5832 ;
    wire new_AGEMA_signal_5833 ;
    wire new_AGEMA_signal_5834 ;
    wire new_AGEMA_signal_5835 ;
    wire new_AGEMA_signal_5836 ;
    wire new_AGEMA_signal_5837 ;
    wire new_AGEMA_signal_5838 ;
    wire new_AGEMA_signal_5839 ;
    wire new_AGEMA_signal_5840 ;
    wire new_AGEMA_signal_5841 ;
    wire new_AGEMA_signal_5842 ;
    wire new_AGEMA_signal_5843 ;
    wire new_AGEMA_signal_5844 ;
    wire new_AGEMA_signal_5845 ;
    wire new_AGEMA_signal_5846 ;
    wire new_AGEMA_signal_5847 ;
    wire new_AGEMA_signal_5848 ;
    wire new_AGEMA_signal_5849 ;
    wire new_AGEMA_signal_5850 ;
    wire new_AGEMA_signal_5851 ;
    wire new_AGEMA_signal_5852 ;
    wire new_AGEMA_signal_5853 ;
    wire new_AGEMA_signal_5854 ;
    wire new_AGEMA_signal_5855 ;
    wire new_AGEMA_signal_5856 ;
    wire new_AGEMA_signal_5857 ;
    wire new_AGEMA_signal_5858 ;
    wire new_AGEMA_signal_5859 ;
    wire new_AGEMA_signal_5860 ;
    wire new_AGEMA_signal_5861 ;
    wire new_AGEMA_signal_5862 ;
    wire new_AGEMA_signal_5863 ;
    wire new_AGEMA_signal_5864 ;
    wire new_AGEMA_signal_5865 ;
    wire new_AGEMA_signal_5866 ;
    wire new_AGEMA_signal_5867 ;
    wire new_AGEMA_signal_5868 ;
    wire new_AGEMA_signal_5869 ;
    wire new_AGEMA_signal_5870 ;
    wire new_AGEMA_signal_5871 ;
    wire new_AGEMA_signal_5872 ;
    wire new_AGEMA_signal_5873 ;
    wire new_AGEMA_signal_5874 ;
    wire new_AGEMA_signal_5875 ;
    wire new_AGEMA_signal_5876 ;
    wire new_AGEMA_signal_5877 ;
    wire new_AGEMA_signal_5878 ;
    wire new_AGEMA_signal_5879 ;
    wire new_AGEMA_signal_5880 ;
    wire new_AGEMA_signal_5881 ;
    wire new_AGEMA_signal_5882 ;
    wire new_AGEMA_signal_5883 ;
    wire new_AGEMA_signal_5884 ;
    wire new_AGEMA_signal_5885 ;
    wire new_AGEMA_signal_5886 ;
    wire new_AGEMA_signal_5887 ;
    wire new_AGEMA_signal_5888 ;
    wire new_AGEMA_signal_5889 ;
    wire new_AGEMA_signal_5890 ;
    wire new_AGEMA_signal_5891 ;
    wire new_AGEMA_signal_5892 ;
    wire new_AGEMA_signal_5893 ;
    wire new_AGEMA_signal_5894 ;
    wire new_AGEMA_signal_5895 ;
    wire new_AGEMA_signal_5896 ;
    wire new_AGEMA_signal_5897 ;
    wire new_AGEMA_signal_5898 ;
    wire new_AGEMA_signal_5899 ;
    wire new_AGEMA_signal_5900 ;
    wire new_AGEMA_signal_5901 ;
    wire new_AGEMA_signal_5902 ;
    wire new_AGEMA_signal_5903 ;
    wire new_AGEMA_signal_5904 ;
    wire new_AGEMA_signal_5905 ;
    wire new_AGEMA_signal_5906 ;
    wire new_AGEMA_signal_5907 ;
    wire new_AGEMA_signal_5908 ;
    wire new_AGEMA_signal_5909 ;
    wire new_AGEMA_signal_5910 ;
    wire new_AGEMA_signal_5911 ;
    wire new_AGEMA_signal_5912 ;
    wire new_AGEMA_signal_5913 ;
    wire new_AGEMA_signal_5914 ;
    wire new_AGEMA_signal_5915 ;
    wire new_AGEMA_signal_5916 ;
    wire new_AGEMA_signal_5917 ;
    wire new_AGEMA_signal_5918 ;
    wire new_AGEMA_signal_5919 ;
    wire new_AGEMA_signal_5920 ;
    wire new_AGEMA_signal_5921 ;
    wire new_AGEMA_signal_5922 ;
    wire new_AGEMA_signal_5923 ;
    wire new_AGEMA_signal_5924 ;
    wire new_AGEMA_signal_5925 ;
    wire new_AGEMA_signal_5926 ;
    wire new_AGEMA_signal_5927 ;
    wire new_AGEMA_signal_5928 ;
    wire new_AGEMA_signal_5929 ;
    wire new_AGEMA_signal_5930 ;
    wire new_AGEMA_signal_5931 ;
    wire new_AGEMA_signal_5932 ;
    wire new_AGEMA_signal_5933 ;
    wire new_AGEMA_signal_5934 ;
    wire new_AGEMA_signal_5935 ;
    wire new_AGEMA_signal_5936 ;
    wire new_AGEMA_signal_5937 ;
    wire new_AGEMA_signal_5938 ;
    wire new_AGEMA_signal_5939 ;
    wire new_AGEMA_signal_5940 ;
    wire new_AGEMA_signal_5941 ;
    wire new_AGEMA_signal_5942 ;
    wire new_AGEMA_signal_5943 ;
    wire new_AGEMA_signal_5944 ;
    wire new_AGEMA_signal_5945 ;
    wire new_AGEMA_signal_5946 ;
    wire new_AGEMA_signal_5947 ;
    wire new_AGEMA_signal_5948 ;
    wire new_AGEMA_signal_5949 ;
    wire new_AGEMA_signal_5950 ;
    wire new_AGEMA_signal_5951 ;
    wire new_AGEMA_signal_5952 ;
    wire new_AGEMA_signal_5953 ;
    wire new_AGEMA_signal_5954 ;
    wire new_AGEMA_signal_5955 ;
    wire new_AGEMA_signal_5956 ;
    wire new_AGEMA_signal_5957 ;
    wire new_AGEMA_signal_5958 ;
    wire new_AGEMA_signal_5959 ;
    wire new_AGEMA_signal_5960 ;
    wire new_AGEMA_signal_5961 ;
    wire new_AGEMA_signal_5962 ;
    wire new_AGEMA_signal_5963 ;
    wire new_AGEMA_signal_5964 ;
    wire new_AGEMA_signal_5965 ;
    wire new_AGEMA_signal_5966 ;
    wire new_AGEMA_signal_5967 ;
    wire new_AGEMA_signal_5968 ;
    wire new_AGEMA_signal_5969 ;
    wire new_AGEMA_signal_5970 ;
    wire new_AGEMA_signal_5971 ;
    wire new_AGEMA_signal_5972 ;
    wire new_AGEMA_signal_5973 ;
    wire new_AGEMA_signal_5974 ;
    wire new_AGEMA_signal_5975 ;
    wire new_AGEMA_signal_5976 ;
    wire new_AGEMA_signal_5977 ;
    wire new_AGEMA_signal_5978 ;
    wire new_AGEMA_signal_5979 ;
    wire new_AGEMA_signal_5980 ;
    wire new_AGEMA_signal_5981 ;
    wire new_AGEMA_signal_5982 ;
    wire new_AGEMA_signal_5983 ;
    wire new_AGEMA_signal_5984 ;
    wire new_AGEMA_signal_5985 ;
    wire new_AGEMA_signal_5986 ;
    wire new_AGEMA_signal_5987 ;
    wire new_AGEMA_signal_5988 ;
    wire new_AGEMA_signal_5989 ;
    wire new_AGEMA_signal_5990 ;
    wire new_AGEMA_signal_5991 ;
    wire new_AGEMA_signal_5992 ;
    wire new_AGEMA_signal_5993 ;
    wire new_AGEMA_signal_5994 ;
    wire new_AGEMA_signal_5995 ;
    wire new_AGEMA_signal_5996 ;
    wire new_AGEMA_signal_5997 ;
    wire new_AGEMA_signal_5998 ;
    wire new_AGEMA_signal_5999 ;
    wire new_AGEMA_signal_6000 ;
    wire new_AGEMA_signal_6001 ;
    wire new_AGEMA_signal_6002 ;
    wire new_AGEMA_signal_6003 ;
    wire new_AGEMA_signal_6004 ;
    wire new_AGEMA_signal_6005 ;
    wire new_AGEMA_signal_6006 ;
    wire new_AGEMA_signal_6007 ;
    wire new_AGEMA_signal_6008 ;
    wire new_AGEMA_signal_6009 ;
    wire new_AGEMA_signal_6010 ;
    wire new_AGEMA_signal_6011 ;
    wire new_AGEMA_signal_6012 ;
    wire new_AGEMA_signal_6013 ;
    wire new_AGEMA_signal_6014 ;
    wire new_AGEMA_signal_6015 ;
    wire new_AGEMA_signal_6016 ;
    wire new_AGEMA_signal_6017 ;
    wire new_AGEMA_signal_6018 ;
    wire new_AGEMA_signal_6019 ;
    wire new_AGEMA_signal_6020 ;
    wire new_AGEMA_signal_6021 ;
    wire new_AGEMA_signal_6022 ;
    wire new_AGEMA_signal_6023 ;
    wire new_AGEMA_signal_6024 ;
    wire new_AGEMA_signal_6025 ;
    wire new_AGEMA_signal_6026 ;
    wire new_AGEMA_signal_6027 ;
    wire new_AGEMA_signal_6028 ;
    wire new_AGEMA_signal_6029 ;
    wire new_AGEMA_signal_6030 ;
    wire new_AGEMA_signal_6031 ;
    wire new_AGEMA_signal_6032 ;
    wire new_AGEMA_signal_6033 ;
    wire new_AGEMA_signal_6034 ;
    wire new_AGEMA_signal_6035 ;
    wire new_AGEMA_signal_6036 ;
    wire new_AGEMA_signal_6037 ;
    wire new_AGEMA_signal_6038 ;
    wire new_AGEMA_signal_6039 ;
    wire new_AGEMA_signal_6040 ;
    wire new_AGEMA_signal_6041 ;
    wire new_AGEMA_signal_6042 ;
    wire new_AGEMA_signal_6043 ;
    wire new_AGEMA_signal_6044 ;
    wire new_AGEMA_signal_6045 ;
    wire new_AGEMA_signal_6046 ;
    wire new_AGEMA_signal_6047 ;
    wire new_AGEMA_signal_6048 ;
    wire new_AGEMA_signal_6049 ;
    wire new_AGEMA_signal_6050 ;
    wire new_AGEMA_signal_6051 ;
    wire new_AGEMA_signal_6052 ;
    wire new_AGEMA_signal_6053 ;
    wire new_AGEMA_signal_6054 ;
    wire new_AGEMA_signal_6055 ;
    wire new_AGEMA_signal_6056 ;
    wire new_AGEMA_signal_6057 ;
    wire new_AGEMA_signal_6058 ;
    wire new_AGEMA_signal_6059 ;
    wire new_AGEMA_signal_6060 ;
    wire new_AGEMA_signal_6061 ;
    wire new_AGEMA_signal_6062 ;
    wire new_AGEMA_signal_6063 ;
    wire new_AGEMA_signal_6064 ;
    wire new_AGEMA_signal_6065 ;
    wire new_AGEMA_signal_6066 ;
    wire new_AGEMA_signal_6067 ;
    wire new_AGEMA_signal_6068 ;
    wire new_AGEMA_signal_6069 ;
    wire new_AGEMA_signal_6070 ;
    wire new_AGEMA_signal_6071 ;
    wire new_AGEMA_signal_6072 ;
    wire new_AGEMA_signal_6073 ;
    wire new_AGEMA_signal_6074 ;
    wire new_AGEMA_signal_6075 ;
    wire new_AGEMA_signal_6076 ;
    wire new_AGEMA_signal_6077 ;
    wire new_AGEMA_signal_6078 ;
    wire new_AGEMA_signal_6079 ;
    wire new_AGEMA_signal_6080 ;
    wire new_AGEMA_signal_6081 ;
    wire new_AGEMA_signal_6082 ;
    wire new_AGEMA_signal_6083 ;
    wire new_AGEMA_signal_6084 ;
    wire new_AGEMA_signal_6085 ;
    wire new_AGEMA_signal_6086 ;
    wire new_AGEMA_signal_6087 ;
    wire new_AGEMA_signal_6088 ;
    wire new_AGEMA_signal_6089 ;
    wire new_AGEMA_signal_6090 ;
    wire new_AGEMA_signal_6091 ;
    wire new_AGEMA_signal_6092 ;
    wire new_AGEMA_signal_6093 ;
    wire new_AGEMA_signal_6094 ;
    wire new_AGEMA_signal_6095 ;
    wire new_AGEMA_signal_6096 ;
    wire new_AGEMA_signal_6097 ;
    wire new_AGEMA_signal_6098 ;
    wire new_AGEMA_signal_6099 ;
    wire new_AGEMA_signal_6100 ;
    wire new_AGEMA_signal_6101 ;
    wire new_AGEMA_signal_6102 ;
    wire new_AGEMA_signal_6103 ;
    wire new_AGEMA_signal_6104 ;
    wire new_AGEMA_signal_6105 ;
    wire new_AGEMA_signal_6106 ;
    wire new_AGEMA_signal_6107 ;
    wire new_AGEMA_signal_6108 ;
    wire new_AGEMA_signal_6109 ;
    wire new_AGEMA_signal_6110 ;
    wire new_AGEMA_signal_6111 ;
    wire new_AGEMA_signal_6112 ;
    wire new_AGEMA_signal_6113 ;
    wire new_AGEMA_signal_6114 ;
    wire new_AGEMA_signal_6115 ;
    wire new_AGEMA_signal_6116 ;
    wire new_AGEMA_signal_6117 ;
    wire new_AGEMA_signal_6118 ;
    wire new_AGEMA_signal_6119 ;
    wire new_AGEMA_signal_6120 ;
    wire new_AGEMA_signal_6121 ;
    wire new_AGEMA_signal_6122 ;
    wire new_AGEMA_signal_6123 ;
    wire new_AGEMA_signal_6124 ;
    wire new_AGEMA_signal_6125 ;
    wire new_AGEMA_signal_6126 ;
    wire new_AGEMA_signal_6127 ;
    wire new_AGEMA_signal_6128 ;
    wire new_AGEMA_signal_6129 ;
    wire new_AGEMA_signal_6130 ;
    wire new_AGEMA_signal_6131 ;
    wire new_AGEMA_signal_6132 ;
    wire new_AGEMA_signal_6133 ;
    wire new_AGEMA_signal_6134 ;
    wire new_AGEMA_signal_6135 ;
    wire new_AGEMA_signal_6136 ;
    wire new_AGEMA_signal_6137 ;
    wire new_AGEMA_signal_6138 ;
    wire new_AGEMA_signal_6139 ;
    wire new_AGEMA_signal_6140 ;
    wire new_AGEMA_signal_6141 ;
    wire new_AGEMA_signal_6142 ;
    wire new_AGEMA_signal_6143 ;
    wire new_AGEMA_signal_6144 ;
    wire new_AGEMA_signal_6145 ;
    wire new_AGEMA_signal_6146 ;
    wire new_AGEMA_signal_6147 ;
    wire new_AGEMA_signal_6148 ;
    wire new_AGEMA_signal_6149 ;
    wire new_AGEMA_signal_6150 ;
    wire new_AGEMA_signal_6151 ;
    wire new_AGEMA_signal_6152 ;
    wire new_AGEMA_signal_6153 ;
    wire new_AGEMA_signal_6154 ;
    wire new_AGEMA_signal_6155 ;
    wire new_AGEMA_signal_6156 ;
    wire new_AGEMA_signal_6157 ;
    wire new_AGEMA_signal_6158 ;
    wire new_AGEMA_signal_6159 ;
    wire new_AGEMA_signal_6160 ;
    wire new_AGEMA_signal_6161 ;
    wire new_AGEMA_signal_6162 ;
    wire new_AGEMA_signal_6163 ;
    wire new_AGEMA_signal_6164 ;
    wire new_AGEMA_signal_6165 ;
    wire new_AGEMA_signal_6166 ;
    wire new_AGEMA_signal_6167 ;
    wire new_AGEMA_signal_6168 ;
    wire new_AGEMA_signal_6169 ;
    wire new_AGEMA_signal_6170 ;
    wire new_AGEMA_signal_6171 ;
    wire new_AGEMA_signal_6172 ;
    wire new_AGEMA_signal_6173 ;
    wire new_AGEMA_signal_6174 ;
    wire new_AGEMA_signal_6175 ;
    wire new_AGEMA_signal_6176 ;
    wire new_AGEMA_signal_6177 ;
    wire new_AGEMA_signal_6178 ;
    wire new_AGEMA_signal_6179 ;
    wire new_AGEMA_signal_6180 ;
    wire new_AGEMA_signal_6181 ;
    wire new_AGEMA_signal_6182 ;
    wire new_AGEMA_signal_6183 ;
    wire new_AGEMA_signal_6184 ;
    wire new_AGEMA_signal_6185 ;
    wire new_AGEMA_signal_6186 ;
    wire new_AGEMA_signal_6187 ;
    wire new_AGEMA_signal_6188 ;
    wire new_AGEMA_signal_6189 ;
    wire new_AGEMA_signal_6190 ;
    wire new_AGEMA_signal_6191 ;
    wire new_AGEMA_signal_6192 ;
    wire new_AGEMA_signal_6193 ;
    wire new_AGEMA_signal_6194 ;
    wire new_AGEMA_signal_6195 ;
    wire new_AGEMA_signal_6196 ;
    wire new_AGEMA_signal_6197 ;
    wire new_AGEMA_signal_6198 ;
    wire new_AGEMA_signal_6199 ;
    wire new_AGEMA_signal_6200 ;
    wire new_AGEMA_signal_6201 ;
    wire new_AGEMA_signal_6202 ;
    wire new_AGEMA_signal_6203 ;
    wire new_AGEMA_signal_6204 ;
    wire new_AGEMA_signal_6205 ;
    wire new_AGEMA_signal_6206 ;
    wire new_AGEMA_signal_6207 ;
    wire new_AGEMA_signal_6208 ;
    wire new_AGEMA_signal_6209 ;
    wire new_AGEMA_signal_6210 ;
    wire new_AGEMA_signal_6211 ;
    wire new_AGEMA_signal_6212 ;
    wire new_AGEMA_signal_6213 ;
    wire new_AGEMA_signal_6214 ;
    wire new_AGEMA_signal_6215 ;
    wire new_AGEMA_signal_6216 ;
    wire new_AGEMA_signal_6217 ;
    wire new_AGEMA_signal_6218 ;
    wire new_AGEMA_signal_6219 ;
    wire new_AGEMA_signal_6220 ;
    wire new_AGEMA_signal_6221 ;
    wire new_AGEMA_signal_6222 ;
    wire new_AGEMA_signal_6223 ;
    wire new_AGEMA_signal_6224 ;
    wire new_AGEMA_signal_6225 ;
    wire new_AGEMA_signal_6226 ;
    wire new_AGEMA_signal_6227 ;
    wire new_AGEMA_signal_6228 ;
    wire new_AGEMA_signal_6229 ;
    wire new_AGEMA_signal_6230 ;
    wire new_AGEMA_signal_6231 ;
    wire new_AGEMA_signal_6232 ;
    wire new_AGEMA_signal_6233 ;
    wire new_AGEMA_signal_6234 ;
    wire new_AGEMA_signal_6235 ;
    wire new_AGEMA_signal_6236 ;
    wire new_AGEMA_signal_6237 ;
    wire new_AGEMA_signal_6238 ;
    wire new_AGEMA_signal_6239 ;
    wire new_AGEMA_signal_6240 ;
    wire new_AGEMA_signal_6241 ;
    wire new_AGEMA_signal_6242 ;
    wire new_AGEMA_signal_6243 ;
    wire new_AGEMA_signal_6244 ;
    wire new_AGEMA_signal_6245 ;
    wire new_AGEMA_signal_6246 ;
    wire new_AGEMA_signal_6247 ;
    wire new_AGEMA_signal_6248 ;
    wire new_AGEMA_signal_6249 ;
    wire new_AGEMA_signal_6250 ;
    wire new_AGEMA_signal_6251 ;
    wire new_AGEMA_signal_6252 ;
    wire new_AGEMA_signal_6253 ;
    wire new_AGEMA_signal_6254 ;
    wire new_AGEMA_signal_6255 ;
    wire new_AGEMA_signal_6256 ;
    wire new_AGEMA_signal_6257 ;
    wire new_AGEMA_signal_6258 ;
    wire new_AGEMA_signal_6259 ;
    wire new_AGEMA_signal_6260 ;
    wire new_AGEMA_signal_6261 ;
    wire new_AGEMA_signal_6262 ;
    wire new_AGEMA_signal_6263 ;
    wire new_AGEMA_signal_6264 ;
    wire new_AGEMA_signal_6265 ;
    wire new_AGEMA_signal_6266 ;
    wire new_AGEMA_signal_6267 ;
    wire new_AGEMA_signal_6268 ;
    wire new_AGEMA_signal_6269 ;
    wire new_AGEMA_signal_6270 ;
    wire new_AGEMA_signal_6271 ;
    wire new_AGEMA_signal_6272 ;
    wire new_AGEMA_signal_6273 ;
    wire new_AGEMA_signal_6274 ;
    wire new_AGEMA_signal_6275 ;
    wire new_AGEMA_signal_6276 ;
    wire new_AGEMA_signal_6277 ;
    wire new_AGEMA_signal_6278 ;
    wire new_AGEMA_signal_6279 ;
    wire new_AGEMA_signal_6280 ;
    wire new_AGEMA_signal_6281 ;
    wire new_AGEMA_signal_6282 ;
    wire new_AGEMA_signal_6283 ;
    wire new_AGEMA_signal_6284 ;
    wire new_AGEMA_signal_6285 ;
    wire new_AGEMA_signal_6286 ;
    wire new_AGEMA_signal_6287 ;
    wire new_AGEMA_signal_6288 ;
    wire new_AGEMA_signal_6289 ;
    wire new_AGEMA_signal_6290 ;
    wire new_AGEMA_signal_6291 ;
    wire new_AGEMA_signal_6292 ;
    wire new_AGEMA_signal_6293 ;
    wire new_AGEMA_signal_6294 ;
    wire new_AGEMA_signal_6295 ;
    wire new_AGEMA_signal_6296 ;
    wire new_AGEMA_signal_6297 ;

    /* cells in depth 0 */
    INV_X1 U28 ( .A (selSR), .ZN (n12) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) U29 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({new_AGEMA_signal_1983, keyStateIn[0]}), .c ({new_AGEMA_signal_1984, StateOutXORroundKey[0]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) U30 ( .a ({ciphertext_s1[121], ciphertext_s0[121]}), .b ({new_AGEMA_signal_1986, keyStateIn[1]}), .c ({new_AGEMA_signal_1987, StateOutXORroundKey[1]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) U31 ( .a ({ciphertext_s1[122], ciphertext_s0[122]}), .b ({new_AGEMA_signal_1989, keyStateIn[2]}), .c ({new_AGEMA_signal_1990, StateOutXORroundKey[2]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) U32 ( .a ({ciphertext_s1[123], ciphertext_s0[123]}), .b ({new_AGEMA_signal_1992, keyStateIn[3]}), .c ({new_AGEMA_signal_1993, StateOutXORroundKey[3]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) U33 ( .a ({ciphertext_s1[124], ciphertext_s0[124]}), .b ({new_AGEMA_signal_1995, keyStateIn[4]}), .c ({new_AGEMA_signal_1996, StateOutXORroundKey[4]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) U34 ( .a ({ciphertext_s1[125], ciphertext_s0[125]}), .b ({new_AGEMA_signal_1998, keyStateIn[5]}), .c ({new_AGEMA_signal_1999, StateOutXORroundKey[5]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) U35 ( .a ({ciphertext_s1[126], ciphertext_s0[126]}), .b ({new_AGEMA_signal_2001, keyStateIn[6]}), .c ({new_AGEMA_signal_2002, StateOutXORroundKey[6]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) U36 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({new_AGEMA_signal_2004, keyStateIn[7]}), .c ({new_AGEMA_signal_2005, StateOutXORroundKey[7]}) ) ;
    NAND2_X1 U37 ( .A1 (intFinal), .A2 (finalStep), .ZN (n13) ) ;
    NOR2_X1 U38 ( .A1 (n10), .A2 (n13), .ZN (done) ) ;
    AND2_X1 U39 ( .A1 (notFirst), .A2 (selXOR), .ZN (intselXOR) ) ;
    INV_X1 U40 ( .A (start), .ZN (n9) ) ;
    NOR2_X1 ctrl_U20 ( .A1 (ctrl_n16), .A2 (ctrl_n4), .ZN (ctrl_nRstSeq4) ) ;
    XNOR2_X1 ctrl_U19 ( .A (ctrl_seq6Out_4_), .B (ctrl_seq6In_1_), .ZN (ctrl_n13) ) ;
    NOR2_X1 ctrl_U18 ( .A1 (ctrl_n15), .A2 (ctrl_n14), .ZN (finalStep) ) ;
    NAND2_X1 ctrl_U17 ( .A1 (ctrl_seq4In_1_), .A2 (ctrl_n2), .ZN (ctrl_n14) ) ;
    INV_X1 ctrl_U16 ( .A (ctrl_n16), .ZN (ctrl_n15) ) ;
    INV_X1 ctrl_U15 ( .A (ctrl_seq4Out_1_), .ZN (ctrl_n2) ) ;
    NAND2_X1 ctrl_U14 ( .A1 (ctrl_n11), .A2 (ctrl_n10), .ZN (ctrl_N14) ) ;
    NAND2_X1 ctrl_U13 ( .A1 (selXOR), .A2 (ctrl_n6), .ZN (ctrl_n11) ) ;
    NOR2_X1 ctrl_U12 ( .A1 (ctrl_seq6In_3_), .A2 (ctrl_seq6Out_4_), .ZN (ctrl_n7) ) ;
    NOR2_X1 ctrl_U11 ( .A1 (ctrl_seq6In_1_), .A2 (ctrl_seq6In_4_), .ZN (ctrl_n8) ) ;
    NOR2_X1 ctrl_U10 ( .A1 (ctrl_n4), .A2 (ctrl_n5), .ZN (selXOR) ) ;
    NOR2_X1 ctrl_U9 ( .A1 (ctrl_seq4Out_1_), .A2 (ctrl_seq4In_1_), .ZN (ctrl_n5) ) ;
    INV_X1 ctrl_U8 ( .A (nReset), .ZN (ctrl_n4) ) ;
    NAND2_X1 ctrl_U7 ( .A1 (ctrl_n8), .A2 (ctrl_n7), .ZN (ctrl_n9) ) ;
    NOR2_X1 ctrl_U6 ( .A1 (ctrl_seq6In_2_), .A2 (ctrl_n9), .ZN (ctrl_n16) ) ;
    NAND2_X1 ctrl_U5 ( .A1 (nReset), .A2 (ctrl_n16), .ZN (ctrl_n10) ) ;
    INV_X1 ctrl_U4 ( .A (ctrl_n10), .ZN (selSR) ) ;
    NOR2_X1 ctrl_U3 ( .A1 (ctrl_n12), .A2 (ctrl_n4), .ZN (selMC) ) ;
    MUX2_X1 ctrl_seq6_SFF_0_MUXInst_U1 ( .S (nReset), .A (1'b1), .B (ctrl_n13), .Z (ctrl_seq6_SFF_0_QD) ) ;
    MUX2_X1 ctrl_seq6_SFF_1_MUXInst_U1 ( .S (nReset), .A (1'b0), .B (ctrl_seq6In_1_), .Z (ctrl_seq6_SFF_1_QD) ) ;
    MUX2_X1 ctrl_seq6_SFF_2_MUXInst_U1 ( .S (nReset), .A (1'b1), .B (ctrl_seq6In_2_), .Z (ctrl_seq6_SFF_2_QD) ) ;
    MUX2_X1 ctrl_seq6_SFF_3_MUXInst_U1 ( .S (nReset), .A (1'b0), .B (ctrl_seq6In_3_), .Z (ctrl_seq6_SFF_3_QD) ) ;
    MUX2_X1 ctrl_seq6_SFF_4_MUXInst_U1 ( .S (nReset), .A (1'b1), .B (ctrl_seq6In_4_), .Z (ctrl_seq6_SFF_4_QD) ) ;
    MUX2_X1 ctrl_seq4_SFF_0_MUXInst_U1 ( .S (ctrl_nRstSeq4), .A (1'b1), .B (ctrl_n2), .Z (ctrl_seq4_SFF_0_QD) ) ;
    MUX2_X1 ctrl_seq4_SFF_1_MUXInst_U1 ( .S (ctrl_nRstSeq4), .A (1'b0), .B (ctrl_seq4In_1_), .Z (ctrl_seq4_SFF_1_QD) ) ;
    INV_X1 ctrl_CSselMC_reg_U1 ( .A (ctrl_n6), .ZN (ctrl_n12) ) ;
    INV_X1 stateArray_U21 ( .A (selMC), .ZN (stateArray_n24) ) ;
    INV_X1 stateArray_U20 ( .A (stateArray_n24), .ZN (stateArray_n22) ) ;
    INV_X1 stateArray_U19 ( .A (nReset), .ZN (stateArray_n33) ) ;
    INV_X1 stateArray_U18 ( .A (stateArray_n33), .ZN (stateArray_n25) ) ;
    INV_X1 stateArray_U17 ( .A (stateArray_n21), .ZN (stateArray_n13) ) ;
    INV_X1 stateArray_U16 ( .A (stateArray_n24), .ZN (stateArray_n23) ) ;
    INV_X1 stateArray_U15 ( .A (stateArray_n33), .ZN (stateArray_n29) ) ;
    INV_X1 stateArray_U14 ( .A (stateArray_n21), .ZN (stateArray_n17) ) ;
    INV_X1 stateArray_U13 ( .A (stateArray_n33), .ZN (stateArray_n31) ) ;
    INV_X1 stateArray_U12 ( .A (stateArray_n21), .ZN (stateArray_n19) ) ;
    INV_X1 stateArray_U11 ( .A (stateArray_n33), .ZN (stateArray_n27) ) ;
    INV_X1 stateArray_U10 ( .A (stateArray_n21), .ZN (stateArray_n15) ) ;
    INV_X1 stateArray_U9 ( .A (stateArray_n33), .ZN (stateArray_n32) ) ;
    INV_X1 stateArray_U8 ( .A (stateArray_n21), .ZN (stateArray_n20) ) ;
    INV_X1 stateArray_U7 ( .A (stateArray_n33), .ZN (stateArray_n30) ) ;
    INV_X1 stateArray_U6 ( .A (stateArray_n21), .ZN (stateArray_n18) ) ;
    INV_X1 stateArray_U5 ( .A (stateArray_n33), .ZN (stateArray_n28) ) ;
    INV_X1 stateArray_U4 ( .A (stateArray_n21), .ZN (stateArray_n16) ) ;
    INV_X1 stateArray_U3 ( .A (stateArray_n33), .ZN (stateArray_n26) ) ;
    INV_X1 stateArray_U2 ( .A (stateArray_n21), .ZN (stateArray_n14) ) ;
    INV_X1 stateArray_U1 ( .A (selSR), .ZN (stateArray_n21) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S00reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2156, stateArray_inS00ser[0]}), .a ({ciphertext_s1[120], ciphertext_s0[120]}), .c ({new_AGEMA_signal_3126, stateArray_S00reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S00reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2159, stateArray_inS00ser[1]}), .a ({ciphertext_s1[121], ciphertext_s0[121]}), .c ({new_AGEMA_signal_3127, stateArray_S00reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S00reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2162, stateArray_inS00ser[2]}), .a ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_3128, stateArray_S00reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S00reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2165, stateArray_inS00ser[3]}), .a ({ciphertext_s1[123], ciphertext_s0[123]}), .c ({new_AGEMA_signal_3129, stateArray_S00reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S00reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2168, stateArray_inS00ser[4]}), .a ({ciphertext_s1[124], ciphertext_s0[124]}), .c ({new_AGEMA_signal_3130, stateArray_S00reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S00reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2171, stateArray_inS00ser[5]}), .a ({ciphertext_s1[125], ciphertext_s0[125]}), .c ({new_AGEMA_signal_3131, stateArray_S00reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S00reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2174, stateArray_inS00ser[6]}), .a ({ciphertext_s1[126], ciphertext_s0[126]}), .c ({new_AGEMA_signal_3132, stateArray_S00reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S00reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2177, stateArray_inS00ser[7]}), .a ({ciphertext_s1[127], ciphertext_s0[127]}), .c ({new_AGEMA_signal_3133, stateArray_S00reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S01reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2180, stateArray_inS01ser[0]}), .a ({ciphertext_s1[112], ciphertext_s0[112]}), .c ({new_AGEMA_signal_3134, stateArray_S01reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S01reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2183, stateArray_inS01ser[1]}), .a ({ciphertext_s1[113], ciphertext_s0[113]}), .c ({new_AGEMA_signal_3135, stateArray_S01reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S01reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2186, stateArray_inS01ser[2]}), .a ({ciphertext_s1[114], ciphertext_s0[114]}), .c ({new_AGEMA_signal_3136, stateArray_S01reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S01reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2189, stateArray_inS01ser[3]}), .a ({ciphertext_s1[115], ciphertext_s0[115]}), .c ({new_AGEMA_signal_3137, stateArray_S01reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S01reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2192, stateArray_inS01ser[4]}), .a ({ciphertext_s1[116], ciphertext_s0[116]}), .c ({new_AGEMA_signal_3138, stateArray_S01reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S01reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2195, stateArray_inS01ser[5]}), .a ({ciphertext_s1[117], ciphertext_s0[117]}), .c ({new_AGEMA_signal_3139, stateArray_S01reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S01reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2198, stateArray_inS01ser[6]}), .a ({ciphertext_s1[118], ciphertext_s0[118]}), .c ({new_AGEMA_signal_3140, stateArray_S01reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S01reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2201, stateArray_inS01ser[7]}), .a ({ciphertext_s1[119], ciphertext_s0[119]}), .c ({new_AGEMA_signal_3141, stateArray_S01reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S02reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_2204, stateArray_inS02ser[0]}), .a ({ciphertext_s1[104], ciphertext_s0[104]}), .c ({new_AGEMA_signal_3142, stateArray_S02reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S02reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_2207, stateArray_inS02ser[1]}), .a ({ciphertext_s1[105], ciphertext_s0[105]}), .c ({new_AGEMA_signal_3143, stateArray_S02reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S02reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_2210, stateArray_inS02ser[2]}), .a ({ciphertext_s1[106], ciphertext_s0[106]}), .c ({new_AGEMA_signal_3144, stateArray_S02reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S02reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_2213, stateArray_inS02ser[3]}), .a ({ciphertext_s1[107], ciphertext_s0[107]}), .c ({new_AGEMA_signal_3145, stateArray_S02reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S02reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_2216, stateArray_inS02ser[4]}), .a ({ciphertext_s1[108], ciphertext_s0[108]}), .c ({new_AGEMA_signal_3146, stateArray_S02reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S02reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_2219, stateArray_inS02ser[5]}), .a ({ciphertext_s1[109], ciphertext_s0[109]}), .c ({new_AGEMA_signal_3147, stateArray_S02reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S02reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_2222, stateArray_inS02ser[6]}), .a ({ciphertext_s1[110], ciphertext_s0[110]}), .c ({new_AGEMA_signal_3148, stateArray_S02reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S02reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_2225, stateArray_inS02ser[7]}), .a ({ciphertext_s1[111], ciphertext_s0[111]}), .c ({new_AGEMA_signal_3149, stateArray_S02reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S03reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_3046, stateArray_inS03ser[0]}), .a ({ciphertext_s1[96], ciphertext_s0[96]}), .c ({new_AGEMA_signal_3150, stateArray_S03reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S03reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_3048, stateArray_inS03ser[1]}), .a ({ciphertext_s1[97], ciphertext_s0[97]}), .c ({new_AGEMA_signal_3151, stateArray_S03reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S03reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_3050, stateArray_inS03ser[2]}), .a ({ciphertext_s1[98], ciphertext_s0[98]}), .c ({new_AGEMA_signal_3152, stateArray_S03reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S03reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_3052, stateArray_inS03ser[3]}), .a ({ciphertext_s1[99], ciphertext_s0[99]}), .c ({new_AGEMA_signal_3153, stateArray_S03reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S03reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_3054, stateArray_inS03ser[4]}), .a ({ciphertext_s1[100], ciphertext_s0[100]}), .c ({new_AGEMA_signal_3154, stateArray_S03reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S03reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_3056, stateArray_inS03ser[5]}), .a ({ciphertext_s1[101], ciphertext_s0[101]}), .c ({new_AGEMA_signal_3155, stateArray_S03reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S03reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_3058, stateArray_inS03ser[6]}), .a ({ciphertext_s1[102], ciphertext_s0[102]}), .c ({new_AGEMA_signal_3156, stateArray_S03reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S03reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_3060, stateArray_inS03ser[7]}), .a ({ciphertext_s1[103], ciphertext_s0[103]}), .c ({new_AGEMA_signal_3157, stateArray_S03reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S10reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2228, stateArray_inS10ser[0]}), .a ({ciphertext_s1[80], ciphertext_s0[80]}), .c ({new_AGEMA_signal_3158, stateArray_S10reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S10reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2231, stateArray_inS10ser[1]}), .a ({ciphertext_s1[81], ciphertext_s0[81]}), .c ({new_AGEMA_signal_3159, stateArray_S10reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S10reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2234, stateArray_inS10ser[2]}), .a ({ciphertext_s1[82], ciphertext_s0[82]}), .c ({new_AGEMA_signal_3160, stateArray_S10reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S10reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2237, stateArray_inS10ser[3]}), .a ({ciphertext_s1[83], ciphertext_s0[83]}), .c ({new_AGEMA_signal_3161, stateArray_S10reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S10reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2240, stateArray_inS10ser[4]}), .a ({ciphertext_s1[84], ciphertext_s0[84]}), .c ({new_AGEMA_signal_3162, stateArray_S10reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S10reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2243, stateArray_inS10ser[5]}), .a ({ciphertext_s1[85], ciphertext_s0[85]}), .c ({new_AGEMA_signal_3163, stateArray_S10reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S10reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2246, stateArray_inS10ser[6]}), .a ({ciphertext_s1[86], ciphertext_s0[86]}), .c ({new_AGEMA_signal_3164, stateArray_S10reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S10reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2249, stateArray_inS10ser[7]}), .a ({ciphertext_s1[87], ciphertext_s0[87]}), .c ({new_AGEMA_signal_3165, stateArray_S10reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S11reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2252, stateArray_inS11ser[0]}), .a ({ciphertext_s1[72], ciphertext_s0[72]}), .c ({new_AGEMA_signal_3166, stateArray_S11reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S11reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2255, stateArray_inS11ser[1]}), .a ({ciphertext_s1[73], ciphertext_s0[73]}), .c ({new_AGEMA_signal_3167, stateArray_S11reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S11reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2258, stateArray_inS11ser[2]}), .a ({ciphertext_s1[74], ciphertext_s0[74]}), .c ({new_AGEMA_signal_3168, stateArray_S11reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S11reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2261, stateArray_inS11ser[3]}), .a ({ciphertext_s1[75], ciphertext_s0[75]}), .c ({new_AGEMA_signal_3169, stateArray_S11reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S11reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2264, stateArray_inS11ser[4]}), .a ({ciphertext_s1[76], ciphertext_s0[76]}), .c ({new_AGEMA_signal_3170, stateArray_S11reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S11reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2267, stateArray_inS11ser[5]}), .a ({ciphertext_s1[77], ciphertext_s0[77]}), .c ({new_AGEMA_signal_3171, stateArray_S11reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S11reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2270, stateArray_inS11ser[6]}), .a ({ciphertext_s1[78], ciphertext_s0[78]}), .c ({new_AGEMA_signal_3172, stateArray_S11reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S11reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2273, stateArray_inS11ser[7]}), .a ({ciphertext_s1[79], ciphertext_s0[79]}), .c ({new_AGEMA_signal_3173, stateArray_S11reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S12reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_2276, stateArray_inS12ser[0]}), .a ({ciphertext_s1[64], ciphertext_s0[64]}), .c ({new_AGEMA_signal_3174, stateArray_S12reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S12reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_2279, stateArray_inS12ser[1]}), .a ({ciphertext_s1[65], ciphertext_s0[65]}), .c ({new_AGEMA_signal_3175, stateArray_S12reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S12reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_2282, stateArray_inS12ser[2]}), .a ({ciphertext_s1[66], ciphertext_s0[66]}), .c ({new_AGEMA_signal_3176, stateArray_S12reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S12reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_2285, stateArray_inS12ser[3]}), .a ({ciphertext_s1[67], ciphertext_s0[67]}), .c ({new_AGEMA_signal_3177, stateArray_S12reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S12reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_2288, stateArray_inS12ser[4]}), .a ({ciphertext_s1[68], ciphertext_s0[68]}), .c ({new_AGEMA_signal_3178, stateArray_S12reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S12reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_2291, stateArray_inS12ser[5]}), .a ({ciphertext_s1[69], ciphertext_s0[69]}), .c ({new_AGEMA_signal_3179, stateArray_S12reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S12reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_2294, stateArray_inS12ser[6]}), .a ({ciphertext_s1[70], ciphertext_s0[70]}), .c ({new_AGEMA_signal_3180, stateArray_S12reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S12reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_2297, stateArray_inS12ser[7]}), .a ({ciphertext_s1[71], ciphertext_s0[71]}), .c ({new_AGEMA_signal_3181, stateArray_S12reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S13reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_3062, stateArray_inS13ser[0]}), .a ({ciphertext_s1[88], ciphertext_s0[88]}), .c ({new_AGEMA_signal_3182, stateArray_S13reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S13reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_3064, stateArray_inS13ser[1]}), .a ({ciphertext_s1[89], ciphertext_s0[89]}), .c ({new_AGEMA_signal_3183, stateArray_S13reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S13reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_3066, stateArray_inS13ser[2]}), .a ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_3184, stateArray_S13reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S13reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_3068, stateArray_inS13ser[3]}), .a ({ciphertext_s1[91], ciphertext_s0[91]}), .c ({new_AGEMA_signal_3185, stateArray_S13reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S13reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_3070, stateArray_inS13ser[4]}), .a ({ciphertext_s1[92], ciphertext_s0[92]}), .c ({new_AGEMA_signal_3186, stateArray_S13reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S13reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_3072, stateArray_inS13ser[5]}), .a ({ciphertext_s1[93], ciphertext_s0[93]}), .c ({new_AGEMA_signal_3187, stateArray_S13reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S13reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_3074, stateArray_inS13ser[6]}), .a ({ciphertext_s1[94], ciphertext_s0[94]}), .c ({new_AGEMA_signal_3188, stateArray_S13reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S13reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_3076, stateArray_inS13ser[7]}), .a ({ciphertext_s1[95], ciphertext_s0[95]}), .c ({new_AGEMA_signal_3189, stateArray_S13reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S20reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2300, stateArray_inS20ser[0]}), .a ({ciphertext_s1[40], ciphertext_s0[40]}), .c ({new_AGEMA_signal_3190, stateArray_S20reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S20reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2303, stateArray_inS20ser[1]}), .a ({ciphertext_s1[41], ciphertext_s0[41]}), .c ({new_AGEMA_signal_3191, stateArray_S20reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S20reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2306, stateArray_inS20ser[2]}), .a ({ciphertext_s1[42], ciphertext_s0[42]}), .c ({new_AGEMA_signal_3192, stateArray_S20reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S20reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2309, stateArray_inS20ser[3]}), .a ({ciphertext_s1[43], ciphertext_s0[43]}), .c ({new_AGEMA_signal_3193, stateArray_S20reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S20reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2312, stateArray_inS20ser[4]}), .a ({ciphertext_s1[44], ciphertext_s0[44]}), .c ({new_AGEMA_signal_3194, stateArray_S20reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S20reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2315, stateArray_inS20ser[5]}), .a ({ciphertext_s1[45], ciphertext_s0[45]}), .c ({new_AGEMA_signal_3195, stateArray_S20reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S20reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2318, stateArray_inS20ser[6]}), .a ({ciphertext_s1[46], ciphertext_s0[46]}), .c ({new_AGEMA_signal_3196, stateArray_S20reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S20reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2321, stateArray_inS20ser[7]}), .a ({ciphertext_s1[47], ciphertext_s0[47]}), .c ({new_AGEMA_signal_3197, stateArray_S20reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S21reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2324, stateArray_inS21ser[0]}), .a ({ciphertext_s1[32], ciphertext_s0[32]}), .c ({new_AGEMA_signal_3198, stateArray_S21reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S21reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2327, stateArray_inS21ser[1]}), .a ({ciphertext_s1[33], ciphertext_s0[33]}), .c ({new_AGEMA_signal_3199, stateArray_S21reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S21reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2330, stateArray_inS21ser[2]}), .a ({ciphertext_s1[34], ciphertext_s0[34]}), .c ({new_AGEMA_signal_3200, stateArray_S21reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S21reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2333, stateArray_inS21ser[3]}), .a ({ciphertext_s1[35], ciphertext_s0[35]}), .c ({new_AGEMA_signal_3201, stateArray_S21reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S21reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2336, stateArray_inS21ser[4]}), .a ({ciphertext_s1[36], ciphertext_s0[36]}), .c ({new_AGEMA_signal_3202, stateArray_S21reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S21reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2339, stateArray_inS21ser[5]}), .a ({ciphertext_s1[37], ciphertext_s0[37]}), .c ({new_AGEMA_signal_3203, stateArray_S21reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S21reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2342, stateArray_inS21ser[6]}), .a ({ciphertext_s1[38], ciphertext_s0[38]}), .c ({new_AGEMA_signal_3204, stateArray_S21reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S21reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2345, stateArray_inS21ser[7]}), .a ({ciphertext_s1[39], ciphertext_s0[39]}), .c ({new_AGEMA_signal_3205, stateArray_S21reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S22reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_2348, stateArray_inS22ser[0]}), .a ({ciphertext_s1[56], ciphertext_s0[56]}), .c ({new_AGEMA_signal_3206, stateArray_S22reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S22reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_2351, stateArray_inS22ser[1]}), .a ({ciphertext_s1[57], ciphertext_s0[57]}), .c ({new_AGEMA_signal_3207, stateArray_S22reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S22reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_2354, stateArray_inS22ser[2]}), .a ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_3208, stateArray_S22reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S22reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_2357, stateArray_inS22ser[3]}), .a ({ciphertext_s1[59], ciphertext_s0[59]}), .c ({new_AGEMA_signal_3209, stateArray_S22reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S22reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_2360, stateArray_inS22ser[4]}), .a ({ciphertext_s1[60], ciphertext_s0[60]}), .c ({new_AGEMA_signal_3210, stateArray_S22reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S22reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_2363, stateArray_inS22ser[5]}), .a ({ciphertext_s1[61], ciphertext_s0[61]}), .c ({new_AGEMA_signal_3211, stateArray_S22reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S22reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_2366, stateArray_inS22ser[6]}), .a ({ciphertext_s1[62], ciphertext_s0[62]}), .c ({new_AGEMA_signal_3212, stateArray_S22reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S22reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_2369, stateArray_inS22ser[7]}), .a ({ciphertext_s1[63], ciphertext_s0[63]}), .c ({new_AGEMA_signal_3213, stateArray_S22reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S23reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_3078, stateArray_inS23ser[0]}), .a ({ciphertext_s1[48], ciphertext_s0[48]}), .c ({new_AGEMA_signal_3214, stateArray_S23reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S23reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_3080, stateArray_inS23ser[1]}), .a ({ciphertext_s1[49], ciphertext_s0[49]}), .c ({new_AGEMA_signal_3215, stateArray_S23reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S23reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_3082, stateArray_inS23ser[2]}), .a ({ciphertext_s1[50], ciphertext_s0[50]}), .c ({new_AGEMA_signal_3216, stateArray_S23reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S23reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_3084, stateArray_inS23ser[3]}), .a ({ciphertext_s1[51], ciphertext_s0[51]}), .c ({new_AGEMA_signal_3217, stateArray_S23reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S23reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_3086, stateArray_inS23ser[4]}), .a ({ciphertext_s1[52], ciphertext_s0[52]}), .c ({new_AGEMA_signal_3218, stateArray_S23reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S23reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_3088, stateArray_inS23ser[5]}), .a ({ciphertext_s1[53], ciphertext_s0[53]}), .c ({new_AGEMA_signal_3219, stateArray_S23reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S23reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_3090, stateArray_inS23ser[6]}), .a ({ciphertext_s1[54], ciphertext_s0[54]}), .c ({new_AGEMA_signal_3220, stateArray_S23reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S23reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_3092, stateArray_inS23ser[7]}), .a ({ciphertext_s1[55], ciphertext_s0[55]}), .c ({new_AGEMA_signal_3221, stateArray_S23reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S30reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_2372, stateArray_inS30ser[0]}), .a ({ciphertext_s1[0], ciphertext_s0[0]}), .c ({new_AGEMA_signal_3222, stateArray_S30reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S30reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_2375, stateArray_inS30ser[1]}), .a ({ciphertext_s1[1], ciphertext_s0[1]}), .c ({new_AGEMA_signal_3223, stateArray_S30reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S30reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_2378, stateArray_inS30ser[2]}), .a ({ciphertext_s1[2], ciphertext_s0[2]}), .c ({new_AGEMA_signal_3224, stateArray_S30reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S30reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_2381, stateArray_inS30ser[3]}), .a ({ciphertext_s1[3], ciphertext_s0[3]}), .c ({new_AGEMA_signal_3225, stateArray_S30reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S30reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_2384, stateArray_inS30ser[4]}), .a ({ciphertext_s1[4], ciphertext_s0[4]}), .c ({new_AGEMA_signal_3226, stateArray_S30reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S30reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_2387, stateArray_inS30ser[5]}), .a ({ciphertext_s1[5], ciphertext_s0[5]}), .c ({new_AGEMA_signal_3227, stateArray_S30reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S30reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_2390, stateArray_inS30ser[6]}), .a ({ciphertext_s1[6], ciphertext_s0[6]}), .c ({new_AGEMA_signal_3228, stateArray_S30reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S30reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_2393, stateArray_inS30ser[7]}), .a ({ciphertext_s1[7], ciphertext_s0[7]}), .c ({new_AGEMA_signal_3229, stateArray_S30reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S31reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_2396, stateArray_inS31ser[0]}), .a ({ciphertext_s1[24], ciphertext_s0[24]}), .c ({new_AGEMA_signal_3230, stateArray_S31reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S31reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_2399, stateArray_inS31ser[1]}), .a ({ciphertext_s1[25], ciphertext_s0[25]}), .c ({new_AGEMA_signal_3231, stateArray_S31reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S31reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_2402, stateArray_inS31ser[2]}), .a ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_3232, stateArray_S31reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S31reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_2405, stateArray_inS31ser[3]}), .a ({ciphertext_s1[27], ciphertext_s0[27]}), .c ({new_AGEMA_signal_3233, stateArray_S31reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S31reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_2408, stateArray_inS31ser[4]}), .a ({ciphertext_s1[28], ciphertext_s0[28]}), .c ({new_AGEMA_signal_3234, stateArray_S31reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S31reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_2411, stateArray_inS31ser[5]}), .a ({ciphertext_s1[29], ciphertext_s0[29]}), .c ({new_AGEMA_signal_3235, stateArray_S31reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S31reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_2414, stateArray_inS31ser[6]}), .a ({ciphertext_s1[30], ciphertext_s0[30]}), .c ({new_AGEMA_signal_3236, stateArray_S31reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S31reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_2417, stateArray_inS31ser[7]}), .a ({ciphertext_s1[31], ciphertext_s0[31]}), .c ({new_AGEMA_signal_3237, stateArray_S31reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S32reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_2420, stateArray_inS32ser[0]}), .a ({ciphertext_s1[16], ciphertext_s0[16]}), .c ({new_AGEMA_signal_3238, stateArray_S32reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S32reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_2423, stateArray_inS32ser[1]}), .a ({ciphertext_s1[17], ciphertext_s0[17]}), .c ({new_AGEMA_signal_3239, stateArray_S32reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S32reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_2426, stateArray_inS32ser[2]}), .a ({ciphertext_s1[18], ciphertext_s0[18]}), .c ({new_AGEMA_signal_3240, stateArray_S32reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S32reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_2429, stateArray_inS32ser[3]}), .a ({ciphertext_s1[19], ciphertext_s0[19]}), .c ({new_AGEMA_signal_3241, stateArray_S32reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S32reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_2432, stateArray_inS32ser[4]}), .a ({ciphertext_s1[20], ciphertext_s0[20]}), .c ({new_AGEMA_signal_3242, stateArray_S32reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S32reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_2435, stateArray_inS32ser[5]}), .a ({ciphertext_s1[21], ciphertext_s0[21]}), .c ({new_AGEMA_signal_3243, stateArray_S32reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S32reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_2438, stateArray_inS32ser[6]}), .a ({ciphertext_s1[22], ciphertext_s0[22]}), .c ({new_AGEMA_signal_3244, stateArray_S32reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S32reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_2441, stateArray_inS32ser[7]}), .a ({ciphertext_s1[23], ciphertext_s0[23]}), .c ({new_AGEMA_signal_3245, stateArray_S32reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS00ser_mux_inst_0_U1 ( .s (stateArray_n32), .b ({plaintext_s1[120], plaintext_s0[120]}), .a ({ciphertext_s1[112], ciphertext_s0[112]}), .c ({new_AGEMA_signal_2156, stateArray_inS00ser[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS00ser_mux_inst_1_U1 ( .s (stateArray_n32), .b ({plaintext_s1[121], plaintext_s0[121]}), .a ({ciphertext_s1[113], ciphertext_s0[113]}), .c ({new_AGEMA_signal_2159, stateArray_inS00ser[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS00ser_mux_inst_2_U1 ( .s (stateArray_n32), .b ({plaintext_s1[122], plaintext_s0[122]}), .a ({ciphertext_s1[114], ciphertext_s0[114]}), .c ({new_AGEMA_signal_2162, stateArray_inS00ser[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS00ser_mux_inst_3_U1 ( .s (stateArray_n32), .b ({plaintext_s1[123], plaintext_s0[123]}), .a ({ciphertext_s1[115], ciphertext_s0[115]}), .c ({new_AGEMA_signal_2165, stateArray_inS00ser[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS00ser_mux_inst_4_U1 ( .s (stateArray_n32), .b ({plaintext_s1[124], plaintext_s0[124]}), .a ({ciphertext_s1[116], ciphertext_s0[116]}), .c ({new_AGEMA_signal_2168, stateArray_inS00ser[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS00ser_mux_inst_5_U1 ( .s (stateArray_n32), .b ({plaintext_s1[125], plaintext_s0[125]}), .a ({ciphertext_s1[117], ciphertext_s0[117]}), .c ({new_AGEMA_signal_2171, stateArray_inS00ser[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS00ser_mux_inst_6_U1 ( .s (stateArray_n32), .b ({plaintext_s1[126], plaintext_s0[126]}), .a ({ciphertext_s1[118], ciphertext_s0[118]}), .c ({new_AGEMA_signal_2174, stateArray_inS00ser[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS00ser_mux_inst_7_U1 ( .s (stateArray_n32), .b ({plaintext_s1[127], plaintext_s0[127]}), .a ({ciphertext_s1[119], ciphertext_s0[119]}), .c ({new_AGEMA_signal_2177, stateArray_inS00ser[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS01ser_mux_inst_0_U1 ( .s (stateArray_n32), .b ({plaintext_s1[112], plaintext_s0[112]}), .a ({ciphertext_s1[104], ciphertext_s0[104]}), .c ({new_AGEMA_signal_2180, stateArray_inS01ser[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS01ser_mux_inst_1_U1 ( .s (stateArray_n32), .b ({plaintext_s1[113], plaintext_s0[113]}), .a ({ciphertext_s1[105], ciphertext_s0[105]}), .c ({new_AGEMA_signal_2183, stateArray_inS01ser[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS01ser_mux_inst_2_U1 ( .s (stateArray_n32), .b ({plaintext_s1[114], plaintext_s0[114]}), .a ({ciphertext_s1[106], ciphertext_s0[106]}), .c ({new_AGEMA_signal_2186, stateArray_inS01ser[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS01ser_mux_inst_3_U1 ( .s (stateArray_n32), .b ({plaintext_s1[115], plaintext_s0[115]}), .a ({ciphertext_s1[107], ciphertext_s0[107]}), .c ({new_AGEMA_signal_2189, stateArray_inS01ser[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS01ser_mux_inst_4_U1 ( .s (stateArray_n32), .b ({plaintext_s1[116], plaintext_s0[116]}), .a ({ciphertext_s1[108], ciphertext_s0[108]}), .c ({new_AGEMA_signal_2192, stateArray_inS01ser[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS01ser_mux_inst_5_U1 ( .s (stateArray_n32), .b ({plaintext_s1[117], plaintext_s0[117]}), .a ({ciphertext_s1[109], ciphertext_s0[109]}), .c ({new_AGEMA_signal_2195, stateArray_inS01ser[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS01ser_mux_inst_6_U1 ( .s (stateArray_n32), .b ({plaintext_s1[118], plaintext_s0[118]}), .a ({ciphertext_s1[110], ciphertext_s0[110]}), .c ({new_AGEMA_signal_2198, stateArray_inS01ser[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS01ser_mux_inst_7_U1 ( .s (stateArray_n32), .b ({plaintext_s1[119], plaintext_s0[119]}), .a ({ciphertext_s1[111], ciphertext_s0[111]}), .c ({new_AGEMA_signal_2201, stateArray_inS01ser[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS02ser_mux_inst_0_U1 ( .s (stateArray_n31), .b ({plaintext_s1[104], plaintext_s0[104]}), .a ({ciphertext_s1[96], ciphertext_s0[96]}), .c ({new_AGEMA_signal_2204, stateArray_inS02ser[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS02ser_mux_inst_1_U1 ( .s (stateArray_n31), .b ({plaintext_s1[105], plaintext_s0[105]}), .a ({ciphertext_s1[97], ciphertext_s0[97]}), .c ({new_AGEMA_signal_2207, stateArray_inS02ser[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS02ser_mux_inst_2_U1 ( .s (stateArray_n31), .b ({plaintext_s1[106], plaintext_s0[106]}), .a ({ciphertext_s1[98], ciphertext_s0[98]}), .c ({new_AGEMA_signal_2210, stateArray_inS02ser[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS02ser_mux_inst_3_U1 ( .s (stateArray_n31), .b ({plaintext_s1[107], plaintext_s0[107]}), .a ({ciphertext_s1[99], ciphertext_s0[99]}), .c ({new_AGEMA_signal_2213, stateArray_inS02ser[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS02ser_mux_inst_4_U1 ( .s (stateArray_n31), .b ({plaintext_s1[108], plaintext_s0[108]}), .a ({ciphertext_s1[100], ciphertext_s0[100]}), .c ({new_AGEMA_signal_2216, stateArray_inS02ser[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS02ser_mux_inst_5_U1 ( .s (stateArray_n31), .b ({plaintext_s1[109], plaintext_s0[109]}), .a ({ciphertext_s1[101], ciphertext_s0[101]}), .c ({new_AGEMA_signal_2219, stateArray_inS02ser[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS02ser_mux_inst_6_U1 ( .s (stateArray_n31), .b ({plaintext_s1[110], plaintext_s0[110]}), .a ({ciphertext_s1[102], ciphertext_s0[102]}), .c ({new_AGEMA_signal_2222, stateArray_inS02ser[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS02ser_mux_inst_7_U1 ( .s (stateArray_n31), .b ({plaintext_s1[111], plaintext_s0[111]}), .a ({ciphertext_s1[103], ciphertext_s0[103]}), .c ({new_AGEMA_signal_2225, stateArray_inS02ser[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_outS10_MC_mux_inst_0_U1 ( .s (stateArray_n23), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .a ({new_AGEMA_signal_2880, StateInMC[24]}), .c ({new_AGEMA_signal_3008, stateArray_outS10ser_MC[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_outS10_MC_mux_inst_1_U1 ( .s (stateArray_n23), .b ({ciphertext_s1[89], ciphertext_s0[89]}), .a ({new_AGEMA_signal_2881, StateInMC[25]}), .c ({new_AGEMA_signal_3009, stateArray_outS10ser_MC[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_outS10_MC_mux_inst_2_U1 ( .s (stateArray_n23), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .a ({new_AGEMA_signal_2882, StateInMC[26]}), .c ({new_AGEMA_signal_3010, stateArray_outS10ser_MC[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_outS10_MC_mux_inst_3_U1 ( .s (stateArray_n23), .b ({ciphertext_s1[91], ciphertext_s0[91]}), .a ({new_AGEMA_signal_2883, StateInMC[27]}), .c ({new_AGEMA_signal_3011, stateArray_outS10ser_MC[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_outS10_MC_mux_inst_4_U1 ( .s (stateArray_n23), .b ({ciphertext_s1[92], ciphertext_s0[92]}), .a ({new_AGEMA_signal_2884, StateInMC[28]}), .c ({new_AGEMA_signal_3012, stateArray_outS10ser_MC[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_outS10_MC_mux_inst_5_U1 ( .s (stateArray_n23), .b ({ciphertext_s1[93], ciphertext_s0[93]}), .a ({new_AGEMA_signal_2885, StateInMC[29]}), .c ({new_AGEMA_signal_3013, stateArray_outS10ser_MC[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_outS10_MC_mux_inst_6_U1 ( .s (stateArray_n23), .b ({ciphertext_s1[94], ciphertext_s0[94]}), .a ({new_AGEMA_signal_2886, StateInMC[30]}), .c ({new_AGEMA_signal_3014, stateArray_outS10ser_MC[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_outS10_MC_mux_inst_7_U1 ( .s (stateArray_n23), .b ({ciphertext_s1[95], ciphertext_s0[95]}), .a ({new_AGEMA_signal_2887, StateInMC[31]}), .c ({new_AGEMA_signal_3015, stateArray_outS10ser_MC[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS03ser_mux_inst_0_U1 ( .s (stateArray_n31), .b ({plaintext_s1[96], plaintext_s0[96]}), .a ({new_AGEMA_signal_3008, stateArray_outS10ser_MC[0]}), .c ({new_AGEMA_signal_3046, stateArray_inS03ser[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS03ser_mux_inst_1_U1 ( .s (stateArray_n31), .b ({plaintext_s1[97], plaintext_s0[97]}), .a ({new_AGEMA_signal_3009, stateArray_outS10ser_MC[1]}), .c ({new_AGEMA_signal_3048, stateArray_inS03ser[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS03ser_mux_inst_2_U1 ( .s (stateArray_n31), .b ({plaintext_s1[98], plaintext_s0[98]}), .a ({new_AGEMA_signal_3010, stateArray_outS10ser_MC[2]}), .c ({new_AGEMA_signal_3050, stateArray_inS03ser[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS03ser_mux_inst_3_U1 ( .s (stateArray_n31), .b ({plaintext_s1[99], plaintext_s0[99]}), .a ({new_AGEMA_signal_3011, stateArray_outS10ser_MC[3]}), .c ({new_AGEMA_signal_3052, stateArray_inS03ser[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS03ser_mux_inst_4_U1 ( .s (stateArray_n31), .b ({plaintext_s1[100], plaintext_s0[100]}), .a ({new_AGEMA_signal_3012, stateArray_outS10ser_MC[4]}), .c ({new_AGEMA_signal_3054, stateArray_inS03ser[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS03ser_mux_inst_5_U1 ( .s (stateArray_n31), .b ({plaintext_s1[101], plaintext_s0[101]}), .a ({new_AGEMA_signal_3013, stateArray_outS10ser_MC[5]}), .c ({new_AGEMA_signal_3056, stateArray_inS03ser[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS03ser_mux_inst_6_U1 ( .s (stateArray_n31), .b ({plaintext_s1[102], plaintext_s0[102]}), .a ({new_AGEMA_signal_3014, stateArray_outS10ser_MC[6]}), .c ({new_AGEMA_signal_3058, stateArray_inS03ser[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS03ser_mux_inst_7_U1 ( .s (stateArray_n31), .b ({plaintext_s1[103], plaintext_s0[103]}), .a ({new_AGEMA_signal_3015, stateArray_outS10ser_MC[7]}), .c ({new_AGEMA_signal_3060, stateArray_inS03ser[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS10ser_mux_inst_0_U1 ( .s (stateArray_n30), .b ({plaintext_s1[88], plaintext_s0[88]}), .a ({ciphertext_s1[80], ciphertext_s0[80]}), .c ({new_AGEMA_signal_2228, stateArray_inS10ser[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS10ser_mux_inst_1_U1 ( .s (stateArray_n30), .b ({plaintext_s1[89], plaintext_s0[89]}), .a ({ciphertext_s1[81], ciphertext_s0[81]}), .c ({new_AGEMA_signal_2231, stateArray_inS10ser[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS10ser_mux_inst_2_U1 ( .s (stateArray_n30), .b ({plaintext_s1[90], plaintext_s0[90]}), .a ({ciphertext_s1[82], ciphertext_s0[82]}), .c ({new_AGEMA_signal_2234, stateArray_inS10ser[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS10ser_mux_inst_3_U1 ( .s (stateArray_n30), .b ({plaintext_s1[91], plaintext_s0[91]}), .a ({ciphertext_s1[83], ciphertext_s0[83]}), .c ({new_AGEMA_signal_2237, stateArray_inS10ser[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS10ser_mux_inst_4_U1 ( .s (stateArray_n30), .b ({plaintext_s1[92], plaintext_s0[92]}), .a ({ciphertext_s1[84], ciphertext_s0[84]}), .c ({new_AGEMA_signal_2240, stateArray_inS10ser[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS10ser_mux_inst_5_U1 ( .s (stateArray_n30), .b ({plaintext_s1[93], plaintext_s0[93]}), .a ({ciphertext_s1[85], ciphertext_s0[85]}), .c ({new_AGEMA_signal_2243, stateArray_inS10ser[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS10ser_mux_inst_6_U1 ( .s (stateArray_n30), .b ({plaintext_s1[94], plaintext_s0[94]}), .a ({ciphertext_s1[86], ciphertext_s0[86]}), .c ({new_AGEMA_signal_2246, stateArray_inS10ser[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS10ser_mux_inst_7_U1 ( .s (stateArray_n30), .b ({plaintext_s1[95], plaintext_s0[95]}), .a ({ciphertext_s1[87], ciphertext_s0[87]}), .c ({new_AGEMA_signal_2249, stateArray_inS10ser[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS11ser_mux_inst_0_U1 ( .s (stateArray_n30), .b ({plaintext_s1[80], plaintext_s0[80]}), .a ({ciphertext_s1[72], ciphertext_s0[72]}), .c ({new_AGEMA_signal_2252, stateArray_inS11ser[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS11ser_mux_inst_1_U1 ( .s (stateArray_n30), .b ({plaintext_s1[81], plaintext_s0[81]}), .a ({ciphertext_s1[73], ciphertext_s0[73]}), .c ({new_AGEMA_signal_2255, stateArray_inS11ser[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS11ser_mux_inst_2_U1 ( .s (stateArray_n30), .b ({plaintext_s1[82], plaintext_s0[82]}), .a ({ciphertext_s1[74], ciphertext_s0[74]}), .c ({new_AGEMA_signal_2258, stateArray_inS11ser[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS11ser_mux_inst_3_U1 ( .s (stateArray_n30), .b ({plaintext_s1[83], plaintext_s0[83]}), .a ({ciphertext_s1[75], ciphertext_s0[75]}), .c ({new_AGEMA_signal_2261, stateArray_inS11ser[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS11ser_mux_inst_4_U1 ( .s (stateArray_n30), .b ({plaintext_s1[84], plaintext_s0[84]}), .a ({ciphertext_s1[76], ciphertext_s0[76]}), .c ({new_AGEMA_signal_2264, stateArray_inS11ser[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS11ser_mux_inst_5_U1 ( .s (stateArray_n30), .b ({plaintext_s1[85], plaintext_s0[85]}), .a ({ciphertext_s1[77], ciphertext_s0[77]}), .c ({new_AGEMA_signal_2267, stateArray_inS11ser[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS11ser_mux_inst_6_U1 ( .s (stateArray_n30), .b ({plaintext_s1[86], plaintext_s0[86]}), .a ({ciphertext_s1[78], ciphertext_s0[78]}), .c ({new_AGEMA_signal_2270, stateArray_inS11ser[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS11ser_mux_inst_7_U1 ( .s (stateArray_n30), .b ({plaintext_s1[87], plaintext_s0[87]}), .a ({ciphertext_s1[79], ciphertext_s0[79]}), .c ({new_AGEMA_signal_2273, stateArray_inS11ser[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS12ser_mux_inst_0_U1 ( .s (stateArray_n29), .b ({plaintext_s1[72], plaintext_s0[72]}), .a ({ciphertext_s1[64], ciphertext_s0[64]}), .c ({new_AGEMA_signal_2276, stateArray_inS12ser[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS12ser_mux_inst_1_U1 ( .s (stateArray_n29), .b ({plaintext_s1[73], plaintext_s0[73]}), .a ({ciphertext_s1[65], ciphertext_s0[65]}), .c ({new_AGEMA_signal_2279, stateArray_inS12ser[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS12ser_mux_inst_2_U1 ( .s (stateArray_n29), .b ({plaintext_s1[74], plaintext_s0[74]}), .a ({ciphertext_s1[66], ciphertext_s0[66]}), .c ({new_AGEMA_signal_2282, stateArray_inS12ser[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS12ser_mux_inst_3_U1 ( .s (stateArray_n29), .b ({plaintext_s1[75], plaintext_s0[75]}), .a ({ciphertext_s1[67], ciphertext_s0[67]}), .c ({new_AGEMA_signal_2285, stateArray_inS12ser[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS12ser_mux_inst_4_U1 ( .s (stateArray_n29), .b ({plaintext_s1[76], plaintext_s0[76]}), .a ({ciphertext_s1[68], ciphertext_s0[68]}), .c ({new_AGEMA_signal_2288, stateArray_inS12ser[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS12ser_mux_inst_5_U1 ( .s (stateArray_n29), .b ({plaintext_s1[77], plaintext_s0[77]}), .a ({ciphertext_s1[69], ciphertext_s0[69]}), .c ({new_AGEMA_signal_2291, stateArray_inS12ser[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS12ser_mux_inst_6_U1 ( .s (stateArray_n29), .b ({plaintext_s1[78], plaintext_s0[78]}), .a ({ciphertext_s1[70], ciphertext_s0[70]}), .c ({new_AGEMA_signal_2294, stateArray_inS12ser[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS12ser_mux_inst_7_U1 ( .s (stateArray_n29), .b ({plaintext_s1[79], plaintext_s0[79]}), .a ({ciphertext_s1[71], ciphertext_s0[71]}), .c ({new_AGEMA_signal_2297, stateArray_inS12ser[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_outS20_MC_mux_inst_0_U1 ( .s (stateArray_n23), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .a ({new_AGEMA_signal_2872, StateInMC[16]}), .c ({new_AGEMA_signal_3016, stateArray_outS20ser_MC[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_outS20_MC_mux_inst_1_U1 ( .s (stateArray_n23), .b ({ciphertext_s1[57], ciphertext_s0[57]}), .a ({new_AGEMA_signal_2873, StateInMC[17]}), .c ({new_AGEMA_signal_3017, stateArray_outS20ser_MC[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_outS20_MC_mux_inst_2_U1 ( .s (stateArray_n23), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .a ({new_AGEMA_signal_2874, StateInMC[18]}), .c ({new_AGEMA_signal_3018, stateArray_outS20ser_MC[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_outS20_MC_mux_inst_3_U1 ( .s (stateArray_n23), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .a ({new_AGEMA_signal_2875, StateInMC[19]}), .c ({new_AGEMA_signal_3019, stateArray_outS20ser_MC[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_outS20_MC_mux_inst_4_U1 ( .s (stateArray_n23), .b ({ciphertext_s1[60], ciphertext_s0[60]}), .a ({new_AGEMA_signal_2876, StateInMC[20]}), .c ({new_AGEMA_signal_3020, stateArray_outS20ser_MC[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_outS20_MC_mux_inst_5_U1 ( .s (stateArray_n23), .b ({ciphertext_s1[61], ciphertext_s0[61]}), .a ({new_AGEMA_signal_2877, StateInMC[21]}), .c ({new_AGEMA_signal_3021, stateArray_outS20ser_MC[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_outS20_MC_mux_inst_6_U1 ( .s (stateArray_n23), .b ({ciphertext_s1[62], ciphertext_s0[62]}), .a ({new_AGEMA_signal_2878, StateInMC[22]}), .c ({new_AGEMA_signal_3022, stateArray_outS20ser_MC[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_outS20_MC_mux_inst_7_U1 ( .s (stateArray_n23), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .a ({new_AGEMA_signal_2879, StateInMC[23]}), .c ({new_AGEMA_signal_3023, stateArray_outS20ser_MC[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS13ser_mux_inst_0_U1 ( .s (stateArray_n29), .b ({plaintext_s1[64], plaintext_s0[64]}), .a ({new_AGEMA_signal_3016, stateArray_outS20ser_MC[0]}), .c ({new_AGEMA_signal_3062, stateArray_inS13ser[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS13ser_mux_inst_1_U1 ( .s (stateArray_n29), .b ({plaintext_s1[65], plaintext_s0[65]}), .a ({new_AGEMA_signal_3017, stateArray_outS20ser_MC[1]}), .c ({new_AGEMA_signal_3064, stateArray_inS13ser[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS13ser_mux_inst_2_U1 ( .s (stateArray_n29), .b ({plaintext_s1[66], plaintext_s0[66]}), .a ({new_AGEMA_signal_3018, stateArray_outS20ser_MC[2]}), .c ({new_AGEMA_signal_3066, stateArray_inS13ser[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS13ser_mux_inst_3_U1 ( .s (stateArray_n29), .b ({plaintext_s1[67], plaintext_s0[67]}), .a ({new_AGEMA_signal_3019, stateArray_outS20ser_MC[3]}), .c ({new_AGEMA_signal_3068, stateArray_inS13ser[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS13ser_mux_inst_4_U1 ( .s (stateArray_n29), .b ({plaintext_s1[68], plaintext_s0[68]}), .a ({new_AGEMA_signal_3020, stateArray_outS20ser_MC[4]}), .c ({new_AGEMA_signal_3070, stateArray_inS13ser[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS13ser_mux_inst_5_U1 ( .s (stateArray_n29), .b ({plaintext_s1[69], plaintext_s0[69]}), .a ({new_AGEMA_signal_3021, stateArray_outS20ser_MC[5]}), .c ({new_AGEMA_signal_3072, stateArray_inS13ser[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS13ser_mux_inst_6_U1 ( .s (stateArray_n29), .b ({plaintext_s1[70], plaintext_s0[70]}), .a ({new_AGEMA_signal_3022, stateArray_outS20ser_MC[6]}), .c ({new_AGEMA_signal_3074, stateArray_inS13ser[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS13ser_mux_inst_7_U1 ( .s (stateArray_n29), .b ({plaintext_s1[71], plaintext_s0[71]}), .a ({new_AGEMA_signal_3023, stateArray_outS20ser_MC[7]}), .c ({new_AGEMA_signal_3076, stateArray_inS13ser[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS20ser_mux_inst_0_U1 ( .s (stateArray_n28), .b ({plaintext_s1[56], plaintext_s0[56]}), .a ({ciphertext_s1[48], ciphertext_s0[48]}), .c ({new_AGEMA_signal_2300, stateArray_inS20ser[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS20ser_mux_inst_1_U1 ( .s (stateArray_n28), .b ({plaintext_s1[57], plaintext_s0[57]}), .a ({ciphertext_s1[49], ciphertext_s0[49]}), .c ({new_AGEMA_signal_2303, stateArray_inS20ser[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS20ser_mux_inst_2_U1 ( .s (stateArray_n28), .b ({plaintext_s1[58], plaintext_s0[58]}), .a ({ciphertext_s1[50], ciphertext_s0[50]}), .c ({new_AGEMA_signal_2306, stateArray_inS20ser[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS20ser_mux_inst_3_U1 ( .s (stateArray_n28), .b ({plaintext_s1[59], plaintext_s0[59]}), .a ({ciphertext_s1[51], ciphertext_s0[51]}), .c ({new_AGEMA_signal_2309, stateArray_inS20ser[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS20ser_mux_inst_4_U1 ( .s (stateArray_n28), .b ({plaintext_s1[60], plaintext_s0[60]}), .a ({ciphertext_s1[52], ciphertext_s0[52]}), .c ({new_AGEMA_signal_2312, stateArray_inS20ser[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS20ser_mux_inst_5_U1 ( .s (stateArray_n28), .b ({plaintext_s1[61], plaintext_s0[61]}), .a ({ciphertext_s1[53], ciphertext_s0[53]}), .c ({new_AGEMA_signal_2315, stateArray_inS20ser[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS20ser_mux_inst_6_U1 ( .s (stateArray_n28), .b ({plaintext_s1[62], plaintext_s0[62]}), .a ({ciphertext_s1[54], ciphertext_s0[54]}), .c ({new_AGEMA_signal_2318, stateArray_inS20ser[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS20ser_mux_inst_7_U1 ( .s (stateArray_n28), .b ({plaintext_s1[63], plaintext_s0[63]}), .a ({ciphertext_s1[55], ciphertext_s0[55]}), .c ({new_AGEMA_signal_2321, stateArray_inS20ser[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS21ser_mux_inst_0_U1 ( .s (stateArray_n28), .b ({plaintext_s1[48], plaintext_s0[48]}), .a ({ciphertext_s1[40], ciphertext_s0[40]}), .c ({new_AGEMA_signal_2324, stateArray_inS21ser[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS21ser_mux_inst_1_U1 ( .s (stateArray_n28), .b ({plaintext_s1[49], plaintext_s0[49]}), .a ({ciphertext_s1[41], ciphertext_s0[41]}), .c ({new_AGEMA_signal_2327, stateArray_inS21ser[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS21ser_mux_inst_2_U1 ( .s (stateArray_n28), .b ({plaintext_s1[50], plaintext_s0[50]}), .a ({ciphertext_s1[42], ciphertext_s0[42]}), .c ({new_AGEMA_signal_2330, stateArray_inS21ser[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS21ser_mux_inst_3_U1 ( .s (stateArray_n28), .b ({plaintext_s1[51], plaintext_s0[51]}), .a ({ciphertext_s1[43], ciphertext_s0[43]}), .c ({new_AGEMA_signal_2333, stateArray_inS21ser[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS21ser_mux_inst_4_U1 ( .s (stateArray_n28), .b ({plaintext_s1[52], plaintext_s0[52]}), .a ({ciphertext_s1[44], ciphertext_s0[44]}), .c ({new_AGEMA_signal_2336, stateArray_inS21ser[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS21ser_mux_inst_5_U1 ( .s (stateArray_n28), .b ({plaintext_s1[53], plaintext_s0[53]}), .a ({ciphertext_s1[45], ciphertext_s0[45]}), .c ({new_AGEMA_signal_2339, stateArray_inS21ser[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS21ser_mux_inst_6_U1 ( .s (stateArray_n28), .b ({plaintext_s1[54], plaintext_s0[54]}), .a ({ciphertext_s1[46], ciphertext_s0[46]}), .c ({new_AGEMA_signal_2342, stateArray_inS21ser[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS21ser_mux_inst_7_U1 ( .s (stateArray_n28), .b ({plaintext_s1[55], plaintext_s0[55]}), .a ({ciphertext_s1[47], ciphertext_s0[47]}), .c ({new_AGEMA_signal_2345, stateArray_inS21ser[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS22ser_mux_inst_0_U1 ( .s (stateArray_n27), .b ({plaintext_s1[40], plaintext_s0[40]}), .a ({ciphertext_s1[32], ciphertext_s0[32]}), .c ({new_AGEMA_signal_2348, stateArray_inS22ser[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS22ser_mux_inst_1_U1 ( .s (stateArray_n27), .b ({plaintext_s1[41], plaintext_s0[41]}), .a ({ciphertext_s1[33], ciphertext_s0[33]}), .c ({new_AGEMA_signal_2351, stateArray_inS22ser[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS22ser_mux_inst_2_U1 ( .s (stateArray_n27), .b ({plaintext_s1[42], plaintext_s0[42]}), .a ({ciphertext_s1[34], ciphertext_s0[34]}), .c ({new_AGEMA_signal_2354, stateArray_inS22ser[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS22ser_mux_inst_3_U1 ( .s (stateArray_n27), .b ({plaintext_s1[43], plaintext_s0[43]}), .a ({ciphertext_s1[35], ciphertext_s0[35]}), .c ({new_AGEMA_signal_2357, stateArray_inS22ser[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS22ser_mux_inst_4_U1 ( .s (stateArray_n27), .b ({plaintext_s1[44], plaintext_s0[44]}), .a ({ciphertext_s1[36], ciphertext_s0[36]}), .c ({new_AGEMA_signal_2360, stateArray_inS22ser[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS22ser_mux_inst_5_U1 ( .s (stateArray_n27), .b ({plaintext_s1[45], plaintext_s0[45]}), .a ({ciphertext_s1[37], ciphertext_s0[37]}), .c ({new_AGEMA_signal_2363, stateArray_inS22ser[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS22ser_mux_inst_6_U1 ( .s (stateArray_n27), .b ({plaintext_s1[46], plaintext_s0[46]}), .a ({ciphertext_s1[38], ciphertext_s0[38]}), .c ({new_AGEMA_signal_2366, stateArray_inS22ser[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS22ser_mux_inst_7_U1 ( .s (stateArray_n27), .b ({plaintext_s1[47], plaintext_s0[47]}), .a ({ciphertext_s1[39], ciphertext_s0[39]}), .c ({new_AGEMA_signal_2369, stateArray_inS22ser[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_outS30_MC_mux_inst_0_U1 ( .s (stateArray_n22), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .a ({new_AGEMA_signal_2864, StateInMC[8]}), .c ({new_AGEMA_signal_3024, stateArray_outS30ser_MC[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_outS30_MC_mux_inst_1_U1 ( .s (stateArray_n22), .b ({ciphertext_s1[25], ciphertext_s0[25]}), .a ({new_AGEMA_signal_2865, StateInMC[9]}), .c ({new_AGEMA_signal_3025, stateArray_outS30ser_MC[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_outS30_MC_mux_inst_2_U1 ( .s (stateArray_n22), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .a ({new_AGEMA_signal_2866, StateInMC[10]}), .c ({new_AGEMA_signal_3026, stateArray_outS30ser_MC[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_outS30_MC_mux_inst_3_U1 ( .s (stateArray_n22), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .a ({new_AGEMA_signal_2867, StateInMC[11]}), .c ({new_AGEMA_signal_3027, stateArray_outS30ser_MC[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_outS30_MC_mux_inst_4_U1 ( .s (stateArray_n22), .b ({ciphertext_s1[28], ciphertext_s0[28]}), .a ({new_AGEMA_signal_2868, StateInMC[12]}), .c ({new_AGEMA_signal_3028, stateArray_outS30ser_MC[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_outS30_MC_mux_inst_5_U1 ( .s (stateArray_n22), .b ({ciphertext_s1[29], ciphertext_s0[29]}), .a ({new_AGEMA_signal_2869, StateInMC[13]}), .c ({new_AGEMA_signal_3029, stateArray_outS30ser_MC[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_outS30_MC_mux_inst_6_U1 ( .s (stateArray_n22), .b ({ciphertext_s1[30], ciphertext_s0[30]}), .a ({new_AGEMA_signal_2870, StateInMC[14]}), .c ({new_AGEMA_signal_3030, stateArray_outS30ser_MC[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_outS30_MC_mux_inst_7_U1 ( .s (stateArray_n22), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .a ({new_AGEMA_signal_2871, StateInMC[15]}), .c ({new_AGEMA_signal_3031, stateArray_outS30ser_MC[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS23ser_mux_inst_0_U1 ( .s (stateArray_n27), .b ({plaintext_s1[32], plaintext_s0[32]}), .a ({new_AGEMA_signal_3024, stateArray_outS30ser_MC[0]}), .c ({new_AGEMA_signal_3078, stateArray_inS23ser[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS23ser_mux_inst_1_U1 ( .s (stateArray_n27), .b ({plaintext_s1[33], plaintext_s0[33]}), .a ({new_AGEMA_signal_3025, stateArray_outS30ser_MC[1]}), .c ({new_AGEMA_signal_3080, stateArray_inS23ser[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS23ser_mux_inst_2_U1 ( .s (stateArray_n27), .b ({plaintext_s1[34], plaintext_s0[34]}), .a ({new_AGEMA_signal_3026, stateArray_outS30ser_MC[2]}), .c ({new_AGEMA_signal_3082, stateArray_inS23ser[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS23ser_mux_inst_3_U1 ( .s (stateArray_n27), .b ({plaintext_s1[35], plaintext_s0[35]}), .a ({new_AGEMA_signal_3027, stateArray_outS30ser_MC[3]}), .c ({new_AGEMA_signal_3084, stateArray_inS23ser[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS23ser_mux_inst_4_U1 ( .s (stateArray_n27), .b ({plaintext_s1[36], plaintext_s0[36]}), .a ({new_AGEMA_signal_3028, stateArray_outS30ser_MC[4]}), .c ({new_AGEMA_signal_3086, stateArray_inS23ser[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS23ser_mux_inst_5_U1 ( .s (stateArray_n27), .b ({plaintext_s1[37], plaintext_s0[37]}), .a ({new_AGEMA_signal_3029, stateArray_outS30ser_MC[5]}), .c ({new_AGEMA_signal_3088, stateArray_inS23ser[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS23ser_mux_inst_6_U1 ( .s (stateArray_n27), .b ({plaintext_s1[38], plaintext_s0[38]}), .a ({new_AGEMA_signal_3030, stateArray_outS30ser_MC[6]}), .c ({new_AGEMA_signal_3090, stateArray_inS23ser[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS23ser_mux_inst_7_U1 ( .s (stateArray_n27), .b ({plaintext_s1[39], plaintext_s0[39]}), .a ({new_AGEMA_signal_3031, stateArray_outS30ser_MC[7]}), .c ({new_AGEMA_signal_3092, stateArray_inS23ser[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS30ser_mux_inst_0_U1 ( .s (stateArray_n26), .b ({plaintext_s1[24], plaintext_s0[24]}), .a ({ciphertext_s1[16], ciphertext_s0[16]}), .c ({new_AGEMA_signal_2372, stateArray_inS30ser[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS30ser_mux_inst_1_U1 ( .s (stateArray_n26), .b ({plaintext_s1[25], plaintext_s0[25]}), .a ({ciphertext_s1[17], ciphertext_s0[17]}), .c ({new_AGEMA_signal_2375, stateArray_inS30ser[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS30ser_mux_inst_2_U1 ( .s (stateArray_n26), .b ({plaintext_s1[26], plaintext_s0[26]}), .a ({ciphertext_s1[18], ciphertext_s0[18]}), .c ({new_AGEMA_signal_2378, stateArray_inS30ser[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS30ser_mux_inst_3_U1 ( .s (stateArray_n26), .b ({plaintext_s1[27], plaintext_s0[27]}), .a ({ciphertext_s1[19], ciphertext_s0[19]}), .c ({new_AGEMA_signal_2381, stateArray_inS30ser[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS30ser_mux_inst_4_U1 ( .s (stateArray_n26), .b ({plaintext_s1[28], plaintext_s0[28]}), .a ({ciphertext_s1[20], ciphertext_s0[20]}), .c ({new_AGEMA_signal_2384, stateArray_inS30ser[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS30ser_mux_inst_5_U1 ( .s (stateArray_n26), .b ({plaintext_s1[29], plaintext_s0[29]}), .a ({ciphertext_s1[21], ciphertext_s0[21]}), .c ({new_AGEMA_signal_2387, stateArray_inS30ser[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS30ser_mux_inst_6_U1 ( .s (stateArray_n26), .b ({plaintext_s1[30], plaintext_s0[30]}), .a ({ciphertext_s1[22], ciphertext_s0[22]}), .c ({new_AGEMA_signal_2390, stateArray_inS30ser[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS30ser_mux_inst_7_U1 ( .s (stateArray_n26), .b ({plaintext_s1[31], plaintext_s0[31]}), .a ({ciphertext_s1[23], ciphertext_s0[23]}), .c ({new_AGEMA_signal_2393, stateArray_inS30ser[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS31ser_mux_inst_0_U1 ( .s (stateArray_n26), .b ({plaintext_s1[16], plaintext_s0[16]}), .a ({ciphertext_s1[8], ciphertext_s0[8]}), .c ({new_AGEMA_signal_2396, stateArray_inS31ser[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS31ser_mux_inst_1_U1 ( .s (stateArray_n26), .b ({plaintext_s1[17], plaintext_s0[17]}), .a ({ciphertext_s1[9], ciphertext_s0[9]}), .c ({new_AGEMA_signal_2399, stateArray_inS31ser[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS31ser_mux_inst_2_U1 ( .s (stateArray_n26), .b ({plaintext_s1[18], plaintext_s0[18]}), .a ({ciphertext_s1[10], ciphertext_s0[10]}), .c ({new_AGEMA_signal_2402, stateArray_inS31ser[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS31ser_mux_inst_3_U1 ( .s (stateArray_n26), .b ({plaintext_s1[19], plaintext_s0[19]}), .a ({ciphertext_s1[11], ciphertext_s0[11]}), .c ({new_AGEMA_signal_2405, stateArray_inS31ser[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS31ser_mux_inst_4_U1 ( .s (stateArray_n26), .b ({plaintext_s1[20], plaintext_s0[20]}), .a ({ciphertext_s1[12], ciphertext_s0[12]}), .c ({new_AGEMA_signal_2408, stateArray_inS31ser[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS31ser_mux_inst_5_U1 ( .s (stateArray_n26), .b ({plaintext_s1[21], plaintext_s0[21]}), .a ({ciphertext_s1[13], ciphertext_s0[13]}), .c ({new_AGEMA_signal_2411, stateArray_inS31ser[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS31ser_mux_inst_6_U1 ( .s (stateArray_n26), .b ({plaintext_s1[22], plaintext_s0[22]}), .a ({ciphertext_s1[14], ciphertext_s0[14]}), .c ({new_AGEMA_signal_2414, stateArray_inS31ser[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS31ser_mux_inst_7_U1 ( .s (stateArray_n26), .b ({plaintext_s1[23], plaintext_s0[23]}), .a ({ciphertext_s1[15], ciphertext_s0[15]}), .c ({new_AGEMA_signal_2417, stateArray_inS31ser[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS32ser_mux_inst_0_U1 ( .s (stateArray_n25), .b ({plaintext_s1[8], plaintext_s0[8]}), .a ({ciphertext_s1[0], ciphertext_s0[0]}), .c ({new_AGEMA_signal_2420, stateArray_inS32ser[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS32ser_mux_inst_1_U1 ( .s (stateArray_n25), .b ({plaintext_s1[9], plaintext_s0[9]}), .a ({ciphertext_s1[1], ciphertext_s0[1]}), .c ({new_AGEMA_signal_2423, stateArray_inS32ser[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS32ser_mux_inst_2_U1 ( .s (stateArray_n25), .b ({plaintext_s1[10], plaintext_s0[10]}), .a ({ciphertext_s1[2], ciphertext_s0[2]}), .c ({new_AGEMA_signal_2426, stateArray_inS32ser[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS32ser_mux_inst_3_U1 ( .s (stateArray_n25), .b ({plaintext_s1[11], plaintext_s0[11]}), .a ({ciphertext_s1[3], ciphertext_s0[3]}), .c ({new_AGEMA_signal_2429, stateArray_inS32ser[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS32ser_mux_inst_4_U1 ( .s (stateArray_n25), .b ({plaintext_s1[12], plaintext_s0[12]}), .a ({ciphertext_s1[4], ciphertext_s0[4]}), .c ({new_AGEMA_signal_2432, stateArray_inS32ser[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS32ser_mux_inst_5_U1 ( .s (stateArray_n25), .b ({plaintext_s1[13], plaintext_s0[13]}), .a ({ciphertext_s1[5], ciphertext_s0[5]}), .c ({new_AGEMA_signal_2435, stateArray_inS32ser[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS32ser_mux_inst_6_U1 ( .s (stateArray_n25), .b ({plaintext_s1[14], plaintext_s0[14]}), .a ({ciphertext_s1[6], ciphertext_s0[6]}), .c ({new_AGEMA_signal_2438, stateArray_inS32ser[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS32ser_mux_inst_7_U1 ( .s (stateArray_n25), .b ({plaintext_s1[15], plaintext_s0[15]}), .a ({ciphertext_s1[7], ciphertext_s0[7]}), .c ({new_AGEMA_signal_2441, stateArray_inS32ser[7]}) ) ;
    INV_X1 MUX_StateInMC_U3 ( .A (intFinal), .ZN (MUX_StateInMC_n7) ) ;
    INV_X1 MUX_StateInMC_U2 ( .A (MUX_StateInMC_n7), .ZN (MUX_StateInMC_n6) ) ;
    INV_X1 MUX_StateInMC_U1 ( .A (MUX_StateInMC_n7), .ZN (MUX_StateInMC_n5) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateInMC_mux_inst_0_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_2825, MCout[0]}), .a ({ciphertext_s1[24], ciphertext_s0[24]}), .c ({new_AGEMA_signal_2860, StateInMC[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateInMC_mux_inst_1_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_2849, MCout[1]}), .a ({ciphertext_s1[25], ciphertext_s0[25]}), .c ({new_AGEMA_signal_2861, StateInMC[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateInMC_mux_inst_2_U1 ( .s (intFinal), .b ({new_AGEMA_signal_2823, MCout[2]}), .a ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_2834, StateInMC[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateInMC_mux_inst_3_U1 ( .s (intFinal), .b ({new_AGEMA_signal_2848, MCout[3]}), .a ({ciphertext_s1[27], ciphertext_s0[27]}), .c ({new_AGEMA_signal_2862, StateInMC[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateInMC_mux_inst_4_U1 ( .s (intFinal), .b ({new_AGEMA_signal_2847, MCout[4]}), .a ({ciphertext_s1[28], ciphertext_s0[28]}), .c ({new_AGEMA_signal_2863, StateInMC[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateInMC_mux_inst_5_U1 ( .s (intFinal), .b ({new_AGEMA_signal_2820, MCout[5]}), .a ({ciphertext_s1[29], ciphertext_s0[29]}), .c ({new_AGEMA_signal_2835, StateInMC[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateInMC_mux_inst_6_U1 ( .s (intFinal), .b ({new_AGEMA_signal_2819, MCout[6]}), .a ({ciphertext_s1[30], ciphertext_s0[30]}), .c ({new_AGEMA_signal_2836, StateInMC[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateInMC_mux_inst_7_U1 ( .s (intFinal), .b ({new_AGEMA_signal_2818, MCout[7]}), .a ({ciphertext_s1[31], ciphertext_s0[31]}), .c ({new_AGEMA_signal_2837, StateInMC[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateInMC_mux_inst_8_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_2817, MCout[8]}), .a ({ciphertext_s1[56], ciphertext_s0[56]}), .c ({new_AGEMA_signal_2864, StateInMC[8]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateInMC_mux_inst_9_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_2846, MCout[9]}), .a ({ciphertext_s1[57], ciphertext_s0[57]}), .c ({new_AGEMA_signal_2865, StateInMC[9]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateInMC_mux_inst_10_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_2815, MCout[10]}), .a ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_2866, StateInMC[10]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateInMC_mux_inst_11_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_2845, MCout[11]}), .a ({ciphertext_s1[59], ciphertext_s0[59]}), .c ({new_AGEMA_signal_2867, StateInMC[11]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateInMC_mux_inst_12_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_2844, MCout[12]}), .a ({ciphertext_s1[60], ciphertext_s0[60]}), .c ({new_AGEMA_signal_2868, StateInMC[12]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateInMC_mux_inst_13_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_2812, MCout[13]}), .a ({ciphertext_s1[61], ciphertext_s0[61]}), .c ({new_AGEMA_signal_2869, StateInMC[13]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateInMC_mux_inst_14_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_2811, MCout[14]}), .a ({ciphertext_s1[62], ciphertext_s0[62]}), .c ({new_AGEMA_signal_2870, StateInMC[14]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateInMC_mux_inst_15_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_2810, MCout[15]}), .a ({ciphertext_s1[63], ciphertext_s0[63]}), .c ({new_AGEMA_signal_2871, StateInMC[15]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateInMC_mux_inst_16_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_2809, MCout[16]}), .a ({ciphertext_s1[88], ciphertext_s0[88]}), .c ({new_AGEMA_signal_2872, StateInMC[16]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateInMC_mux_inst_17_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_2843, MCout[17]}), .a ({ciphertext_s1[89], ciphertext_s0[89]}), .c ({new_AGEMA_signal_2873, StateInMC[17]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateInMC_mux_inst_18_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_2807, MCout[18]}), .a ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_2874, StateInMC[18]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateInMC_mux_inst_19_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_2842, MCout[19]}), .a ({ciphertext_s1[91], ciphertext_s0[91]}), .c ({new_AGEMA_signal_2875, StateInMC[19]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateInMC_mux_inst_20_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_2841, MCout[20]}), .a ({ciphertext_s1[92], ciphertext_s0[92]}), .c ({new_AGEMA_signal_2876, StateInMC[20]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateInMC_mux_inst_21_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_2804, MCout[21]}), .a ({ciphertext_s1[93], ciphertext_s0[93]}), .c ({new_AGEMA_signal_2877, StateInMC[21]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateInMC_mux_inst_22_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_2803, MCout[22]}), .a ({ciphertext_s1[94], ciphertext_s0[94]}), .c ({new_AGEMA_signal_2878, StateInMC[22]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateInMC_mux_inst_23_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_2802, MCout[23]}), .a ({ciphertext_s1[95], ciphertext_s0[95]}), .c ({new_AGEMA_signal_2879, StateInMC[23]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateInMC_mux_inst_24_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_2801, MCout[24]}), .a ({ciphertext_s1[120], ciphertext_s0[120]}), .c ({new_AGEMA_signal_2880, StateInMC[24]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateInMC_mux_inst_25_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_2840, MCout[25]}), .a ({ciphertext_s1[121], ciphertext_s0[121]}), .c ({new_AGEMA_signal_2881, StateInMC[25]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateInMC_mux_inst_26_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_2799, MCout[26]}), .a ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_2882, StateInMC[26]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateInMC_mux_inst_27_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_2839, MCout[27]}), .a ({ciphertext_s1[123], ciphertext_s0[123]}), .c ({new_AGEMA_signal_2883, StateInMC[27]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateInMC_mux_inst_28_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_2838, MCout[28]}), .a ({ciphertext_s1[124], ciphertext_s0[124]}), .c ({new_AGEMA_signal_2884, StateInMC[28]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateInMC_mux_inst_29_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_2796, MCout[29]}), .a ({ciphertext_s1[125], ciphertext_s0[125]}), .c ({new_AGEMA_signal_2885, StateInMC[29]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateInMC_mux_inst_30_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_2795, MCout[30]}), .a ({ciphertext_s1[126], ciphertext_s0[126]}), .c ({new_AGEMA_signal_2886, StateInMC[30]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateInMC_mux_inst_31_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_2794, MCout[31]}), .a ({ciphertext_s1[127], ciphertext_s0[127]}), .c ({new_AGEMA_signal_2887, StateInMC[31]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) KeyArray_U50 ( .a ({new_AGEMA_signal_2006, KeyArray_outS01ser_7_}), .b ({new_AGEMA_signal_2004, keyStateIn[7]}), .c ({new_AGEMA_signal_2007, KeyArray_outS01ser_XOR_00[7]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) KeyArray_U49 ( .a ({new_AGEMA_signal_2008, KeyArray_outS01ser_6_}), .b ({new_AGEMA_signal_2001, keyStateIn[6]}), .c ({new_AGEMA_signal_2009, KeyArray_outS01ser_XOR_00[6]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) KeyArray_U48 ( .a ({new_AGEMA_signal_2010, KeyArray_outS01ser_5_}), .b ({new_AGEMA_signal_1998, keyStateIn[5]}), .c ({new_AGEMA_signal_2011, KeyArray_outS01ser_XOR_00[5]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) KeyArray_U47 ( .a ({new_AGEMA_signal_2012, KeyArray_outS01ser_4_}), .b ({new_AGEMA_signal_1995, keyStateIn[4]}), .c ({new_AGEMA_signal_2013, KeyArray_outS01ser_XOR_00[4]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) KeyArray_U46 ( .a ({new_AGEMA_signal_2014, KeyArray_outS01ser_3_}), .b ({new_AGEMA_signal_1992, keyStateIn[3]}), .c ({new_AGEMA_signal_2015, KeyArray_outS01ser_XOR_00[3]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) KeyArray_U45 ( .a ({new_AGEMA_signal_2016, KeyArray_outS01ser_2_}), .b ({new_AGEMA_signal_1989, keyStateIn[2]}), .c ({new_AGEMA_signal_2017, KeyArray_outS01ser_XOR_00[2]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) KeyArray_U44 ( .a ({new_AGEMA_signal_2018, KeyArray_outS01ser_1_}), .b ({new_AGEMA_signal_1986, keyStateIn[1]}), .c ({new_AGEMA_signal_2019, KeyArray_outS01ser_XOR_00[1]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) KeyArray_U43 ( .a ({new_AGEMA_signal_2020, KeyArray_outS01ser_0_}), .b ({new_AGEMA_signal_1983, keyStateIn[0]}), .c ({new_AGEMA_signal_2021, KeyArray_outS01ser_XOR_00[0]}) ) ;
    INV_X1 KeyArray_U26 ( .A (KeyArray_n47), .ZN (KeyArray_n46) ) ;
    INV_X1 KeyArray_U25 ( .A (KeyArray_n47), .ZN (KeyArray_n45) ) ;
    INV_X1 KeyArray_U24 ( .A (KeyArray_n47), .ZN (KeyArray_n44) ) ;
    INV_X1 KeyArray_U23 ( .A (KeyArray_n47), .ZN (KeyArray_n43) ) ;
    INV_X1 KeyArray_U22 ( .A (KeyArray_n47), .ZN (KeyArray_n42) ) ;
    INV_X1 KeyArray_U21 ( .A (KeyArray_n47), .ZN (KeyArray_n41) ) ;
    INV_X1 KeyArray_U20 ( .A (KeyArray_n47), .ZN (KeyArray_n40) ) ;
    INV_X1 KeyArray_U19 ( .A (KeyArray_n47), .ZN (KeyArray_n39) ) ;
    INV_X1 KeyArray_U18 ( .A (nReset), .ZN (KeyArray_n47) ) ;
    INV_X1 KeyArray_U17 ( .A (KeyArray_n38), .ZN (KeyArray_n31) ) ;
    INV_X1 KeyArray_U16 ( .A (KeyArray_n29), .ZN (KeyArray_n23) ) ;
    INV_X1 KeyArray_U15 ( .A (KeyArray_n38), .ZN (KeyArray_n37) ) ;
    INV_X1 KeyArray_U14 ( .A (KeyArray_n29), .ZN (KeyArray_n28) ) ;
    INV_X1 KeyArray_U13 ( .A (KeyArray_n38), .ZN (KeyArray_n36) ) ;
    INV_X1 KeyArray_U12 ( .A (KeyArray_n29), .ZN (KeyArray_n27) ) ;
    INV_X1 KeyArray_U11 ( .A (KeyArray_n38), .ZN (KeyArray_n35) ) ;
    INV_X1 KeyArray_U10 ( .A (KeyArray_n29), .ZN (KeyArray_n26) ) ;
    INV_X1 KeyArray_U9 ( .A (KeyArray_n38), .ZN (KeyArray_n32) ) ;
    INV_X1 KeyArray_U8 ( .A (KeyArray_n29), .ZN (KeyArray_n24) ) ;
    INV_X1 KeyArray_U7 ( .A (KeyArray_n38), .ZN (KeyArray_n33) ) ;
    INV_X1 KeyArray_U6 ( .A (KeyArray_n29), .ZN (KeyArray_n25) ) ;
    INV_X1 KeyArray_U5 ( .A (KeyArray_n38), .ZN (KeyArray_n30) ) ;
    INV_X1 KeyArray_U4 ( .A (KeyArray_n29), .ZN (KeyArray_n22) ) ;
    INV_X1 KeyArray_U3 ( .A (KeyArray_n38), .ZN (KeyArray_n34) ) ;
    INV_X1 KeyArray_U2 ( .A (selMC), .ZN (KeyArray_n38) ) ;
    INV_X1 KeyArray_U1 ( .A (n12), .ZN (KeyArray_n29) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S00reg_gff_1_SFF_0_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_1983, keyStateIn[0]}), .a ({new_AGEMA_signal_3267, KeyArray_S00reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_3375, KeyArray_S00reg_gff_1_SFF_0_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_3247, KeyArray_inS00ser[0]}), .a ({new_AGEMA_signal_2491, KeyArray_outS10ser[0]}), .c ({new_AGEMA_signal_3267, KeyArray_S00reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S00reg_gff_1_SFF_1_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_1986, keyStateIn[1]}), .a ({new_AGEMA_signal_3268, KeyArray_S00reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_3376, KeyArray_S00reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_3249, KeyArray_inS00ser[1]}), .a ({new_AGEMA_signal_2494, KeyArray_outS10ser[1]}), .c ({new_AGEMA_signal_3268, KeyArray_S00reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S00reg_gff_1_SFF_2_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_1989, keyStateIn[2]}), .a ({new_AGEMA_signal_3269, KeyArray_S00reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_3377, KeyArray_S00reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_3251, KeyArray_inS00ser[2]}), .a ({new_AGEMA_signal_2497, KeyArray_outS10ser[2]}), .c ({new_AGEMA_signal_3269, KeyArray_S00reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S00reg_gff_1_SFF_3_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_1992, keyStateIn[3]}), .a ({new_AGEMA_signal_3270, KeyArray_S00reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_3378, KeyArray_S00reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_3253, KeyArray_inS00ser[3]}), .a ({new_AGEMA_signal_2500, KeyArray_outS10ser[3]}), .c ({new_AGEMA_signal_3270, KeyArray_S00reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S00reg_gff_1_SFF_4_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_1995, keyStateIn[4]}), .a ({new_AGEMA_signal_3271, KeyArray_S00reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_3379, KeyArray_S00reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_3255, KeyArray_inS00ser[4]}), .a ({new_AGEMA_signal_2503, KeyArray_outS10ser[4]}), .c ({new_AGEMA_signal_3271, KeyArray_S00reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S00reg_gff_1_SFF_5_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_1998, keyStateIn[5]}), .a ({new_AGEMA_signal_3272, KeyArray_S00reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_3380, KeyArray_S00reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_3257, KeyArray_inS00ser[5]}), .a ({new_AGEMA_signal_2506, KeyArray_outS10ser[5]}), .c ({new_AGEMA_signal_3272, KeyArray_S00reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S00reg_gff_1_SFF_6_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2001, keyStateIn[6]}), .a ({new_AGEMA_signal_3273, KeyArray_S00reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_3381, KeyArray_S00reg_gff_1_SFF_6_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_3259, KeyArray_inS00ser[6]}), .a ({new_AGEMA_signal_2509, KeyArray_outS10ser[6]}), .c ({new_AGEMA_signal_3273, KeyArray_S00reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S00reg_gff_1_SFF_7_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2004, keyStateIn[7]}), .a ({new_AGEMA_signal_3274, KeyArray_S00reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_3382, KeyArray_S00reg_gff_1_SFF_7_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_3261, KeyArray_inS00ser[7]}), .a ({new_AGEMA_signal_2512, KeyArray_outS10ser[7]}), .c ({new_AGEMA_signal_3274, KeyArray_S00reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S01reg_gff_1_SFF_0_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2020, KeyArray_outS01ser_0_}), .a ({new_AGEMA_signal_2888, KeyArray_S01reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_3275, KeyArray_S01reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_2444, KeyArray_inS01ser[0]}), .a ({new_AGEMA_signal_2515, KeyArray_outS11ser[0]}), .c ({new_AGEMA_signal_2888, KeyArray_S01reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S01reg_gff_1_SFF_1_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2018, KeyArray_outS01ser_1_}), .a ({new_AGEMA_signal_2889, KeyArray_S01reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_3276, KeyArray_S01reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_2447, KeyArray_inS01ser[1]}), .a ({new_AGEMA_signal_2518, KeyArray_outS11ser[1]}), .c ({new_AGEMA_signal_2889, KeyArray_S01reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S01reg_gff_1_SFF_2_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2016, KeyArray_outS01ser_2_}), .a ({new_AGEMA_signal_2890, KeyArray_S01reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_3277, KeyArray_S01reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_2450, KeyArray_inS01ser[2]}), .a ({new_AGEMA_signal_2521, KeyArray_outS11ser[2]}), .c ({new_AGEMA_signal_2890, KeyArray_S01reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S01reg_gff_1_SFF_3_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2014, KeyArray_outS01ser_3_}), .a ({new_AGEMA_signal_2891, KeyArray_S01reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_3278, KeyArray_S01reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_2453, KeyArray_inS01ser[3]}), .a ({new_AGEMA_signal_2524, KeyArray_outS11ser[3]}), .c ({new_AGEMA_signal_2891, KeyArray_S01reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S01reg_gff_1_SFF_4_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2012, KeyArray_outS01ser_4_}), .a ({new_AGEMA_signal_2892, KeyArray_S01reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_3279, KeyArray_S01reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_2456, KeyArray_inS01ser[4]}), .a ({new_AGEMA_signal_2527, KeyArray_outS11ser[4]}), .c ({new_AGEMA_signal_2892, KeyArray_S01reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S01reg_gff_1_SFF_5_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2010, KeyArray_outS01ser_5_}), .a ({new_AGEMA_signal_2893, KeyArray_S01reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_3280, KeyArray_S01reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_2459, KeyArray_inS01ser[5]}), .a ({new_AGEMA_signal_2530, KeyArray_outS11ser[5]}), .c ({new_AGEMA_signal_2893, KeyArray_S01reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S01reg_gff_1_SFF_6_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2008, KeyArray_outS01ser_6_}), .a ({new_AGEMA_signal_2894, KeyArray_S01reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_3281, KeyArray_S01reg_gff_1_SFF_6_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_2462, KeyArray_inS01ser[6]}), .a ({new_AGEMA_signal_2533, KeyArray_outS11ser[6]}), .c ({new_AGEMA_signal_2894, KeyArray_S01reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S01reg_gff_1_SFF_7_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2006, KeyArray_outS01ser_7_}), .a ({new_AGEMA_signal_2895, KeyArray_S01reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_3282, KeyArray_S01reg_gff_1_SFF_7_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_2465, KeyArray_inS01ser[7]}), .a ({new_AGEMA_signal_2536, KeyArray_outS11ser[7]}), .c ({new_AGEMA_signal_2895, KeyArray_S01reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S02reg_gff_1_SFF_0_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_2443, KeyArray_outS02ser[0]}), .a ({new_AGEMA_signal_2896, KeyArray_S02reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_3283, KeyArray_S02reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_2468, KeyArray_inS02ser[0]}), .a ({new_AGEMA_signal_2539, KeyArray_outS12ser[0]}), .c ({new_AGEMA_signal_2896, KeyArray_S02reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S02reg_gff_1_SFF_1_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_2446, KeyArray_outS02ser[1]}), .a ({new_AGEMA_signal_2897, KeyArray_S02reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_3284, KeyArray_S02reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_2471, KeyArray_inS02ser[1]}), .a ({new_AGEMA_signal_2542, KeyArray_outS12ser[1]}), .c ({new_AGEMA_signal_2897, KeyArray_S02reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S02reg_gff_1_SFF_2_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_2449, KeyArray_outS02ser[2]}), .a ({new_AGEMA_signal_2898, KeyArray_S02reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_3285, KeyArray_S02reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_2474, KeyArray_inS02ser[2]}), .a ({new_AGEMA_signal_2545, KeyArray_outS12ser[2]}), .c ({new_AGEMA_signal_2898, KeyArray_S02reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S02reg_gff_1_SFF_3_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_2452, KeyArray_outS02ser[3]}), .a ({new_AGEMA_signal_2899, KeyArray_S02reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_3286, KeyArray_S02reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_2477, KeyArray_inS02ser[3]}), .a ({new_AGEMA_signal_2548, KeyArray_outS12ser[3]}), .c ({new_AGEMA_signal_2899, KeyArray_S02reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S02reg_gff_1_SFF_4_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_2455, KeyArray_outS02ser[4]}), .a ({new_AGEMA_signal_2900, KeyArray_S02reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_3287, KeyArray_S02reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_2480, KeyArray_inS02ser[4]}), .a ({new_AGEMA_signal_2551, KeyArray_outS12ser[4]}), .c ({new_AGEMA_signal_2900, KeyArray_S02reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S02reg_gff_1_SFF_5_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_2458, KeyArray_outS02ser[5]}), .a ({new_AGEMA_signal_2901, KeyArray_S02reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_3288, KeyArray_S02reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_2483, KeyArray_inS02ser[5]}), .a ({new_AGEMA_signal_2554, KeyArray_outS12ser[5]}), .c ({new_AGEMA_signal_2901, KeyArray_S02reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S02reg_gff_1_SFF_6_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_2461, KeyArray_outS02ser[6]}), .a ({new_AGEMA_signal_2902, KeyArray_S02reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_3289, KeyArray_S02reg_gff_1_SFF_6_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_2486, KeyArray_inS02ser[6]}), .a ({new_AGEMA_signal_2557, KeyArray_outS12ser[6]}), .c ({new_AGEMA_signal_2902, KeyArray_S02reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S02reg_gff_1_SFF_7_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_2464, KeyArray_outS02ser[7]}), .a ({new_AGEMA_signal_2903, KeyArray_S02reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_3290, KeyArray_S02reg_gff_1_SFF_7_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_2489, KeyArray_inS02ser[7]}), .a ({new_AGEMA_signal_2560, KeyArray_outS12ser[7]}), .c ({new_AGEMA_signal_2903, KeyArray_S02reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S03reg_gff_1_SFF_0_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_2467, KeyArray_outS03ser[0]}), .a ({new_AGEMA_signal_2904, KeyArray_S03reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_3291, KeyArray_S03reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_2492, KeyArray_inS03ser[0]}), .a ({new_AGEMA_signal_2563, keySBIn[0]}), .c ({new_AGEMA_signal_2904, KeyArray_S03reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S03reg_gff_1_SFF_1_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_2470, KeyArray_outS03ser[1]}), .a ({new_AGEMA_signal_2905, KeyArray_S03reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_3292, KeyArray_S03reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_2495, KeyArray_inS03ser[1]}), .a ({new_AGEMA_signal_2566, keySBIn[1]}), .c ({new_AGEMA_signal_2905, KeyArray_S03reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S03reg_gff_1_SFF_2_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_2473, KeyArray_outS03ser[2]}), .a ({new_AGEMA_signal_2906, KeyArray_S03reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_3293, KeyArray_S03reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_2498, KeyArray_inS03ser[2]}), .a ({new_AGEMA_signal_2569, keySBIn[2]}), .c ({new_AGEMA_signal_2906, KeyArray_S03reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S03reg_gff_1_SFF_3_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_2476, KeyArray_outS03ser[3]}), .a ({new_AGEMA_signal_2907, KeyArray_S03reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_3294, KeyArray_S03reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_2501, KeyArray_inS03ser[3]}), .a ({new_AGEMA_signal_2572, keySBIn[3]}), .c ({new_AGEMA_signal_2907, KeyArray_S03reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S03reg_gff_1_SFF_4_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_2479, KeyArray_outS03ser[4]}), .a ({new_AGEMA_signal_2908, KeyArray_S03reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_3295, KeyArray_S03reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_2504, KeyArray_inS03ser[4]}), .a ({new_AGEMA_signal_2575, keySBIn[4]}), .c ({new_AGEMA_signal_2908, KeyArray_S03reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S03reg_gff_1_SFF_5_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_2482, KeyArray_outS03ser[5]}), .a ({new_AGEMA_signal_2909, KeyArray_S03reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_3296, KeyArray_S03reg_gff_1_SFF_5_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_2507, KeyArray_inS03ser[5]}), .a ({new_AGEMA_signal_2578, keySBIn[5]}), .c ({new_AGEMA_signal_2909, KeyArray_S03reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S03reg_gff_1_SFF_6_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_2485, KeyArray_outS03ser[6]}), .a ({new_AGEMA_signal_2910, KeyArray_S03reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_3297, KeyArray_S03reg_gff_1_SFF_6_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_2510, KeyArray_inS03ser[6]}), .a ({new_AGEMA_signal_2581, keySBIn[6]}), .c ({new_AGEMA_signal_2910, KeyArray_S03reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S03reg_gff_1_SFF_7_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_2488, KeyArray_outS03ser[7]}), .a ({new_AGEMA_signal_2911, KeyArray_S03reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_3298, KeyArray_S03reg_gff_1_SFF_7_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_2513, KeyArray_inS03ser[7]}), .a ({new_AGEMA_signal_2584, keySBIn[7]}), .c ({new_AGEMA_signal_2911, KeyArray_S03reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S10reg_gff_1_SFF_0_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_2491, KeyArray_outS10ser[0]}), .a ({new_AGEMA_signal_2912, KeyArray_S10reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_3299, KeyArray_S10reg_gff_1_SFF_0_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_2516, KeyArray_inS10ser[0]}), .a ({new_AGEMA_signal_2587, KeyArray_outS20ser[0]}), .c ({new_AGEMA_signal_2912, KeyArray_S10reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S10reg_gff_1_SFF_1_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_2494, KeyArray_outS10ser[1]}), .a ({new_AGEMA_signal_2913, KeyArray_S10reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_3300, KeyArray_S10reg_gff_1_SFF_1_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_2519, KeyArray_inS10ser[1]}), .a ({new_AGEMA_signal_2590, KeyArray_outS20ser[1]}), .c ({new_AGEMA_signal_2913, KeyArray_S10reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S10reg_gff_1_SFF_2_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_2497, KeyArray_outS10ser[2]}), .a ({new_AGEMA_signal_2914, KeyArray_S10reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_3301, KeyArray_S10reg_gff_1_SFF_2_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_2522, KeyArray_inS10ser[2]}), .a ({new_AGEMA_signal_2593, KeyArray_outS20ser[2]}), .c ({new_AGEMA_signal_2914, KeyArray_S10reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S10reg_gff_1_SFF_3_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_2500, KeyArray_outS10ser[3]}), .a ({new_AGEMA_signal_2915, KeyArray_S10reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_3302, KeyArray_S10reg_gff_1_SFF_3_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_2525, KeyArray_inS10ser[3]}), .a ({new_AGEMA_signal_2596, KeyArray_outS20ser[3]}), .c ({new_AGEMA_signal_2915, KeyArray_S10reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S10reg_gff_1_SFF_4_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_2503, KeyArray_outS10ser[4]}), .a ({new_AGEMA_signal_2916, KeyArray_S10reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_3303, KeyArray_S10reg_gff_1_SFF_4_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_2528, KeyArray_inS10ser[4]}), .a ({new_AGEMA_signal_2599, KeyArray_outS20ser[4]}), .c ({new_AGEMA_signal_2916, KeyArray_S10reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S10reg_gff_1_SFF_5_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_2506, KeyArray_outS10ser[5]}), .a ({new_AGEMA_signal_2917, KeyArray_S10reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_3304, KeyArray_S10reg_gff_1_SFF_5_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_2531, KeyArray_inS10ser[5]}), .a ({new_AGEMA_signal_2602, KeyArray_outS20ser[5]}), .c ({new_AGEMA_signal_2917, KeyArray_S10reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S10reg_gff_1_SFF_6_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_2509, KeyArray_outS10ser[6]}), .a ({new_AGEMA_signal_2918, KeyArray_S10reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_3305, KeyArray_S10reg_gff_1_SFF_6_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_2534, KeyArray_inS10ser[6]}), .a ({new_AGEMA_signal_2605, KeyArray_outS20ser[6]}), .c ({new_AGEMA_signal_2918, KeyArray_S10reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S10reg_gff_1_SFF_7_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_2512, KeyArray_outS10ser[7]}), .a ({new_AGEMA_signal_2919, KeyArray_S10reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_3306, KeyArray_S10reg_gff_1_SFF_7_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_2537, KeyArray_inS10ser[7]}), .a ({new_AGEMA_signal_2608, KeyArray_outS20ser[7]}), .c ({new_AGEMA_signal_2919, KeyArray_S10reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S11reg_gff_1_SFF_0_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_2515, KeyArray_outS11ser[0]}), .a ({new_AGEMA_signal_2920, KeyArray_S11reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_3307, KeyArray_S11reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_2540, KeyArray_inS11ser[0]}), .a ({new_AGEMA_signal_2611, KeyArray_outS21ser[0]}), .c ({new_AGEMA_signal_2920, KeyArray_S11reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S11reg_gff_1_SFF_1_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_2518, KeyArray_outS11ser[1]}), .a ({new_AGEMA_signal_2921, KeyArray_S11reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_3308, KeyArray_S11reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_2543, KeyArray_inS11ser[1]}), .a ({new_AGEMA_signal_2614, KeyArray_outS21ser[1]}), .c ({new_AGEMA_signal_2921, KeyArray_S11reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S11reg_gff_1_SFF_2_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_2521, KeyArray_outS11ser[2]}), .a ({new_AGEMA_signal_2922, KeyArray_S11reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_3309, KeyArray_S11reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_2546, KeyArray_inS11ser[2]}), .a ({new_AGEMA_signal_2617, KeyArray_outS21ser[2]}), .c ({new_AGEMA_signal_2922, KeyArray_S11reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S11reg_gff_1_SFF_3_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_2524, KeyArray_outS11ser[3]}), .a ({new_AGEMA_signal_2923, KeyArray_S11reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_3310, KeyArray_S11reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_2549, KeyArray_inS11ser[3]}), .a ({new_AGEMA_signal_2620, KeyArray_outS21ser[3]}), .c ({new_AGEMA_signal_2923, KeyArray_S11reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S11reg_gff_1_SFF_4_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_2527, KeyArray_outS11ser[4]}), .a ({new_AGEMA_signal_2924, KeyArray_S11reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_3311, KeyArray_S11reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_2552, KeyArray_inS11ser[4]}), .a ({new_AGEMA_signal_2623, KeyArray_outS21ser[4]}), .c ({new_AGEMA_signal_2924, KeyArray_S11reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S11reg_gff_1_SFF_5_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_2530, KeyArray_outS11ser[5]}), .a ({new_AGEMA_signal_2925, KeyArray_S11reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_3312, KeyArray_S11reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_2555, KeyArray_inS11ser[5]}), .a ({new_AGEMA_signal_2626, KeyArray_outS21ser[5]}), .c ({new_AGEMA_signal_2925, KeyArray_S11reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S11reg_gff_1_SFF_6_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_2533, KeyArray_outS11ser[6]}), .a ({new_AGEMA_signal_2926, KeyArray_S11reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_3313, KeyArray_S11reg_gff_1_SFF_6_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_2558, KeyArray_inS11ser[6]}), .a ({new_AGEMA_signal_2629, KeyArray_outS21ser[6]}), .c ({new_AGEMA_signal_2926, KeyArray_S11reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S11reg_gff_1_SFF_7_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_2536, KeyArray_outS11ser[7]}), .a ({new_AGEMA_signal_2927, KeyArray_S11reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_3314, KeyArray_S11reg_gff_1_SFF_7_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_2561, KeyArray_inS11ser[7]}), .a ({new_AGEMA_signal_2632, KeyArray_outS21ser[7]}), .c ({new_AGEMA_signal_2927, KeyArray_S11reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S12reg_gff_1_SFF_0_U1 ( .s (n12), .b ({new_AGEMA_signal_2539, KeyArray_outS12ser[0]}), .a ({new_AGEMA_signal_2928, KeyArray_S12reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_3093, KeyArray_S12reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_2564, KeyArray_inS12ser[0]}), .a ({new_AGEMA_signal_2635, KeyArray_outS22ser[0]}), .c ({new_AGEMA_signal_2928, KeyArray_S12reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S12reg_gff_1_SFF_1_U1 ( .s (n12), .b ({new_AGEMA_signal_2542, KeyArray_outS12ser[1]}), .a ({new_AGEMA_signal_2929, KeyArray_S12reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_3094, KeyArray_S12reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_2567, KeyArray_inS12ser[1]}), .a ({new_AGEMA_signal_2638, KeyArray_outS22ser[1]}), .c ({new_AGEMA_signal_2929, KeyArray_S12reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S12reg_gff_1_SFF_2_U1 ( .s (n12), .b ({new_AGEMA_signal_2545, KeyArray_outS12ser[2]}), .a ({new_AGEMA_signal_2930, KeyArray_S12reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_3095, KeyArray_S12reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_2570, KeyArray_inS12ser[2]}), .a ({new_AGEMA_signal_2641, KeyArray_outS22ser[2]}), .c ({new_AGEMA_signal_2930, KeyArray_S12reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S12reg_gff_1_SFF_3_U1 ( .s (n12), .b ({new_AGEMA_signal_2548, KeyArray_outS12ser[3]}), .a ({new_AGEMA_signal_2931, KeyArray_S12reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_3096, KeyArray_S12reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_2573, KeyArray_inS12ser[3]}), .a ({new_AGEMA_signal_2644, KeyArray_outS22ser[3]}), .c ({new_AGEMA_signal_2931, KeyArray_S12reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S12reg_gff_1_SFF_4_U1 ( .s (n12), .b ({new_AGEMA_signal_2551, KeyArray_outS12ser[4]}), .a ({new_AGEMA_signal_2932, KeyArray_S12reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_3097, KeyArray_S12reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_2576, KeyArray_inS12ser[4]}), .a ({new_AGEMA_signal_2647, KeyArray_outS22ser[4]}), .c ({new_AGEMA_signal_2932, KeyArray_S12reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S12reg_gff_1_SFF_5_U1 ( .s (n12), .b ({new_AGEMA_signal_2554, KeyArray_outS12ser[5]}), .a ({new_AGEMA_signal_2933, KeyArray_S12reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_3098, KeyArray_S12reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_2579, KeyArray_inS12ser[5]}), .a ({new_AGEMA_signal_2650, KeyArray_outS22ser[5]}), .c ({new_AGEMA_signal_2933, KeyArray_S12reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S12reg_gff_1_SFF_6_U1 ( .s (n12), .b ({new_AGEMA_signal_2557, KeyArray_outS12ser[6]}), .a ({new_AGEMA_signal_2934, KeyArray_S12reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_3099, KeyArray_S12reg_gff_1_SFF_6_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_2582, KeyArray_inS12ser[6]}), .a ({new_AGEMA_signal_2653, KeyArray_outS22ser[6]}), .c ({new_AGEMA_signal_2934, KeyArray_S12reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S12reg_gff_1_SFF_7_U1 ( .s (n12), .b ({new_AGEMA_signal_2560, KeyArray_outS12ser[7]}), .a ({new_AGEMA_signal_2935, KeyArray_S12reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_3100, KeyArray_S12reg_gff_1_SFF_7_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_2585, KeyArray_inS12ser[7]}), .a ({new_AGEMA_signal_2656, KeyArray_outS22ser[7]}), .c ({new_AGEMA_signal_2935, KeyArray_S12reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S13reg_gff_1_SFF_0_U1 ( .s (n12), .b ({new_AGEMA_signal_2563, keySBIn[0]}), .a ({new_AGEMA_signal_2936, KeyArray_S13reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_3101, KeyArray_S13reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_2588, KeyArray_inS13ser[0]}), .a ({new_AGEMA_signal_2659, KeyArray_outS23ser[0]}), .c ({new_AGEMA_signal_2936, KeyArray_S13reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S13reg_gff_1_SFF_1_U1 ( .s (n12), .b ({new_AGEMA_signal_2566, keySBIn[1]}), .a ({new_AGEMA_signal_2937, KeyArray_S13reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_3102, KeyArray_S13reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_2591, KeyArray_inS13ser[1]}), .a ({new_AGEMA_signal_2662, KeyArray_outS23ser[1]}), .c ({new_AGEMA_signal_2937, KeyArray_S13reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S13reg_gff_1_SFF_2_U1 ( .s (n12), .b ({new_AGEMA_signal_2569, keySBIn[2]}), .a ({new_AGEMA_signal_2938, KeyArray_S13reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_3103, KeyArray_S13reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_2594, KeyArray_inS13ser[2]}), .a ({new_AGEMA_signal_2665, KeyArray_outS23ser[2]}), .c ({new_AGEMA_signal_2938, KeyArray_S13reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S13reg_gff_1_SFF_3_U1 ( .s (n12), .b ({new_AGEMA_signal_2572, keySBIn[3]}), .a ({new_AGEMA_signal_2939, KeyArray_S13reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_3104, KeyArray_S13reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_2597, KeyArray_inS13ser[3]}), .a ({new_AGEMA_signal_2668, KeyArray_outS23ser[3]}), .c ({new_AGEMA_signal_2939, KeyArray_S13reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S13reg_gff_1_SFF_4_U1 ( .s (n12), .b ({new_AGEMA_signal_2575, keySBIn[4]}), .a ({new_AGEMA_signal_2940, KeyArray_S13reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_3105, KeyArray_S13reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_2600, KeyArray_inS13ser[4]}), .a ({new_AGEMA_signal_2671, KeyArray_outS23ser[4]}), .c ({new_AGEMA_signal_2940, KeyArray_S13reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S13reg_gff_1_SFF_5_U1 ( .s (n12), .b ({new_AGEMA_signal_2578, keySBIn[5]}), .a ({new_AGEMA_signal_2941, KeyArray_S13reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_3106, KeyArray_S13reg_gff_1_SFF_5_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_2603, KeyArray_inS13ser[5]}), .a ({new_AGEMA_signal_2674, KeyArray_outS23ser[5]}), .c ({new_AGEMA_signal_2941, KeyArray_S13reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S13reg_gff_1_SFF_6_U1 ( .s (n12), .b ({new_AGEMA_signal_2581, keySBIn[6]}), .a ({new_AGEMA_signal_2942, KeyArray_S13reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_3107, KeyArray_S13reg_gff_1_SFF_6_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_2606, KeyArray_inS13ser[6]}), .a ({new_AGEMA_signal_2677, KeyArray_outS23ser[6]}), .c ({new_AGEMA_signal_2942, KeyArray_S13reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S13reg_gff_1_SFF_7_U1 ( .s (n12), .b ({new_AGEMA_signal_2584, keySBIn[7]}), .a ({new_AGEMA_signal_2943, KeyArray_S13reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_3108, KeyArray_S13reg_gff_1_SFF_7_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_2609, KeyArray_inS13ser[7]}), .a ({new_AGEMA_signal_2680, KeyArray_outS23ser[7]}), .c ({new_AGEMA_signal_2943, KeyArray_S13reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S20reg_gff_1_SFF_0_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_2587, KeyArray_outS20ser[0]}), .a ({new_AGEMA_signal_2944, KeyArray_S20reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_3315, KeyArray_S20reg_gff_1_SFF_0_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_2612, KeyArray_inS20ser[0]}), .a ({new_AGEMA_signal_2683, KeyArray_outS30ser[0]}), .c ({new_AGEMA_signal_2944, KeyArray_S20reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S20reg_gff_1_SFF_1_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_2590, KeyArray_outS20ser[1]}), .a ({new_AGEMA_signal_2945, KeyArray_S20reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_3316, KeyArray_S20reg_gff_1_SFF_1_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_2615, KeyArray_inS20ser[1]}), .a ({new_AGEMA_signal_2686, KeyArray_outS30ser[1]}), .c ({new_AGEMA_signal_2945, KeyArray_S20reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S20reg_gff_1_SFF_2_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_2593, KeyArray_outS20ser[2]}), .a ({new_AGEMA_signal_2946, KeyArray_S20reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_3317, KeyArray_S20reg_gff_1_SFF_2_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_2618, KeyArray_inS20ser[2]}), .a ({new_AGEMA_signal_2689, KeyArray_outS30ser[2]}), .c ({new_AGEMA_signal_2946, KeyArray_S20reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S20reg_gff_1_SFF_3_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_2596, KeyArray_outS20ser[3]}), .a ({new_AGEMA_signal_2947, KeyArray_S20reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_3318, KeyArray_S20reg_gff_1_SFF_3_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_2621, KeyArray_inS20ser[3]}), .a ({new_AGEMA_signal_2692, KeyArray_outS30ser[3]}), .c ({new_AGEMA_signal_2947, KeyArray_S20reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S20reg_gff_1_SFF_4_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_2599, KeyArray_outS20ser[4]}), .a ({new_AGEMA_signal_2948, KeyArray_S20reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_3319, KeyArray_S20reg_gff_1_SFF_4_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_2624, KeyArray_inS20ser[4]}), .a ({new_AGEMA_signal_2695, KeyArray_outS30ser[4]}), .c ({new_AGEMA_signal_2948, KeyArray_S20reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S20reg_gff_1_SFF_5_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_2602, KeyArray_outS20ser[5]}), .a ({new_AGEMA_signal_2949, KeyArray_S20reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_3320, KeyArray_S20reg_gff_1_SFF_5_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_2627, KeyArray_inS20ser[5]}), .a ({new_AGEMA_signal_2698, KeyArray_outS30ser[5]}), .c ({new_AGEMA_signal_2949, KeyArray_S20reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S20reg_gff_1_SFF_6_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_2605, KeyArray_outS20ser[6]}), .a ({new_AGEMA_signal_2950, KeyArray_S20reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_3321, KeyArray_S20reg_gff_1_SFF_6_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_2630, KeyArray_inS20ser[6]}), .a ({new_AGEMA_signal_2701, KeyArray_outS30ser[6]}), .c ({new_AGEMA_signal_2950, KeyArray_S20reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S20reg_gff_1_SFF_7_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_2608, KeyArray_outS20ser[7]}), .a ({new_AGEMA_signal_2951, KeyArray_S20reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_3322, KeyArray_S20reg_gff_1_SFF_7_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_2633, KeyArray_inS20ser[7]}), .a ({new_AGEMA_signal_2704, KeyArray_outS30ser[7]}), .c ({new_AGEMA_signal_2951, KeyArray_S20reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S21reg_gff_1_SFF_0_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_2611, KeyArray_outS21ser[0]}), .a ({new_AGEMA_signal_2952, KeyArray_S21reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_3323, KeyArray_S21reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_2636, KeyArray_inS21ser[0]}), .a ({new_AGEMA_signal_2707, KeyArray_outS31ser[0]}), .c ({new_AGEMA_signal_2952, KeyArray_S21reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S21reg_gff_1_SFF_1_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_2614, KeyArray_outS21ser[1]}), .a ({new_AGEMA_signal_2953, KeyArray_S21reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_3324, KeyArray_S21reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_2639, KeyArray_inS21ser[1]}), .a ({new_AGEMA_signal_2710, KeyArray_outS31ser[1]}), .c ({new_AGEMA_signal_2953, KeyArray_S21reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S21reg_gff_1_SFF_2_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_2617, KeyArray_outS21ser[2]}), .a ({new_AGEMA_signal_2954, KeyArray_S21reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_3325, KeyArray_S21reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_2642, KeyArray_inS21ser[2]}), .a ({new_AGEMA_signal_2713, KeyArray_outS31ser[2]}), .c ({new_AGEMA_signal_2954, KeyArray_S21reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S21reg_gff_1_SFF_3_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_2620, KeyArray_outS21ser[3]}), .a ({new_AGEMA_signal_2955, KeyArray_S21reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_3326, KeyArray_S21reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_2645, KeyArray_inS21ser[3]}), .a ({new_AGEMA_signal_2716, KeyArray_outS31ser[3]}), .c ({new_AGEMA_signal_2955, KeyArray_S21reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S21reg_gff_1_SFF_4_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_2623, KeyArray_outS21ser[4]}), .a ({new_AGEMA_signal_2956, KeyArray_S21reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_3327, KeyArray_S21reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_2648, KeyArray_inS21ser[4]}), .a ({new_AGEMA_signal_2719, KeyArray_outS31ser[4]}), .c ({new_AGEMA_signal_2956, KeyArray_S21reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S21reg_gff_1_SFF_5_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_2626, KeyArray_outS21ser[5]}), .a ({new_AGEMA_signal_2957, KeyArray_S21reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_3328, KeyArray_S21reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_2651, KeyArray_inS21ser[5]}), .a ({new_AGEMA_signal_2722, KeyArray_outS31ser[5]}), .c ({new_AGEMA_signal_2957, KeyArray_S21reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S21reg_gff_1_SFF_6_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_2629, KeyArray_outS21ser[6]}), .a ({new_AGEMA_signal_2958, KeyArray_S21reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_3329, KeyArray_S21reg_gff_1_SFF_6_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_2654, KeyArray_inS21ser[6]}), .a ({new_AGEMA_signal_2725, KeyArray_outS31ser[6]}), .c ({new_AGEMA_signal_2958, KeyArray_S21reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S21reg_gff_1_SFF_7_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_2632, KeyArray_outS21ser[7]}), .a ({new_AGEMA_signal_2959, KeyArray_S21reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_3330, KeyArray_S21reg_gff_1_SFF_7_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_2657, KeyArray_inS21ser[7]}), .a ({new_AGEMA_signal_2728, KeyArray_outS31ser[7]}), .c ({new_AGEMA_signal_2959, KeyArray_S21reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S22reg_gff_1_SFF_0_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_2635, KeyArray_outS22ser[0]}), .a ({new_AGEMA_signal_2960, KeyArray_S22reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_3331, KeyArray_S22reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_2660, KeyArray_inS22ser[0]}), .a ({new_AGEMA_signal_2731, KeyArray_outS32ser[0]}), .c ({new_AGEMA_signal_2960, KeyArray_S22reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S22reg_gff_1_SFF_1_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_2638, KeyArray_outS22ser[1]}), .a ({new_AGEMA_signal_2961, KeyArray_S22reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_3332, KeyArray_S22reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_2663, KeyArray_inS22ser[1]}), .a ({new_AGEMA_signal_2734, KeyArray_outS32ser[1]}), .c ({new_AGEMA_signal_2961, KeyArray_S22reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S22reg_gff_1_SFF_2_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_2641, KeyArray_outS22ser[2]}), .a ({new_AGEMA_signal_2962, KeyArray_S22reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_3333, KeyArray_S22reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_2666, KeyArray_inS22ser[2]}), .a ({new_AGEMA_signal_2737, KeyArray_outS32ser[2]}), .c ({new_AGEMA_signal_2962, KeyArray_S22reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S22reg_gff_1_SFF_3_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_2644, KeyArray_outS22ser[3]}), .a ({new_AGEMA_signal_2963, KeyArray_S22reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_3334, KeyArray_S22reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_2669, KeyArray_inS22ser[3]}), .a ({new_AGEMA_signal_2740, KeyArray_outS32ser[3]}), .c ({new_AGEMA_signal_2963, KeyArray_S22reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S22reg_gff_1_SFF_4_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_2647, KeyArray_outS22ser[4]}), .a ({new_AGEMA_signal_2964, KeyArray_S22reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_3335, KeyArray_S22reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_2672, KeyArray_inS22ser[4]}), .a ({new_AGEMA_signal_2743, KeyArray_outS32ser[4]}), .c ({new_AGEMA_signal_2964, KeyArray_S22reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S22reg_gff_1_SFF_5_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_2650, KeyArray_outS22ser[5]}), .a ({new_AGEMA_signal_2965, KeyArray_S22reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_3336, KeyArray_S22reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_2675, KeyArray_inS22ser[5]}), .a ({new_AGEMA_signal_2746, KeyArray_outS32ser[5]}), .c ({new_AGEMA_signal_2965, KeyArray_S22reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S22reg_gff_1_SFF_6_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_2653, KeyArray_outS22ser[6]}), .a ({new_AGEMA_signal_2966, KeyArray_S22reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_3337, KeyArray_S22reg_gff_1_SFF_6_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_2678, KeyArray_inS22ser[6]}), .a ({new_AGEMA_signal_2749, KeyArray_outS32ser[6]}), .c ({new_AGEMA_signal_2966, KeyArray_S22reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S22reg_gff_1_SFF_7_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_2656, KeyArray_outS22ser[7]}), .a ({new_AGEMA_signal_2967, KeyArray_S22reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_3338, KeyArray_S22reg_gff_1_SFF_7_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_2681, KeyArray_inS22ser[7]}), .a ({new_AGEMA_signal_2752, KeyArray_outS32ser[7]}), .c ({new_AGEMA_signal_2967, KeyArray_S22reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S23reg_gff_1_SFF_0_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_2659, KeyArray_outS23ser[0]}), .a ({new_AGEMA_signal_2968, KeyArray_S23reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_3339, KeyArray_S23reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_2684, KeyArray_inS23ser[0]}), .a ({new_AGEMA_signal_2755, KeyArray_outS33ser[0]}), .c ({new_AGEMA_signal_2968, KeyArray_S23reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S23reg_gff_1_SFF_1_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_2662, KeyArray_outS23ser[1]}), .a ({new_AGEMA_signal_2969, KeyArray_S23reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_3340, KeyArray_S23reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_2687, KeyArray_inS23ser[1]}), .a ({new_AGEMA_signal_2758, KeyArray_outS33ser[1]}), .c ({new_AGEMA_signal_2969, KeyArray_S23reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S23reg_gff_1_SFF_2_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_2665, KeyArray_outS23ser[2]}), .a ({new_AGEMA_signal_2970, KeyArray_S23reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_3341, KeyArray_S23reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_2690, KeyArray_inS23ser[2]}), .a ({new_AGEMA_signal_2761, KeyArray_outS33ser[2]}), .c ({new_AGEMA_signal_2970, KeyArray_S23reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S23reg_gff_1_SFF_3_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_2668, KeyArray_outS23ser[3]}), .a ({new_AGEMA_signal_2971, KeyArray_S23reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_3342, KeyArray_S23reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_2693, KeyArray_inS23ser[3]}), .a ({new_AGEMA_signal_2764, KeyArray_outS33ser[3]}), .c ({new_AGEMA_signal_2971, KeyArray_S23reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S23reg_gff_1_SFF_4_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_2671, KeyArray_outS23ser[4]}), .a ({new_AGEMA_signal_2972, KeyArray_S23reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_3343, KeyArray_S23reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_2696, KeyArray_inS23ser[4]}), .a ({new_AGEMA_signal_2767, KeyArray_outS33ser[4]}), .c ({new_AGEMA_signal_2972, KeyArray_S23reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S23reg_gff_1_SFF_5_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_2674, KeyArray_outS23ser[5]}), .a ({new_AGEMA_signal_2973, KeyArray_S23reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_3344, KeyArray_S23reg_gff_1_SFF_5_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_2699, KeyArray_inS23ser[5]}), .a ({new_AGEMA_signal_2770, KeyArray_outS33ser[5]}), .c ({new_AGEMA_signal_2973, KeyArray_S23reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S23reg_gff_1_SFF_6_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_2677, KeyArray_outS23ser[6]}), .a ({new_AGEMA_signal_2974, KeyArray_S23reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_3345, KeyArray_S23reg_gff_1_SFF_6_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_2702, KeyArray_inS23ser[6]}), .a ({new_AGEMA_signal_2773, KeyArray_outS33ser[6]}), .c ({new_AGEMA_signal_2974, KeyArray_S23reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S23reg_gff_1_SFF_7_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_2680, KeyArray_outS23ser[7]}), .a ({new_AGEMA_signal_2975, KeyArray_S23reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_3346, KeyArray_S23reg_gff_1_SFF_7_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_2705, KeyArray_inS23ser[7]}), .a ({new_AGEMA_signal_2776, KeyArray_outS33ser[7]}), .c ({new_AGEMA_signal_2975, KeyArray_S23reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S31reg_gff_1_SFF_0_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_2707, KeyArray_outS31ser[0]}), .a ({new_AGEMA_signal_2976, KeyArray_S31reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_3347, KeyArray_S31reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_2732, KeyArray_inS31ser[0]}), .a ({new_AGEMA_signal_2020, KeyArray_outS01ser_0_}), .c ({new_AGEMA_signal_2976, KeyArray_S31reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S31reg_gff_1_SFF_1_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_2710, KeyArray_outS31ser[1]}), .a ({new_AGEMA_signal_2977, KeyArray_S31reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_3348, KeyArray_S31reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_2735, KeyArray_inS31ser[1]}), .a ({new_AGEMA_signal_2018, KeyArray_outS01ser_1_}), .c ({new_AGEMA_signal_2977, KeyArray_S31reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S31reg_gff_1_SFF_2_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_2713, KeyArray_outS31ser[2]}), .a ({new_AGEMA_signal_2978, KeyArray_S31reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_3349, KeyArray_S31reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_2738, KeyArray_inS31ser[2]}), .a ({new_AGEMA_signal_2016, KeyArray_outS01ser_2_}), .c ({new_AGEMA_signal_2978, KeyArray_S31reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S31reg_gff_1_SFF_3_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_2716, KeyArray_outS31ser[3]}), .a ({new_AGEMA_signal_2979, KeyArray_S31reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_3350, KeyArray_S31reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_2741, KeyArray_inS31ser[3]}), .a ({new_AGEMA_signal_2014, KeyArray_outS01ser_3_}), .c ({new_AGEMA_signal_2979, KeyArray_S31reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S31reg_gff_1_SFF_4_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_2719, KeyArray_outS31ser[4]}), .a ({new_AGEMA_signal_2980, KeyArray_S31reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_3351, KeyArray_S31reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_2744, KeyArray_inS31ser[4]}), .a ({new_AGEMA_signal_2012, KeyArray_outS01ser_4_}), .c ({new_AGEMA_signal_2980, KeyArray_S31reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S31reg_gff_1_SFF_5_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_2722, KeyArray_outS31ser[5]}), .a ({new_AGEMA_signal_2981, KeyArray_S31reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_3352, KeyArray_S31reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_2747, KeyArray_inS31ser[5]}), .a ({new_AGEMA_signal_2010, KeyArray_outS01ser_5_}), .c ({new_AGEMA_signal_2981, KeyArray_S31reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S31reg_gff_1_SFF_6_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_2725, KeyArray_outS31ser[6]}), .a ({new_AGEMA_signal_2982, KeyArray_S31reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_3353, KeyArray_S31reg_gff_1_SFF_6_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_2750, KeyArray_inS31ser[6]}), .a ({new_AGEMA_signal_2008, KeyArray_outS01ser_6_}), .c ({new_AGEMA_signal_2982, KeyArray_S31reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S31reg_gff_1_SFF_7_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_2728, KeyArray_outS31ser[7]}), .a ({new_AGEMA_signal_2983, KeyArray_S31reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_3354, KeyArray_S31reg_gff_1_SFF_7_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_2753, KeyArray_inS31ser[7]}), .a ({new_AGEMA_signal_2006, KeyArray_outS01ser_7_}), .c ({new_AGEMA_signal_2983, KeyArray_S31reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S32reg_gff_1_SFF_0_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_2731, KeyArray_outS32ser[0]}), .a ({new_AGEMA_signal_2984, KeyArray_S32reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_3355, KeyArray_S32reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_2756, KeyArray_inS32ser[0]}), .a ({new_AGEMA_signal_2443, KeyArray_outS02ser[0]}), .c ({new_AGEMA_signal_2984, KeyArray_S32reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S32reg_gff_1_SFF_1_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_2734, KeyArray_outS32ser[1]}), .a ({new_AGEMA_signal_2985, KeyArray_S32reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_3356, KeyArray_S32reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_2759, KeyArray_inS32ser[1]}), .a ({new_AGEMA_signal_2446, KeyArray_outS02ser[1]}), .c ({new_AGEMA_signal_2985, KeyArray_S32reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S32reg_gff_1_SFF_2_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_2737, KeyArray_outS32ser[2]}), .a ({new_AGEMA_signal_2986, KeyArray_S32reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_3357, KeyArray_S32reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_2762, KeyArray_inS32ser[2]}), .a ({new_AGEMA_signal_2449, KeyArray_outS02ser[2]}), .c ({new_AGEMA_signal_2986, KeyArray_S32reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S32reg_gff_1_SFF_3_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_2740, KeyArray_outS32ser[3]}), .a ({new_AGEMA_signal_2987, KeyArray_S32reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_3358, KeyArray_S32reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_2765, KeyArray_inS32ser[3]}), .a ({new_AGEMA_signal_2452, KeyArray_outS02ser[3]}), .c ({new_AGEMA_signal_2987, KeyArray_S32reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S32reg_gff_1_SFF_4_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_2743, KeyArray_outS32ser[4]}), .a ({new_AGEMA_signal_2988, KeyArray_S32reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_3359, KeyArray_S32reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_2768, KeyArray_inS32ser[4]}), .a ({new_AGEMA_signal_2455, KeyArray_outS02ser[4]}), .c ({new_AGEMA_signal_2988, KeyArray_S32reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S32reg_gff_1_SFF_5_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_2746, KeyArray_outS32ser[5]}), .a ({new_AGEMA_signal_2989, KeyArray_S32reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_3360, KeyArray_S32reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_2771, KeyArray_inS32ser[5]}), .a ({new_AGEMA_signal_2458, KeyArray_outS02ser[5]}), .c ({new_AGEMA_signal_2989, KeyArray_S32reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S32reg_gff_1_SFF_6_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_2749, KeyArray_outS32ser[6]}), .a ({new_AGEMA_signal_2990, KeyArray_S32reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_3361, KeyArray_S32reg_gff_1_SFF_6_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_2774, KeyArray_inS32ser[6]}), .a ({new_AGEMA_signal_2461, KeyArray_outS02ser[6]}), .c ({new_AGEMA_signal_2990, KeyArray_S32reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S32reg_gff_1_SFF_7_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_2752, KeyArray_outS32ser[7]}), .a ({new_AGEMA_signal_2991, KeyArray_S32reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_3362, KeyArray_S32reg_gff_1_SFF_7_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_2777, KeyArray_inS32ser[7]}), .a ({new_AGEMA_signal_2464, KeyArray_outS02ser[7]}), .c ({new_AGEMA_signal_2991, KeyArray_S32reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S33reg_gff_1_SFF_0_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_2755, KeyArray_outS33ser[0]}), .a ({new_AGEMA_signal_2992, KeyArray_S33reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_3363, KeyArray_S33reg_gff_1_SFF_0_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_2779, KeyArray_inS33ser[0]}), .a ({new_AGEMA_signal_2467, KeyArray_outS03ser[0]}), .c ({new_AGEMA_signal_2992, KeyArray_S33reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S33reg_gff_1_SFF_1_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_2758, KeyArray_outS33ser[1]}), .a ({new_AGEMA_signal_2993, KeyArray_S33reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_3364, KeyArray_S33reg_gff_1_SFF_1_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_2781, KeyArray_inS33ser[1]}), .a ({new_AGEMA_signal_2470, KeyArray_outS03ser[1]}), .c ({new_AGEMA_signal_2993, KeyArray_S33reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S33reg_gff_1_SFF_2_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_2761, KeyArray_outS33ser[2]}), .a ({new_AGEMA_signal_2994, KeyArray_S33reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_3365, KeyArray_S33reg_gff_1_SFF_2_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_2783, KeyArray_inS33ser[2]}), .a ({new_AGEMA_signal_2473, KeyArray_outS03ser[2]}), .c ({new_AGEMA_signal_2994, KeyArray_S33reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S33reg_gff_1_SFF_3_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_2764, KeyArray_outS33ser[3]}), .a ({new_AGEMA_signal_2995, KeyArray_S33reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_3366, KeyArray_S33reg_gff_1_SFF_3_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_2785, KeyArray_inS33ser[3]}), .a ({new_AGEMA_signal_2476, KeyArray_outS03ser[3]}), .c ({new_AGEMA_signal_2995, KeyArray_S33reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S33reg_gff_1_SFF_4_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_2767, KeyArray_outS33ser[4]}), .a ({new_AGEMA_signal_2996, KeyArray_S33reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_3367, KeyArray_S33reg_gff_1_SFF_4_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_2787, KeyArray_inS33ser[4]}), .a ({new_AGEMA_signal_2479, KeyArray_outS03ser[4]}), .c ({new_AGEMA_signal_2996, KeyArray_S33reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S33reg_gff_1_SFF_5_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_2770, KeyArray_outS33ser[5]}), .a ({new_AGEMA_signal_2997, KeyArray_S33reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_3368, KeyArray_S33reg_gff_1_SFF_5_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_2789, KeyArray_inS33ser[5]}), .a ({new_AGEMA_signal_2482, KeyArray_outS03ser[5]}), .c ({new_AGEMA_signal_2997, KeyArray_S33reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S33reg_gff_1_SFF_6_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_2773, KeyArray_outS33ser[6]}), .a ({new_AGEMA_signal_2998, KeyArray_S33reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_3369, KeyArray_S33reg_gff_1_SFF_6_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_2791, KeyArray_inS33ser[6]}), .a ({new_AGEMA_signal_2485, KeyArray_outS03ser[6]}), .c ({new_AGEMA_signal_2998, KeyArray_S33reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S33reg_gff_1_SFF_7_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_2776, KeyArray_outS33ser[7]}), .a ({new_AGEMA_signal_2999, KeyArray_S33reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_3370, KeyArray_S33reg_gff_1_SFF_7_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_2793, KeyArray_inS33ser[7]}), .a ({new_AGEMA_signal_2488, KeyArray_outS03ser[7]}), .c ({new_AGEMA_signal_2999, KeyArray_S33reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_selXOR_mux_inst_0_U1 ( .s (intselXOR), .b ({new_AGEMA_signal_2020, KeyArray_outS01ser_0_}), .a ({new_AGEMA_signal_2021, KeyArray_outS01ser_XOR_00[0]}), .c ({new_AGEMA_signal_3109, KeyArray_outS01ser_p[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_selXOR_mux_inst_1_U1 ( .s (intselXOR), .b ({new_AGEMA_signal_2018, KeyArray_outS01ser_1_}), .a ({new_AGEMA_signal_2019, KeyArray_outS01ser_XOR_00[1]}), .c ({new_AGEMA_signal_3110, KeyArray_outS01ser_p[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_selXOR_mux_inst_2_U1 ( .s (intselXOR), .b ({new_AGEMA_signal_2016, KeyArray_outS01ser_2_}), .a ({new_AGEMA_signal_2017, KeyArray_outS01ser_XOR_00[2]}), .c ({new_AGEMA_signal_3111, KeyArray_outS01ser_p[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_selXOR_mux_inst_3_U1 ( .s (intselXOR), .b ({new_AGEMA_signal_2014, KeyArray_outS01ser_3_}), .a ({new_AGEMA_signal_2015, KeyArray_outS01ser_XOR_00[3]}), .c ({new_AGEMA_signal_3112, KeyArray_outS01ser_p[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_selXOR_mux_inst_4_U1 ( .s (intselXOR), .b ({new_AGEMA_signal_2012, KeyArray_outS01ser_4_}), .a ({new_AGEMA_signal_2013, KeyArray_outS01ser_XOR_00[4]}), .c ({new_AGEMA_signal_3113, KeyArray_outS01ser_p[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_selXOR_mux_inst_5_U1 ( .s (intselXOR), .b ({new_AGEMA_signal_2010, KeyArray_outS01ser_5_}), .a ({new_AGEMA_signal_2011, KeyArray_outS01ser_XOR_00[5]}), .c ({new_AGEMA_signal_3114, KeyArray_outS01ser_p[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_selXOR_mux_inst_6_U1 ( .s (intselXOR), .b ({new_AGEMA_signal_2008, KeyArray_outS01ser_6_}), .a ({new_AGEMA_signal_2009, KeyArray_outS01ser_XOR_00[6]}), .c ({new_AGEMA_signal_3115, KeyArray_outS01ser_p[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_selXOR_mux_inst_7_U1 ( .s (intselXOR), .b ({new_AGEMA_signal_2006, KeyArray_outS01ser_7_}), .a ({new_AGEMA_signal_2007, KeyArray_outS01ser_XOR_00[7]}), .c ({new_AGEMA_signal_3116, KeyArray_outS01ser_p[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS00ser_mux_inst_0_U1 ( .s (KeyArray_n46), .b ({key_s1[120], key_s0[120]}), .a ({new_AGEMA_signal_3109, KeyArray_outS01ser_p[0]}), .c ({new_AGEMA_signal_3247, KeyArray_inS00ser[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS00ser_mux_inst_1_U1 ( .s (KeyArray_n46), .b ({key_s1[121], key_s0[121]}), .a ({new_AGEMA_signal_3110, KeyArray_outS01ser_p[1]}), .c ({new_AGEMA_signal_3249, KeyArray_inS00ser[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS00ser_mux_inst_2_U1 ( .s (KeyArray_n46), .b ({key_s1[122], key_s0[122]}), .a ({new_AGEMA_signal_3111, KeyArray_outS01ser_p[2]}), .c ({new_AGEMA_signal_3251, KeyArray_inS00ser[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS00ser_mux_inst_3_U1 ( .s (KeyArray_n46), .b ({key_s1[123], key_s0[123]}), .a ({new_AGEMA_signal_3112, KeyArray_outS01ser_p[3]}), .c ({new_AGEMA_signal_3253, KeyArray_inS00ser[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS00ser_mux_inst_4_U1 ( .s (KeyArray_n46), .b ({key_s1[124], key_s0[124]}), .a ({new_AGEMA_signal_3113, KeyArray_outS01ser_p[4]}), .c ({new_AGEMA_signal_3255, KeyArray_inS00ser[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS00ser_mux_inst_5_U1 ( .s (KeyArray_n46), .b ({key_s1[125], key_s0[125]}), .a ({new_AGEMA_signal_3114, KeyArray_outS01ser_p[5]}), .c ({new_AGEMA_signal_3257, KeyArray_inS00ser[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS00ser_mux_inst_6_U1 ( .s (KeyArray_n46), .b ({key_s1[126], key_s0[126]}), .a ({new_AGEMA_signal_3115, KeyArray_outS01ser_p[6]}), .c ({new_AGEMA_signal_3259, KeyArray_inS00ser[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS00ser_mux_inst_7_U1 ( .s (KeyArray_n46), .b ({key_s1[127], key_s0[127]}), .a ({new_AGEMA_signal_3116, KeyArray_outS01ser_p[7]}), .c ({new_AGEMA_signal_3261, KeyArray_inS00ser[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS01ser_mux_inst_0_U1 ( .s (KeyArray_n46), .b ({key_s1[112], key_s0[112]}), .a ({new_AGEMA_signal_2443, KeyArray_outS02ser[0]}), .c ({new_AGEMA_signal_2444, KeyArray_inS01ser[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS01ser_mux_inst_1_U1 ( .s (KeyArray_n46), .b ({key_s1[113], key_s0[113]}), .a ({new_AGEMA_signal_2446, KeyArray_outS02ser[1]}), .c ({new_AGEMA_signal_2447, KeyArray_inS01ser[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS01ser_mux_inst_2_U1 ( .s (KeyArray_n46), .b ({key_s1[114], key_s0[114]}), .a ({new_AGEMA_signal_2449, KeyArray_outS02ser[2]}), .c ({new_AGEMA_signal_2450, KeyArray_inS01ser[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS01ser_mux_inst_3_U1 ( .s (KeyArray_n46), .b ({key_s1[115], key_s0[115]}), .a ({new_AGEMA_signal_2452, KeyArray_outS02ser[3]}), .c ({new_AGEMA_signal_2453, KeyArray_inS01ser[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS01ser_mux_inst_4_U1 ( .s (KeyArray_n46), .b ({key_s1[116], key_s0[116]}), .a ({new_AGEMA_signal_2455, KeyArray_outS02ser[4]}), .c ({new_AGEMA_signal_2456, KeyArray_inS01ser[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS01ser_mux_inst_5_U1 ( .s (KeyArray_n46), .b ({key_s1[117], key_s0[117]}), .a ({new_AGEMA_signal_2458, KeyArray_outS02ser[5]}), .c ({new_AGEMA_signal_2459, KeyArray_inS01ser[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS01ser_mux_inst_6_U1 ( .s (KeyArray_n46), .b ({key_s1[118], key_s0[118]}), .a ({new_AGEMA_signal_2461, KeyArray_outS02ser[6]}), .c ({new_AGEMA_signal_2462, KeyArray_inS01ser[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS01ser_mux_inst_7_U1 ( .s (KeyArray_n46), .b ({key_s1[119], key_s0[119]}), .a ({new_AGEMA_signal_2464, KeyArray_outS02ser[7]}), .c ({new_AGEMA_signal_2465, KeyArray_inS01ser[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS02ser_mux_inst_0_U1 ( .s (KeyArray_n45), .b ({key_s1[104], key_s0[104]}), .a ({new_AGEMA_signal_2467, KeyArray_outS03ser[0]}), .c ({new_AGEMA_signal_2468, KeyArray_inS02ser[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS02ser_mux_inst_1_U1 ( .s (KeyArray_n45), .b ({key_s1[105], key_s0[105]}), .a ({new_AGEMA_signal_2470, KeyArray_outS03ser[1]}), .c ({new_AGEMA_signal_2471, KeyArray_inS02ser[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS02ser_mux_inst_2_U1 ( .s (KeyArray_n45), .b ({key_s1[106], key_s0[106]}), .a ({new_AGEMA_signal_2473, KeyArray_outS03ser[2]}), .c ({new_AGEMA_signal_2474, KeyArray_inS02ser[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS02ser_mux_inst_3_U1 ( .s (KeyArray_n45), .b ({key_s1[107], key_s0[107]}), .a ({new_AGEMA_signal_2476, KeyArray_outS03ser[3]}), .c ({new_AGEMA_signal_2477, KeyArray_inS02ser[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS02ser_mux_inst_4_U1 ( .s (KeyArray_n45), .b ({key_s1[108], key_s0[108]}), .a ({new_AGEMA_signal_2479, KeyArray_outS03ser[4]}), .c ({new_AGEMA_signal_2480, KeyArray_inS02ser[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS02ser_mux_inst_5_U1 ( .s (KeyArray_n45), .b ({key_s1[109], key_s0[109]}), .a ({new_AGEMA_signal_2482, KeyArray_outS03ser[5]}), .c ({new_AGEMA_signal_2483, KeyArray_inS02ser[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS02ser_mux_inst_6_U1 ( .s (KeyArray_n45), .b ({key_s1[110], key_s0[110]}), .a ({new_AGEMA_signal_2485, KeyArray_outS03ser[6]}), .c ({new_AGEMA_signal_2486, KeyArray_inS02ser[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS02ser_mux_inst_7_U1 ( .s (KeyArray_n45), .b ({key_s1[111], key_s0[111]}), .a ({new_AGEMA_signal_2488, KeyArray_outS03ser[7]}), .c ({new_AGEMA_signal_2489, KeyArray_inS02ser[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS03ser_mux_inst_0_U1 ( .s (KeyArray_n45), .b ({key_s1[96], key_s0[96]}), .a ({new_AGEMA_signal_2491, KeyArray_outS10ser[0]}), .c ({new_AGEMA_signal_2492, KeyArray_inS03ser[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS03ser_mux_inst_1_U1 ( .s (KeyArray_n45), .b ({key_s1[97], key_s0[97]}), .a ({new_AGEMA_signal_2494, KeyArray_outS10ser[1]}), .c ({new_AGEMA_signal_2495, KeyArray_inS03ser[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS03ser_mux_inst_2_U1 ( .s (KeyArray_n45), .b ({key_s1[98], key_s0[98]}), .a ({new_AGEMA_signal_2497, KeyArray_outS10ser[2]}), .c ({new_AGEMA_signal_2498, KeyArray_inS03ser[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS03ser_mux_inst_3_U1 ( .s (KeyArray_n45), .b ({key_s1[99], key_s0[99]}), .a ({new_AGEMA_signal_2500, KeyArray_outS10ser[3]}), .c ({new_AGEMA_signal_2501, KeyArray_inS03ser[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS03ser_mux_inst_4_U1 ( .s (KeyArray_n45), .b ({key_s1[100], key_s0[100]}), .a ({new_AGEMA_signal_2503, KeyArray_outS10ser[4]}), .c ({new_AGEMA_signal_2504, KeyArray_inS03ser[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS03ser_mux_inst_5_U1 ( .s (KeyArray_n45), .b ({key_s1[101], key_s0[101]}), .a ({new_AGEMA_signal_2506, KeyArray_outS10ser[5]}), .c ({new_AGEMA_signal_2507, KeyArray_inS03ser[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS03ser_mux_inst_6_U1 ( .s (KeyArray_n45), .b ({key_s1[102], key_s0[102]}), .a ({new_AGEMA_signal_2509, KeyArray_outS10ser[6]}), .c ({new_AGEMA_signal_2510, KeyArray_inS03ser[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS03ser_mux_inst_7_U1 ( .s (KeyArray_n45), .b ({key_s1[103], key_s0[103]}), .a ({new_AGEMA_signal_2512, KeyArray_outS10ser[7]}), .c ({new_AGEMA_signal_2513, KeyArray_inS03ser[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS10ser_mux_inst_0_U1 ( .s (KeyArray_n44), .b ({key_s1[88], key_s0[88]}), .a ({new_AGEMA_signal_2515, KeyArray_outS11ser[0]}), .c ({new_AGEMA_signal_2516, KeyArray_inS10ser[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS10ser_mux_inst_1_U1 ( .s (KeyArray_n44), .b ({key_s1[89], key_s0[89]}), .a ({new_AGEMA_signal_2518, KeyArray_outS11ser[1]}), .c ({new_AGEMA_signal_2519, KeyArray_inS10ser[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS10ser_mux_inst_2_U1 ( .s (KeyArray_n44), .b ({key_s1[90], key_s0[90]}), .a ({new_AGEMA_signal_2521, KeyArray_outS11ser[2]}), .c ({new_AGEMA_signal_2522, KeyArray_inS10ser[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS10ser_mux_inst_3_U1 ( .s (KeyArray_n44), .b ({key_s1[91], key_s0[91]}), .a ({new_AGEMA_signal_2524, KeyArray_outS11ser[3]}), .c ({new_AGEMA_signal_2525, KeyArray_inS10ser[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS10ser_mux_inst_4_U1 ( .s (KeyArray_n44), .b ({key_s1[92], key_s0[92]}), .a ({new_AGEMA_signal_2527, KeyArray_outS11ser[4]}), .c ({new_AGEMA_signal_2528, KeyArray_inS10ser[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS10ser_mux_inst_5_U1 ( .s (KeyArray_n44), .b ({key_s1[93], key_s0[93]}), .a ({new_AGEMA_signal_2530, KeyArray_outS11ser[5]}), .c ({new_AGEMA_signal_2531, KeyArray_inS10ser[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS10ser_mux_inst_6_U1 ( .s (KeyArray_n44), .b ({key_s1[94], key_s0[94]}), .a ({new_AGEMA_signal_2533, KeyArray_outS11ser[6]}), .c ({new_AGEMA_signal_2534, KeyArray_inS10ser[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS10ser_mux_inst_7_U1 ( .s (KeyArray_n44), .b ({key_s1[95], key_s0[95]}), .a ({new_AGEMA_signal_2536, KeyArray_outS11ser[7]}), .c ({new_AGEMA_signal_2537, KeyArray_inS10ser[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS11ser_mux_inst_0_U1 ( .s (KeyArray_n44), .b ({key_s1[80], key_s0[80]}), .a ({new_AGEMA_signal_2539, KeyArray_outS12ser[0]}), .c ({new_AGEMA_signal_2540, KeyArray_inS11ser[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS11ser_mux_inst_1_U1 ( .s (KeyArray_n44), .b ({key_s1[81], key_s0[81]}), .a ({new_AGEMA_signal_2542, KeyArray_outS12ser[1]}), .c ({new_AGEMA_signal_2543, KeyArray_inS11ser[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS11ser_mux_inst_2_U1 ( .s (KeyArray_n44), .b ({key_s1[82], key_s0[82]}), .a ({new_AGEMA_signal_2545, KeyArray_outS12ser[2]}), .c ({new_AGEMA_signal_2546, KeyArray_inS11ser[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS11ser_mux_inst_3_U1 ( .s (KeyArray_n44), .b ({key_s1[83], key_s0[83]}), .a ({new_AGEMA_signal_2548, KeyArray_outS12ser[3]}), .c ({new_AGEMA_signal_2549, KeyArray_inS11ser[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS11ser_mux_inst_4_U1 ( .s (KeyArray_n44), .b ({key_s1[84], key_s0[84]}), .a ({new_AGEMA_signal_2551, KeyArray_outS12ser[4]}), .c ({new_AGEMA_signal_2552, KeyArray_inS11ser[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS11ser_mux_inst_5_U1 ( .s (KeyArray_n44), .b ({key_s1[85], key_s0[85]}), .a ({new_AGEMA_signal_2554, KeyArray_outS12ser[5]}), .c ({new_AGEMA_signal_2555, KeyArray_inS11ser[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS11ser_mux_inst_6_U1 ( .s (KeyArray_n44), .b ({key_s1[86], key_s0[86]}), .a ({new_AGEMA_signal_2557, KeyArray_outS12ser[6]}), .c ({new_AGEMA_signal_2558, KeyArray_inS11ser[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS11ser_mux_inst_7_U1 ( .s (KeyArray_n44), .b ({key_s1[87], key_s0[87]}), .a ({new_AGEMA_signal_2560, KeyArray_outS12ser[7]}), .c ({new_AGEMA_signal_2561, KeyArray_inS11ser[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS12ser_mux_inst_0_U1 ( .s (KeyArray_n43), .b ({key_s1[72], key_s0[72]}), .a ({new_AGEMA_signal_2563, keySBIn[0]}), .c ({new_AGEMA_signal_2564, KeyArray_inS12ser[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS12ser_mux_inst_1_U1 ( .s (KeyArray_n43), .b ({key_s1[73], key_s0[73]}), .a ({new_AGEMA_signal_2566, keySBIn[1]}), .c ({new_AGEMA_signal_2567, KeyArray_inS12ser[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS12ser_mux_inst_2_U1 ( .s (KeyArray_n43), .b ({key_s1[74], key_s0[74]}), .a ({new_AGEMA_signal_2569, keySBIn[2]}), .c ({new_AGEMA_signal_2570, KeyArray_inS12ser[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS12ser_mux_inst_3_U1 ( .s (KeyArray_n43), .b ({key_s1[75], key_s0[75]}), .a ({new_AGEMA_signal_2572, keySBIn[3]}), .c ({new_AGEMA_signal_2573, KeyArray_inS12ser[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS12ser_mux_inst_4_U1 ( .s (KeyArray_n43), .b ({key_s1[76], key_s0[76]}), .a ({new_AGEMA_signal_2575, keySBIn[4]}), .c ({new_AGEMA_signal_2576, KeyArray_inS12ser[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS12ser_mux_inst_5_U1 ( .s (KeyArray_n43), .b ({key_s1[77], key_s0[77]}), .a ({new_AGEMA_signal_2578, keySBIn[5]}), .c ({new_AGEMA_signal_2579, KeyArray_inS12ser[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS12ser_mux_inst_6_U1 ( .s (KeyArray_n43), .b ({key_s1[78], key_s0[78]}), .a ({new_AGEMA_signal_2581, keySBIn[6]}), .c ({new_AGEMA_signal_2582, KeyArray_inS12ser[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS12ser_mux_inst_7_U1 ( .s (KeyArray_n43), .b ({key_s1[79], key_s0[79]}), .a ({new_AGEMA_signal_2584, keySBIn[7]}), .c ({new_AGEMA_signal_2585, KeyArray_inS12ser[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS13ser_mux_inst_0_U1 ( .s (KeyArray_n43), .b ({key_s1[64], key_s0[64]}), .a ({new_AGEMA_signal_2587, KeyArray_outS20ser[0]}), .c ({new_AGEMA_signal_2588, KeyArray_inS13ser[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS13ser_mux_inst_1_U1 ( .s (KeyArray_n43), .b ({key_s1[65], key_s0[65]}), .a ({new_AGEMA_signal_2590, KeyArray_outS20ser[1]}), .c ({new_AGEMA_signal_2591, KeyArray_inS13ser[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS13ser_mux_inst_2_U1 ( .s (KeyArray_n43), .b ({key_s1[66], key_s0[66]}), .a ({new_AGEMA_signal_2593, KeyArray_outS20ser[2]}), .c ({new_AGEMA_signal_2594, KeyArray_inS13ser[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS13ser_mux_inst_3_U1 ( .s (KeyArray_n43), .b ({key_s1[67], key_s0[67]}), .a ({new_AGEMA_signal_2596, KeyArray_outS20ser[3]}), .c ({new_AGEMA_signal_2597, KeyArray_inS13ser[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS13ser_mux_inst_4_U1 ( .s (KeyArray_n43), .b ({key_s1[68], key_s0[68]}), .a ({new_AGEMA_signal_2599, KeyArray_outS20ser[4]}), .c ({new_AGEMA_signal_2600, KeyArray_inS13ser[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS13ser_mux_inst_5_U1 ( .s (KeyArray_n43), .b ({key_s1[69], key_s0[69]}), .a ({new_AGEMA_signal_2602, KeyArray_outS20ser[5]}), .c ({new_AGEMA_signal_2603, KeyArray_inS13ser[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS13ser_mux_inst_6_U1 ( .s (KeyArray_n43), .b ({key_s1[70], key_s0[70]}), .a ({new_AGEMA_signal_2605, KeyArray_outS20ser[6]}), .c ({new_AGEMA_signal_2606, KeyArray_inS13ser[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS13ser_mux_inst_7_U1 ( .s (KeyArray_n43), .b ({key_s1[71], key_s0[71]}), .a ({new_AGEMA_signal_2608, KeyArray_outS20ser[7]}), .c ({new_AGEMA_signal_2609, KeyArray_inS13ser[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS20ser_mux_inst_0_U1 ( .s (KeyArray_n42), .b ({key_s1[56], key_s0[56]}), .a ({new_AGEMA_signal_2611, KeyArray_outS21ser[0]}), .c ({new_AGEMA_signal_2612, KeyArray_inS20ser[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS20ser_mux_inst_1_U1 ( .s (KeyArray_n42), .b ({key_s1[57], key_s0[57]}), .a ({new_AGEMA_signal_2614, KeyArray_outS21ser[1]}), .c ({new_AGEMA_signal_2615, KeyArray_inS20ser[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS20ser_mux_inst_2_U1 ( .s (KeyArray_n42), .b ({key_s1[58], key_s0[58]}), .a ({new_AGEMA_signal_2617, KeyArray_outS21ser[2]}), .c ({new_AGEMA_signal_2618, KeyArray_inS20ser[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS20ser_mux_inst_3_U1 ( .s (KeyArray_n42), .b ({key_s1[59], key_s0[59]}), .a ({new_AGEMA_signal_2620, KeyArray_outS21ser[3]}), .c ({new_AGEMA_signal_2621, KeyArray_inS20ser[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS20ser_mux_inst_4_U1 ( .s (KeyArray_n42), .b ({key_s1[60], key_s0[60]}), .a ({new_AGEMA_signal_2623, KeyArray_outS21ser[4]}), .c ({new_AGEMA_signal_2624, KeyArray_inS20ser[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS20ser_mux_inst_5_U1 ( .s (KeyArray_n42), .b ({key_s1[61], key_s0[61]}), .a ({new_AGEMA_signal_2626, KeyArray_outS21ser[5]}), .c ({new_AGEMA_signal_2627, KeyArray_inS20ser[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS20ser_mux_inst_6_U1 ( .s (KeyArray_n42), .b ({key_s1[62], key_s0[62]}), .a ({new_AGEMA_signal_2629, KeyArray_outS21ser[6]}), .c ({new_AGEMA_signal_2630, KeyArray_inS20ser[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS20ser_mux_inst_7_U1 ( .s (KeyArray_n42), .b ({key_s1[63], key_s0[63]}), .a ({new_AGEMA_signal_2632, KeyArray_outS21ser[7]}), .c ({new_AGEMA_signal_2633, KeyArray_inS20ser[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS21ser_mux_inst_0_U1 ( .s (KeyArray_n42), .b ({key_s1[48], key_s0[48]}), .a ({new_AGEMA_signal_2635, KeyArray_outS22ser[0]}), .c ({new_AGEMA_signal_2636, KeyArray_inS21ser[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS21ser_mux_inst_1_U1 ( .s (KeyArray_n42), .b ({key_s1[49], key_s0[49]}), .a ({new_AGEMA_signal_2638, KeyArray_outS22ser[1]}), .c ({new_AGEMA_signal_2639, KeyArray_inS21ser[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS21ser_mux_inst_2_U1 ( .s (KeyArray_n42), .b ({key_s1[50], key_s0[50]}), .a ({new_AGEMA_signal_2641, KeyArray_outS22ser[2]}), .c ({new_AGEMA_signal_2642, KeyArray_inS21ser[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS21ser_mux_inst_3_U1 ( .s (KeyArray_n42), .b ({key_s1[51], key_s0[51]}), .a ({new_AGEMA_signal_2644, KeyArray_outS22ser[3]}), .c ({new_AGEMA_signal_2645, KeyArray_inS21ser[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS21ser_mux_inst_4_U1 ( .s (KeyArray_n42), .b ({key_s1[52], key_s0[52]}), .a ({new_AGEMA_signal_2647, KeyArray_outS22ser[4]}), .c ({new_AGEMA_signal_2648, KeyArray_inS21ser[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS21ser_mux_inst_5_U1 ( .s (KeyArray_n42), .b ({key_s1[53], key_s0[53]}), .a ({new_AGEMA_signal_2650, KeyArray_outS22ser[5]}), .c ({new_AGEMA_signal_2651, KeyArray_inS21ser[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS21ser_mux_inst_6_U1 ( .s (KeyArray_n42), .b ({key_s1[54], key_s0[54]}), .a ({new_AGEMA_signal_2653, KeyArray_outS22ser[6]}), .c ({new_AGEMA_signal_2654, KeyArray_inS21ser[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS21ser_mux_inst_7_U1 ( .s (KeyArray_n42), .b ({key_s1[55], key_s0[55]}), .a ({new_AGEMA_signal_2656, KeyArray_outS22ser[7]}), .c ({new_AGEMA_signal_2657, KeyArray_inS21ser[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS22ser_mux_inst_0_U1 ( .s (KeyArray_n41), .b ({key_s1[40], key_s0[40]}), .a ({new_AGEMA_signal_2659, KeyArray_outS23ser[0]}), .c ({new_AGEMA_signal_2660, KeyArray_inS22ser[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS22ser_mux_inst_1_U1 ( .s (KeyArray_n41), .b ({key_s1[41], key_s0[41]}), .a ({new_AGEMA_signal_2662, KeyArray_outS23ser[1]}), .c ({new_AGEMA_signal_2663, KeyArray_inS22ser[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS22ser_mux_inst_2_U1 ( .s (KeyArray_n41), .b ({key_s1[42], key_s0[42]}), .a ({new_AGEMA_signal_2665, KeyArray_outS23ser[2]}), .c ({new_AGEMA_signal_2666, KeyArray_inS22ser[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS22ser_mux_inst_3_U1 ( .s (KeyArray_n41), .b ({key_s1[43], key_s0[43]}), .a ({new_AGEMA_signal_2668, KeyArray_outS23ser[3]}), .c ({new_AGEMA_signal_2669, KeyArray_inS22ser[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS22ser_mux_inst_4_U1 ( .s (KeyArray_n41), .b ({key_s1[44], key_s0[44]}), .a ({new_AGEMA_signal_2671, KeyArray_outS23ser[4]}), .c ({new_AGEMA_signal_2672, KeyArray_inS22ser[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS22ser_mux_inst_5_U1 ( .s (KeyArray_n41), .b ({key_s1[45], key_s0[45]}), .a ({new_AGEMA_signal_2674, KeyArray_outS23ser[5]}), .c ({new_AGEMA_signal_2675, KeyArray_inS22ser[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS22ser_mux_inst_6_U1 ( .s (KeyArray_n41), .b ({key_s1[46], key_s0[46]}), .a ({new_AGEMA_signal_2677, KeyArray_outS23ser[6]}), .c ({new_AGEMA_signal_2678, KeyArray_inS22ser[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS22ser_mux_inst_7_U1 ( .s (KeyArray_n41), .b ({key_s1[47], key_s0[47]}), .a ({new_AGEMA_signal_2680, KeyArray_outS23ser[7]}), .c ({new_AGEMA_signal_2681, KeyArray_inS22ser[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS23ser_mux_inst_0_U1 ( .s (KeyArray_n41), .b ({key_s1[32], key_s0[32]}), .a ({new_AGEMA_signal_2683, KeyArray_outS30ser[0]}), .c ({new_AGEMA_signal_2684, KeyArray_inS23ser[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS23ser_mux_inst_1_U1 ( .s (KeyArray_n41), .b ({key_s1[33], key_s0[33]}), .a ({new_AGEMA_signal_2686, KeyArray_outS30ser[1]}), .c ({new_AGEMA_signal_2687, KeyArray_inS23ser[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS23ser_mux_inst_2_U1 ( .s (KeyArray_n41), .b ({key_s1[34], key_s0[34]}), .a ({new_AGEMA_signal_2689, KeyArray_outS30ser[2]}), .c ({new_AGEMA_signal_2690, KeyArray_inS23ser[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS23ser_mux_inst_3_U1 ( .s (KeyArray_n41), .b ({key_s1[35], key_s0[35]}), .a ({new_AGEMA_signal_2692, KeyArray_outS30ser[3]}), .c ({new_AGEMA_signal_2693, KeyArray_inS23ser[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS23ser_mux_inst_4_U1 ( .s (KeyArray_n41), .b ({key_s1[36], key_s0[36]}), .a ({new_AGEMA_signal_2695, KeyArray_outS30ser[4]}), .c ({new_AGEMA_signal_2696, KeyArray_inS23ser[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS23ser_mux_inst_5_U1 ( .s (KeyArray_n41), .b ({key_s1[37], key_s0[37]}), .a ({new_AGEMA_signal_2698, KeyArray_outS30ser[5]}), .c ({new_AGEMA_signal_2699, KeyArray_inS23ser[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS23ser_mux_inst_6_U1 ( .s (KeyArray_n41), .b ({key_s1[38], key_s0[38]}), .a ({new_AGEMA_signal_2701, KeyArray_outS30ser[6]}), .c ({new_AGEMA_signal_2702, KeyArray_inS23ser[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS23ser_mux_inst_7_U1 ( .s (KeyArray_n41), .b ({key_s1[39], key_s0[39]}), .a ({new_AGEMA_signal_2704, KeyArray_outS30ser[7]}), .c ({new_AGEMA_signal_2705, KeyArray_inS23ser[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS30ser_mux_inst_0_U1 ( .s (KeyArray_n40), .b ({key_s1[24], key_s0[24]}), .a ({new_AGEMA_signal_2707, KeyArray_outS31ser[0]}), .c ({new_AGEMA_signal_2708, KeyArray_inS30ser[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS30ser_mux_inst_1_U1 ( .s (KeyArray_n40), .b ({key_s1[25], key_s0[25]}), .a ({new_AGEMA_signal_2710, KeyArray_outS31ser[1]}), .c ({new_AGEMA_signal_2711, KeyArray_inS30ser[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS30ser_mux_inst_2_U1 ( .s (KeyArray_n40), .b ({key_s1[26], key_s0[26]}), .a ({new_AGEMA_signal_2713, KeyArray_outS31ser[2]}), .c ({new_AGEMA_signal_2714, KeyArray_inS30ser[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS30ser_mux_inst_3_U1 ( .s (KeyArray_n40), .b ({key_s1[27], key_s0[27]}), .a ({new_AGEMA_signal_2716, KeyArray_outS31ser[3]}), .c ({new_AGEMA_signal_2717, KeyArray_inS30ser[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS30ser_mux_inst_4_U1 ( .s (KeyArray_n40), .b ({key_s1[28], key_s0[28]}), .a ({new_AGEMA_signal_2719, KeyArray_outS31ser[4]}), .c ({new_AGEMA_signal_2720, KeyArray_inS30ser[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS30ser_mux_inst_5_U1 ( .s (KeyArray_n40), .b ({key_s1[29], key_s0[29]}), .a ({new_AGEMA_signal_2722, KeyArray_outS31ser[5]}), .c ({new_AGEMA_signal_2723, KeyArray_inS30ser[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS30ser_mux_inst_6_U1 ( .s (KeyArray_n40), .b ({key_s1[30], key_s0[30]}), .a ({new_AGEMA_signal_2725, KeyArray_outS31ser[6]}), .c ({new_AGEMA_signal_2726, KeyArray_inS30ser[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS30ser_mux_inst_7_U1 ( .s (KeyArray_n40), .b ({key_s1[31], key_s0[31]}), .a ({new_AGEMA_signal_2728, KeyArray_outS31ser[7]}), .c ({new_AGEMA_signal_2729, KeyArray_inS30ser[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS31ser_mux_inst_0_U1 ( .s (KeyArray_n40), .b ({key_s1[16], key_s0[16]}), .a ({new_AGEMA_signal_2731, KeyArray_outS32ser[0]}), .c ({new_AGEMA_signal_2732, KeyArray_inS31ser[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS31ser_mux_inst_1_U1 ( .s (KeyArray_n40), .b ({key_s1[17], key_s0[17]}), .a ({new_AGEMA_signal_2734, KeyArray_outS32ser[1]}), .c ({new_AGEMA_signal_2735, KeyArray_inS31ser[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS31ser_mux_inst_2_U1 ( .s (KeyArray_n40), .b ({key_s1[18], key_s0[18]}), .a ({new_AGEMA_signal_2737, KeyArray_outS32ser[2]}), .c ({new_AGEMA_signal_2738, KeyArray_inS31ser[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS31ser_mux_inst_3_U1 ( .s (KeyArray_n40), .b ({key_s1[19], key_s0[19]}), .a ({new_AGEMA_signal_2740, KeyArray_outS32ser[3]}), .c ({new_AGEMA_signal_2741, KeyArray_inS31ser[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS31ser_mux_inst_4_U1 ( .s (KeyArray_n40), .b ({key_s1[20], key_s0[20]}), .a ({new_AGEMA_signal_2743, KeyArray_outS32ser[4]}), .c ({new_AGEMA_signal_2744, KeyArray_inS31ser[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS31ser_mux_inst_5_U1 ( .s (KeyArray_n40), .b ({key_s1[21], key_s0[21]}), .a ({new_AGEMA_signal_2746, KeyArray_outS32ser[5]}), .c ({new_AGEMA_signal_2747, KeyArray_inS31ser[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS31ser_mux_inst_6_U1 ( .s (KeyArray_n40), .b ({key_s1[22], key_s0[22]}), .a ({new_AGEMA_signal_2749, KeyArray_outS32ser[6]}), .c ({new_AGEMA_signal_2750, KeyArray_inS31ser[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS31ser_mux_inst_7_U1 ( .s (KeyArray_n40), .b ({key_s1[23], key_s0[23]}), .a ({new_AGEMA_signal_2752, KeyArray_outS32ser[7]}), .c ({new_AGEMA_signal_2753, KeyArray_inS31ser[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS32ser_mux_inst_0_U1 ( .s (KeyArray_n39), .b ({key_s1[8], key_s0[8]}), .a ({new_AGEMA_signal_2755, KeyArray_outS33ser[0]}), .c ({new_AGEMA_signal_2756, KeyArray_inS32ser[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS32ser_mux_inst_1_U1 ( .s (KeyArray_n39), .b ({key_s1[9], key_s0[9]}), .a ({new_AGEMA_signal_2758, KeyArray_outS33ser[1]}), .c ({new_AGEMA_signal_2759, KeyArray_inS32ser[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS32ser_mux_inst_2_U1 ( .s (KeyArray_n39), .b ({key_s1[10], key_s0[10]}), .a ({new_AGEMA_signal_2761, KeyArray_outS33ser[2]}), .c ({new_AGEMA_signal_2762, KeyArray_inS32ser[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS32ser_mux_inst_3_U1 ( .s (KeyArray_n39), .b ({key_s1[11], key_s0[11]}), .a ({new_AGEMA_signal_2764, KeyArray_outS33ser[3]}), .c ({new_AGEMA_signal_2765, KeyArray_inS32ser[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS32ser_mux_inst_4_U1 ( .s (KeyArray_n39), .b ({key_s1[12], key_s0[12]}), .a ({new_AGEMA_signal_2767, KeyArray_outS33ser[4]}), .c ({new_AGEMA_signal_2768, KeyArray_inS32ser[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS32ser_mux_inst_5_U1 ( .s (KeyArray_n39), .b ({key_s1[13], key_s0[13]}), .a ({new_AGEMA_signal_2770, KeyArray_outS33ser[5]}), .c ({new_AGEMA_signal_2771, KeyArray_inS32ser[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS32ser_mux_inst_6_U1 ( .s (KeyArray_n39), .b ({key_s1[14], key_s0[14]}), .a ({new_AGEMA_signal_2773, KeyArray_outS33ser[6]}), .c ({new_AGEMA_signal_2774, KeyArray_inS32ser[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS32ser_mux_inst_7_U1 ( .s (KeyArray_n39), .b ({key_s1[15], key_s0[15]}), .a ({new_AGEMA_signal_2776, KeyArray_outS33ser[7]}), .c ({new_AGEMA_signal_2777, KeyArray_inS32ser[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS33ser_mux_inst_0_U1 ( .s (KeyArray_n39), .b ({key_s1[0], key_s0[0]}), .a ({new_AGEMA_signal_1983, keyStateIn[0]}), .c ({new_AGEMA_signal_2779, KeyArray_inS33ser[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS33ser_mux_inst_1_U1 ( .s (KeyArray_n39), .b ({key_s1[1], key_s0[1]}), .a ({new_AGEMA_signal_1986, keyStateIn[1]}), .c ({new_AGEMA_signal_2781, KeyArray_inS33ser[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS33ser_mux_inst_2_U1 ( .s (KeyArray_n39), .b ({key_s1[2], key_s0[2]}), .a ({new_AGEMA_signal_1989, keyStateIn[2]}), .c ({new_AGEMA_signal_2783, KeyArray_inS33ser[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS33ser_mux_inst_3_U1 ( .s (KeyArray_n39), .b ({key_s1[3], key_s0[3]}), .a ({new_AGEMA_signal_1992, keyStateIn[3]}), .c ({new_AGEMA_signal_2785, KeyArray_inS33ser[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS33ser_mux_inst_4_U1 ( .s (KeyArray_n39), .b ({key_s1[4], key_s0[4]}), .a ({new_AGEMA_signal_1995, keyStateIn[4]}), .c ({new_AGEMA_signal_2787, KeyArray_inS33ser[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS33ser_mux_inst_5_U1 ( .s (KeyArray_n39), .b ({key_s1[5], key_s0[5]}), .a ({new_AGEMA_signal_1998, keyStateIn[5]}), .c ({new_AGEMA_signal_2789, KeyArray_inS33ser[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS33ser_mux_inst_6_U1 ( .s (KeyArray_n39), .b ({key_s1[6], key_s0[6]}), .a ({new_AGEMA_signal_2001, keyStateIn[6]}), .c ({new_AGEMA_signal_2791, KeyArray_inS33ser[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_MUX_inS33ser_mux_inst_7_U1 ( .s (KeyArray_n39), .b ({key_s1[7], key_s0[7]}), .a ({new_AGEMA_signal_2004, keyStateIn[7]}), .c ({new_AGEMA_signal_2793, KeyArray_inS33ser[7]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_U24 ( .a ({new_AGEMA_signal_2122, MixColumns_line0_n16}), .b ({new_AGEMA_signal_2024, MixColumns_line0_n15}), .c ({new_AGEMA_signal_2794, MCout[31]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_U23 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .c ({new_AGEMA_signal_2024, MixColumns_line0_n15}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_U22 ( .a ({ciphertext_s1[126], ciphertext_s0[126]}), .b ({new_AGEMA_signal_2051, MixColumns_line0_S13[7]}), .c ({new_AGEMA_signal_2122, MixColumns_line0_n16}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_U21 ( .a ({new_AGEMA_signal_2123, MixColumns_line0_n14}), .b ({new_AGEMA_signal_2027, MixColumns_line0_n13}), .c ({new_AGEMA_signal_2795, MCout[30]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_U20 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({ciphertext_s1[30], ciphertext_s0[30]}), .c ({new_AGEMA_signal_2027, MixColumns_line0_n13}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_U19 ( .a ({ciphertext_s1[125], ciphertext_s0[125]}), .b ({new_AGEMA_signal_2053, MixColumns_line0_S13[6]}), .c ({new_AGEMA_signal_2123, MixColumns_line0_n14}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_U18 ( .a ({new_AGEMA_signal_2124, MixColumns_line0_n12}), .b ({new_AGEMA_signal_2030, MixColumns_line0_n11}), .c ({new_AGEMA_signal_2796, MCout[29]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_U17 ( .a ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({ciphertext_s1[29], ciphertext_s0[29]}), .c ({new_AGEMA_signal_2030, MixColumns_line0_n11}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_U16 ( .a ({ciphertext_s1[124], ciphertext_s0[124]}), .b ({new_AGEMA_signal_2055, MixColumns_line0_S13[5]}), .c ({new_AGEMA_signal_2124, MixColumns_line0_n12}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_U15 ( .a ({new_AGEMA_signal_2797, MixColumns_line0_n10}), .b ({new_AGEMA_signal_2033, MixColumns_line0_n9}), .c ({new_AGEMA_signal_2838, MCout[28]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_U14 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({ciphertext_s1[28], ciphertext_s0[28]}), .c ({new_AGEMA_signal_2033, MixColumns_line0_n9}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_U13 ( .a ({new_AGEMA_signal_2046, MixColumns_line0_S02[4]}), .b ({new_AGEMA_signal_2127, MixColumns_line0_S13[4]}), .c ({new_AGEMA_signal_2797, MixColumns_line0_n10}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_U12 ( .a ({new_AGEMA_signal_2798, MixColumns_line0_n8}), .b ({new_AGEMA_signal_2036, MixColumns_line0_n7}), .c ({new_AGEMA_signal_2839, MCout[27]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_U11 ( .a ({ciphertext_s1[59], ciphertext_s0[59]}), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .c ({new_AGEMA_signal_2036, MixColumns_line0_n7}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_U10 ( .a ({new_AGEMA_signal_2047, MixColumns_line0_S02[3]}), .b ({new_AGEMA_signal_2128, MixColumns_line0_S13[3]}), .c ({new_AGEMA_signal_2798, MixColumns_line0_n8}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_U9 ( .a ({new_AGEMA_signal_2125, MixColumns_line0_n6}), .b ({new_AGEMA_signal_2039, MixColumns_line0_n5}), .c ({new_AGEMA_signal_2799, MCout[26]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_U8 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_2039, MixColumns_line0_n5}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_U7 ( .a ({ciphertext_s1[121], ciphertext_s0[121]}), .b ({new_AGEMA_signal_2058, MixColumns_line0_S13[2]}), .c ({new_AGEMA_signal_2125, MixColumns_line0_n6}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_U6 ( .a ({new_AGEMA_signal_2800, MixColumns_line0_n4}), .b ({new_AGEMA_signal_2042, MixColumns_line0_n3}), .c ({new_AGEMA_signal_2840, MCout[25]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_U5 ( .a ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({ciphertext_s1[57], ciphertext_s0[57]}), .c ({new_AGEMA_signal_2042, MixColumns_line0_n3}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_U4 ( .a ({new_AGEMA_signal_2048, MixColumns_line0_S02[1]}), .b ({new_AGEMA_signal_2129, MixColumns_line0_S13[1]}), .c ({new_AGEMA_signal_2800, MixColumns_line0_n4}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_U3 ( .a ({new_AGEMA_signal_2126, MixColumns_line0_n2}), .b ({new_AGEMA_signal_2045, MixColumns_line0_n1}), .c ({new_AGEMA_signal_2801, MCout[24]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_U2 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .c ({new_AGEMA_signal_2045, MixColumns_line0_n1}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_U1 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({new_AGEMA_signal_2060, MixColumns_line0_S13[0]}), .c ({new_AGEMA_signal_2126, MixColumns_line0_n2}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_timesTWO_U3 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[123], ciphertext_s0[123]}), .c ({new_AGEMA_signal_2046, MixColumns_line0_S02[4]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_timesTWO_U2 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_2047, MixColumns_line0_S02[3]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_timesTWO_U1 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[120], ciphertext_s0[120]}), .c ({new_AGEMA_signal_2048, MixColumns_line0_S02[1]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_timesTHREE_U8 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[94], ciphertext_s0[94]}), .c ({new_AGEMA_signal_2051, MixColumns_line0_S13[7]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_timesTHREE_U7 ( .a ({ciphertext_s1[94], ciphertext_s0[94]}), .b ({ciphertext_s1[93], ciphertext_s0[93]}), .c ({new_AGEMA_signal_2053, MixColumns_line0_S13[6]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_timesTHREE_U6 ( .a ({ciphertext_s1[93], ciphertext_s0[93]}), .b ({ciphertext_s1[92], ciphertext_s0[92]}), .c ({new_AGEMA_signal_2055, MixColumns_line0_S13[5]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_timesTHREE_U5 ( .a ({ciphertext_s1[92], ciphertext_s0[92]}), .b ({new_AGEMA_signal_2062, MixColumns_line0_timesTHREE_input2[4]}), .c ({new_AGEMA_signal_2127, MixColumns_line0_S13[4]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_timesTHREE_U4 ( .a ({ciphertext_s1[91], ciphertext_s0[91]}), .b ({new_AGEMA_signal_2063, MixColumns_line0_timesTHREE_input2[3]}), .c ({new_AGEMA_signal_2128, MixColumns_line0_S13[3]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_timesTHREE_U3 ( .a ({ciphertext_s1[90], ciphertext_s0[90]}), .b ({ciphertext_s1[89], ciphertext_s0[89]}), .c ({new_AGEMA_signal_2058, MixColumns_line0_S13[2]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_timesTHREE_U2 ( .a ({ciphertext_s1[89], ciphertext_s0[89]}), .b ({new_AGEMA_signal_2064, MixColumns_line0_timesTHREE_input2[1]}), .c ({new_AGEMA_signal_2129, MixColumns_line0_S13[1]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_timesTHREE_U1 ( .a ({ciphertext_s1[88], ciphertext_s0[88]}), .b ({ciphertext_s1[95], ciphertext_s0[95]}), .c ({new_AGEMA_signal_2060, MixColumns_line0_S13[0]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_timesTHREE_timesTWO_U3 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[91], ciphertext_s0[91]}), .c ({new_AGEMA_signal_2062, MixColumns_line0_timesTHREE_input2[4]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_timesTHREE_timesTWO_U2 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_2063, MixColumns_line0_timesTHREE_input2[3]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line0_timesTHREE_timesTWO_U1 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .c ({new_AGEMA_signal_2064, MixColumns_line0_timesTHREE_input2[1]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_U24 ( .a ({new_AGEMA_signal_2130, MixColumns_line1_n16}), .b ({new_AGEMA_signal_2065, MixColumns_line1_n15}), .c ({new_AGEMA_signal_2802, MCout[23]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_U23 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[127], ciphertext_s0[127]}), .c ({new_AGEMA_signal_2065, MixColumns_line1_n15}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_U22 ( .a ({ciphertext_s1[94], ciphertext_s0[94]}), .b ({new_AGEMA_signal_2076, MixColumns_line1_S13[7]}), .c ({new_AGEMA_signal_2130, MixColumns_line1_n16}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_U21 ( .a ({new_AGEMA_signal_2131, MixColumns_line1_n14}), .b ({new_AGEMA_signal_2066, MixColumns_line1_n13}), .c ({new_AGEMA_signal_2803, MCout[22]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_U20 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({ciphertext_s1[126], ciphertext_s0[126]}), .c ({new_AGEMA_signal_2066, MixColumns_line1_n13}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_U19 ( .a ({ciphertext_s1[93], ciphertext_s0[93]}), .b ({new_AGEMA_signal_2077, MixColumns_line1_S13[6]}), .c ({new_AGEMA_signal_2131, MixColumns_line1_n14}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_U18 ( .a ({new_AGEMA_signal_2132, MixColumns_line1_n12}), .b ({new_AGEMA_signal_2067, MixColumns_line1_n11}), .c ({new_AGEMA_signal_2804, MCout[21]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_U17 ( .a ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({ciphertext_s1[125], ciphertext_s0[125]}), .c ({new_AGEMA_signal_2067, MixColumns_line1_n11}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_U16 ( .a ({ciphertext_s1[92], ciphertext_s0[92]}), .b ({new_AGEMA_signal_2078, MixColumns_line1_S13[5]}), .c ({new_AGEMA_signal_2132, MixColumns_line1_n12}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_U15 ( .a ({new_AGEMA_signal_2805, MixColumns_line1_n10}), .b ({new_AGEMA_signal_2068, MixColumns_line1_n9}), .c ({new_AGEMA_signal_2841, MCout[20]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_U14 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({ciphertext_s1[124], ciphertext_s0[124]}), .c ({new_AGEMA_signal_2068, MixColumns_line1_n9}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_U13 ( .a ({new_AGEMA_signal_2073, MixColumns_line1_S02_4_}), .b ({new_AGEMA_signal_2135, MixColumns_line1_S13[4]}), .c ({new_AGEMA_signal_2805, MixColumns_line1_n10}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_U12 ( .a ({new_AGEMA_signal_2806, MixColumns_line1_n8}), .b ({new_AGEMA_signal_2069, MixColumns_line1_n7}), .c ({new_AGEMA_signal_2842, MCout[19]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_U11 ( .a ({ciphertext_s1[27], ciphertext_s0[27]}), .b ({ciphertext_s1[123], ciphertext_s0[123]}), .c ({new_AGEMA_signal_2069, MixColumns_line1_n7}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_U10 ( .a ({new_AGEMA_signal_2074, MixColumns_line1_S02_3_}), .b ({new_AGEMA_signal_2136, MixColumns_line1_S13[3]}), .c ({new_AGEMA_signal_2806, MixColumns_line1_n8}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_U9 ( .a ({new_AGEMA_signal_2133, MixColumns_line1_n6}), .b ({new_AGEMA_signal_2070, MixColumns_line1_n5}), .c ({new_AGEMA_signal_2807, MCout[18]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_U8 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_2070, MixColumns_line1_n5}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_U7 ( .a ({ciphertext_s1[89], ciphertext_s0[89]}), .b ({new_AGEMA_signal_2079, MixColumns_line1_S13[2]}), .c ({new_AGEMA_signal_2133, MixColumns_line1_n6}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_U6 ( .a ({new_AGEMA_signal_2808, MixColumns_line1_n4}), .b ({new_AGEMA_signal_2071, MixColumns_line1_n3}), .c ({new_AGEMA_signal_2843, MCout[17]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_U5 ( .a ({ciphertext_s1[121], ciphertext_s0[121]}), .b ({ciphertext_s1[25], ciphertext_s0[25]}), .c ({new_AGEMA_signal_2071, MixColumns_line1_n3}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_U4 ( .a ({new_AGEMA_signal_2075, MixColumns_line1_S02_1_}), .b ({new_AGEMA_signal_2137, MixColumns_line1_S13[1]}), .c ({new_AGEMA_signal_2808, MixColumns_line1_n4}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_U3 ( .a ({new_AGEMA_signal_2134, MixColumns_line1_n2}), .b ({new_AGEMA_signal_2072, MixColumns_line1_n1}), .c ({new_AGEMA_signal_2809, MCout[16]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_U2 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .c ({new_AGEMA_signal_2072, MixColumns_line1_n1}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_U1 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({new_AGEMA_signal_2080, MixColumns_line1_S13[0]}), .c ({new_AGEMA_signal_2134, MixColumns_line1_n2}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_timesTWO_U3 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[91], ciphertext_s0[91]}), .c ({new_AGEMA_signal_2073, MixColumns_line1_S02_4_}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_timesTWO_U2 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_2074, MixColumns_line1_S02_3_}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_timesTWO_U1 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .c ({new_AGEMA_signal_2075, MixColumns_line1_S02_1_}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_timesTHREE_U8 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[62], ciphertext_s0[62]}), .c ({new_AGEMA_signal_2076, MixColumns_line1_S13[7]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_timesTHREE_U7 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({ciphertext_s1[61], ciphertext_s0[61]}), .c ({new_AGEMA_signal_2077, MixColumns_line1_S13[6]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_timesTHREE_U6 ( .a ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({ciphertext_s1[60], ciphertext_s0[60]}), .c ({new_AGEMA_signal_2078, MixColumns_line1_S13[5]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_timesTHREE_U5 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({new_AGEMA_signal_2081, MixColumns_line1_timesTHREE_input2[4]}), .c ({new_AGEMA_signal_2135, MixColumns_line1_S13[4]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_timesTHREE_U4 ( .a ({ciphertext_s1[59], ciphertext_s0[59]}), .b ({new_AGEMA_signal_2082, MixColumns_line1_timesTHREE_input2[3]}), .c ({new_AGEMA_signal_2136, MixColumns_line1_S13[3]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_timesTHREE_U3 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({ciphertext_s1[57], ciphertext_s0[57]}), .c ({new_AGEMA_signal_2079, MixColumns_line1_S13[2]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_timesTHREE_U2 ( .a ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({new_AGEMA_signal_2083, MixColumns_line1_timesTHREE_input2[1]}), .c ({new_AGEMA_signal_2137, MixColumns_line1_S13[1]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_timesTHREE_U1 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .c ({new_AGEMA_signal_2080, MixColumns_line1_S13[0]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_timesTHREE_timesTWO_U3 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .c ({new_AGEMA_signal_2081, MixColumns_line1_timesTHREE_input2[4]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_timesTHREE_timesTWO_U2 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_2082, MixColumns_line1_timesTHREE_input2[3]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line1_timesTHREE_timesTWO_U1 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .c ({new_AGEMA_signal_2083, MixColumns_line1_timesTHREE_input2[1]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_U24 ( .a ({new_AGEMA_signal_2138, MixColumns_line2_n16}), .b ({new_AGEMA_signal_2084, MixColumns_line2_n15}), .c ({new_AGEMA_signal_2810, MCout[15]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_U23 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[95], ciphertext_s0[95]}), .c ({new_AGEMA_signal_2084, MixColumns_line2_n15}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_U22 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({new_AGEMA_signal_2095, MixColumns_line2_S13[7]}), .c ({new_AGEMA_signal_2138, MixColumns_line2_n16}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_U21 ( .a ({new_AGEMA_signal_2139, MixColumns_line2_n14}), .b ({new_AGEMA_signal_2085, MixColumns_line2_n13}), .c ({new_AGEMA_signal_2811, MCout[14]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_U20 ( .a ({ciphertext_s1[126], ciphertext_s0[126]}), .b ({ciphertext_s1[94], ciphertext_s0[94]}), .c ({new_AGEMA_signal_2085, MixColumns_line2_n13}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_U19 ( .a ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({new_AGEMA_signal_2096, MixColumns_line2_S13[6]}), .c ({new_AGEMA_signal_2139, MixColumns_line2_n14}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_U18 ( .a ({new_AGEMA_signal_2140, MixColumns_line2_n12}), .b ({new_AGEMA_signal_2086, MixColumns_line2_n11}), .c ({new_AGEMA_signal_2812, MCout[13]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_U17 ( .a ({ciphertext_s1[125], ciphertext_s0[125]}), .b ({ciphertext_s1[93], ciphertext_s0[93]}), .c ({new_AGEMA_signal_2086, MixColumns_line2_n11}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_U16 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({new_AGEMA_signal_2097, MixColumns_line2_S13[5]}), .c ({new_AGEMA_signal_2140, MixColumns_line2_n12}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_U15 ( .a ({new_AGEMA_signal_2813, MixColumns_line2_n10}), .b ({new_AGEMA_signal_2087, MixColumns_line2_n9}), .c ({new_AGEMA_signal_2844, MCout[12]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_U14 ( .a ({ciphertext_s1[124], ciphertext_s0[124]}), .b ({ciphertext_s1[92], ciphertext_s0[92]}), .c ({new_AGEMA_signal_2087, MixColumns_line2_n9}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_U13 ( .a ({new_AGEMA_signal_2092, MixColumns_line2_S02_4_}), .b ({new_AGEMA_signal_2143, MixColumns_line2_S13[4]}), .c ({new_AGEMA_signal_2813, MixColumns_line2_n10}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_U12 ( .a ({new_AGEMA_signal_2814, MixColumns_line2_n8}), .b ({new_AGEMA_signal_2088, MixColumns_line2_n7}), .c ({new_AGEMA_signal_2845, MCout[11]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_U11 ( .a ({ciphertext_s1[123], ciphertext_s0[123]}), .b ({ciphertext_s1[91], ciphertext_s0[91]}), .c ({new_AGEMA_signal_2088, MixColumns_line2_n7}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_U10 ( .a ({new_AGEMA_signal_2093, MixColumns_line2_S02_3_}), .b ({new_AGEMA_signal_2144, MixColumns_line2_S13[3]}), .c ({new_AGEMA_signal_2814, MixColumns_line2_n8}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_U9 ( .a ({new_AGEMA_signal_2141, MixColumns_line2_n6}), .b ({new_AGEMA_signal_2089, MixColumns_line2_n5}), .c ({new_AGEMA_signal_2815, MCout[10]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_U8 ( .a ({ciphertext_s1[122], ciphertext_s0[122]}), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_2089, MixColumns_line2_n5}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_U7 ( .a ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({new_AGEMA_signal_2098, MixColumns_line2_S13[2]}), .c ({new_AGEMA_signal_2141, MixColumns_line2_n6}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_U6 ( .a ({new_AGEMA_signal_2816, MixColumns_line2_n4}), .b ({new_AGEMA_signal_2090, MixColumns_line2_n3}), .c ({new_AGEMA_signal_2846, MCout[9]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_U5 ( .a ({ciphertext_s1[89], ciphertext_s0[89]}), .b ({ciphertext_s1[121], ciphertext_s0[121]}), .c ({new_AGEMA_signal_2090, MixColumns_line2_n3}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_U4 ( .a ({new_AGEMA_signal_2094, MixColumns_line2_S02_1_}), .b ({new_AGEMA_signal_2145, MixColumns_line2_S13[1]}), .c ({new_AGEMA_signal_2816, MixColumns_line2_n4}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_U3 ( .a ({new_AGEMA_signal_2142, MixColumns_line2_n2}), .b ({new_AGEMA_signal_2091, MixColumns_line2_n1}), .c ({new_AGEMA_signal_2817, MCout[8]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_U2 ( .a ({ciphertext_s1[88], ciphertext_s0[88]}), .b ({ciphertext_s1[120], ciphertext_s0[120]}), .c ({new_AGEMA_signal_2091, MixColumns_line2_n1}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_U1 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({new_AGEMA_signal_2099, MixColumns_line2_S13[0]}), .c ({new_AGEMA_signal_2142, MixColumns_line2_n2}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_timesTWO_U3 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .c ({new_AGEMA_signal_2092, MixColumns_line2_S02_4_}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_timesTWO_U2 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_2093, MixColumns_line2_S02_3_}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_timesTWO_U1 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .c ({new_AGEMA_signal_2094, MixColumns_line2_S02_1_}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_timesTHREE_U8 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[30], ciphertext_s0[30]}), .c ({new_AGEMA_signal_2095, MixColumns_line2_S13[7]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_timesTHREE_U7 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({ciphertext_s1[29], ciphertext_s0[29]}), .c ({new_AGEMA_signal_2096, MixColumns_line2_S13[6]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_timesTHREE_U6 ( .a ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({ciphertext_s1[28], ciphertext_s0[28]}), .c ({new_AGEMA_signal_2097, MixColumns_line2_S13[5]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_timesTHREE_U5 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({new_AGEMA_signal_2100, MixColumns_line2_timesTHREE_input2[4]}), .c ({new_AGEMA_signal_2143, MixColumns_line2_S13[4]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_timesTHREE_U4 ( .a ({ciphertext_s1[27], ciphertext_s0[27]}), .b ({new_AGEMA_signal_2101, MixColumns_line2_timesTHREE_input2[3]}), .c ({new_AGEMA_signal_2144, MixColumns_line2_S13[3]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_timesTHREE_U3 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({ciphertext_s1[25], ciphertext_s0[25]}), .c ({new_AGEMA_signal_2098, MixColumns_line2_S13[2]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_timesTHREE_U2 ( .a ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({new_AGEMA_signal_2102, MixColumns_line2_timesTHREE_input2[1]}), .c ({new_AGEMA_signal_2145, MixColumns_line2_S13[1]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_timesTHREE_U1 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .c ({new_AGEMA_signal_2099, MixColumns_line2_S13[0]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_timesTHREE_timesTWO_U3 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .c ({new_AGEMA_signal_2100, MixColumns_line2_timesTHREE_input2[4]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_timesTHREE_timesTWO_U2 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_2101, MixColumns_line2_timesTHREE_input2[3]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line2_timesTHREE_timesTWO_U1 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .c ({new_AGEMA_signal_2102, MixColumns_line2_timesTHREE_input2[1]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_U24 ( .a ({new_AGEMA_signal_2146, MixColumns_line3_n16}), .b ({new_AGEMA_signal_2103, MixColumns_line3_n15}), .c ({new_AGEMA_signal_2818, MCout[7]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_U23 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .c ({new_AGEMA_signal_2103, MixColumns_line3_n15}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_U22 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({new_AGEMA_signal_2114, MixColumns_line3_S13[7]}), .c ({new_AGEMA_signal_2146, MixColumns_line3_n16}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_U21 ( .a ({new_AGEMA_signal_2147, MixColumns_line3_n14}), .b ({new_AGEMA_signal_2104, MixColumns_line3_n13}), .c ({new_AGEMA_signal_2819, MCout[6]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_U20 ( .a ({ciphertext_s1[94], ciphertext_s0[94]}), .b ({ciphertext_s1[62], ciphertext_s0[62]}), .c ({new_AGEMA_signal_2104, MixColumns_line3_n13}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_U19 ( .a ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({new_AGEMA_signal_2115, MixColumns_line3_S13[6]}), .c ({new_AGEMA_signal_2147, MixColumns_line3_n14}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_U18 ( .a ({new_AGEMA_signal_2148, MixColumns_line3_n12}), .b ({new_AGEMA_signal_2105, MixColumns_line3_n11}), .c ({new_AGEMA_signal_2820, MCout[5]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_U17 ( .a ({ciphertext_s1[93], ciphertext_s0[93]}), .b ({ciphertext_s1[61], ciphertext_s0[61]}), .c ({new_AGEMA_signal_2105, MixColumns_line3_n11}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_U16 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({new_AGEMA_signal_2116, MixColumns_line3_S13[5]}), .c ({new_AGEMA_signal_2148, MixColumns_line3_n12}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_U15 ( .a ({new_AGEMA_signal_2821, MixColumns_line3_n10}), .b ({new_AGEMA_signal_2106, MixColumns_line3_n9}), .c ({new_AGEMA_signal_2847, MCout[4]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_U14 ( .a ({ciphertext_s1[92], ciphertext_s0[92]}), .b ({ciphertext_s1[60], ciphertext_s0[60]}), .c ({new_AGEMA_signal_2106, MixColumns_line3_n9}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_U13 ( .a ({new_AGEMA_signal_2111, MixColumns_line3_S02_4_}), .b ({new_AGEMA_signal_2151, MixColumns_line3_S13[4]}), .c ({new_AGEMA_signal_2821, MixColumns_line3_n10}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_U12 ( .a ({new_AGEMA_signal_2822, MixColumns_line3_n8}), .b ({new_AGEMA_signal_2107, MixColumns_line3_n7}), .c ({new_AGEMA_signal_2848, MCout[3]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_U11 ( .a ({ciphertext_s1[91], ciphertext_s0[91]}), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .c ({new_AGEMA_signal_2107, MixColumns_line3_n7}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_U10 ( .a ({new_AGEMA_signal_2112, MixColumns_line3_S02_3_}), .b ({new_AGEMA_signal_2152, MixColumns_line3_S13[3]}), .c ({new_AGEMA_signal_2822, MixColumns_line3_n8}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_U9 ( .a ({new_AGEMA_signal_2149, MixColumns_line3_n6}), .b ({new_AGEMA_signal_2108, MixColumns_line3_n5}), .c ({new_AGEMA_signal_2823, MCout[2]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_U8 ( .a ({ciphertext_s1[90], ciphertext_s0[90]}), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_2108, MixColumns_line3_n5}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_U7 ( .a ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({new_AGEMA_signal_2117, MixColumns_line3_S13[2]}), .c ({new_AGEMA_signal_2149, MixColumns_line3_n6}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_U6 ( .a ({new_AGEMA_signal_2824, MixColumns_line3_n4}), .b ({new_AGEMA_signal_2109, MixColumns_line3_n3}), .c ({new_AGEMA_signal_2849, MCout[1]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_U5 ( .a ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({ciphertext_s1[89], ciphertext_s0[89]}), .c ({new_AGEMA_signal_2109, MixColumns_line3_n3}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_U4 ( .a ({new_AGEMA_signal_2113, MixColumns_line3_S02_1_}), .b ({new_AGEMA_signal_2153, MixColumns_line3_S13[1]}), .c ({new_AGEMA_signal_2824, MixColumns_line3_n4}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_U3 ( .a ({new_AGEMA_signal_2150, MixColumns_line3_n2}), .b ({new_AGEMA_signal_2110, MixColumns_line3_n1}), .c ({new_AGEMA_signal_2825, MCout[0]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_U2 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .c ({new_AGEMA_signal_2110, MixColumns_line3_n1}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_U1 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({new_AGEMA_signal_2118, MixColumns_line3_S13[0]}), .c ({new_AGEMA_signal_2150, MixColumns_line3_n2}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_timesTWO_U3 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .c ({new_AGEMA_signal_2111, MixColumns_line3_S02_4_}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_timesTWO_U2 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_2112, MixColumns_line3_S02_3_}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_timesTWO_U1 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .c ({new_AGEMA_signal_2113, MixColumns_line3_S02_1_}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_timesTHREE_U8 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[126], ciphertext_s0[126]}), .c ({new_AGEMA_signal_2114, MixColumns_line3_S13[7]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_timesTHREE_U7 ( .a ({ciphertext_s1[126], ciphertext_s0[126]}), .b ({ciphertext_s1[125], ciphertext_s0[125]}), .c ({new_AGEMA_signal_2115, MixColumns_line3_S13[6]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_timesTHREE_U6 ( .a ({ciphertext_s1[125], ciphertext_s0[125]}), .b ({ciphertext_s1[124], ciphertext_s0[124]}), .c ({new_AGEMA_signal_2116, MixColumns_line3_S13[5]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_timesTHREE_U5 ( .a ({ciphertext_s1[124], ciphertext_s0[124]}), .b ({new_AGEMA_signal_2119, MixColumns_line3_timesTHREE_input2_4_}), .c ({new_AGEMA_signal_2151, MixColumns_line3_S13[4]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_timesTHREE_U4 ( .a ({ciphertext_s1[123], ciphertext_s0[123]}), .b ({new_AGEMA_signal_2120, MixColumns_line3_timesTHREE_input2_3_}), .c ({new_AGEMA_signal_2152, MixColumns_line3_S13[3]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_timesTHREE_U3 ( .a ({ciphertext_s1[122], ciphertext_s0[122]}), .b ({ciphertext_s1[121], ciphertext_s0[121]}), .c ({new_AGEMA_signal_2117, MixColumns_line3_S13[2]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_timesTHREE_U2 ( .a ({ciphertext_s1[121], ciphertext_s0[121]}), .b ({new_AGEMA_signal_2121, MixColumns_line3_timesTHREE_input2_1_}), .c ({new_AGEMA_signal_2153, MixColumns_line3_S13[1]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_timesTHREE_U1 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({ciphertext_s1[127], ciphertext_s0[127]}), .c ({new_AGEMA_signal_2118, MixColumns_line3_S13[0]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_timesTHREE_timesTWO_U3 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[123], ciphertext_s0[123]}), .c ({new_AGEMA_signal_2119, MixColumns_line3_timesTHREE_input2_4_}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_timesTHREE_timesTWO_U2 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_2120, MixColumns_line3_timesTHREE_input2_3_}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) MixColumns_line3_timesTHREE_timesTWO_U1 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[120], ciphertext_s0[120]}), .c ({new_AGEMA_signal_2121, MixColumns_line3_timesTHREE_input2_1_}) ) ;
    NOR2_X1 calcRCon_U46 ( .A1 (calcRCon_n11), .A2 (calcRCon_n38), .ZN (roundConstant[7]) ) ;
    NOR2_X1 calcRCon_U45 ( .A1 (calcRCon_n16), .A2 (calcRCon_n38), .ZN (roundConstant[6]) ) ;
    AND2_X1 calcRCon_U44 ( .A1 (calcRCon_s_current_state_5_), .A2 (enRCon), .ZN (roundConstant[5]) ) ;
    AND2_X1 calcRCon_U43 ( .A1 (calcRCon_s_current_state_4_), .A2 (enRCon), .ZN (roundConstant[4]) ) ;
    NOR2_X1 calcRCon_U42 ( .A1 (calcRCon_n15), .A2 (calcRCon_n38), .ZN (roundConstant[3]) ) ;
    NOR2_X1 calcRCon_U41 ( .A1 (calcRCon_n12), .A2 (calcRCon_n38), .ZN (roundConstant[2]) ) ;
    NOR2_X1 calcRCon_U40 ( .A1 (calcRCon_n14), .A2 (calcRCon_n38), .ZN (roundConstant[1]) ) ;
    NOR2_X1 calcRCon_U39 ( .A1 (calcRCon_n13), .A2 (calcRCon_n38), .ZN (roundConstant[0]) ) ;
    INV_X1 calcRCon_U38 ( .A (enRCon), .ZN (calcRCon_n38) ) ;
    NAND2_X1 calcRCon_U37 ( .A1 (calcRCon_n37), .A2 (calcRCon_n36), .ZN (notFirst) ) ;
    NOR2_X1 calcRCon_U36 ( .A1 (calcRCon_n35), .A2 (calcRCon_n34), .ZN (calcRCon_n36) ) ;
    NAND2_X1 calcRCon_U35 ( .A1 (calcRCon_n33), .A2 (calcRCon_n32), .ZN (calcRCon_n34) ) ;
    NOR2_X1 calcRCon_U34 ( .A1 (calcRCon_s_current_state_1_), .A2 (calcRCon_n15), .ZN (calcRCon_n32) ) ;
    NOR2_X1 calcRCon_U33 ( .A1 (calcRCon_s_current_state_6_), .A2 (calcRCon_n13), .ZN (calcRCon_n33) ) ;
    NAND2_X1 calcRCon_U32 ( .A1 (calcRCon_s_current_state_2_), .A2 (calcRCon_n3), .ZN (calcRCon_n35) ) ;
    NOR2_X1 calcRCon_U31 ( .A1 (calcRCon_s_current_state_4_), .A2 (calcRCon_s_current_state_5_), .ZN (calcRCon_n37) ) ;
    NAND2_X1 calcRCon_U30 ( .A1 (nReset), .A2 (calcRCon_n31), .ZN (calcRCon_n51) ) ;
    MUX2_X1 calcRCon_U29 ( .S (calcRCon_n5), .A (calcRCon_n11), .B (calcRCon_n13), .Z (calcRCon_n31) ) ;
    NAND2_X1 calcRCon_U28 ( .A1 (calcRCon_n30), .A2 (calcRCon_n29), .ZN (calcRCon_n50) ) ;
    NAND2_X1 calcRCon_U27 ( .A1 (calcRCon_n28), .A2 (calcRCon_s_current_state_1_), .ZN (calcRCon_n29) ) ;
    NAND2_X1 calcRCon_U26 ( .A1 (calcRCon_n27), .A2 (calcRCon_n26), .ZN (calcRCon_n30) ) ;
    XOR2_X1 calcRCon_U25 ( .A (calcRCon_s_current_state_0_), .B (calcRCon_n3), .Z (calcRCon_n27) ) ;
    NAND2_X1 calcRCon_U24 ( .A1 (nReset), .A2 (calcRCon_n25), .ZN (calcRCon_n49) ) ;
    MUX2_X1 calcRCon_U23 ( .S (calcRCon_n5), .A (calcRCon_n14), .B (calcRCon_n12), .Z (calcRCon_n25) ) ;
    NAND2_X1 calcRCon_U22 ( .A1 (nReset), .A2 (calcRCon_n24), .ZN (calcRCon_n48) ) ;
    MUX2_X1 calcRCon_U21 ( .S (calcRCon_n5), .A (calcRCon_n23), .B (calcRCon_n15), .Z (calcRCon_n24) ) ;
    XNOR2_X1 calcRCon_U20 ( .A (calcRCon_n3), .B (calcRCon_s_current_state_2_), .ZN (calcRCon_n23) ) ;
    NAND2_X1 calcRCon_U19 ( .A1 (calcRCon_n22), .A2 (calcRCon_n21), .ZN (calcRCon_n47) ) ;
    NAND2_X1 calcRCon_U18 ( .A1 (calcRCon_s_current_state_4_), .A2 (calcRCon_n28), .ZN (calcRCon_n21) ) ;
    NAND2_X1 calcRCon_U17 ( .A1 (calcRCon_n20), .A2 (calcRCon_n26), .ZN (calcRCon_n22) ) ;
    XOR2_X1 calcRCon_U16 ( .A (calcRCon_n15), .B (calcRCon_n11), .Z (calcRCon_n20) ) ;
    NAND2_X1 calcRCon_U15 ( .A1 (calcRCon_n19), .A2 (calcRCon_n18), .ZN (calcRCon_n46) ) ;
    NAND2_X1 calcRCon_U14 ( .A1 (calcRCon_s_current_state_4_), .A2 (calcRCon_n26), .ZN (calcRCon_n18) ) ;
    NAND2_X1 calcRCon_U13 ( .A1 (calcRCon_s_current_state_5_), .A2 (calcRCon_n28), .ZN (calcRCon_n19) ) ;
    NAND2_X1 calcRCon_U12 ( .A1 (calcRCon_n17), .A2 (calcRCon_n10), .ZN (calcRCon_n45) ) ;
    NAND2_X1 calcRCon_U11 ( .A1 (calcRCon_s_current_state_5_), .A2 (calcRCon_n26), .ZN (calcRCon_n10) ) ;
    NOR2_X1 calcRCon_U10 ( .A1 (calcRCon_n5), .A2 (calcRCon_n6), .ZN (calcRCon_n26) ) ;
    NAND2_X1 calcRCon_U9 ( .A1 (calcRCon_s_current_state_6_), .A2 (calcRCon_n28), .ZN (calcRCon_n17) ) ;
    NOR2_X1 calcRCon_U8 ( .A1 (selSR), .A2 (calcRCon_n6), .ZN (calcRCon_n28) ) ;
    NAND2_X1 calcRCon_U7 ( .A1 (nReset), .A2 (calcRCon_n9), .ZN (calcRCon_n44) ) ;
    MUX2_X1 calcRCon_U6 ( .S (calcRCon_n5), .A (calcRCon_n16), .B (calcRCon_n11), .Z (calcRCon_n9) ) ;
    NAND2_X1 calcRCon_U5 ( .A1 (calcRCon_s_current_state_4_), .A2 (calcRCon_s_current_state_2_), .ZN (calcRCon_n7) ) ;
    NAND2_X1 calcRCon_U4 ( .A1 (calcRCon_s_current_state_1_), .A2 (calcRCon_s_current_state_5_), .ZN (calcRCon_n8) ) ;
    INV_X1 calcRCon_U3 ( .A (nReset), .ZN (calcRCon_n6) ) ;
    INV_X1 calcRCon_U2 ( .A (selSR), .ZN (calcRCon_n5) ) ;
    NOR2_X1 calcRCon_U1 ( .A1 (calcRCon_n8), .A2 (calcRCon_n7), .ZN (intFinal) ) ;
    INV_X1 calcRCon_s_current_state_reg_0__U1 ( .A (calcRCon_s_current_state_0_), .ZN (calcRCon_n13) ) ;
    INV_X1 calcRCon_s_current_state_reg_1__U1 ( .A (calcRCon_s_current_state_1_), .ZN (calcRCon_n14) ) ;
    INV_X1 calcRCon_s_current_state_reg_2__U1 ( .A (calcRCon_s_current_state_2_), .ZN (calcRCon_n12) ) ;
    INV_X1 calcRCon_s_current_state_reg_3__U1 ( .A (calcRCon_s_current_state_3_), .ZN (calcRCon_n15) ) ;
    INV_X1 calcRCon_s_current_state_reg_6__U1 ( .A (calcRCon_s_current_state_6_), .ZN (calcRCon_n16) ) ;
    INV_X1 calcRCon_s_current_state_reg_7__U1 ( .A (calcRCon_n3), .ZN (calcRCon_n11) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_SboxIn_mux_inst_0_U1 ( .s (selMC), .b ({new_AGEMA_signal_1984, StateOutXORroundKey[0]}), .a ({new_AGEMA_signal_2563, keySBIn[0]}), .c ({new_AGEMA_signal_2826, SboxIn[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_SboxIn_mux_inst_1_U1 ( .s (selMC), .b ({new_AGEMA_signal_1987, StateOutXORroundKey[1]}), .a ({new_AGEMA_signal_2566, keySBIn[1]}), .c ({new_AGEMA_signal_2827, SboxIn[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_SboxIn_mux_inst_2_U1 ( .s (selMC), .b ({new_AGEMA_signal_1990, StateOutXORroundKey[2]}), .a ({new_AGEMA_signal_2569, keySBIn[2]}), .c ({new_AGEMA_signal_2828, SboxIn[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_SboxIn_mux_inst_3_U1 ( .s (selMC), .b ({new_AGEMA_signal_1993, StateOutXORroundKey[3]}), .a ({new_AGEMA_signal_2572, keySBIn[3]}), .c ({new_AGEMA_signal_2829, SboxIn[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_SboxIn_mux_inst_4_U1 ( .s (selMC), .b ({new_AGEMA_signal_1996, StateOutXORroundKey[4]}), .a ({new_AGEMA_signal_2575, keySBIn[4]}), .c ({new_AGEMA_signal_2830, SboxIn[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_SboxIn_mux_inst_5_U1 ( .s (selMC), .b ({new_AGEMA_signal_1999, StateOutXORroundKey[5]}), .a ({new_AGEMA_signal_2578, keySBIn[5]}), .c ({new_AGEMA_signal_2831, SboxIn[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_SboxIn_mux_inst_6_U1 ( .s (selMC), .b ({new_AGEMA_signal_2002, StateOutXORroundKey[6]}), .a ({new_AGEMA_signal_2581, keySBIn[6]}), .c ({new_AGEMA_signal_2832, SboxIn[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_SboxIn_mux_inst_7_U1 ( .s (selMC), .b ({new_AGEMA_signal_2005, StateOutXORroundKey[7]}), .a ({new_AGEMA_signal_2584, keySBIn[7]}), .c ({new_AGEMA_signal_2833, SboxIn[7]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_T1_U1 ( .a ({new_AGEMA_signal_2833, SboxIn[7]}), .b ({new_AGEMA_signal_2830, SboxIn[4]}), .c ({new_AGEMA_signal_2850, Inst_bSbox_T1}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_T2_U1 ( .a ({new_AGEMA_signal_2833, SboxIn[7]}), .b ({new_AGEMA_signal_2828, SboxIn[2]}), .c ({new_AGEMA_signal_2851, Inst_bSbox_T2}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_T3_U1 ( .a ({new_AGEMA_signal_2833, SboxIn[7]}), .b ({new_AGEMA_signal_2827, SboxIn[1]}), .c ({new_AGEMA_signal_2852, Inst_bSbox_T3}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_T4_U1 ( .a ({new_AGEMA_signal_2830, SboxIn[4]}), .b ({new_AGEMA_signal_2828, SboxIn[2]}), .c ({new_AGEMA_signal_2853, Inst_bSbox_T4}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_T5_U1 ( .a ({new_AGEMA_signal_2829, SboxIn[3]}), .b ({new_AGEMA_signal_2827, SboxIn[1]}), .c ({new_AGEMA_signal_2854, Inst_bSbox_T5}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_T6_U1 ( .a ({new_AGEMA_signal_2850, Inst_bSbox_T1}), .b ({new_AGEMA_signal_2854, Inst_bSbox_T5}), .c ({new_AGEMA_signal_3000, Inst_bSbox_T6}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_T7_U1 ( .a ({new_AGEMA_signal_2832, SboxIn[6]}), .b ({new_AGEMA_signal_2831, SboxIn[5]}), .c ({new_AGEMA_signal_2855, Inst_bSbox_T7}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_T8_U1 ( .a ({new_AGEMA_signal_2826, SboxIn[0]}), .b ({new_AGEMA_signal_3000, Inst_bSbox_T6}), .c ({new_AGEMA_signal_3032, Inst_bSbox_T8}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_T9_U1 ( .a ({new_AGEMA_signal_2826, SboxIn[0]}), .b ({new_AGEMA_signal_2855, Inst_bSbox_T7}), .c ({new_AGEMA_signal_3001, Inst_bSbox_T9}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_T10_U1 ( .a ({new_AGEMA_signal_3000, Inst_bSbox_T6}), .b ({new_AGEMA_signal_2855, Inst_bSbox_T7}), .c ({new_AGEMA_signal_3033, Inst_bSbox_T10}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_T11_U1 ( .a ({new_AGEMA_signal_2832, SboxIn[6]}), .b ({new_AGEMA_signal_2828, SboxIn[2]}), .c ({new_AGEMA_signal_2856, Inst_bSbox_T11}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_T12_U1 ( .a ({new_AGEMA_signal_2831, SboxIn[5]}), .b ({new_AGEMA_signal_2828, SboxIn[2]}), .c ({new_AGEMA_signal_2857, Inst_bSbox_T12}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_T13_U1 ( .a ({new_AGEMA_signal_2852, Inst_bSbox_T3}), .b ({new_AGEMA_signal_2853, Inst_bSbox_T4}), .c ({new_AGEMA_signal_3002, Inst_bSbox_T13}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_T14_U1 ( .a ({new_AGEMA_signal_3000, Inst_bSbox_T6}), .b ({new_AGEMA_signal_2856, Inst_bSbox_T11}), .c ({new_AGEMA_signal_3034, Inst_bSbox_T14}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_T15_U1 ( .a ({new_AGEMA_signal_2854, Inst_bSbox_T5}), .b ({new_AGEMA_signal_2856, Inst_bSbox_T11}), .c ({new_AGEMA_signal_3003, Inst_bSbox_T15}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_T16_U1 ( .a ({new_AGEMA_signal_2854, Inst_bSbox_T5}), .b ({new_AGEMA_signal_2857, Inst_bSbox_T12}), .c ({new_AGEMA_signal_3004, Inst_bSbox_T16}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_T17_U1 ( .a ({new_AGEMA_signal_3001, Inst_bSbox_T9}), .b ({new_AGEMA_signal_3004, Inst_bSbox_T16}), .c ({new_AGEMA_signal_3035, Inst_bSbox_T17}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_T18_U1 ( .a ({new_AGEMA_signal_2830, SboxIn[4]}), .b ({new_AGEMA_signal_2826, SboxIn[0]}), .c ({new_AGEMA_signal_2858, Inst_bSbox_T18}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_T19_U1 ( .a ({new_AGEMA_signal_2855, Inst_bSbox_T7}), .b ({new_AGEMA_signal_2858, Inst_bSbox_T18}), .c ({new_AGEMA_signal_3005, Inst_bSbox_T19}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_T20_U1 ( .a ({new_AGEMA_signal_2850, Inst_bSbox_T1}), .b ({new_AGEMA_signal_3005, Inst_bSbox_T19}), .c ({new_AGEMA_signal_3036, Inst_bSbox_T20}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_T21_U1 ( .a ({new_AGEMA_signal_2827, SboxIn[1]}), .b ({new_AGEMA_signal_2826, SboxIn[0]}), .c ({new_AGEMA_signal_2859, Inst_bSbox_T21}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_T22_U1 ( .a ({new_AGEMA_signal_2855, Inst_bSbox_T7}), .b ({new_AGEMA_signal_2859, Inst_bSbox_T21}), .c ({new_AGEMA_signal_3006, Inst_bSbox_T22}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_T23_U1 ( .a ({new_AGEMA_signal_2851, Inst_bSbox_T2}), .b ({new_AGEMA_signal_3006, Inst_bSbox_T22}), .c ({new_AGEMA_signal_3037, Inst_bSbox_T23}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_T24_U1 ( .a ({new_AGEMA_signal_2851, Inst_bSbox_T2}), .b ({new_AGEMA_signal_3033, Inst_bSbox_T10}), .c ({new_AGEMA_signal_3117, Inst_bSbox_T24}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_T25_U1 ( .a ({new_AGEMA_signal_3036, Inst_bSbox_T20}), .b ({new_AGEMA_signal_3035, Inst_bSbox_T17}), .c ({new_AGEMA_signal_3118, Inst_bSbox_T25}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_T26_U1 ( .a ({new_AGEMA_signal_2852, Inst_bSbox_T3}), .b ({new_AGEMA_signal_3004, Inst_bSbox_T16}), .c ({new_AGEMA_signal_3038, Inst_bSbox_T26}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_T27_U1 ( .a ({new_AGEMA_signal_2850, Inst_bSbox_T1}), .b ({new_AGEMA_signal_2857, Inst_bSbox_T12}), .c ({new_AGEMA_signal_3007, Inst_bSbox_T27}) ) ;
    INV_X1 nReset_reg_U1 ( .A (nReset), .ZN (n10) ) ;

    /* cells in depth 1 */
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M1_U1 ( .a ({new_AGEMA_signal_3002, Inst_bSbox_T13}), .b ({new_AGEMA_signal_3000, Inst_bSbox_T6}), .clk (clk), .r ({Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_3039, Inst_bSbox_M1}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M2_U1 ( .a ({new_AGEMA_signal_3037, Inst_bSbox_T23}), .b ({new_AGEMA_signal_3032, Inst_bSbox_T8}), .clk (clk), .r ({Fresh[7], Fresh[6], Fresh[5], Fresh[4]}), .c ({new_AGEMA_signal_3119, Inst_bSbox_M2}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_M3_U1 ( .a ({new_AGEMA_signal_3671, new_AGEMA_signal_3670}), .b ({new_AGEMA_signal_3039, Inst_bSbox_M1}), .c ({new_AGEMA_signal_3120, Inst_bSbox_M3}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M4_U1 ( .a ({new_AGEMA_signal_3005, Inst_bSbox_T19}), .b ({new_AGEMA_signal_2826, SboxIn[0]}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8]}), .c ({new_AGEMA_signal_3040, Inst_bSbox_M4}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_M5_U1 ( .a ({new_AGEMA_signal_3040, Inst_bSbox_M4}), .b ({new_AGEMA_signal_3039, Inst_bSbox_M1}), .c ({new_AGEMA_signal_3121, Inst_bSbox_M5}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M6_U1 ( .a ({new_AGEMA_signal_2852, Inst_bSbox_T3}), .b ({new_AGEMA_signal_3004, Inst_bSbox_T16}), .clk (clk), .r ({Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_3041, Inst_bSbox_M6}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M7_U1 ( .a ({new_AGEMA_signal_3006, Inst_bSbox_T22}), .b ({new_AGEMA_signal_3001, Inst_bSbox_T9}), .clk (clk), .r ({Fresh[19], Fresh[18], Fresh[17], Fresh[16]}), .c ({new_AGEMA_signal_3042, Inst_bSbox_M7}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_M8_U1 ( .a ({new_AGEMA_signal_3673, new_AGEMA_signal_3672}), .b ({new_AGEMA_signal_3041, Inst_bSbox_M6}), .c ({new_AGEMA_signal_3122, Inst_bSbox_M8}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M9_U1 ( .a ({new_AGEMA_signal_3036, Inst_bSbox_T20}), .b ({new_AGEMA_signal_3035, Inst_bSbox_T17}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20]}), .c ({new_AGEMA_signal_3123, Inst_bSbox_M9}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_M10_U1 ( .a ({new_AGEMA_signal_3123, Inst_bSbox_M9}), .b ({new_AGEMA_signal_3041, Inst_bSbox_M6}), .c ({new_AGEMA_signal_3262, Inst_bSbox_M10}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M11_U1 ( .a ({new_AGEMA_signal_2850, Inst_bSbox_T1}), .b ({new_AGEMA_signal_3003, Inst_bSbox_T15}), .clk (clk), .r ({Fresh[27], Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_3043, Inst_bSbox_M11}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M12_U1 ( .a ({new_AGEMA_signal_2853, Inst_bSbox_T4}), .b ({new_AGEMA_signal_3007, Inst_bSbox_T27}), .clk (clk), .r ({Fresh[31], Fresh[30], Fresh[29], Fresh[28]}), .c ({new_AGEMA_signal_3044, Inst_bSbox_M12}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_M13_U1 ( .a ({new_AGEMA_signal_3044, Inst_bSbox_M12}), .b ({new_AGEMA_signal_3043, Inst_bSbox_M11}), .c ({new_AGEMA_signal_3124, Inst_bSbox_M13}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M14_U1 ( .a ({new_AGEMA_signal_2851, Inst_bSbox_T2}), .b ({new_AGEMA_signal_3033, Inst_bSbox_T10}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33], Fresh[32]}), .c ({new_AGEMA_signal_3125, Inst_bSbox_M14}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_M15_U1 ( .a ({new_AGEMA_signal_3125, Inst_bSbox_M14}), .b ({new_AGEMA_signal_3043, Inst_bSbox_M11}), .c ({new_AGEMA_signal_3263, Inst_bSbox_M15}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_M16_U1 ( .a ({new_AGEMA_signal_3120, Inst_bSbox_M3}), .b ({new_AGEMA_signal_3119, Inst_bSbox_M2}), .c ({new_AGEMA_signal_3264, Inst_bSbox_M16}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_M17_U1 ( .a ({new_AGEMA_signal_3121, Inst_bSbox_M5}), .b ({new_AGEMA_signal_3675, new_AGEMA_signal_3674}), .c ({new_AGEMA_signal_3265, Inst_bSbox_M17}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_M18_U1 ( .a ({new_AGEMA_signal_3122, Inst_bSbox_M8}), .b ({new_AGEMA_signal_3042, Inst_bSbox_M7}), .c ({new_AGEMA_signal_3266, Inst_bSbox_M18}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_M19_U1 ( .a ({new_AGEMA_signal_3262, Inst_bSbox_M10}), .b ({new_AGEMA_signal_3263, Inst_bSbox_M15}), .c ({new_AGEMA_signal_3371, Inst_bSbox_M19}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_M20_U1 ( .a ({new_AGEMA_signal_3264, Inst_bSbox_M16}), .b ({new_AGEMA_signal_3124, Inst_bSbox_M13}), .c ({new_AGEMA_signal_3372, Inst_bSbox_M20}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_M21_U1 ( .a ({new_AGEMA_signal_3265, Inst_bSbox_M17}), .b ({new_AGEMA_signal_3263, Inst_bSbox_M15}), .c ({new_AGEMA_signal_3373, Inst_bSbox_M21}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_M22_U1 ( .a ({new_AGEMA_signal_3266, Inst_bSbox_M18}), .b ({new_AGEMA_signal_3124, Inst_bSbox_M13}), .c ({new_AGEMA_signal_3374, Inst_bSbox_M22}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_M23_U1 ( .a ({new_AGEMA_signal_3371, Inst_bSbox_M19}), .b ({new_AGEMA_signal_3677, new_AGEMA_signal_3676}), .c ({new_AGEMA_signal_3383, Inst_bSbox_M23}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_M24_U1 ( .a ({new_AGEMA_signal_3374, Inst_bSbox_M22}), .b ({new_AGEMA_signal_3383, Inst_bSbox_M23}), .c ({new_AGEMA_signal_3387, Inst_bSbox_M24}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_M27_U1 ( .a ({new_AGEMA_signal_3372, Inst_bSbox_M20}), .b ({new_AGEMA_signal_3373, Inst_bSbox_M21}), .c ({new_AGEMA_signal_3385, Inst_bSbox_M27}) ) ;
    buf_clk new_AGEMA_reg_buffer_1714 ( .C (clk), .D (Inst_bSbox_T14), .Q (new_AGEMA_signal_3670) ) ;
    buf_clk new_AGEMA_reg_buffer_1715 ( .C (clk), .D (new_AGEMA_signal_3034), .Q (new_AGEMA_signal_3671) ) ;
    buf_clk new_AGEMA_reg_buffer_1716 ( .C (clk), .D (Inst_bSbox_T26), .Q (new_AGEMA_signal_3672) ) ;
    buf_clk new_AGEMA_reg_buffer_1717 ( .C (clk), .D (new_AGEMA_signal_3038), .Q (new_AGEMA_signal_3673) ) ;
    buf_clk new_AGEMA_reg_buffer_1718 ( .C (clk), .D (Inst_bSbox_T24), .Q (new_AGEMA_signal_3674) ) ;
    buf_clk new_AGEMA_reg_buffer_1719 ( .C (clk), .D (new_AGEMA_signal_3117), .Q (new_AGEMA_signal_3675) ) ;
    buf_clk new_AGEMA_reg_buffer_1720 ( .C (clk), .D (Inst_bSbox_T25), .Q (new_AGEMA_signal_3676) ) ;
    buf_clk new_AGEMA_reg_buffer_1721 ( .C (clk), .D (new_AGEMA_signal_3118), .Q (new_AGEMA_signal_3677) ) ;
    buf_clk new_AGEMA_reg_buffer_1738 ( .C (clk), .D (intFinal), .Q (new_AGEMA_signal_3694) ) ;
    buf_clk new_AGEMA_reg_buffer_1742 ( .C (clk), .D (StateOutXORroundKey[0]), .Q (new_AGEMA_signal_3698) ) ;
    buf_clk new_AGEMA_reg_buffer_1746 ( .C (clk), .D (new_AGEMA_signal_1984), .Q (new_AGEMA_signal_3702) ) ;
    buf_clk new_AGEMA_reg_buffer_1750 ( .C (clk), .D (StateOutXORroundKey[1]), .Q (new_AGEMA_signal_3706) ) ;
    buf_clk new_AGEMA_reg_buffer_1754 ( .C (clk), .D (new_AGEMA_signal_1987), .Q (new_AGEMA_signal_3710) ) ;
    buf_clk new_AGEMA_reg_buffer_1758 ( .C (clk), .D (StateOutXORroundKey[2]), .Q (new_AGEMA_signal_3714) ) ;
    buf_clk new_AGEMA_reg_buffer_1762 ( .C (clk), .D (new_AGEMA_signal_1990), .Q (new_AGEMA_signal_3718) ) ;
    buf_clk new_AGEMA_reg_buffer_1766 ( .C (clk), .D (StateOutXORroundKey[3]), .Q (new_AGEMA_signal_3722) ) ;
    buf_clk new_AGEMA_reg_buffer_1770 ( .C (clk), .D (new_AGEMA_signal_1993), .Q (new_AGEMA_signal_3726) ) ;
    buf_clk new_AGEMA_reg_buffer_1774 ( .C (clk), .D (StateOutXORroundKey[4]), .Q (new_AGEMA_signal_3730) ) ;
    buf_clk new_AGEMA_reg_buffer_1778 ( .C (clk), .D (new_AGEMA_signal_1996), .Q (new_AGEMA_signal_3734) ) ;
    buf_clk new_AGEMA_reg_buffer_1782 ( .C (clk), .D (StateOutXORroundKey[5]), .Q (new_AGEMA_signal_3738) ) ;
    buf_clk new_AGEMA_reg_buffer_1786 ( .C (clk), .D (new_AGEMA_signal_1999), .Q (new_AGEMA_signal_3742) ) ;
    buf_clk new_AGEMA_reg_buffer_1790 ( .C (clk), .D (StateOutXORroundKey[6]), .Q (new_AGEMA_signal_3746) ) ;
    buf_clk new_AGEMA_reg_buffer_1794 ( .C (clk), .D (new_AGEMA_signal_2002), .Q (new_AGEMA_signal_3750) ) ;
    buf_clk new_AGEMA_reg_buffer_1798 ( .C (clk), .D (StateOutXORroundKey[7]), .Q (new_AGEMA_signal_3754) ) ;
    buf_clk new_AGEMA_reg_buffer_1802 ( .C (clk), .D (new_AGEMA_signal_2005), .Q (new_AGEMA_signal_3758) ) ;
    buf_clk new_AGEMA_reg_buffer_1806 ( .C (clk), .D (stateArray_n13), .Q (new_AGEMA_signal_3762) ) ;
    buf_clk new_AGEMA_reg_buffer_1810 ( .C (clk), .D (ciphertext_s0[8]), .Q (new_AGEMA_signal_3766) ) ;
    buf_clk new_AGEMA_reg_buffer_1814 ( .C (clk), .D (ciphertext_s1[8]), .Q (new_AGEMA_signal_3770) ) ;
    buf_clk new_AGEMA_reg_buffer_1818 ( .C (clk), .D (ciphertext_s0[9]), .Q (new_AGEMA_signal_3774) ) ;
    buf_clk new_AGEMA_reg_buffer_1822 ( .C (clk), .D (ciphertext_s1[9]), .Q (new_AGEMA_signal_3778) ) ;
    buf_clk new_AGEMA_reg_buffer_1826 ( .C (clk), .D (ciphertext_s0[10]), .Q (new_AGEMA_signal_3782) ) ;
    buf_clk new_AGEMA_reg_buffer_1830 ( .C (clk), .D (ciphertext_s1[10]), .Q (new_AGEMA_signal_3786) ) ;
    buf_clk new_AGEMA_reg_buffer_1834 ( .C (clk), .D (ciphertext_s0[11]), .Q (new_AGEMA_signal_3790) ) ;
    buf_clk new_AGEMA_reg_buffer_1838 ( .C (clk), .D (ciphertext_s1[11]), .Q (new_AGEMA_signal_3794) ) ;
    buf_clk new_AGEMA_reg_buffer_1842 ( .C (clk), .D (ciphertext_s0[12]), .Q (new_AGEMA_signal_3798) ) ;
    buf_clk new_AGEMA_reg_buffer_1846 ( .C (clk), .D (ciphertext_s1[12]), .Q (new_AGEMA_signal_3802) ) ;
    buf_clk new_AGEMA_reg_buffer_1850 ( .C (clk), .D (ciphertext_s0[13]), .Q (new_AGEMA_signal_3806) ) ;
    buf_clk new_AGEMA_reg_buffer_1854 ( .C (clk), .D (ciphertext_s1[13]), .Q (new_AGEMA_signal_3810) ) ;
    buf_clk new_AGEMA_reg_buffer_1858 ( .C (clk), .D (ciphertext_s0[14]), .Q (new_AGEMA_signal_3814) ) ;
    buf_clk new_AGEMA_reg_buffer_1862 ( .C (clk), .D (ciphertext_s1[14]), .Q (new_AGEMA_signal_3818) ) ;
    buf_clk new_AGEMA_reg_buffer_1866 ( .C (clk), .D (ciphertext_s0[15]), .Q (new_AGEMA_signal_3822) ) ;
    buf_clk new_AGEMA_reg_buffer_1870 ( .C (clk), .D (ciphertext_s1[15]), .Q (new_AGEMA_signal_3826) ) ;
    buf_clk new_AGEMA_reg_buffer_1874 ( .C (clk), .D (stateArray_n22), .Q (new_AGEMA_signal_3830) ) ;
    buf_clk new_AGEMA_reg_buffer_1878 ( .C (clk), .D (StateInMC[0]), .Q (new_AGEMA_signal_3834) ) ;
    buf_clk new_AGEMA_reg_buffer_1882 ( .C (clk), .D (new_AGEMA_signal_2860), .Q (new_AGEMA_signal_3838) ) ;
    buf_clk new_AGEMA_reg_buffer_1886 ( .C (clk), .D (StateInMC[1]), .Q (new_AGEMA_signal_3842) ) ;
    buf_clk new_AGEMA_reg_buffer_1890 ( .C (clk), .D (new_AGEMA_signal_2861), .Q (new_AGEMA_signal_3846) ) ;
    buf_clk new_AGEMA_reg_buffer_1894 ( .C (clk), .D (StateInMC[2]), .Q (new_AGEMA_signal_3850) ) ;
    buf_clk new_AGEMA_reg_buffer_1898 ( .C (clk), .D (new_AGEMA_signal_2834), .Q (new_AGEMA_signal_3854) ) ;
    buf_clk new_AGEMA_reg_buffer_1902 ( .C (clk), .D (StateInMC[3]), .Q (new_AGEMA_signal_3858) ) ;
    buf_clk new_AGEMA_reg_buffer_1906 ( .C (clk), .D (new_AGEMA_signal_2862), .Q (new_AGEMA_signal_3862) ) ;
    buf_clk new_AGEMA_reg_buffer_1910 ( .C (clk), .D (StateInMC[4]), .Q (new_AGEMA_signal_3866) ) ;
    buf_clk new_AGEMA_reg_buffer_1914 ( .C (clk), .D (new_AGEMA_signal_2863), .Q (new_AGEMA_signal_3870) ) ;
    buf_clk new_AGEMA_reg_buffer_1918 ( .C (clk), .D (StateInMC[5]), .Q (new_AGEMA_signal_3874) ) ;
    buf_clk new_AGEMA_reg_buffer_1922 ( .C (clk), .D (new_AGEMA_signal_2835), .Q (new_AGEMA_signal_3878) ) ;
    buf_clk new_AGEMA_reg_buffer_1926 ( .C (clk), .D (StateInMC[6]), .Q (new_AGEMA_signal_3882) ) ;
    buf_clk new_AGEMA_reg_buffer_1930 ( .C (clk), .D (new_AGEMA_signal_2836), .Q (new_AGEMA_signal_3886) ) ;
    buf_clk new_AGEMA_reg_buffer_1934 ( .C (clk), .D (StateInMC[7]), .Q (new_AGEMA_signal_3890) ) ;
    buf_clk new_AGEMA_reg_buffer_1938 ( .C (clk), .D (new_AGEMA_signal_2837), .Q (new_AGEMA_signal_3894) ) ;
    buf_clk new_AGEMA_reg_buffer_1942 ( .C (clk), .D (stateArray_n25), .Q (new_AGEMA_signal_3898) ) ;
    buf_clk new_AGEMA_reg_buffer_1946 ( .C (clk), .D (plaintext_s0[0]), .Q (new_AGEMA_signal_3902) ) ;
    buf_clk new_AGEMA_reg_buffer_1950 ( .C (clk), .D (plaintext_s1[0]), .Q (new_AGEMA_signal_3906) ) ;
    buf_clk new_AGEMA_reg_buffer_1954 ( .C (clk), .D (plaintext_s0[1]), .Q (new_AGEMA_signal_3910) ) ;
    buf_clk new_AGEMA_reg_buffer_1958 ( .C (clk), .D (plaintext_s1[1]), .Q (new_AGEMA_signal_3914) ) ;
    buf_clk new_AGEMA_reg_buffer_1962 ( .C (clk), .D (plaintext_s0[2]), .Q (new_AGEMA_signal_3918) ) ;
    buf_clk new_AGEMA_reg_buffer_1966 ( .C (clk), .D (plaintext_s1[2]), .Q (new_AGEMA_signal_3922) ) ;
    buf_clk new_AGEMA_reg_buffer_1970 ( .C (clk), .D (plaintext_s0[3]), .Q (new_AGEMA_signal_3926) ) ;
    buf_clk new_AGEMA_reg_buffer_1974 ( .C (clk), .D (plaintext_s1[3]), .Q (new_AGEMA_signal_3930) ) ;
    buf_clk new_AGEMA_reg_buffer_1978 ( .C (clk), .D (plaintext_s0[4]), .Q (new_AGEMA_signal_3934) ) ;
    buf_clk new_AGEMA_reg_buffer_1982 ( .C (clk), .D (plaintext_s1[4]), .Q (new_AGEMA_signal_3938) ) ;
    buf_clk new_AGEMA_reg_buffer_1986 ( .C (clk), .D (plaintext_s0[5]), .Q (new_AGEMA_signal_3942) ) ;
    buf_clk new_AGEMA_reg_buffer_1990 ( .C (clk), .D (plaintext_s1[5]), .Q (new_AGEMA_signal_3946) ) ;
    buf_clk new_AGEMA_reg_buffer_1994 ( .C (clk), .D (plaintext_s0[6]), .Q (new_AGEMA_signal_3950) ) ;
    buf_clk new_AGEMA_reg_buffer_1998 ( .C (clk), .D (plaintext_s1[6]), .Q (new_AGEMA_signal_3954) ) ;
    buf_clk new_AGEMA_reg_buffer_2002 ( .C (clk), .D (plaintext_s0[7]), .Q (new_AGEMA_signal_3958) ) ;
    buf_clk new_AGEMA_reg_buffer_2006 ( .C (clk), .D (plaintext_s1[7]), .Q (new_AGEMA_signal_3962) ) ;
    buf_clk new_AGEMA_reg_buffer_2010 ( .C (clk), .D (keyStateIn[7]), .Q (new_AGEMA_signal_3966) ) ;
    buf_clk new_AGEMA_reg_buffer_2014 ( .C (clk), .D (new_AGEMA_signal_2004), .Q (new_AGEMA_signal_3970) ) ;
    buf_clk new_AGEMA_reg_buffer_2018 ( .C (clk), .D (roundConstant[7]), .Q (new_AGEMA_signal_3974) ) ;
    buf_clk new_AGEMA_reg_buffer_2022 ( .C (clk), .D (keyStateIn[6]), .Q (new_AGEMA_signal_3978) ) ;
    buf_clk new_AGEMA_reg_buffer_2026 ( .C (clk), .D (new_AGEMA_signal_2001), .Q (new_AGEMA_signal_3982) ) ;
    buf_clk new_AGEMA_reg_buffer_2030 ( .C (clk), .D (roundConstant[6]), .Q (new_AGEMA_signal_3986) ) ;
    buf_clk new_AGEMA_reg_buffer_2034 ( .C (clk), .D (keyStateIn[5]), .Q (new_AGEMA_signal_3990) ) ;
    buf_clk new_AGEMA_reg_buffer_2038 ( .C (clk), .D (new_AGEMA_signal_1998), .Q (new_AGEMA_signal_3994) ) ;
    buf_clk new_AGEMA_reg_buffer_2042 ( .C (clk), .D (roundConstant[5]), .Q (new_AGEMA_signal_3998) ) ;
    buf_clk new_AGEMA_reg_buffer_2046 ( .C (clk), .D (keyStateIn[4]), .Q (new_AGEMA_signal_4002) ) ;
    buf_clk new_AGEMA_reg_buffer_2050 ( .C (clk), .D (new_AGEMA_signal_1995), .Q (new_AGEMA_signal_4006) ) ;
    buf_clk new_AGEMA_reg_buffer_2054 ( .C (clk), .D (roundConstant[4]), .Q (new_AGEMA_signal_4010) ) ;
    buf_clk new_AGEMA_reg_buffer_2058 ( .C (clk), .D (keyStateIn[3]), .Q (new_AGEMA_signal_4014) ) ;
    buf_clk new_AGEMA_reg_buffer_2062 ( .C (clk), .D (new_AGEMA_signal_1992), .Q (new_AGEMA_signal_4018) ) ;
    buf_clk new_AGEMA_reg_buffer_2066 ( .C (clk), .D (roundConstant[3]), .Q (new_AGEMA_signal_4022) ) ;
    buf_clk new_AGEMA_reg_buffer_2070 ( .C (clk), .D (keyStateIn[2]), .Q (new_AGEMA_signal_4026) ) ;
    buf_clk new_AGEMA_reg_buffer_2074 ( .C (clk), .D (new_AGEMA_signal_1989), .Q (new_AGEMA_signal_4030) ) ;
    buf_clk new_AGEMA_reg_buffer_2078 ( .C (clk), .D (roundConstant[2]), .Q (new_AGEMA_signal_4034) ) ;
    buf_clk new_AGEMA_reg_buffer_2082 ( .C (clk), .D (keyStateIn[1]), .Q (new_AGEMA_signal_4038) ) ;
    buf_clk new_AGEMA_reg_buffer_2086 ( .C (clk), .D (new_AGEMA_signal_1986), .Q (new_AGEMA_signal_4042) ) ;
    buf_clk new_AGEMA_reg_buffer_2090 ( .C (clk), .D (roundConstant[1]), .Q (new_AGEMA_signal_4046) ) ;
    buf_clk new_AGEMA_reg_buffer_2094 ( .C (clk), .D (keyStateIn[0]), .Q (new_AGEMA_signal_4050) ) ;
    buf_clk new_AGEMA_reg_buffer_2098 ( .C (clk), .D (new_AGEMA_signal_1983), .Q (new_AGEMA_signal_4054) ) ;
    buf_clk new_AGEMA_reg_buffer_2102 ( .C (clk), .D (roundConstant[0]), .Q (new_AGEMA_signal_4058) ) ;
    buf_clk new_AGEMA_reg_buffer_2106 ( .C (clk), .D (KeyArray_n23), .Q (new_AGEMA_signal_4062) ) ;
    buf_clk new_AGEMA_reg_buffer_2110 ( .C (clk), .D (KeyArray_outS30ser[0]), .Q (new_AGEMA_signal_4066) ) ;
    buf_clk new_AGEMA_reg_buffer_2114 ( .C (clk), .D (new_AGEMA_signal_2683), .Q (new_AGEMA_signal_4070) ) ;
    buf_clk new_AGEMA_reg_buffer_2118 ( .C (clk), .D (KeyArray_n31), .Q (new_AGEMA_signal_4074) ) ;
    buf_clk new_AGEMA_reg_buffer_2122 ( .C (clk), .D (KeyArray_inS30ser[0]), .Q (new_AGEMA_signal_4078) ) ;
    buf_clk new_AGEMA_reg_buffer_2126 ( .C (clk), .D (new_AGEMA_signal_2708), .Q (new_AGEMA_signal_4082) ) ;
    buf_clk new_AGEMA_reg_buffer_2130 ( .C (clk), .D (KeyArray_outS30ser[1]), .Q (new_AGEMA_signal_4086) ) ;
    buf_clk new_AGEMA_reg_buffer_2134 ( .C (clk), .D (new_AGEMA_signal_2686), .Q (new_AGEMA_signal_4090) ) ;
    buf_clk new_AGEMA_reg_buffer_2138 ( .C (clk), .D (KeyArray_inS30ser[1]), .Q (new_AGEMA_signal_4094) ) ;
    buf_clk new_AGEMA_reg_buffer_2142 ( .C (clk), .D (new_AGEMA_signal_2711), .Q (new_AGEMA_signal_4098) ) ;
    buf_clk new_AGEMA_reg_buffer_2146 ( .C (clk), .D (KeyArray_outS30ser[2]), .Q (new_AGEMA_signal_4102) ) ;
    buf_clk new_AGEMA_reg_buffer_2150 ( .C (clk), .D (new_AGEMA_signal_2689), .Q (new_AGEMA_signal_4106) ) ;
    buf_clk new_AGEMA_reg_buffer_2154 ( .C (clk), .D (KeyArray_inS30ser[2]), .Q (new_AGEMA_signal_4110) ) ;
    buf_clk new_AGEMA_reg_buffer_2158 ( .C (clk), .D (new_AGEMA_signal_2714), .Q (new_AGEMA_signal_4114) ) ;
    buf_clk new_AGEMA_reg_buffer_2162 ( .C (clk), .D (KeyArray_outS30ser[3]), .Q (new_AGEMA_signal_4118) ) ;
    buf_clk new_AGEMA_reg_buffer_2166 ( .C (clk), .D (new_AGEMA_signal_2692), .Q (new_AGEMA_signal_4122) ) ;
    buf_clk new_AGEMA_reg_buffer_2170 ( .C (clk), .D (KeyArray_inS30ser[3]), .Q (new_AGEMA_signal_4126) ) ;
    buf_clk new_AGEMA_reg_buffer_2174 ( .C (clk), .D (new_AGEMA_signal_2717), .Q (new_AGEMA_signal_4130) ) ;
    buf_clk new_AGEMA_reg_buffer_2178 ( .C (clk), .D (KeyArray_outS30ser[4]), .Q (new_AGEMA_signal_4134) ) ;
    buf_clk new_AGEMA_reg_buffer_2182 ( .C (clk), .D (new_AGEMA_signal_2695), .Q (new_AGEMA_signal_4138) ) ;
    buf_clk new_AGEMA_reg_buffer_2186 ( .C (clk), .D (KeyArray_inS30ser[4]), .Q (new_AGEMA_signal_4142) ) ;
    buf_clk new_AGEMA_reg_buffer_2190 ( .C (clk), .D (new_AGEMA_signal_2720), .Q (new_AGEMA_signal_4146) ) ;
    buf_clk new_AGEMA_reg_buffer_2194 ( .C (clk), .D (KeyArray_outS30ser[5]), .Q (new_AGEMA_signal_4150) ) ;
    buf_clk new_AGEMA_reg_buffer_2198 ( .C (clk), .D (new_AGEMA_signal_2698), .Q (new_AGEMA_signal_4154) ) ;
    buf_clk new_AGEMA_reg_buffer_2202 ( .C (clk), .D (KeyArray_inS30ser[5]), .Q (new_AGEMA_signal_4158) ) ;
    buf_clk new_AGEMA_reg_buffer_2206 ( .C (clk), .D (new_AGEMA_signal_2723), .Q (new_AGEMA_signal_4162) ) ;
    buf_clk new_AGEMA_reg_buffer_2210 ( .C (clk), .D (KeyArray_outS30ser[6]), .Q (new_AGEMA_signal_4166) ) ;
    buf_clk new_AGEMA_reg_buffer_2214 ( .C (clk), .D (new_AGEMA_signal_2701), .Q (new_AGEMA_signal_4170) ) ;
    buf_clk new_AGEMA_reg_buffer_2218 ( .C (clk), .D (KeyArray_inS30ser[6]), .Q (new_AGEMA_signal_4174) ) ;
    buf_clk new_AGEMA_reg_buffer_2222 ( .C (clk), .D (new_AGEMA_signal_2726), .Q (new_AGEMA_signal_4178) ) ;
    buf_clk new_AGEMA_reg_buffer_2226 ( .C (clk), .D (KeyArray_outS30ser[7]), .Q (new_AGEMA_signal_4182) ) ;
    buf_clk new_AGEMA_reg_buffer_2230 ( .C (clk), .D (new_AGEMA_signal_2704), .Q (new_AGEMA_signal_4186) ) ;
    buf_clk new_AGEMA_reg_buffer_2234 ( .C (clk), .D (KeyArray_inS30ser[7]), .Q (new_AGEMA_signal_4190) ) ;
    buf_clk new_AGEMA_reg_buffer_2238 ( .C (clk), .D (new_AGEMA_signal_2729), .Q (new_AGEMA_signal_4194) ) ;
    buf_clk new_AGEMA_reg_buffer_2242 ( .C (clk), .D (Inst_bSbox_T6), .Q (new_AGEMA_signal_4198) ) ;
    buf_clk new_AGEMA_reg_buffer_2245 ( .C (clk), .D (new_AGEMA_signal_3000), .Q (new_AGEMA_signal_4201) ) ;
    buf_clk new_AGEMA_reg_buffer_2248 ( .C (clk), .D (Inst_bSbox_T8), .Q (new_AGEMA_signal_4204) ) ;
    buf_clk new_AGEMA_reg_buffer_2251 ( .C (clk), .D (new_AGEMA_signal_3032), .Q (new_AGEMA_signal_4207) ) ;
    buf_clk new_AGEMA_reg_buffer_2254 ( .C (clk), .D (SboxIn[0]), .Q (new_AGEMA_signal_4210) ) ;
    buf_clk new_AGEMA_reg_buffer_2257 ( .C (clk), .D (new_AGEMA_signal_2826), .Q (new_AGEMA_signal_4213) ) ;
    buf_clk new_AGEMA_reg_buffer_2260 ( .C (clk), .D (Inst_bSbox_T16), .Q (new_AGEMA_signal_4216) ) ;
    buf_clk new_AGEMA_reg_buffer_2263 ( .C (clk), .D (new_AGEMA_signal_3004), .Q (new_AGEMA_signal_4219) ) ;
    buf_clk new_AGEMA_reg_buffer_2266 ( .C (clk), .D (Inst_bSbox_T9), .Q (new_AGEMA_signal_4222) ) ;
    buf_clk new_AGEMA_reg_buffer_2269 ( .C (clk), .D (new_AGEMA_signal_3001), .Q (new_AGEMA_signal_4225) ) ;
    buf_clk new_AGEMA_reg_buffer_2272 ( .C (clk), .D (Inst_bSbox_T17), .Q (new_AGEMA_signal_4228) ) ;
    buf_clk new_AGEMA_reg_buffer_2275 ( .C (clk), .D (new_AGEMA_signal_3035), .Q (new_AGEMA_signal_4231) ) ;
    buf_clk new_AGEMA_reg_buffer_2278 ( .C (clk), .D (Inst_bSbox_T15), .Q (new_AGEMA_signal_4234) ) ;
    buf_clk new_AGEMA_reg_buffer_2281 ( .C (clk), .D (new_AGEMA_signal_3003), .Q (new_AGEMA_signal_4237) ) ;
    buf_clk new_AGEMA_reg_buffer_2284 ( .C (clk), .D (Inst_bSbox_T27), .Q (new_AGEMA_signal_4240) ) ;
    buf_clk new_AGEMA_reg_buffer_2287 ( .C (clk), .D (new_AGEMA_signal_3007), .Q (new_AGEMA_signal_4243) ) ;
    buf_clk new_AGEMA_reg_buffer_2290 ( .C (clk), .D (Inst_bSbox_T10), .Q (new_AGEMA_signal_4246) ) ;
    buf_clk new_AGEMA_reg_buffer_2293 ( .C (clk), .D (new_AGEMA_signal_3033), .Q (new_AGEMA_signal_4249) ) ;
    buf_clk new_AGEMA_reg_buffer_2296 ( .C (clk), .D (Inst_bSbox_T13), .Q (new_AGEMA_signal_4252) ) ;
    buf_clk new_AGEMA_reg_buffer_2299 ( .C (clk), .D (new_AGEMA_signal_3002), .Q (new_AGEMA_signal_4255) ) ;
    buf_clk new_AGEMA_reg_buffer_2302 ( .C (clk), .D (Inst_bSbox_T23), .Q (new_AGEMA_signal_4258) ) ;
    buf_clk new_AGEMA_reg_buffer_2305 ( .C (clk), .D (new_AGEMA_signal_3037), .Q (new_AGEMA_signal_4261) ) ;
    buf_clk new_AGEMA_reg_buffer_2308 ( .C (clk), .D (Inst_bSbox_T19), .Q (new_AGEMA_signal_4264) ) ;
    buf_clk new_AGEMA_reg_buffer_2311 ( .C (clk), .D (new_AGEMA_signal_3005), .Q (new_AGEMA_signal_4267) ) ;
    buf_clk new_AGEMA_reg_buffer_2314 ( .C (clk), .D (Inst_bSbox_T3), .Q (new_AGEMA_signal_4270) ) ;
    buf_clk new_AGEMA_reg_buffer_2317 ( .C (clk), .D (new_AGEMA_signal_2852), .Q (new_AGEMA_signal_4273) ) ;
    buf_clk new_AGEMA_reg_buffer_2320 ( .C (clk), .D (Inst_bSbox_T22), .Q (new_AGEMA_signal_4276) ) ;
    buf_clk new_AGEMA_reg_buffer_2323 ( .C (clk), .D (new_AGEMA_signal_3006), .Q (new_AGEMA_signal_4279) ) ;
    buf_clk new_AGEMA_reg_buffer_2326 ( .C (clk), .D (Inst_bSbox_T20), .Q (new_AGEMA_signal_4282) ) ;
    buf_clk new_AGEMA_reg_buffer_2329 ( .C (clk), .D (new_AGEMA_signal_3036), .Q (new_AGEMA_signal_4285) ) ;
    buf_clk new_AGEMA_reg_buffer_2332 ( .C (clk), .D (Inst_bSbox_T1), .Q (new_AGEMA_signal_4288) ) ;
    buf_clk new_AGEMA_reg_buffer_2335 ( .C (clk), .D (new_AGEMA_signal_2850), .Q (new_AGEMA_signal_4291) ) ;
    buf_clk new_AGEMA_reg_buffer_2338 ( .C (clk), .D (Inst_bSbox_T4), .Q (new_AGEMA_signal_4294) ) ;
    buf_clk new_AGEMA_reg_buffer_2341 ( .C (clk), .D (new_AGEMA_signal_2853), .Q (new_AGEMA_signal_4297) ) ;
    buf_clk new_AGEMA_reg_buffer_2344 ( .C (clk), .D (Inst_bSbox_T2), .Q (new_AGEMA_signal_4300) ) ;
    buf_clk new_AGEMA_reg_buffer_2347 ( .C (clk), .D (new_AGEMA_signal_2851), .Q (new_AGEMA_signal_4303) ) ;
    buf_clk new_AGEMA_reg_buffer_2350 ( .C (clk), .D (ctrl_seq6_SFF_0_QD), .Q (new_AGEMA_signal_4306) ) ;
    buf_clk new_AGEMA_reg_buffer_2354 ( .C (clk), .D (ctrl_seq6_SFF_1_QD), .Q (new_AGEMA_signal_4310) ) ;
    buf_clk new_AGEMA_reg_buffer_2358 ( .C (clk), .D (ctrl_seq6_SFF_2_QD), .Q (new_AGEMA_signal_4314) ) ;
    buf_clk new_AGEMA_reg_buffer_2362 ( .C (clk), .D (ctrl_seq6_SFF_3_QD), .Q (new_AGEMA_signal_4318) ) ;
    buf_clk new_AGEMA_reg_buffer_2366 ( .C (clk), .D (ctrl_seq6_SFF_4_QD), .Q (new_AGEMA_signal_4322) ) ;
    buf_clk new_AGEMA_reg_buffer_2370 ( .C (clk), .D (ctrl_seq4_SFF_0_QD), .Q (new_AGEMA_signal_4326) ) ;
    buf_clk new_AGEMA_reg_buffer_2374 ( .C (clk), .D (ctrl_seq4_SFF_1_QD), .Q (new_AGEMA_signal_4330) ) ;
    buf_clk new_AGEMA_reg_buffer_2378 ( .C (clk), .D (ctrl_N14), .Q (new_AGEMA_signal_4334) ) ;
    buf_clk new_AGEMA_reg_buffer_2382 ( .C (clk), .D (selSR), .Q (new_AGEMA_signal_4338) ) ;
    buf_clk new_AGEMA_reg_buffer_2386 ( .C (clk), .D (stateArray_S00reg_gff_1_SFF_0_QD), .Q (new_AGEMA_signal_4342) ) ;
    buf_clk new_AGEMA_reg_buffer_2390 ( .C (clk), .D (new_AGEMA_signal_3126), .Q (new_AGEMA_signal_4346) ) ;
    buf_clk new_AGEMA_reg_buffer_2394 ( .C (clk), .D (stateArray_S00reg_gff_1_SFF_1_QD), .Q (new_AGEMA_signal_4350) ) ;
    buf_clk new_AGEMA_reg_buffer_2398 ( .C (clk), .D (new_AGEMA_signal_3127), .Q (new_AGEMA_signal_4354) ) ;
    buf_clk new_AGEMA_reg_buffer_2402 ( .C (clk), .D (stateArray_S00reg_gff_1_SFF_2_QD), .Q (new_AGEMA_signal_4358) ) ;
    buf_clk new_AGEMA_reg_buffer_2406 ( .C (clk), .D (new_AGEMA_signal_3128), .Q (new_AGEMA_signal_4362) ) ;
    buf_clk new_AGEMA_reg_buffer_2410 ( .C (clk), .D (stateArray_S00reg_gff_1_SFF_3_QD), .Q (new_AGEMA_signal_4366) ) ;
    buf_clk new_AGEMA_reg_buffer_2414 ( .C (clk), .D (new_AGEMA_signal_3129), .Q (new_AGEMA_signal_4370) ) ;
    buf_clk new_AGEMA_reg_buffer_2418 ( .C (clk), .D (stateArray_S00reg_gff_1_SFF_4_QD), .Q (new_AGEMA_signal_4374) ) ;
    buf_clk new_AGEMA_reg_buffer_2422 ( .C (clk), .D (new_AGEMA_signal_3130), .Q (new_AGEMA_signal_4378) ) ;
    buf_clk new_AGEMA_reg_buffer_2426 ( .C (clk), .D (stateArray_S00reg_gff_1_SFF_5_QD), .Q (new_AGEMA_signal_4382) ) ;
    buf_clk new_AGEMA_reg_buffer_2430 ( .C (clk), .D (new_AGEMA_signal_3131), .Q (new_AGEMA_signal_4386) ) ;
    buf_clk new_AGEMA_reg_buffer_2434 ( .C (clk), .D (stateArray_S00reg_gff_1_SFF_6_QD), .Q (new_AGEMA_signal_4390) ) ;
    buf_clk new_AGEMA_reg_buffer_2438 ( .C (clk), .D (new_AGEMA_signal_3132), .Q (new_AGEMA_signal_4394) ) ;
    buf_clk new_AGEMA_reg_buffer_2442 ( .C (clk), .D (stateArray_S00reg_gff_1_SFF_7_QD), .Q (new_AGEMA_signal_4398) ) ;
    buf_clk new_AGEMA_reg_buffer_2446 ( .C (clk), .D (new_AGEMA_signal_3133), .Q (new_AGEMA_signal_4402) ) ;
    buf_clk new_AGEMA_reg_buffer_2450 ( .C (clk), .D (stateArray_S01reg_gff_1_SFF_0_QD), .Q (new_AGEMA_signal_4406) ) ;
    buf_clk new_AGEMA_reg_buffer_2454 ( .C (clk), .D (new_AGEMA_signal_3134), .Q (new_AGEMA_signal_4410) ) ;
    buf_clk new_AGEMA_reg_buffer_2458 ( .C (clk), .D (stateArray_S01reg_gff_1_SFF_1_QD), .Q (new_AGEMA_signal_4414) ) ;
    buf_clk new_AGEMA_reg_buffer_2462 ( .C (clk), .D (new_AGEMA_signal_3135), .Q (new_AGEMA_signal_4418) ) ;
    buf_clk new_AGEMA_reg_buffer_2466 ( .C (clk), .D (stateArray_S01reg_gff_1_SFF_2_QD), .Q (new_AGEMA_signal_4422) ) ;
    buf_clk new_AGEMA_reg_buffer_2470 ( .C (clk), .D (new_AGEMA_signal_3136), .Q (new_AGEMA_signal_4426) ) ;
    buf_clk new_AGEMA_reg_buffer_2474 ( .C (clk), .D (stateArray_S01reg_gff_1_SFF_3_QD), .Q (new_AGEMA_signal_4430) ) ;
    buf_clk new_AGEMA_reg_buffer_2478 ( .C (clk), .D (new_AGEMA_signal_3137), .Q (new_AGEMA_signal_4434) ) ;
    buf_clk new_AGEMA_reg_buffer_2482 ( .C (clk), .D (stateArray_S01reg_gff_1_SFF_4_QD), .Q (new_AGEMA_signal_4438) ) ;
    buf_clk new_AGEMA_reg_buffer_2486 ( .C (clk), .D (new_AGEMA_signal_3138), .Q (new_AGEMA_signal_4442) ) ;
    buf_clk new_AGEMA_reg_buffer_2490 ( .C (clk), .D (stateArray_S01reg_gff_1_SFF_5_QD), .Q (new_AGEMA_signal_4446) ) ;
    buf_clk new_AGEMA_reg_buffer_2494 ( .C (clk), .D (new_AGEMA_signal_3139), .Q (new_AGEMA_signal_4450) ) ;
    buf_clk new_AGEMA_reg_buffer_2498 ( .C (clk), .D (stateArray_S01reg_gff_1_SFF_6_QD), .Q (new_AGEMA_signal_4454) ) ;
    buf_clk new_AGEMA_reg_buffer_2502 ( .C (clk), .D (new_AGEMA_signal_3140), .Q (new_AGEMA_signal_4458) ) ;
    buf_clk new_AGEMA_reg_buffer_2506 ( .C (clk), .D (stateArray_S01reg_gff_1_SFF_7_QD), .Q (new_AGEMA_signal_4462) ) ;
    buf_clk new_AGEMA_reg_buffer_2510 ( .C (clk), .D (new_AGEMA_signal_3141), .Q (new_AGEMA_signal_4466) ) ;
    buf_clk new_AGEMA_reg_buffer_2514 ( .C (clk), .D (stateArray_S02reg_gff_1_SFF_0_QD), .Q (new_AGEMA_signal_4470) ) ;
    buf_clk new_AGEMA_reg_buffer_2518 ( .C (clk), .D (new_AGEMA_signal_3142), .Q (new_AGEMA_signal_4474) ) ;
    buf_clk new_AGEMA_reg_buffer_2522 ( .C (clk), .D (stateArray_S02reg_gff_1_SFF_1_QD), .Q (new_AGEMA_signal_4478) ) ;
    buf_clk new_AGEMA_reg_buffer_2526 ( .C (clk), .D (new_AGEMA_signal_3143), .Q (new_AGEMA_signal_4482) ) ;
    buf_clk new_AGEMA_reg_buffer_2530 ( .C (clk), .D (stateArray_S02reg_gff_1_SFF_2_QD), .Q (new_AGEMA_signal_4486) ) ;
    buf_clk new_AGEMA_reg_buffer_2534 ( .C (clk), .D (new_AGEMA_signal_3144), .Q (new_AGEMA_signal_4490) ) ;
    buf_clk new_AGEMA_reg_buffer_2538 ( .C (clk), .D (stateArray_S02reg_gff_1_SFF_3_QD), .Q (new_AGEMA_signal_4494) ) ;
    buf_clk new_AGEMA_reg_buffer_2542 ( .C (clk), .D (new_AGEMA_signal_3145), .Q (new_AGEMA_signal_4498) ) ;
    buf_clk new_AGEMA_reg_buffer_2546 ( .C (clk), .D (stateArray_S02reg_gff_1_SFF_4_QD), .Q (new_AGEMA_signal_4502) ) ;
    buf_clk new_AGEMA_reg_buffer_2550 ( .C (clk), .D (new_AGEMA_signal_3146), .Q (new_AGEMA_signal_4506) ) ;
    buf_clk new_AGEMA_reg_buffer_2554 ( .C (clk), .D (stateArray_S02reg_gff_1_SFF_5_QD), .Q (new_AGEMA_signal_4510) ) ;
    buf_clk new_AGEMA_reg_buffer_2558 ( .C (clk), .D (new_AGEMA_signal_3147), .Q (new_AGEMA_signal_4514) ) ;
    buf_clk new_AGEMA_reg_buffer_2562 ( .C (clk), .D (stateArray_S02reg_gff_1_SFF_6_QD), .Q (new_AGEMA_signal_4518) ) ;
    buf_clk new_AGEMA_reg_buffer_2566 ( .C (clk), .D (new_AGEMA_signal_3148), .Q (new_AGEMA_signal_4522) ) ;
    buf_clk new_AGEMA_reg_buffer_2570 ( .C (clk), .D (stateArray_S02reg_gff_1_SFF_7_QD), .Q (new_AGEMA_signal_4526) ) ;
    buf_clk new_AGEMA_reg_buffer_2574 ( .C (clk), .D (new_AGEMA_signal_3149), .Q (new_AGEMA_signal_4530) ) ;
    buf_clk new_AGEMA_reg_buffer_2578 ( .C (clk), .D (stateArray_S03reg_gff_1_SFF_0_QD), .Q (new_AGEMA_signal_4534) ) ;
    buf_clk new_AGEMA_reg_buffer_2582 ( .C (clk), .D (new_AGEMA_signal_3150), .Q (new_AGEMA_signal_4538) ) ;
    buf_clk new_AGEMA_reg_buffer_2586 ( .C (clk), .D (stateArray_S03reg_gff_1_SFF_1_QD), .Q (new_AGEMA_signal_4542) ) ;
    buf_clk new_AGEMA_reg_buffer_2590 ( .C (clk), .D (new_AGEMA_signal_3151), .Q (new_AGEMA_signal_4546) ) ;
    buf_clk new_AGEMA_reg_buffer_2594 ( .C (clk), .D (stateArray_S03reg_gff_1_SFF_2_QD), .Q (new_AGEMA_signal_4550) ) ;
    buf_clk new_AGEMA_reg_buffer_2598 ( .C (clk), .D (new_AGEMA_signal_3152), .Q (new_AGEMA_signal_4554) ) ;
    buf_clk new_AGEMA_reg_buffer_2602 ( .C (clk), .D (stateArray_S03reg_gff_1_SFF_3_QD), .Q (new_AGEMA_signal_4558) ) ;
    buf_clk new_AGEMA_reg_buffer_2606 ( .C (clk), .D (new_AGEMA_signal_3153), .Q (new_AGEMA_signal_4562) ) ;
    buf_clk new_AGEMA_reg_buffer_2610 ( .C (clk), .D (stateArray_S03reg_gff_1_SFF_4_QD), .Q (new_AGEMA_signal_4566) ) ;
    buf_clk new_AGEMA_reg_buffer_2614 ( .C (clk), .D (new_AGEMA_signal_3154), .Q (new_AGEMA_signal_4570) ) ;
    buf_clk new_AGEMA_reg_buffer_2618 ( .C (clk), .D (stateArray_S03reg_gff_1_SFF_5_QD), .Q (new_AGEMA_signal_4574) ) ;
    buf_clk new_AGEMA_reg_buffer_2622 ( .C (clk), .D (new_AGEMA_signal_3155), .Q (new_AGEMA_signal_4578) ) ;
    buf_clk new_AGEMA_reg_buffer_2626 ( .C (clk), .D (stateArray_S03reg_gff_1_SFF_6_QD), .Q (new_AGEMA_signal_4582) ) ;
    buf_clk new_AGEMA_reg_buffer_2630 ( .C (clk), .D (new_AGEMA_signal_3156), .Q (new_AGEMA_signal_4586) ) ;
    buf_clk new_AGEMA_reg_buffer_2634 ( .C (clk), .D (stateArray_S03reg_gff_1_SFF_7_QD), .Q (new_AGEMA_signal_4590) ) ;
    buf_clk new_AGEMA_reg_buffer_2638 ( .C (clk), .D (new_AGEMA_signal_3157), .Q (new_AGEMA_signal_4594) ) ;
    buf_clk new_AGEMA_reg_buffer_2642 ( .C (clk), .D (stateArray_S10reg_gff_1_SFF_0_QD), .Q (new_AGEMA_signal_4598) ) ;
    buf_clk new_AGEMA_reg_buffer_2646 ( .C (clk), .D (new_AGEMA_signal_3158), .Q (new_AGEMA_signal_4602) ) ;
    buf_clk new_AGEMA_reg_buffer_2650 ( .C (clk), .D (stateArray_S10reg_gff_1_SFF_1_QD), .Q (new_AGEMA_signal_4606) ) ;
    buf_clk new_AGEMA_reg_buffer_2654 ( .C (clk), .D (new_AGEMA_signal_3159), .Q (new_AGEMA_signal_4610) ) ;
    buf_clk new_AGEMA_reg_buffer_2658 ( .C (clk), .D (stateArray_S10reg_gff_1_SFF_2_QD), .Q (new_AGEMA_signal_4614) ) ;
    buf_clk new_AGEMA_reg_buffer_2662 ( .C (clk), .D (new_AGEMA_signal_3160), .Q (new_AGEMA_signal_4618) ) ;
    buf_clk new_AGEMA_reg_buffer_2666 ( .C (clk), .D (stateArray_S10reg_gff_1_SFF_3_QD), .Q (new_AGEMA_signal_4622) ) ;
    buf_clk new_AGEMA_reg_buffer_2670 ( .C (clk), .D (new_AGEMA_signal_3161), .Q (new_AGEMA_signal_4626) ) ;
    buf_clk new_AGEMA_reg_buffer_2674 ( .C (clk), .D (stateArray_S10reg_gff_1_SFF_4_QD), .Q (new_AGEMA_signal_4630) ) ;
    buf_clk new_AGEMA_reg_buffer_2678 ( .C (clk), .D (new_AGEMA_signal_3162), .Q (new_AGEMA_signal_4634) ) ;
    buf_clk new_AGEMA_reg_buffer_2682 ( .C (clk), .D (stateArray_S10reg_gff_1_SFF_5_QD), .Q (new_AGEMA_signal_4638) ) ;
    buf_clk new_AGEMA_reg_buffer_2686 ( .C (clk), .D (new_AGEMA_signal_3163), .Q (new_AGEMA_signal_4642) ) ;
    buf_clk new_AGEMA_reg_buffer_2690 ( .C (clk), .D (stateArray_S10reg_gff_1_SFF_6_QD), .Q (new_AGEMA_signal_4646) ) ;
    buf_clk new_AGEMA_reg_buffer_2694 ( .C (clk), .D (new_AGEMA_signal_3164), .Q (new_AGEMA_signal_4650) ) ;
    buf_clk new_AGEMA_reg_buffer_2698 ( .C (clk), .D (stateArray_S10reg_gff_1_SFF_7_QD), .Q (new_AGEMA_signal_4654) ) ;
    buf_clk new_AGEMA_reg_buffer_2702 ( .C (clk), .D (new_AGEMA_signal_3165), .Q (new_AGEMA_signal_4658) ) ;
    buf_clk new_AGEMA_reg_buffer_2706 ( .C (clk), .D (stateArray_S11reg_gff_1_SFF_0_QD), .Q (new_AGEMA_signal_4662) ) ;
    buf_clk new_AGEMA_reg_buffer_2710 ( .C (clk), .D (new_AGEMA_signal_3166), .Q (new_AGEMA_signal_4666) ) ;
    buf_clk new_AGEMA_reg_buffer_2714 ( .C (clk), .D (stateArray_S11reg_gff_1_SFF_1_QD), .Q (new_AGEMA_signal_4670) ) ;
    buf_clk new_AGEMA_reg_buffer_2718 ( .C (clk), .D (new_AGEMA_signal_3167), .Q (new_AGEMA_signal_4674) ) ;
    buf_clk new_AGEMA_reg_buffer_2722 ( .C (clk), .D (stateArray_S11reg_gff_1_SFF_2_QD), .Q (new_AGEMA_signal_4678) ) ;
    buf_clk new_AGEMA_reg_buffer_2726 ( .C (clk), .D (new_AGEMA_signal_3168), .Q (new_AGEMA_signal_4682) ) ;
    buf_clk new_AGEMA_reg_buffer_2730 ( .C (clk), .D (stateArray_S11reg_gff_1_SFF_3_QD), .Q (new_AGEMA_signal_4686) ) ;
    buf_clk new_AGEMA_reg_buffer_2734 ( .C (clk), .D (new_AGEMA_signal_3169), .Q (new_AGEMA_signal_4690) ) ;
    buf_clk new_AGEMA_reg_buffer_2738 ( .C (clk), .D (stateArray_S11reg_gff_1_SFF_4_QD), .Q (new_AGEMA_signal_4694) ) ;
    buf_clk new_AGEMA_reg_buffer_2742 ( .C (clk), .D (new_AGEMA_signal_3170), .Q (new_AGEMA_signal_4698) ) ;
    buf_clk new_AGEMA_reg_buffer_2746 ( .C (clk), .D (stateArray_S11reg_gff_1_SFF_5_QD), .Q (new_AGEMA_signal_4702) ) ;
    buf_clk new_AGEMA_reg_buffer_2750 ( .C (clk), .D (new_AGEMA_signal_3171), .Q (new_AGEMA_signal_4706) ) ;
    buf_clk new_AGEMA_reg_buffer_2754 ( .C (clk), .D (stateArray_S11reg_gff_1_SFF_6_QD), .Q (new_AGEMA_signal_4710) ) ;
    buf_clk new_AGEMA_reg_buffer_2758 ( .C (clk), .D (new_AGEMA_signal_3172), .Q (new_AGEMA_signal_4714) ) ;
    buf_clk new_AGEMA_reg_buffer_2762 ( .C (clk), .D (stateArray_S11reg_gff_1_SFF_7_QD), .Q (new_AGEMA_signal_4718) ) ;
    buf_clk new_AGEMA_reg_buffer_2766 ( .C (clk), .D (new_AGEMA_signal_3173), .Q (new_AGEMA_signal_4722) ) ;
    buf_clk new_AGEMA_reg_buffer_2770 ( .C (clk), .D (stateArray_S12reg_gff_1_SFF_0_QD), .Q (new_AGEMA_signal_4726) ) ;
    buf_clk new_AGEMA_reg_buffer_2774 ( .C (clk), .D (new_AGEMA_signal_3174), .Q (new_AGEMA_signal_4730) ) ;
    buf_clk new_AGEMA_reg_buffer_2778 ( .C (clk), .D (stateArray_S12reg_gff_1_SFF_1_QD), .Q (new_AGEMA_signal_4734) ) ;
    buf_clk new_AGEMA_reg_buffer_2782 ( .C (clk), .D (new_AGEMA_signal_3175), .Q (new_AGEMA_signal_4738) ) ;
    buf_clk new_AGEMA_reg_buffer_2786 ( .C (clk), .D (stateArray_S12reg_gff_1_SFF_2_QD), .Q (new_AGEMA_signal_4742) ) ;
    buf_clk new_AGEMA_reg_buffer_2790 ( .C (clk), .D (new_AGEMA_signal_3176), .Q (new_AGEMA_signal_4746) ) ;
    buf_clk new_AGEMA_reg_buffer_2794 ( .C (clk), .D (stateArray_S12reg_gff_1_SFF_3_QD), .Q (new_AGEMA_signal_4750) ) ;
    buf_clk new_AGEMA_reg_buffer_2798 ( .C (clk), .D (new_AGEMA_signal_3177), .Q (new_AGEMA_signal_4754) ) ;
    buf_clk new_AGEMA_reg_buffer_2802 ( .C (clk), .D (stateArray_S12reg_gff_1_SFF_4_QD), .Q (new_AGEMA_signal_4758) ) ;
    buf_clk new_AGEMA_reg_buffer_2806 ( .C (clk), .D (new_AGEMA_signal_3178), .Q (new_AGEMA_signal_4762) ) ;
    buf_clk new_AGEMA_reg_buffer_2810 ( .C (clk), .D (stateArray_S12reg_gff_1_SFF_5_QD), .Q (new_AGEMA_signal_4766) ) ;
    buf_clk new_AGEMA_reg_buffer_2814 ( .C (clk), .D (new_AGEMA_signal_3179), .Q (new_AGEMA_signal_4770) ) ;
    buf_clk new_AGEMA_reg_buffer_2818 ( .C (clk), .D (stateArray_S12reg_gff_1_SFF_6_QD), .Q (new_AGEMA_signal_4774) ) ;
    buf_clk new_AGEMA_reg_buffer_2822 ( .C (clk), .D (new_AGEMA_signal_3180), .Q (new_AGEMA_signal_4778) ) ;
    buf_clk new_AGEMA_reg_buffer_2826 ( .C (clk), .D (stateArray_S12reg_gff_1_SFF_7_QD), .Q (new_AGEMA_signal_4782) ) ;
    buf_clk new_AGEMA_reg_buffer_2830 ( .C (clk), .D (new_AGEMA_signal_3181), .Q (new_AGEMA_signal_4786) ) ;
    buf_clk new_AGEMA_reg_buffer_2834 ( .C (clk), .D (stateArray_S13reg_gff_1_SFF_0_QD), .Q (new_AGEMA_signal_4790) ) ;
    buf_clk new_AGEMA_reg_buffer_2838 ( .C (clk), .D (new_AGEMA_signal_3182), .Q (new_AGEMA_signal_4794) ) ;
    buf_clk new_AGEMA_reg_buffer_2842 ( .C (clk), .D (stateArray_S13reg_gff_1_SFF_1_QD), .Q (new_AGEMA_signal_4798) ) ;
    buf_clk new_AGEMA_reg_buffer_2846 ( .C (clk), .D (new_AGEMA_signal_3183), .Q (new_AGEMA_signal_4802) ) ;
    buf_clk new_AGEMA_reg_buffer_2850 ( .C (clk), .D (stateArray_S13reg_gff_1_SFF_2_QD), .Q (new_AGEMA_signal_4806) ) ;
    buf_clk new_AGEMA_reg_buffer_2854 ( .C (clk), .D (new_AGEMA_signal_3184), .Q (new_AGEMA_signal_4810) ) ;
    buf_clk new_AGEMA_reg_buffer_2858 ( .C (clk), .D (stateArray_S13reg_gff_1_SFF_3_QD), .Q (new_AGEMA_signal_4814) ) ;
    buf_clk new_AGEMA_reg_buffer_2862 ( .C (clk), .D (new_AGEMA_signal_3185), .Q (new_AGEMA_signal_4818) ) ;
    buf_clk new_AGEMA_reg_buffer_2866 ( .C (clk), .D (stateArray_S13reg_gff_1_SFF_4_QD), .Q (new_AGEMA_signal_4822) ) ;
    buf_clk new_AGEMA_reg_buffer_2870 ( .C (clk), .D (new_AGEMA_signal_3186), .Q (new_AGEMA_signal_4826) ) ;
    buf_clk new_AGEMA_reg_buffer_2874 ( .C (clk), .D (stateArray_S13reg_gff_1_SFF_5_QD), .Q (new_AGEMA_signal_4830) ) ;
    buf_clk new_AGEMA_reg_buffer_2878 ( .C (clk), .D (new_AGEMA_signal_3187), .Q (new_AGEMA_signal_4834) ) ;
    buf_clk new_AGEMA_reg_buffer_2882 ( .C (clk), .D (stateArray_S13reg_gff_1_SFF_6_QD), .Q (new_AGEMA_signal_4838) ) ;
    buf_clk new_AGEMA_reg_buffer_2886 ( .C (clk), .D (new_AGEMA_signal_3188), .Q (new_AGEMA_signal_4842) ) ;
    buf_clk new_AGEMA_reg_buffer_2890 ( .C (clk), .D (stateArray_S13reg_gff_1_SFF_7_QD), .Q (new_AGEMA_signal_4846) ) ;
    buf_clk new_AGEMA_reg_buffer_2894 ( .C (clk), .D (new_AGEMA_signal_3189), .Q (new_AGEMA_signal_4850) ) ;
    buf_clk new_AGEMA_reg_buffer_2898 ( .C (clk), .D (stateArray_S20reg_gff_1_SFF_0_QD), .Q (new_AGEMA_signal_4854) ) ;
    buf_clk new_AGEMA_reg_buffer_2902 ( .C (clk), .D (new_AGEMA_signal_3190), .Q (new_AGEMA_signal_4858) ) ;
    buf_clk new_AGEMA_reg_buffer_2906 ( .C (clk), .D (stateArray_S20reg_gff_1_SFF_1_QD), .Q (new_AGEMA_signal_4862) ) ;
    buf_clk new_AGEMA_reg_buffer_2910 ( .C (clk), .D (new_AGEMA_signal_3191), .Q (new_AGEMA_signal_4866) ) ;
    buf_clk new_AGEMA_reg_buffer_2914 ( .C (clk), .D (stateArray_S20reg_gff_1_SFF_2_QD), .Q (new_AGEMA_signal_4870) ) ;
    buf_clk new_AGEMA_reg_buffer_2918 ( .C (clk), .D (new_AGEMA_signal_3192), .Q (new_AGEMA_signal_4874) ) ;
    buf_clk new_AGEMA_reg_buffer_2922 ( .C (clk), .D (stateArray_S20reg_gff_1_SFF_3_QD), .Q (new_AGEMA_signal_4878) ) ;
    buf_clk new_AGEMA_reg_buffer_2926 ( .C (clk), .D (new_AGEMA_signal_3193), .Q (new_AGEMA_signal_4882) ) ;
    buf_clk new_AGEMA_reg_buffer_2930 ( .C (clk), .D (stateArray_S20reg_gff_1_SFF_4_QD), .Q (new_AGEMA_signal_4886) ) ;
    buf_clk new_AGEMA_reg_buffer_2934 ( .C (clk), .D (new_AGEMA_signal_3194), .Q (new_AGEMA_signal_4890) ) ;
    buf_clk new_AGEMA_reg_buffer_2938 ( .C (clk), .D (stateArray_S20reg_gff_1_SFF_5_QD), .Q (new_AGEMA_signal_4894) ) ;
    buf_clk new_AGEMA_reg_buffer_2942 ( .C (clk), .D (new_AGEMA_signal_3195), .Q (new_AGEMA_signal_4898) ) ;
    buf_clk new_AGEMA_reg_buffer_2946 ( .C (clk), .D (stateArray_S20reg_gff_1_SFF_6_QD), .Q (new_AGEMA_signal_4902) ) ;
    buf_clk new_AGEMA_reg_buffer_2950 ( .C (clk), .D (new_AGEMA_signal_3196), .Q (new_AGEMA_signal_4906) ) ;
    buf_clk new_AGEMA_reg_buffer_2954 ( .C (clk), .D (stateArray_S20reg_gff_1_SFF_7_QD), .Q (new_AGEMA_signal_4910) ) ;
    buf_clk new_AGEMA_reg_buffer_2958 ( .C (clk), .D (new_AGEMA_signal_3197), .Q (new_AGEMA_signal_4914) ) ;
    buf_clk new_AGEMA_reg_buffer_2962 ( .C (clk), .D (stateArray_S21reg_gff_1_SFF_0_QD), .Q (new_AGEMA_signal_4918) ) ;
    buf_clk new_AGEMA_reg_buffer_2966 ( .C (clk), .D (new_AGEMA_signal_3198), .Q (new_AGEMA_signal_4922) ) ;
    buf_clk new_AGEMA_reg_buffer_2970 ( .C (clk), .D (stateArray_S21reg_gff_1_SFF_1_QD), .Q (new_AGEMA_signal_4926) ) ;
    buf_clk new_AGEMA_reg_buffer_2974 ( .C (clk), .D (new_AGEMA_signal_3199), .Q (new_AGEMA_signal_4930) ) ;
    buf_clk new_AGEMA_reg_buffer_2978 ( .C (clk), .D (stateArray_S21reg_gff_1_SFF_2_QD), .Q (new_AGEMA_signal_4934) ) ;
    buf_clk new_AGEMA_reg_buffer_2982 ( .C (clk), .D (new_AGEMA_signal_3200), .Q (new_AGEMA_signal_4938) ) ;
    buf_clk new_AGEMA_reg_buffer_2986 ( .C (clk), .D (stateArray_S21reg_gff_1_SFF_3_QD), .Q (new_AGEMA_signal_4942) ) ;
    buf_clk new_AGEMA_reg_buffer_2990 ( .C (clk), .D (new_AGEMA_signal_3201), .Q (new_AGEMA_signal_4946) ) ;
    buf_clk new_AGEMA_reg_buffer_2994 ( .C (clk), .D (stateArray_S21reg_gff_1_SFF_4_QD), .Q (new_AGEMA_signal_4950) ) ;
    buf_clk new_AGEMA_reg_buffer_2998 ( .C (clk), .D (new_AGEMA_signal_3202), .Q (new_AGEMA_signal_4954) ) ;
    buf_clk new_AGEMA_reg_buffer_3002 ( .C (clk), .D (stateArray_S21reg_gff_1_SFF_5_QD), .Q (new_AGEMA_signal_4958) ) ;
    buf_clk new_AGEMA_reg_buffer_3006 ( .C (clk), .D (new_AGEMA_signal_3203), .Q (new_AGEMA_signal_4962) ) ;
    buf_clk new_AGEMA_reg_buffer_3010 ( .C (clk), .D (stateArray_S21reg_gff_1_SFF_6_QD), .Q (new_AGEMA_signal_4966) ) ;
    buf_clk new_AGEMA_reg_buffer_3014 ( .C (clk), .D (new_AGEMA_signal_3204), .Q (new_AGEMA_signal_4970) ) ;
    buf_clk new_AGEMA_reg_buffer_3018 ( .C (clk), .D (stateArray_S21reg_gff_1_SFF_7_QD), .Q (new_AGEMA_signal_4974) ) ;
    buf_clk new_AGEMA_reg_buffer_3022 ( .C (clk), .D (new_AGEMA_signal_3205), .Q (new_AGEMA_signal_4978) ) ;
    buf_clk new_AGEMA_reg_buffer_3026 ( .C (clk), .D (stateArray_S22reg_gff_1_SFF_0_QD), .Q (new_AGEMA_signal_4982) ) ;
    buf_clk new_AGEMA_reg_buffer_3030 ( .C (clk), .D (new_AGEMA_signal_3206), .Q (new_AGEMA_signal_4986) ) ;
    buf_clk new_AGEMA_reg_buffer_3034 ( .C (clk), .D (stateArray_S22reg_gff_1_SFF_1_QD), .Q (new_AGEMA_signal_4990) ) ;
    buf_clk new_AGEMA_reg_buffer_3038 ( .C (clk), .D (new_AGEMA_signal_3207), .Q (new_AGEMA_signal_4994) ) ;
    buf_clk new_AGEMA_reg_buffer_3042 ( .C (clk), .D (stateArray_S22reg_gff_1_SFF_2_QD), .Q (new_AGEMA_signal_4998) ) ;
    buf_clk new_AGEMA_reg_buffer_3046 ( .C (clk), .D (new_AGEMA_signal_3208), .Q (new_AGEMA_signal_5002) ) ;
    buf_clk new_AGEMA_reg_buffer_3050 ( .C (clk), .D (stateArray_S22reg_gff_1_SFF_3_QD), .Q (new_AGEMA_signal_5006) ) ;
    buf_clk new_AGEMA_reg_buffer_3054 ( .C (clk), .D (new_AGEMA_signal_3209), .Q (new_AGEMA_signal_5010) ) ;
    buf_clk new_AGEMA_reg_buffer_3058 ( .C (clk), .D (stateArray_S22reg_gff_1_SFF_4_QD), .Q (new_AGEMA_signal_5014) ) ;
    buf_clk new_AGEMA_reg_buffer_3062 ( .C (clk), .D (new_AGEMA_signal_3210), .Q (new_AGEMA_signal_5018) ) ;
    buf_clk new_AGEMA_reg_buffer_3066 ( .C (clk), .D (stateArray_S22reg_gff_1_SFF_5_QD), .Q (new_AGEMA_signal_5022) ) ;
    buf_clk new_AGEMA_reg_buffer_3070 ( .C (clk), .D (new_AGEMA_signal_3211), .Q (new_AGEMA_signal_5026) ) ;
    buf_clk new_AGEMA_reg_buffer_3074 ( .C (clk), .D (stateArray_S22reg_gff_1_SFF_6_QD), .Q (new_AGEMA_signal_5030) ) ;
    buf_clk new_AGEMA_reg_buffer_3078 ( .C (clk), .D (new_AGEMA_signal_3212), .Q (new_AGEMA_signal_5034) ) ;
    buf_clk new_AGEMA_reg_buffer_3082 ( .C (clk), .D (stateArray_S22reg_gff_1_SFF_7_QD), .Q (new_AGEMA_signal_5038) ) ;
    buf_clk new_AGEMA_reg_buffer_3086 ( .C (clk), .D (new_AGEMA_signal_3213), .Q (new_AGEMA_signal_5042) ) ;
    buf_clk new_AGEMA_reg_buffer_3090 ( .C (clk), .D (stateArray_S23reg_gff_1_SFF_0_QD), .Q (new_AGEMA_signal_5046) ) ;
    buf_clk new_AGEMA_reg_buffer_3094 ( .C (clk), .D (new_AGEMA_signal_3214), .Q (new_AGEMA_signal_5050) ) ;
    buf_clk new_AGEMA_reg_buffer_3098 ( .C (clk), .D (stateArray_S23reg_gff_1_SFF_1_QD), .Q (new_AGEMA_signal_5054) ) ;
    buf_clk new_AGEMA_reg_buffer_3102 ( .C (clk), .D (new_AGEMA_signal_3215), .Q (new_AGEMA_signal_5058) ) ;
    buf_clk new_AGEMA_reg_buffer_3106 ( .C (clk), .D (stateArray_S23reg_gff_1_SFF_2_QD), .Q (new_AGEMA_signal_5062) ) ;
    buf_clk new_AGEMA_reg_buffer_3110 ( .C (clk), .D (new_AGEMA_signal_3216), .Q (new_AGEMA_signal_5066) ) ;
    buf_clk new_AGEMA_reg_buffer_3114 ( .C (clk), .D (stateArray_S23reg_gff_1_SFF_3_QD), .Q (new_AGEMA_signal_5070) ) ;
    buf_clk new_AGEMA_reg_buffer_3118 ( .C (clk), .D (new_AGEMA_signal_3217), .Q (new_AGEMA_signal_5074) ) ;
    buf_clk new_AGEMA_reg_buffer_3122 ( .C (clk), .D (stateArray_S23reg_gff_1_SFF_4_QD), .Q (new_AGEMA_signal_5078) ) ;
    buf_clk new_AGEMA_reg_buffer_3126 ( .C (clk), .D (new_AGEMA_signal_3218), .Q (new_AGEMA_signal_5082) ) ;
    buf_clk new_AGEMA_reg_buffer_3130 ( .C (clk), .D (stateArray_S23reg_gff_1_SFF_5_QD), .Q (new_AGEMA_signal_5086) ) ;
    buf_clk new_AGEMA_reg_buffer_3134 ( .C (clk), .D (new_AGEMA_signal_3219), .Q (new_AGEMA_signal_5090) ) ;
    buf_clk new_AGEMA_reg_buffer_3138 ( .C (clk), .D (stateArray_S23reg_gff_1_SFF_6_QD), .Q (new_AGEMA_signal_5094) ) ;
    buf_clk new_AGEMA_reg_buffer_3142 ( .C (clk), .D (new_AGEMA_signal_3220), .Q (new_AGEMA_signal_5098) ) ;
    buf_clk new_AGEMA_reg_buffer_3146 ( .C (clk), .D (stateArray_S23reg_gff_1_SFF_7_QD), .Q (new_AGEMA_signal_5102) ) ;
    buf_clk new_AGEMA_reg_buffer_3150 ( .C (clk), .D (new_AGEMA_signal_3221), .Q (new_AGEMA_signal_5106) ) ;
    buf_clk new_AGEMA_reg_buffer_3154 ( .C (clk), .D (stateArray_S30reg_gff_1_SFF_0_QD), .Q (new_AGEMA_signal_5110) ) ;
    buf_clk new_AGEMA_reg_buffer_3158 ( .C (clk), .D (new_AGEMA_signal_3222), .Q (new_AGEMA_signal_5114) ) ;
    buf_clk new_AGEMA_reg_buffer_3162 ( .C (clk), .D (stateArray_S30reg_gff_1_SFF_1_QD), .Q (new_AGEMA_signal_5118) ) ;
    buf_clk new_AGEMA_reg_buffer_3166 ( .C (clk), .D (new_AGEMA_signal_3223), .Q (new_AGEMA_signal_5122) ) ;
    buf_clk new_AGEMA_reg_buffer_3170 ( .C (clk), .D (stateArray_S30reg_gff_1_SFF_2_QD), .Q (new_AGEMA_signal_5126) ) ;
    buf_clk new_AGEMA_reg_buffer_3174 ( .C (clk), .D (new_AGEMA_signal_3224), .Q (new_AGEMA_signal_5130) ) ;
    buf_clk new_AGEMA_reg_buffer_3178 ( .C (clk), .D (stateArray_S30reg_gff_1_SFF_3_QD), .Q (new_AGEMA_signal_5134) ) ;
    buf_clk new_AGEMA_reg_buffer_3182 ( .C (clk), .D (new_AGEMA_signal_3225), .Q (new_AGEMA_signal_5138) ) ;
    buf_clk new_AGEMA_reg_buffer_3186 ( .C (clk), .D (stateArray_S30reg_gff_1_SFF_4_QD), .Q (new_AGEMA_signal_5142) ) ;
    buf_clk new_AGEMA_reg_buffer_3190 ( .C (clk), .D (new_AGEMA_signal_3226), .Q (new_AGEMA_signal_5146) ) ;
    buf_clk new_AGEMA_reg_buffer_3194 ( .C (clk), .D (stateArray_S30reg_gff_1_SFF_5_QD), .Q (new_AGEMA_signal_5150) ) ;
    buf_clk new_AGEMA_reg_buffer_3198 ( .C (clk), .D (new_AGEMA_signal_3227), .Q (new_AGEMA_signal_5154) ) ;
    buf_clk new_AGEMA_reg_buffer_3202 ( .C (clk), .D (stateArray_S30reg_gff_1_SFF_6_QD), .Q (new_AGEMA_signal_5158) ) ;
    buf_clk new_AGEMA_reg_buffer_3206 ( .C (clk), .D (new_AGEMA_signal_3228), .Q (new_AGEMA_signal_5162) ) ;
    buf_clk new_AGEMA_reg_buffer_3210 ( .C (clk), .D (stateArray_S30reg_gff_1_SFF_7_QD), .Q (new_AGEMA_signal_5166) ) ;
    buf_clk new_AGEMA_reg_buffer_3214 ( .C (clk), .D (new_AGEMA_signal_3229), .Q (new_AGEMA_signal_5170) ) ;
    buf_clk new_AGEMA_reg_buffer_3218 ( .C (clk), .D (stateArray_S31reg_gff_1_SFF_0_QD), .Q (new_AGEMA_signal_5174) ) ;
    buf_clk new_AGEMA_reg_buffer_3222 ( .C (clk), .D (new_AGEMA_signal_3230), .Q (new_AGEMA_signal_5178) ) ;
    buf_clk new_AGEMA_reg_buffer_3226 ( .C (clk), .D (stateArray_S31reg_gff_1_SFF_1_QD), .Q (new_AGEMA_signal_5182) ) ;
    buf_clk new_AGEMA_reg_buffer_3230 ( .C (clk), .D (new_AGEMA_signal_3231), .Q (new_AGEMA_signal_5186) ) ;
    buf_clk new_AGEMA_reg_buffer_3234 ( .C (clk), .D (stateArray_S31reg_gff_1_SFF_2_QD), .Q (new_AGEMA_signal_5190) ) ;
    buf_clk new_AGEMA_reg_buffer_3238 ( .C (clk), .D (new_AGEMA_signal_3232), .Q (new_AGEMA_signal_5194) ) ;
    buf_clk new_AGEMA_reg_buffer_3242 ( .C (clk), .D (stateArray_S31reg_gff_1_SFF_3_QD), .Q (new_AGEMA_signal_5198) ) ;
    buf_clk new_AGEMA_reg_buffer_3246 ( .C (clk), .D (new_AGEMA_signal_3233), .Q (new_AGEMA_signal_5202) ) ;
    buf_clk new_AGEMA_reg_buffer_3250 ( .C (clk), .D (stateArray_S31reg_gff_1_SFF_4_QD), .Q (new_AGEMA_signal_5206) ) ;
    buf_clk new_AGEMA_reg_buffer_3254 ( .C (clk), .D (new_AGEMA_signal_3234), .Q (new_AGEMA_signal_5210) ) ;
    buf_clk new_AGEMA_reg_buffer_3258 ( .C (clk), .D (stateArray_S31reg_gff_1_SFF_5_QD), .Q (new_AGEMA_signal_5214) ) ;
    buf_clk new_AGEMA_reg_buffer_3262 ( .C (clk), .D (new_AGEMA_signal_3235), .Q (new_AGEMA_signal_5218) ) ;
    buf_clk new_AGEMA_reg_buffer_3266 ( .C (clk), .D (stateArray_S31reg_gff_1_SFF_6_QD), .Q (new_AGEMA_signal_5222) ) ;
    buf_clk new_AGEMA_reg_buffer_3270 ( .C (clk), .D (new_AGEMA_signal_3236), .Q (new_AGEMA_signal_5226) ) ;
    buf_clk new_AGEMA_reg_buffer_3274 ( .C (clk), .D (stateArray_S31reg_gff_1_SFF_7_QD), .Q (new_AGEMA_signal_5230) ) ;
    buf_clk new_AGEMA_reg_buffer_3278 ( .C (clk), .D (new_AGEMA_signal_3237), .Q (new_AGEMA_signal_5234) ) ;
    buf_clk new_AGEMA_reg_buffer_3282 ( .C (clk), .D (stateArray_S32reg_gff_1_SFF_0_QD), .Q (new_AGEMA_signal_5238) ) ;
    buf_clk new_AGEMA_reg_buffer_3286 ( .C (clk), .D (new_AGEMA_signal_3238), .Q (new_AGEMA_signal_5242) ) ;
    buf_clk new_AGEMA_reg_buffer_3290 ( .C (clk), .D (stateArray_S32reg_gff_1_SFF_1_QD), .Q (new_AGEMA_signal_5246) ) ;
    buf_clk new_AGEMA_reg_buffer_3294 ( .C (clk), .D (new_AGEMA_signal_3239), .Q (new_AGEMA_signal_5250) ) ;
    buf_clk new_AGEMA_reg_buffer_3298 ( .C (clk), .D (stateArray_S32reg_gff_1_SFF_2_QD), .Q (new_AGEMA_signal_5254) ) ;
    buf_clk new_AGEMA_reg_buffer_3302 ( .C (clk), .D (new_AGEMA_signal_3240), .Q (new_AGEMA_signal_5258) ) ;
    buf_clk new_AGEMA_reg_buffer_3306 ( .C (clk), .D (stateArray_S32reg_gff_1_SFF_3_QD), .Q (new_AGEMA_signal_5262) ) ;
    buf_clk new_AGEMA_reg_buffer_3310 ( .C (clk), .D (new_AGEMA_signal_3241), .Q (new_AGEMA_signal_5266) ) ;
    buf_clk new_AGEMA_reg_buffer_3314 ( .C (clk), .D (stateArray_S32reg_gff_1_SFF_4_QD), .Q (new_AGEMA_signal_5270) ) ;
    buf_clk new_AGEMA_reg_buffer_3318 ( .C (clk), .D (new_AGEMA_signal_3242), .Q (new_AGEMA_signal_5274) ) ;
    buf_clk new_AGEMA_reg_buffer_3322 ( .C (clk), .D (stateArray_S32reg_gff_1_SFF_5_QD), .Q (new_AGEMA_signal_5278) ) ;
    buf_clk new_AGEMA_reg_buffer_3326 ( .C (clk), .D (new_AGEMA_signal_3243), .Q (new_AGEMA_signal_5282) ) ;
    buf_clk new_AGEMA_reg_buffer_3330 ( .C (clk), .D (stateArray_S32reg_gff_1_SFF_6_QD), .Q (new_AGEMA_signal_5286) ) ;
    buf_clk new_AGEMA_reg_buffer_3334 ( .C (clk), .D (new_AGEMA_signal_3244), .Q (new_AGEMA_signal_5290) ) ;
    buf_clk new_AGEMA_reg_buffer_3338 ( .C (clk), .D (stateArray_S32reg_gff_1_SFF_7_QD), .Q (new_AGEMA_signal_5294) ) ;
    buf_clk new_AGEMA_reg_buffer_3342 ( .C (clk), .D (new_AGEMA_signal_3245), .Q (new_AGEMA_signal_5298) ) ;
    buf_clk new_AGEMA_reg_buffer_3346 ( .C (clk), .D (KeyArray_S00reg_gff_1_SFF_0_n5), .Q (new_AGEMA_signal_5302) ) ;
    buf_clk new_AGEMA_reg_buffer_3350 ( .C (clk), .D (new_AGEMA_signal_3375), .Q (new_AGEMA_signal_5306) ) ;
    buf_clk new_AGEMA_reg_buffer_3354 ( .C (clk), .D (KeyArray_S00reg_gff_1_SFF_1_n6), .Q (new_AGEMA_signal_5310) ) ;
    buf_clk new_AGEMA_reg_buffer_3358 ( .C (clk), .D (new_AGEMA_signal_3376), .Q (new_AGEMA_signal_5314) ) ;
    buf_clk new_AGEMA_reg_buffer_3362 ( .C (clk), .D (KeyArray_S00reg_gff_1_SFF_2_n6), .Q (new_AGEMA_signal_5318) ) ;
    buf_clk new_AGEMA_reg_buffer_3366 ( .C (clk), .D (new_AGEMA_signal_3377), .Q (new_AGEMA_signal_5322) ) ;
    buf_clk new_AGEMA_reg_buffer_3370 ( .C (clk), .D (KeyArray_S00reg_gff_1_SFF_3_n6), .Q (new_AGEMA_signal_5326) ) ;
    buf_clk new_AGEMA_reg_buffer_3374 ( .C (clk), .D (new_AGEMA_signal_3378), .Q (new_AGEMA_signal_5330) ) ;
    buf_clk new_AGEMA_reg_buffer_3378 ( .C (clk), .D (KeyArray_S00reg_gff_1_SFF_4_n6), .Q (new_AGEMA_signal_5334) ) ;
    buf_clk new_AGEMA_reg_buffer_3382 ( .C (clk), .D (new_AGEMA_signal_3379), .Q (new_AGEMA_signal_5338) ) ;
    buf_clk new_AGEMA_reg_buffer_3386 ( .C (clk), .D (KeyArray_S00reg_gff_1_SFF_5_n6), .Q (new_AGEMA_signal_5342) ) ;
    buf_clk new_AGEMA_reg_buffer_3390 ( .C (clk), .D (new_AGEMA_signal_3380), .Q (new_AGEMA_signal_5346) ) ;
    buf_clk new_AGEMA_reg_buffer_3394 ( .C (clk), .D (KeyArray_S00reg_gff_1_SFF_6_n6), .Q (new_AGEMA_signal_5350) ) ;
    buf_clk new_AGEMA_reg_buffer_3398 ( .C (clk), .D (new_AGEMA_signal_3381), .Q (new_AGEMA_signal_5354) ) ;
    buf_clk new_AGEMA_reg_buffer_3402 ( .C (clk), .D (KeyArray_S00reg_gff_1_SFF_7_n6), .Q (new_AGEMA_signal_5358) ) ;
    buf_clk new_AGEMA_reg_buffer_3406 ( .C (clk), .D (new_AGEMA_signal_3382), .Q (new_AGEMA_signal_5362) ) ;
    buf_clk new_AGEMA_reg_buffer_3410 ( .C (clk), .D (KeyArray_S01reg_gff_1_SFF_0_n6), .Q (new_AGEMA_signal_5366) ) ;
    buf_clk new_AGEMA_reg_buffer_3414 ( .C (clk), .D (new_AGEMA_signal_3275), .Q (new_AGEMA_signal_5370) ) ;
    buf_clk new_AGEMA_reg_buffer_3418 ( .C (clk), .D (KeyArray_S01reg_gff_1_SFF_1_n6), .Q (new_AGEMA_signal_5374) ) ;
    buf_clk new_AGEMA_reg_buffer_3422 ( .C (clk), .D (new_AGEMA_signal_3276), .Q (new_AGEMA_signal_5378) ) ;
    buf_clk new_AGEMA_reg_buffer_3426 ( .C (clk), .D (KeyArray_S01reg_gff_1_SFF_2_n6), .Q (new_AGEMA_signal_5382) ) ;
    buf_clk new_AGEMA_reg_buffer_3430 ( .C (clk), .D (new_AGEMA_signal_3277), .Q (new_AGEMA_signal_5386) ) ;
    buf_clk new_AGEMA_reg_buffer_3434 ( .C (clk), .D (KeyArray_S01reg_gff_1_SFF_3_n6), .Q (new_AGEMA_signal_5390) ) ;
    buf_clk new_AGEMA_reg_buffer_3438 ( .C (clk), .D (new_AGEMA_signal_3278), .Q (new_AGEMA_signal_5394) ) ;
    buf_clk new_AGEMA_reg_buffer_3442 ( .C (clk), .D (KeyArray_S01reg_gff_1_SFF_4_n6), .Q (new_AGEMA_signal_5398) ) ;
    buf_clk new_AGEMA_reg_buffer_3446 ( .C (clk), .D (new_AGEMA_signal_3279), .Q (new_AGEMA_signal_5402) ) ;
    buf_clk new_AGEMA_reg_buffer_3450 ( .C (clk), .D (KeyArray_S01reg_gff_1_SFF_5_n6), .Q (new_AGEMA_signal_5406) ) ;
    buf_clk new_AGEMA_reg_buffer_3454 ( .C (clk), .D (new_AGEMA_signal_3280), .Q (new_AGEMA_signal_5410) ) ;
    buf_clk new_AGEMA_reg_buffer_3458 ( .C (clk), .D (KeyArray_S01reg_gff_1_SFF_6_n6), .Q (new_AGEMA_signal_5414) ) ;
    buf_clk new_AGEMA_reg_buffer_3462 ( .C (clk), .D (new_AGEMA_signal_3281), .Q (new_AGEMA_signal_5418) ) ;
    buf_clk new_AGEMA_reg_buffer_3466 ( .C (clk), .D (KeyArray_S01reg_gff_1_SFF_7_n6), .Q (new_AGEMA_signal_5422) ) ;
    buf_clk new_AGEMA_reg_buffer_3470 ( .C (clk), .D (new_AGEMA_signal_3282), .Q (new_AGEMA_signal_5426) ) ;
    buf_clk new_AGEMA_reg_buffer_3474 ( .C (clk), .D (KeyArray_S02reg_gff_1_SFF_0_n6), .Q (new_AGEMA_signal_5430) ) ;
    buf_clk new_AGEMA_reg_buffer_3478 ( .C (clk), .D (new_AGEMA_signal_3283), .Q (new_AGEMA_signal_5434) ) ;
    buf_clk new_AGEMA_reg_buffer_3482 ( .C (clk), .D (KeyArray_S02reg_gff_1_SFF_1_n6), .Q (new_AGEMA_signal_5438) ) ;
    buf_clk new_AGEMA_reg_buffer_3486 ( .C (clk), .D (new_AGEMA_signal_3284), .Q (new_AGEMA_signal_5442) ) ;
    buf_clk new_AGEMA_reg_buffer_3490 ( .C (clk), .D (KeyArray_S02reg_gff_1_SFF_2_n6), .Q (new_AGEMA_signal_5446) ) ;
    buf_clk new_AGEMA_reg_buffer_3494 ( .C (clk), .D (new_AGEMA_signal_3285), .Q (new_AGEMA_signal_5450) ) ;
    buf_clk new_AGEMA_reg_buffer_3498 ( .C (clk), .D (KeyArray_S02reg_gff_1_SFF_3_n6), .Q (new_AGEMA_signal_5454) ) ;
    buf_clk new_AGEMA_reg_buffer_3502 ( .C (clk), .D (new_AGEMA_signal_3286), .Q (new_AGEMA_signal_5458) ) ;
    buf_clk new_AGEMA_reg_buffer_3506 ( .C (clk), .D (KeyArray_S02reg_gff_1_SFF_4_n6), .Q (new_AGEMA_signal_5462) ) ;
    buf_clk new_AGEMA_reg_buffer_3510 ( .C (clk), .D (new_AGEMA_signal_3287), .Q (new_AGEMA_signal_5466) ) ;
    buf_clk new_AGEMA_reg_buffer_3514 ( .C (clk), .D (KeyArray_S02reg_gff_1_SFF_5_n6), .Q (new_AGEMA_signal_5470) ) ;
    buf_clk new_AGEMA_reg_buffer_3518 ( .C (clk), .D (new_AGEMA_signal_3288), .Q (new_AGEMA_signal_5474) ) ;
    buf_clk new_AGEMA_reg_buffer_3522 ( .C (clk), .D (KeyArray_S02reg_gff_1_SFF_6_n6), .Q (new_AGEMA_signal_5478) ) ;
    buf_clk new_AGEMA_reg_buffer_3526 ( .C (clk), .D (new_AGEMA_signal_3289), .Q (new_AGEMA_signal_5482) ) ;
    buf_clk new_AGEMA_reg_buffer_3530 ( .C (clk), .D (KeyArray_S02reg_gff_1_SFF_7_n6), .Q (new_AGEMA_signal_5486) ) ;
    buf_clk new_AGEMA_reg_buffer_3534 ( .C (clk), .D (new_AGEMA_signal_3290), .Q (new_AGEMA_signal_5490) ) ;
    buf_clk new_AGEMA_reg_buffer_3538 ( .C (clk), .D (KeyArray_S03reg_gff_1_SFF_0_n6), .Q (new_AGEMA_signal_5494) ) ;
    buf_clk new_AGEMA_reg_buffer_3542 ( .C (clk), .D (new_AGEMA_signal_3291), .Q (new_AGEMA_signal_5498) ) ;
    buf_clk new_AGEMA_reg_buffer_3546 ( .C (clk), .D (KeyArray_S03reg_gff_1_SFF_1_n6), .Q (new_AGEMA_signal_5502) ) ;
    buf_clk new_AGEMA_reg_buffer_3550 ( .C (clk), .D (new_AGEMA_signal_3292), .Q (new_AGEMA_signal_5506) ) ;
    buf_clk new_AGEMA_reg_buffer_3554 ( .C (clk), .D (KeyArray_S03reg_gff_1_SFF_2_n6), .Q (new_AGEMA_signal_5510) ) ;
    buf_clk new_AGEMA_reg_buffer_3558 ( .C (clk), .D (new_AGEMA_signal_3293), .Q (new_AGEMA_signal_5514) ) ;
    buf_clk new_AGEMA_reg_buffer_3562 ( .C (clk), .D (KeyArray_S03reg_gff_1_SFF_3_n6), .Q (new_AGEMA_signal_5518) ) ;
    buf_clk new_AGEMA_reg_buffer_3566 ( .C (clk), .D (new_AGEMA_signal_3294), .Q (new_AGEMA_signal_5522) ) ;
    buf_clk new_AGEMA_reg_buffer_3570 ( .C (clk), .D (KeyArray_S03reg_gff_1_SFF_4_n6), .Q (new_AGEMA_signal_5526) ) ;
    buf_clk new_AGEMA_reg_buffer_3574 ( .C (clk), .D (new_AGEMA_signal_3295), .Q (new_AGEMA_signal_5530) ) ;
    buf_clk new_AGEMA_reg_buffer_3578 ( .C (clk), .D (KeyArray_S03reg_gff_1_SFF_5_n5), .Q (new_AGEMA_signal_5534) ) ;
    buf_clk new_AGEMA_reg_buffer_3582 ( .C (clk), .D (new_AGEMA_signal_3296), .Q (new_AGEMA_signal_5538) ) ;
    buf_clk new_AGEMA_reg_buffer_3586 ( .C (clk), .D (KeyArray_S03reg_gff_1_SFF_6_n5), .Q (new_AGEMA_signal_5542) ) ;
    buf_clk new_AGEMA_reg_buffer_3590 ( .C (clk), .D (new_AGEMA_signal_3297), .Q (new_AGEMA_signal_5546) ) ;
    buf_clk new_AGEMA_reg_buffer_3594 ( .C (clk), .D (KeyArray_S03reg_gff_1_SFF_7_n5), .Q (new_AGEMA_signal_5550) ) ;
    buf_clk new_AGEMA_reg_buffer_3598 ( .C (clk), .D (new_AGEMA_signal_3298), .Q (new_AGEMA_signal_5554) ) ;
    buf_clk new_AGEMA_reg_buffer_3602 ( .C (clk), .D (KeyArray_S10reg_gff_1_SFF_0_n5), .Q (new_AGEMA_signal_5558) ) ;
    buf_clk new_AGEMA_reg_buffer_3606 ( .C (clk), .D (new_AGEMA_signal_3299), .Q (new_AGEMA_signal_5562) ) ;
    buf_clk new_AGEMA_reg_buffer_3610 ( .C (clk), .D (KeyArray_S10reg_gff_1_SFF_1_n5), .Q (new_AGEMA_signal_5566) ) ;
    buf_clk new_AGEMA_reg_buffer_3614 ( .C (clk), .D (new_AGEMA_signal_3300), .Q (new_AGEMA_signal_5570) ) ;
    buf_clk new_AGEMA_reg_buffer_3618 ( .C (clk), .D (KeyArray_S10reg_gff_1_SFF_2_n5), .Q (new_AGEMA_signal_5574) ) ;
    buf_clk new_AGEMA_reg_buffer_3622 ( .C (clk), .D (new_AGEMA_signal_3301), .Q (new_AGEMA_signal_5578) ) ;
    buf_clk new_AGEMA_reg_buffer_3626 ( .C (clk), .D (KeyArray_S10reg_gff_1_SFF_3_n5), .Q (new_AGEMA_signal_5582) ) ;
    buf_clk new_AGEMA_reg_buffer_3630 ( .C (clk), .D (new_AGEMA_signal_3302), .Q (new_AGEMA_signal_5586) ) ;
    buf_clk new_AGEMA_reg_buffer_3634 ( .C (clk), .D (KeyArray_S10reg_gff_1_SFF_4_n5), .Q (new_AGEMA_signal_5590) ) ;
    buf_clk new_AGEMA_reg_buffer_3638 ( .C (clk), .D (new_AGEMA_signal_3303), .Q (new_AGEMA_signal_5594) ) ;
    buf_clk new_AGEMA_reg_buffer_3642 ( .C (clk), .D (KeyArray_S10reg_gff_1_SFF_5_n5), .Q (new_AGEMA_signal_5598) ) ;
    buf_clk new_AGEMA_reg_buffer_3646 ( .C (clk), .D (new_AGEMA_signal_3304), .Q (new_AGEMA_signal_5602) ) ;
    buf_clk new_AGEMA_reg_buffer_3650 ( .C (clk), .D (KeyArray_S10reg_gff_1_SFF_6_n5), .Q (new_AGEMA_signal_5606) ) ;
    buf_clk new_AGEMA_reg_buffer_3654 ( .C (clk), .D (new_AGEMA_signal_3305), .Q (new_AGEMA_signal_5610) ) ;
    buf_clk new_AGEMA_reg_buffer_3658 ( .C (clk), .D (KeyArray_S10reg_gff_1_SFF_7_n5), .Q (new_AGEMA_signal_5614) ) ;
    buf_clk new_AGEMA_reg_buffer_3662 ( .C (clk), .D (new_AGEMA_signal_3306), .Q (new_AGEMA_signal_5618) ) ;
    buf_clk new_AGEMA_reg_buffer_3666 ( .C (clk), .D (KeyArray_S11reg_gff_1_SFF_0_n6), .Q (new_AGEMA_signal_5622) ) ;
    buf_clk new_AGEMA_reg_buffer_3670 ( .C (clk), .D (new_AGEMA_signal_3307), .Q (new_AGEMA_signal_5626) ) ;
    buf_clk new_AGEMA_reg_buffer_3674 ( .C (clk), .D (KeyArray_S11reg_gff_1_SFF_1_n6), .Q (new_AGEMA_signal_5630) ) ;
    buf_clk new_AGEMA_reg_buffer_3678 ( .C (clk), .D (new_AGEMA_signal_3308), .Q (new_AGEMA_signal_5634) ) ;
    buf_clk new_AGEMA_reg_buffer_3682 ( .C (clk), .D (KeyArray_S11reg_gff_1_SFF_2_n6), .Q (new_AGEMA_signal_5638) ) ;
    buf_clk new_AGEMA_reg_buffer_3686 ( .C (clk), .D (new_AGEMA_signal_3309), .Q (new_AGEMA_signal_5642) ) ;
    buf_clk new_AGEMA_reg_buffer_3690 ( .C (clk), .D (KeyArray_S11reg_gff_1_SFF_3_n6), .Q (new_AGEMA_signal_5646) ) ;
    buf_clk new_AGEMA_reg_buffer_3694 ( .C (clk), .D (new_AGEMA_signal_3310), .Q (new_AGEMA_signal_5650) ) ;
    buf_clk new_AGEMA_reg_buffer_3698 ( .C (clk), .D (KeyArray_S11reg_gff_1_SFF_4_n6), .Q (new_AGEMA_signal_5654) ) ;
    buf_clk new_AGEMA_reg_buffer_3702 ( .C (clk), .D (new_AGEMA_signal_3311), .Q (new_AGEMA_signal_5658) ) ;
    buf_clk new_AGEMA_reg_buffer_3706 ( .C (clk), .D (KeyArray_S11reg_gff_1_SFF_5_n6), .Q (new_AGEMA_signal_5662) ) ;
    buf_clk new_AGEMA_reg_buffer_3710 ( .C (clk), .D (new_AGEMA_signal_3312), .Q (new_AGEMA_signal_5666) ) ;
    buf_clk new_AGEMA_reg_buffer_3714 ( .C (clk), .D (KeyArray_S11reg_gff_1_SFF_6_n6), .Q (new_AGEMA_signal_5670) ) ;
    buf_clk new_AGEMA_reg_buffer_3718 ( .C (clk), .D (new_AGEMA_signal_3313), .Q (new_AGEMA_signal_5674) ) ;
    buf_clk new_AGEMA_reg_buffer_3722 ( .C (clk), .D (KeyArray_S11reg_gff_1_SFF_7_n6), .Q (new_AGEMA_signal_5678) ) ;
    buf_clk new_AGEMA_reg_buffer_3726 ( .C (clk), .D (new_AGEMA_signal_3314), .Q (new_AGEMA_signal_5682) ) ;
    buf_clk new_AGEMA_reg_buffer_3730 ( .C (clk), .D (KeyArray_S12reg_gff_1_SFF_0_n6), .Q (new_AGEMA_signal_5686) ) ;
    buf_clk new_AGEMA_reg_buffer_3734 ( .C (clk), .D (new_AGEMA_signal_3093), .Q (new_AGEMA_signal_5690) ) ;
    buf_clk new_AGEMA_reg_buffer_3738 ( .C (clk), .D (KeyArray_S12reg_gff_1_SFF_1_n6), .Q (new_AGEMA_signal_5694) ) ;
    buf_clk new_AGEMA_reg_buffer_3742 ( .C (clk), .D (new_AGEMA_signal_3094), .Q (new_AGEMA_signal_5698) ) ;
    buf_clk new_AGEMA_reg_buffer_3746 ( .C (clk), .D (KeyArray_S12reg_gff_1_SFF_2_n6), .Q (new_AGEMA_signal_5702) ) ;
    buf_clk new_AGEMA_reg_buffer_3750 ( .C (clk), .D (new_AGEMA_signal_3095), .Q (new_AGEMA_signal_5706) ) ;
    buf_clk new_AGEMA_reg_buffer_3754 ( .C (clk), .D (KeyArray_S12reg_gff_1_SFF_3_n6), .Q (new_AGEMA_signal_5710) ) ;
    buf_clk new_AGEMA_reg_buffer_3758 ( .C (clk), .D (new_AGEMA_signal_3096), .Q (new_AGEMA_signal_5714) ) ;
    buf_clk new_AGEMA_reg_buffer_3762 ( .C (clk), .D (KeyArray_S12reg_gff_1_SFF_4_n6), .Q (new_AGEMA_signal_5718) ) ;
    buf_clk new_AGEMA_reg_buffer_3766 ( .C (clk), .D (new_AGEMA_signal_3097), .Q (new_AGEMA_signal_5722) ) ;
    buf_clk new_AGEMA_reg_buffer_3770 ( .C (clk), .D (KeyArray_S12reg_gff_1_SFF_5_n6), .Q (new_AGEMA_signal_5726) ) ;
    buf_clk new_AGEMA_reg_buffer_3774 ( .C (clk), .D (new_AGEMA_signal_3098), .Q (new_AGEMA_signal_5730) ) ;
    buf_clk new_AGEMA_reg_buffer_3778 ( .C (clk), .D (KeyArray_S12reg_gff_1_SFF_6_n6), .Q (new_AGEMA_signal_5734) ) ;
    buf_clk new_AGEMA_reg_buffer_3782 ( .C (clk), .D (new_AGEMA_signal_3099), .Q (new_AGEMA_signal_5738) ) ;
    buf_clk new_AGEMA_reg_buffer_3786 ( .C (clk), .D (KeyArray_S12reg_gff_1_SFF_7_n6), .Q (new_AGEMA_signal_5742) ) ;
    buf_clk new_AGEMA_reg_buffer_3790 ( .C (clk), .D (new_AGEMA_signal_3100), .Q (new_AGEMA_signal_5746) ) ;
    buf_clk new_AGEMA_reg_buffer_3794 ( .C (clk), .D (KeyArray_S13reg_gff_1_SFF_0_n6), .Q (new_AGEMA_signal_5750) ) ;
    buf_clk new_AGEMA_reg_buffer_3798 ( .C (clk), .D (new_AGEMA_signal_3101), .Q (new_AGEMA_signal_5754) ) ;
    buf_clk new_AGEMA_reg_buffer_3802 ( .C (clk), .D (KeyArray_S13reg_gff_1_SFF_1_n6), .Q (new_AGEMA_signal_5758) ) ;
    buf_clk new_AGEMA_reg_buffer_3806 ( .C (clk), .D (new_AGEMA_signal_3102), .Q (new_AGEMA_signal_5762) ) ;
    buf_clk new_AGEMA_reg_buffer_3810 ( .C (clk), .D (KeyArray_S13reg_gff_1_SFF_2_n6), .Q (new_AGEMA_signal_5766) ) ;
    buf_clk new_AGEMA_reg_buffer_3814 ( .C (clk), .D (new_AGEMA_signal_3103), .Q (new_AGEMA_signal_5770) ) ;
    buf_clk new_AGEMA_reg_buffer_3818 ( .C (clk), .D (KeyArray_S13reg_gff_1_SFF_3_n6), .Q (new_AGEMA_signal_5774) ) ;
    buf_clk new_AGEMA_reg_buffer_3822 ( .C (clk), .D (new_AGEMA_signal_3104), .Q (new_AGEMA_signal_5778) ) ;
    buf_clk new_AGEMA_reg_buffer_3826 ( .C (clk), .D (KeyArray_S13reg_gff_1_SFF_4_n6), .Q (new_AGEMA_signal_5782) ) ;
    buf_clk new_AGEMA_reg_buffer_3830 ( .C (clk), .D (new_AGEMA_signal_3105), .Q (new_AGEMA_signal_5786) ) ;
    buf_clk new_AGEMA_reg_buffer_3834 ( .C (clk), .D (KeyArray_S13reg_gff_1_SFF_5_n5), .Q (new_AGEMA_signal_5790) ) ;
    buf_clk new_AGEMA_reg_buffer_3838 ( .C (clk), .D (new_AGEMA_signal_3106), .Q (new_AGEMA_signal_5794) ) ;
    buf_clk new_AGEMA_reg_buffer_3842 ( .C (clk), .D (KeyArray_S13reg_gff_1_SFF_6_n5), .Q (new_AGEMA_signal_5798) ) ;
    buf_clk new_AGEMA_reg_buffer_3846 ( .C (clk), .D (new_AGEMA_signal_3107), .Q (new_AGEMA_signal_5802) ) ;
    buf_clk new_AGEMA_reg_buffer_3850 ( .C (clk), .D (KeyArray_S13reg_gff_1_SFF_7_n5), .Q (new_AGEMA_signal_5806) ) ;
    buf_clk new_AGEMA_reg_buffer_3854 ( .C (clk), .D (new_AGEMA_signal_3108), .Q (new_AGEMA_signal_5810) ) ;
    buf_clk new_AGEMA_reg_buffer_3858 ( .C (clk), .D (KeyArray_S20reg_gff_1_SFF_0_n5), .Q (new_AGEMA_signal_5814) ) ;
    buf_clk new_AGEMA_reg_buffer_3862 ( .C (clk), .D (new_AGEMA_signal_3315), .Q (new_AGEMA_signal_5818) ) ;
    buf_clk new_AGEMA_reg_buffer_3866 ( .C (clk), .D (KeyArray_S20reg_gff_1_SFF_1_n5), .Q (new_AGEMA_signal_5822) ) ;
    buf_clk new_AGEMA_reg_buffer_3870 ( .C (clk), .D (new_AGEMA_signal_3316), .Q (new_AGEMA_signal_5826) ) ;
    buf_clk new_AGEMA_reg_buffer_3874 ( .C (clk), .D (KeyArray_S20reg_gff_1_SFF_2_n5), .Q (new_AGEMA_signal_5830) ) ;
    buf_clk new_AGEMA_reg_buffer_3878 ( .C (clk), .D (new_AGEMA_signal_3317), .Q (new_AGEMA_signal_5834) ) ;
    buf_clk new_AGEMA_reg_buffer_3882 ( .C (clk), .D (KeyArray_S20reg_gff_1_SFF_3_n5), .Q (new_AGEMA_signal_5838) ) ;
    buf_clk new_AGEMA_reg_buffer_3886 ( .C (clk), .D (new_AGEMA_signal_3318), .Q (new_AGEMA_signal_5842) ) ;
    buf_clk new_AGEMA_reg_buffer_3890 ( .C (clk), .D (KeyArray_S20reg_gff_1_SFF_4_n5), .Q (new_AGEMA_signal_5846) ) ;
    buf_clk new_AGEMA_reg_buffer_3894 ( .C (clk), .D (new_AGEMA_signal_3319), .Q (new_AGEMA_signal_5850) ) ;
    buf_clk new_AGEMA_reg_buffer_3898 ( .C (clk), .D (KeyArray_S20reg_gff_1_SFF_5_n5), .Q (new_AGEMA_signal_5854) ) ;
    buf_clk new_AGEMA_reg_buffer_3902 ( .C (clk), .D (new_AGEMA_signal_3320), .Q (new_AGEMA_signal_5858) ) ;
    buf_clk new_AGEMA_reg_buffer_3906 ( .C (clk), .D (KeyArray_S20reg_gff_1_SFF_6_n5), .Q (new_AGEMA_signal_5862) ) ;
    buf_clk new_AGEMA_reg_buffer_3910 ( .C (clk), .D (new_AGEMA_signal_3321), .Q (new_AGEMA_signal_5866) ) ;
    buf_clk new_AGEMA_reg_buffer_3914 ( .C (clk), .D (KeyArray_S20reg_gff_1_SFF_7_n5), .Q (new_AGEMA_signal_5870) ) ;
    buf_clk new_AGEMA_reg_buffer_3918 ( .C (clk), .D (new_AGEMA_signal_3322), .Q (new_AGEMA_signal_5874) ) ;
    buf_clk new_AGEMA_reg_buffer_3922 ( .C (clk), .D (KeyArray_S21reg_gff_1_SFF_0_n6), .Q (new_AGEMA_signal_5878) ) ;
    buf_clk new_AGEMA_reg_buffer_3926 ( .C (clk), .D (new_AGEMA_signal_3323), .Q (new_AGEMA_signal_5882) ) ;
    buf_clk new_AGEMA_reg_buffer_3930 ( .C (clk), .D (KeyArray_S21reg_gff_1_SFF_1_n6), .Q (new_AGEMA_signal_5886) ) ;
    buf_clk new_AGEMA_reg_buffer_3934 ( .C (clk), .D (new_AGEMA_signal_3324), .Q (new_AGEMA_signal_5890) ) ;
    buf_clk new_AGEMA_reg_buffer_3938 ( .C (clk), .D (KeyArray_S21reg_gff_1_SFF_2_n6), .Q (new_AGEMA_signal_5894) ) ;
    buf_clk new_AGEMA_reg_buffer_3942 ( .C (clk), .D (new_AGEMA_signal_3325), .Q (new_AGEMA_signal_5898) ) ;
    buf_clk new_AGEMA_reg_buffer_3946 ( .C (clk), .D (KeyArray_S21reg_gff_1_SFF_3_n6), .Q (new_AGEMA_signal_5902) ) ;
    buf_clk new_AGEMA_reg_buffer_3950 ( .C (clk), .D (new_AGEMA_signal_3326), .Q (new_AGEMA_signal_5906) ) ;
    buf_clk new_AGEMA_reg_buffer_3954 ( .C (clk), .D (KeyArray_S21reg_gff_1_SFF_4_n6), .Q (new_AGEMA_signal_5910) ) ;
    buf_clk new_AGEMA_reg_buffer_3958 ( .C (clk), .D (new_AGEMA_signal_3327), .Q (new_AGEMA_signal_5914) ) ;
    buf_clk new_AGEMA_reg_buffer_3962 ( .C (clk), .D (KeyArray_S21reg_gff_1_SFF_5_n6), .Q (new_AGEMA_signal_5918) ) ;
    buf_clk new_AGEMA_reg_buffer_3966 ( .C (clk), .D (new_AGEMA_signal_3328), .Q (new_AGEMA_signal_5922) ) ;
    buf_clk new_AGEMA_reg_buffer_3970 ( .C (clk), .D (KeyArray_S21reg_gff_1_SFF_6_n6), .Q (new_AGEMA_signal_5926) ) ;
    buf_clk new_AGEMA_reg_buffer_3974 ( .C (clk), .D (new_AGEMA_signal_3329), .Q (new_AGEMA_signal_5930) ) ;
    buf_clk new_AGEMA_reg_buffer_3978 ( .C (clk), .D (KeyArray_S21reg_gff_1_SFF_7_n6), .Q (new_AGEMA_signal_5934) ) ;
    buf_clk new_AGEMA_reg_buffer_3982 ( .C (clk), .D (new_AGEMA_signal_3330), .Q (new_AGEMA_signal_5938) ) ;
    buf_clk new_AGEMA_reg_buffer_3986 ( .C (clk), .D (KeyArray_S22reg_gff_1_SFF_0_n6), .Q (new_AGEMA_signal_5942) ) ;
    buf_clk new_AGEMA_reg_buffer_3990 ( .C (clk), .D (new_AGEMA_signal_3331), .Q (new_AGEMA_signal_5946) ) ;
    buf_clk new_AGEMA_reg_buffer_3994 ( .C (clk), .D (KeyArray_S22reg_gff_1_SFF_1_n6), .Q (new_AGEMA_signal_5950) ) ;
    buf_clk new_AGEMA_reg_buffer_3998 ( .C (clk), .D (new_AGEMA_signal_3332), .Q (new_AGEMA_signal_5954) ) ;
    buf_clk new_AGEMA_reg_buffer_4002 ( .C (clk), .D (KeyArray_S22reg_gff_1_SFF_2_n6), .Q (new_AGEMA_signal_5958) ) ;
    buf_clk new_AGEMA_reg_buffer_4006 ( .C (clk), .D (new_AGEMA_signal_3333), .Q (new_AGEMA_signal_5962) ) ;
    buf_clk new_AGEMA_reg_buffer_4010 ( .C (clk), .D (KeyArray_S22reg_gff_1_SFF_3_n6), .Q (new_AGEMA_signal_5966) ) ;
    buf_clk new_AGEMA_reg_buffer_4014 ( .C (clk), .D (new_AGEMA_signal_3334), .Q (new_AGEMA_signal_5970) ) ;
    buf_clk new_AGEMA_reg_buffer_4018 ( .C (clk), .D (KeyArray_S22reg_gff_1_SFF_4_n6), .Q (new_AGEMA_signal_5974) ) ;
    buf_clk new_AGEMA_reg_buffer_4022 ( .C (clk), .D (new_AGEMA_signal_3335), .Q (new_AGEMA_signal_5978) ) ;
    buf_clk new_AGEMA_reg_buffer_4026 ( .C (clk), .D (KeyArray_S22reg_gff_1_SFF_5_n6), .Q (new_AGEMA_signal_5982) ) ;
    buf_clk new_AGEMA_reg_buffer_4030 ( .C (clk), .D (new_AGEMA_signal_3336), .Q (new_AGEMA_signal_5986) ) ;
    buf_clk new_AGEMA_reg_buffer_4034 ( .C (clk), .D (KeyArray_S22reg_gff_1_SFF_6_n6), .Q (new_AGEMA_signal_5990) ) ;
    buf_clk new_AGEMA_reg_buffer_4038 ( .C (clk), .D (new_AGEMA_signal_3337), .Q (new_AGEMA_signal_5994) ) ;
    buf_clk new_AGEMA_reg_buffer_4042 ( .C (clk), .D (KeyArray_S22reg_gff_1_SFF_7_n6), .Q (new_AGEMA_signal_5998) ) ;
    buf_clk new_AGEMA_reg_buffer_4046 ( .C (clk), .D (new_AGEMA_signal_3338), .Q (new_AGEMA_signal_6002) ) ;
    buf_clk new_AGEMA_reg_buffer_4050 ( .C (clk), .D (KeyArray_S23reg_gff_1_SFF_0_n6), .Q (new_AGEMA_signal_6006) ) ;
    buf_clk new_AGEMA_reg_buffer_4054 ( .C (clk), .D (new_AGEMA_signal_3339), .Q (new_AGEMA_signal_6010) ) ;
    buf_clk new_AGEMA_reg_buffer_4058 ( .C (clk), .D (KeyArray_S23reg_gff_1_SFF_1_n6), .Q (new_AGEMA_signal_6014) ) ;
    buf_clk new_AGEMA_reg_buffer_4062 ( .C (clk), .D (new_AGEMA_signal_3340), .Q (new_AGEMA_signal_6018) ) ;
    buf_clk new_AGEMA_reg_buffer_4066 ( .C (clk), .D (KeyArray_S23reg_gff_1_SFF_2_n6), .Q (new_AGEMA_signal_6022) ) ;
    buf_clk new_AGEMA_reg_buffer_4070 ( .C (clk), .D (new_AGEMA_signal_3341), .Q (new_AGEMA_signal_6026) ) ;
    buf_clk new_AGEMA_reg_buffer_4074 ( .C (clk), .D (KeyArray_S23reg_gff_1_SFF_3_n6), .Q (new_AGEMA_signal_6030) ) ;
    buf_clk new_AGEMA_reg_buffer_4078 ( .C (clk), .D (new_AGEMA_signal_3342), .Q (new_AGEMA_signal_6034) ) ;
    buf_clk new_AGEMA_reg_buffer_4082 ( .C (clk), .D (KeyArray_S23reg_gff_1_SFF_4_n6), .Q (new_AGEMA_signal_6038) ) ;
    buf_clk new_AGEMA_reg_buffer_4086 ( .C (clk), .D (new_AGEMA_signal_3343), .Q (new_AGEMA_signal_6042) ) ;
    buf_clk new_AGEMA_reg_buffer_4090 ( .C (clk), .D (KeyArray_S23reg_gff_1_SFF_5_n5), .Q (new_AGEMA_signal_6046) ) ;
    buf_clk new_AGEMA_reg_buffer_4094 ( .C (clk), .D (new_AGEMA_signal_3344), .Q (new_AGEMA_signal_6050) ) ;
    buf_clk new_AGEMA_reg_buffer_4098 ( .C (clk), .D (KeyArray_S23reg_gff_1_SFF_6_n5), .Q (new_AGEMA_signal_6054) ) ;
    buf_clk new_AGEMA_reg_buffer_4102 ( .C (clk), .D (new_AGEMA_signal_3345), .Q (new_AGEMA_signal_6058) ) ;
    buf_clk new_AGEMA_reg_buffer_4106 ( .C (clk), .D (KeyArray_S23reg_gff_1_SFF_7_n5), .Q (new_AGEMA_signal_6062) ) ;
    buf_clk new_AGEMA_reg_buffer_4110 ( .C (clk), .D (new_AGEMA_signal_3346), .Q (new_AGEMA_signal_6066) ) ;
    buf_clk new_AGEMA_reg_buffer_4114 ( .C (clk), .D (KeyArray_S31reg_gff_1_SFF_0_n6), .Q (new_AGEMA_signal_6070) ) ;
    buf_clk new_AGEMA_reg_buffer_4118 ( .C (clk), .D (new_AGEMA_signal_3347), .Q (new_AGEMA_signal_6074) ) ;
    buf_clk new_AGEMA_reg_buffer_4122 ( .C (clk), .D (KeyArray_S31reg_gff_1_SFF_1_n6), .Q (new_AGEMA_signal_6078) ) ;
    buf_clk new_AGEMA_reg_buffer_4126 ( .C (clk), .D (new_AGEMA_signal_3348), .Q (new_AGEMA_signal_6082) ) ;
    buf_clk new_AGEMA_reg_buffer_4130 ( .C (clk), .D (KeyArray_S31reg_gff_1_SFF_2_n6), .Q (new_AGEMA_signal_6086) ) ;
    buf_clk new_AGEMA_reg_buffer_4134 ( .C (clk), .D (new_AGEMA_signal_3349), .Q (new_AGEMA_signal_6090) ) ;
    buf_clk new_AGEMA_reg_buffer_4138 ( .C (clk), .D (KeyArray_S31reg_gff_1_SFF_3_n6), .Q (new_AGEMA_signal_6094) ) ;
    buf_clk new_AGEMA_reg_buffer_4142 ( .C (clk), .D (new_AGEMA_signal_3350), .Q (new_AGEMA_signal_6098) ) ;
    buf_clk new_AGEMA_reg_buffer_4146 ( .C (clk), .D (KeyArray_S31reg_gff_1_SFF_4_n6), .Q (new_AGEMA_signal_6102) ) ;
    buf_clk new_AGEMA_reg_buffer_4150 ( .C (clk), .D (new_AGEMA_signal_3351), .Q (new_AGEMA_signal_6106) ) ;
    buf_clk new_AGEMA_reg_buffer_4154 ( .C (clk), .D (KeyArray_S31reg_gff_1_SFF_5_n6), .Q (new_AGEMA_signal_6110) ) ;
    buf_clk new_AGEMA_reg_buffer_4158 ( .C (clk), .D (new_AGEMA_signal_3352), .Q (new_AGEMA_signal_6114) ) ;
    buf_clk new_AGEMA_reg_buffer_4162 ( .C (clk), .D (KeyArray_S31reg_gff_1_SFF_6_n6), .Q (new_AGEMA_signal_6118) ) ;
    buf_clk new_AGEMA_reg_buffer_4166 ( .C (clk), .D (new_AGEMA_signal_3353), .Q (new_AGEMA_signal_6122) ) ;
    buf_clk new_AGEMA_reg_buffer_4170 ( .C (clk), .D (KeyArray_S31reg_gff_1_SFF_7_n6), .Q (new_AGEMA_signal_6126) ) ;
    buf_clk new_AGEMA_reg_buffer_4174 ( .C (clk), .D (new_AGEMA_signal_3354), .Q (new_AGEMA_signal_6130) ) ;
    buf_clk new_AGEMA_reg_buffer_4178 ( .C (clk), .D (KeyArray_S32reg_gff_1_SFF_0_n6), .Q (new_AGEMA_signal_6134) ) ;
    buf_clk new_AGEMA_reg_buffer_4182 ( .C (clk), .D (new_AGEMA_signal_3355), .Q (new_AGEMA_signal_6138) ) ;
    buf_clk new_AGEMA_reg_buffer_4186 ( .C (clk), .D (KeyArray_S32reg_gff_1_SFF_1_n6), .Q (new_AGEMA_signal_6142) ) ;
    buf_clk new_AGEMA_reg_buffer_4190 ( .C (clk), .D (new_AGEMA_signal_3356), .Q (new_AGEMA_signal_6146) ) ;
    buf_clk new_AGEMA_reg_buffer_4194 ( .C (clk), .D (KeyArray_S32reg_gff_1_SFF_2_n6), .Q (new_AGEMA_signal_6150) ) ;
    buf_clk new_AGEMA_reg_buffer_4198 ( .C (clk), .D (new_AGEMA_signal_3357), .Q (new_AGEMA_signal_6154) ) ;
    buf_clk new_AGEMA_reg_buffer_4202 ( .C (clk), .D (KeyArray_S32reg_gff_1_SFF_3_n6), .Q (new_AGEMA_signal_6158) ) ;
    buf_clk new_AGEMA_reg_buffer_4206 ( .C (clk), .D (new_AGEMA_signal_3358), .Q (new_AGEMA_signal_6162) ) ;
    buf_clk new_AGEMA_reg_buffer_4210 ( .C (clk), .D (KeyArray_S32reg_gff_1_SFF_4_n6), .Q (new_AGEMA_signal_6166) ) ;
    buf_clk new_AGEMA_reg_buffer_4214 ( .C (clk), .D (new_AGEMA_signal_3359), .Q (new_AGEMA_signal_6170) ) ;
    buf_clk new_AGEMA_reg_buffer_4218 ( .C (clk), .D (KeyArray_S32reg_gff_1_SFF_5_n6), .Q (new_AGEMA_signal_6174) ) ;
    buf_clk new_AGEMA_reg_buffer_4222 ( .C (clk), .D (new_AGEMA_signal_3360), .Q (new_AGEMA_signal_6178) ) ;
    buf_clk new_AGEMA_reg_buffer_4226 ( .C (clk), .D (KeyArray_S32reg_gff_1_SFF_6_n5), .Q (new_AGEMA_signal_6182) ) ;
    buf_clk new_AGEMA_reg_buffer_4230 ( .C (clk), .D (new_AGEMA_signal_3361), .Q (new_AGEMA_signal_6186) ) ;
    buf_clk new_AGEMA_reg_buffer_4234 ( .C (clk), .D (KeyArray_S32reg_gff_1_SFF_7_n5), .Q (new_AGEMA_signal_6190) ) ;
    buf_clk new_AGEMA_reg_buffer_4238 ( .C (clk), .D (new_AGEMA_signal_3362), .Q (new_AGEMA_signal_6194) ) ;
    buf_clk new_AGEMA_reg_buffer_4242 ( .C (clk), .D (KeyArray_S33reg_gff_1_SFF_0_n5), .Q (new_AGEMA_signal_6198) ) ;
    buf_clk new_AGEMA_reg_buffer_4246 ( .C (clk), .D (new_AGEMA_signal_3363), .Q (new_AGEMA_signal_6202) ) ;
    buf_clk new_AGEMA_reg_buffer_4250 ( .C (clk), .D (KeyArray_S33reg_gff_1_SFF_1_n5), .Q (new_AGEMA_signal_6206) ) ;
    buf_clk new_AGEMA_reg_buffer_4254 ( .C (clk), .D (new_AGEMA_signal_3364), .Q (new_AGEMA_signal_6210) ) ;
    buf_clk new_AGEMA_reg_buffer_4258 ( .C (clk), .D (KeyArray_S33reg_gff_1_SFF_2_n5), .Q (new_AGEMA_signal_6214) ) ;
    buf_clk new_AGEMA_reg_buffer_4262 ( .C (clk), .D (new_AGEMA_signal_3365), .Q (new_AGEMA_signal_6218) ) ;
    buf_clk new_AGEMA_reg_buffer_4266 ( .C (clk), .D (KeyArray_S33reg_gff_1_SFF_3_n5), .Q (new_AGEMA_signal_6222) ) ;
    buf_clk new_AGEMA_reg_buffer_4270 ( .C (clk), .D (new_AGEMA_signal_3366), .Q (new_AGEMA_signal_6226) ) ;
    buf_clk new_AGEMA_reg_buffer_4274 ( .C (clk), .D (KeyArray_S33reg_gff_1_SFF_4_n5), .Q (new_AGEMA_signal_6230) ) ;
    buf_clk new_AGEMA_reg_buffer_4278 ( .C (clk), .D (new_AGEMA_signal_3367), .Q (new_AGEMA_signal_6234) ) ;
    buf_clk new_AGEMA_reg_buffer_4282 ( .C (clk), .D (KeyArray_S33reg_gff_1_SFF_5_n5), .Q (new_AGEMA_signal_6238) ) ;
    buf_clk new_AGEMA_reg_buffer_4286 ( .C (clk), .D (new_AGEMA_signal_3368), .Q (new_AGEMA_signal_6242) ) ;
    buf_clk new_AGEMA_reg_buffer_4290 ( .C (clk), .D (KeyArray_S33reg_gff_1_SFF_6_n5), .Q (new_AGEMA_signal_6246) ) ;
    buf_clk new_AGEMA_reg_buffer_4294 ( .C (clk), .D (new_AGEMA_signal_3369), .Q (new_AGEMA_signal_6250) ) ;
    buf_clk new_AGEMA_reg_buffer_4298 ( .C (clk), .D (KeyArray_S33reg_gff_1_SFF_7_n5), .Q (new_AGEMA_signal_6254) ) ;
    buf_clk new_AGEMA_reg_buffer_4302 ( .C (clk), .D (new_AGEMA_signal_3370), .Q (new_AGEMA_signal_6258) ) ;
    buf_clk new_AGEMA_reg_buffer_4306 ( .C (clk), .D (calcRCon_n51), .Q (new_AGEMA_signal_6262) ) ;
    buf_clk new_AGEMA_reg_buffer_4310 ( .C (clk), .D (calcRCon_n50), .Q (new_AGEMA_signal_6266) ) ;
    buf_clk new_AGEMA_reg_buffer_4314 ( .C (clk), .D (calcRCon_n49), .Q (new_AGEMA_signal_6270) ) ;
    buf_clk new_AGEMA_reg_buffer_4318 ( .C (clk), .D (calcRCon_n48), .Q (new_AGEMA_signal_6274) ) ;
    buf_clk new_AGEMA_reg_buffer_4322 ( .C (clk), .D (calcRCon_n47), .Q (new_AGEMA_signal_6278) ) ;
    buf_clk new_AGEMA_reg_buffer_4326 ( .C (clk), .D (calcRCon_n46), .Q (new_AGEMA_signal_6282) ) ;
    buf_clk new_AGEMA_reg_buffer_4330 ( .C (clk), .D (calcRCon_n45), .Q (new_AGEMA_signal_6286) ) ;
    buf_clk new_AGEMA_reg_buffer_4334 ( .C (clk), .D (calcRCon_n44), .Q (new_AGEMA_signal_6290) ) ;
    buf_clk new_AGEMA_reg_buffer_4338 ( .C (clk), .D (n9), .Q (new_AGEMA_signal_6294) ) ;

    /* cells in depth 2 */
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M25_U1 ( .a ({new_AGEMA_signal_3374, Inst_bSbox_M22}), .b ({new_AGEMA_signal_3372, Inst_bSbox_M20}), .clk (clk), .r ({Fresh[39], Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_3384, Inst_bSbox_M25}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_M26_U1 ( .a ({new_AGEMA_signal_3679, new_AGEMA_signal_3678}), .b ({new_AGEMA_signal_3384, Inst_bSbox_M25}), .c ({new_AGEMA_signal_3388, Inst_bSbox_M26}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_M28_U1 ( .a ({new_AGEMA_signal_3681, new_AGEMA_signal_3680}), .b ({new_AGEMA_signal_3384, Inst_bSbox_M25}), .c ({new_AGEMA_signal_3389, Inst_bSbox_M28}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M31_U1 ( .a ({new_AGEMA_signal_3372, Inst_bSbox_M20}), .b ({new_AGEMA_signal_3383, Inst_bSbox_M23}), .clk (clk), .r ({Fresh[43], Fresh[42], Fresh[41], Fresh[40]}), .c ({new_AGEMA_signal_3390, Inst_bSbox_M31}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_M33_U1 ( .a ({new_AGEMA_signal_3683, new_AGEMA_signal_3682}), .b ({new_AGEMA_signal_3384, Inst_bSbox_M25}), .c ({new_AGEMA_signal_3391, Inst_bSbox_M33}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M34_U1 ( .a ({new_AGEMA_signal_3373, Inst_bSbox_M21}), .b ({new_AGEMA_signal_3374, Inst_bSbox_M22}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44]}), .c ({new_AGEMA_signal_3386, Inst_bSbox_M34}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_M36_U1 ( .a ({new_AGEMA_signal_3685, new_AGEMA_signal_3684}), .b ({new_AGEMA_signal_3384, Inst_bSbox_M25}), .c ({new_AGEMA_signal_3396, Inst_bSbox_M36}) ) ;
    buf_clk new_AGEMA_reg_buffer_1722 ( .C (clk), .D (Inst_bSbox_M21), .Q (new_AGEMA_signal_3678) ) ;
    buf_clk new_AGEMA_reg_buffer_1723 ( .C (clk), .D (new_AGEMA_signal_3373), .Q (new_AGEMA_signal_3679) ) ;
    buf_clk new_AGEMA_reg_buffer_1724 ( .C (clk), .D (Inst_bSbox_M23), .Q (new_AGEMA_signal_3680) ) ;
    buf_clk new_AGEMA_reg_buffer_1725 ( .C (clk), .D (new_AGEMA_signal_3383), .Q (new_AGEMA_signal_3681) ) ;
    buf_clk new_AGEMA_reg_buffer_1726 ( .C (clk), .D (Inst_bSbox_M27), .Q (new_AGEMA_signal_3682) ) ;
    buf_clk new_AGEMA_reg_buffer_1727 ( .C (clk), .D (new_AGEMA_signal_3385), .Q (new_AGEMA_signal_3683) ) ;
    buf_clk new_AGEMA_reg_buffer_1728 ( .C (clk), .D (Inst_bSbox_M24), .Q (new_AGEMA_signal_3684) ) ;
    buf_clk new_AGEMA_reg_buffer_1729 ( .C (clk), .D (new_AGEMA_signal_3387), .Q (new_AGEMA_signal_3685) ) ;
    buf_clk new_AGEMA_reg_buffer_1739 ( .C (clk), .D (new_AGEMA_signal_3694), .Q (new_AGEMA_signal_3695) ) ;
    buf_clk new_AGEMA_reg_buffer_1743 ( .C (clk), .D (new_AGEMA_signal_3698), .Q (new_AGEMA_signal_3699) ) ;
    buf_clk new_AGEMA_reg_buffer_1747 ( .C (clk), .D (new_AGEMA_signal_3702), .Q (new_AGEMA_signal_3703) ) ;
    buf_clk new_AGEMA_reg_buffer_1751 ( .C (clk), .D (new_AGEMA_signal_3706), .Q (new_AGEMA_signal_3707) ) ;
    buf_clk new_AGEMA_reg_buffer_1755 ( .C (clk), .D (new_AGEMA_signal_3710), .Q (new_AGEMA_signal_3711) ) ;
    buf_clk new_AGEMA_reg_buffer_1759 ( .C (clk), .D (new_AGEMA_signal_3714), .Q (new_AGEMA_signal_3715) ) ;
    buf_clk new_AGEMA_reg_buffer_1763 ( .C (clk), .D (new_AGEMA_signal_3718), .Q (new_AGEMA_signal_3719) ) ;
    buf_clk new_AGEMA_reg_buffer_1767 ( .C (clk), .D (new_AGEMA_signal_3722), .Q (new_AGEMA_signal_3723) ) ;
    buf_clk new_AGEMA_reg_buffer_1771 ( .C (clk), .D (new_AGEMA_signal_3726), .Q (new_AGEMA_signal_3727) ) ;
    buf_clk new_AGEMA_reg_buffer_1775 ( .C (clk), .D (new_AGEMA_signal_3730), .Q (new_AGEMA_signal_3731) ) ;
    buf_clk new_AGEMA_reg_buffer_1779 ( .C (clk), .D (new_AGEMA_signal_3734), .Q (new_AGEMA_signal_3735) ) ;
    buf_clk new_AGEMA_reg_buffer_1783 ( .C (clk), .D (new_AGEMA_signal_3738), .Q (new_AGEMA_signal_3739) ) ;
    buf_clk new_AGEMA_reg_buffer_1787 ( .C (clk), .D (new_AGEMA_signal_3742), .Q (new_AGEMA_signal_3743) ) ;
    buf_clk new_AGEMA_reg_buffer_1791 ( .C (clk), .D (new_AGEMA_signal_3746), .Q (new_AGEMA_signal_3747) ) ;
    buf_clk new_AGEMA_reg_buffer_1795 ( .C (clk), .D (new_AGEMA_signal_3750), .Q (new_AGEMA_signal_3751) ) ;
    buf_clk new_AGEMA_reg_buffer_1799 ( .C (clk), .D (new_AGEMA_signal_3754), .Q (new_AGEMA_signal_3755) ) ;
    buf_clk new_AGEMA_reg_buffer_1803 ( .C (clk), .D (new_AGEMA_signal_3758), .Q (new_AGEMA_signal_3759) ) ;
    buf_clk new_AGEMA_reg_buffer_1807 ( .C (clk), .D (new_AGEMA_signal_3762), .Q (new_AGEMA_signal_3763) ) ;
    buf_clk new_AGEMA_reg_buffer_1811 ( .C (clk), .D (new_AGEMA_signal_3766), .Q (new_AGEMA_signal_3767) ) ;
    buf_clk new_AGEMA_reg_buffer_1815 ( .C (clk), .D (new_AGEMA_signal_3770), .Q (new_AGEMA_signal_3771) ) ;
    buf_clk new_AGEMA_reg_buffer_1819 ( .C (clk), .D (new_AGEMA_signal_3774), .Q (new_AGEMA_signal_3775) ) ;
    buf_clk new_AGEMA_reg_buffer_1823 ( .C (clk), .D (new_AGEMA_signal_3778), .Q (new_AGEMA_signal_3779) ) ;
    buf_clk new_AGEMA_reg_buffer_1827 ( .C (clk), .D (new_AGEMA_signal_3782), .Q (new_AGEMA_signal_3783) ) ;
    buf_clk new_AGEMA_reg_buffer_1831 ( .C (clk), .D (new_AGEMA_signal_3786), .Q (new_AGEMA_signal_3787) ) ;
    buf_clk new_AGEMA_reg_buffer_1835 ( .C (clk), .D (new_AGEMA_signal_3790), .Q (new_AGEMA_signal_3791) ) ;
    buf_clk new_AGEMA_reg_buffer_1839 ( .C (clk), .D (new_AGEMA_signal_3794), .Q (new_AGEMA_signal_3795) ) ;
    buf_clk new_AGEMA_reg_buffer_1843 ( .C (clk), .D (new_AGEMA_signal_3798), .Q (new_AGEMA_signal_3799) ) ;
    buf_clk new_AGEMA_reg_buffer_1847 ( .C (clk), .D (new_AGEMA_signal_3802), .Q (new_AGEMA_signal_3803) ) ;
    buf_clk new_AGEMA_reg_buffer_1851 ( .C (clk), .D (new_AGEMA_signal_3806), .Q (new_AGEMA_signal_3807) ) ;
    buf_clk new_AGEMA_reg_buffer_1855 ( .C (clk), .D (new_AGEMA_signal_3810), .Q (new_AGEMA_signal_3811) ) ;
    buf_clk new_AGEMA_reg_buffer_1859 ( .C (clk), .D (new_AGEMA_signal_3814), .Q (new_AGEMA_signal_3815) ) ;
    buf_clk new_AGEMA_reg_buffer_1863 ( .C (clk), .D (new_AGEMA_signal_3818), .Q (new_AGEMA_signal_3819) ) ;
    buf_clk new_AGEMA_reg_buffer_1867 ( .C (clk), .D (new_AGEMA_signal_3822), .Q (new_AGEMA_signal_3823) ) ;
    buf_clk new_AGEMA_reg_buffer_1871 ( .C (clk), .D (new_AGEMA_signal_3826), .Q (new_AGEMA_signal_3827) ) ;
    buf_clk new_AGEMA_reg_buffer_1875 ( .C (clk), .D (new_AGEMA_signal_3830), .Q (new_AGEMA_signal_3831) ) ;
    buf_clk new_AGEMA_reg_buffer_1879 ( .C (clk), .D (new_AGEMA_signal_3834), .Q (new_AGEMA_signal_3835) ) ;
    buf_clk new_AGEMA_reg_buffer_1883 ( .C (clk), .D (new_AGEMA_signal_3838), .Q (new_AGEMA_signal_3839) ) ;
    buf_clk new_AGEMA_reg_buffer_1887 ( .C (clk), .D (new_AGEMA_signal_3842), .Q (new_AGEMA_signal_3843) ) ;
    buf_clk new_AGEMA_reg_buffer_1891 ( .C (clk), .D (new_AGEMA_signal_3846), .Q (new_AGEMA_signal_3847) ) ;
    buf_clk new_AGEMA_reg_buffer_1895 ( .C (clk), .D (new_AGEMA_signal_3850), .Q (new_AGEMA_signal_3851) ) ;
    buf_clk new_AGEMA_reg_buffer_1899 ( .C (clk), .D (new_AGEMA_signal_3854), .Q (new_AGEMA_signal_3855) ) ;
    buf_clk new_AGEMA_reg_buffer_1903 ( .C (clk), .D (new_AGEMA_signal_3858), .Q (new_AGEMA_signal_3859) ) ;
    buf_clk new_AGEMA_reg_buffer_1907 ( .C (clk), .D (new_AGEMA_signal_3862), .Q (new_AGEMA_signal_3863) ) ;
    buf_clk new_AGEMA_reg_buffer_1911 ( .C (clk), .D (new_AGEMA_signal_3866), .Q (new_AGEMA_signal_3867) ) ;
    buf_clk new_AGEMA_reg_buffer_1915 ( .C (clk), .D (new_AGEMA_signal_3870), .Q (new_AGEMA_signal_3871) ) ;
    buf_clk new_AGEMA_reg_buffer_1919 ( .C (clk), .D (new_AGEMA_signal_3874), .Q (new_AGEMA_signal_3875) ) ;
    buf_clk new_AGEMA_reg_buffer_1923 ( .C (clk), .D (new_AGEMA_signal_3878), .Q (new_AGEMA_signal_3879) ) ;
    buf_clk new_AGEMA_reg_buffer_1927 ( .C (clk), .D (new_AGEMA_signal_3882), .Q (new_AGEMA_signal_3883) ) ;
    buf_clk new_AGEMA_reg_buffer_1931 ( .C (clk), .D (new_AGEMA_signal_3886), .Q (new_AGEMA_signal_3887) ) ;
    buf_clk new_AGEMA_reg_buffer_1935 ( .C (clk), .D (new_AGEMA_signal_3890), .Q (new_AGEMA_signal_3891) ) ;
    buf_clk new_AGEMA_reg_buffer_1939 ( .C (clk), .D (new_AGEMA_signal_3894), .Q (new_AGEMA_signal_3895) ) ;
    buf_clk new_AGEMA_reg_buffer_1943 ( .C (clk), .D (new_AGEMA_signal_3898), .Q (new_AGEMA_signal_3899) ) ;
    buf_clk new_AGEMA_reg_buffer_1947 ( .C (clk), .D (new_AGEMA_signal_3902), .Q (new_AGEMA_signal_3903) ) ;
    buf_clk new_AGEMA_reg_buffer_1951 ( .C (clk), .D (new_AGEMA_signal_3906), .Q (new_AGEMA_signal_3907) ) ;
    buf_clk new_AGEMA_reg_buffer_1955 ( .C (clk), .D (new_AGEMA_signal_3910), .Q (new_AGEMA_signal_3911) ) ;
    buf_clk new_AGEMA_reg_buffer_1959 ( .C (clk), .D (new_AGEMA_signal_3914), .Q (new_AGEMA_signal_3915) ) ;
    buf_clk new_AGEMA_reg_buffer_1963 ( .C (clk), .D (new_AGEMA_signal_3918), .Q (new_AGEMA_signal_3919) ) ;
    buf_clk new_AGEMA_reg_buffer_1967 ( .C (clk), .D (new_AGEMA_signal_3922), .Q (new_AGEMA_signal_3923) ) ;
    buf_clk new_AGEMA_reg_buffer_1971 ( .C (clk), .D (new_AGEMA_signal_3926), .Q (new_AGEMA_signal_3927) ) ;
    buf_clk new_AGEMA_reg_buffer_1975 ( .C (clk), .D (new_AGEMA_signal_3930), .Q (new_AGEMA_signal_3931) ) ;
    buf_clk new_AGEMA_reg_buffer_1979 ( .C (clk), .D (new_AGEMA_signal_3934), .Q (new_AGEMA_signal_3935) ) ;
    buf_clk new_AGEMA_reg_buffer_1983 ( .C (clk), .D (new_AGEMA_signal_3938), .Q (new_AGEMA_signal_3939) ) ;
    buf_clk new_AGEMA_reg_buffer_1987 ( .C (clk), .D (new_AGEMA_signal_3942), .Q (new_AGEMA_signal_3943) ) ;
    buf_clk new_AGEMA_reg_buffer_1991 ( .C (clk), .D (new_AGEMA_signal_3946), .Q (new_AGEMA_signal_3947) ) ;
    buf_clk new_AGEMA_reg_buffer_1995 ( .C (clk), .D (new_AGEMA_signal_3950), .Q (new_AGEMA_signal_3951) ) ;
    buf_clk new_AGEMA_reg_buffer_1999 ( .C (clk), .D (new_AGEMA_signal_3954), .Q (new_AGEMA_signal_3955) ) ;
    buf_clk new_AGEMA_reg_buffer_2003 ( .C (clk), .D (new_AGEMA_signal_3958), .Q (new_AGEMA_signal_3959) ) ;
    buf_clk new_AGEMA_reg_buffer_2007 ( .C (clk), .D (new_AGEMA_signal_3962), .Q (new_AGEMA_signal_3963) ) ;
    buf_clk new_AGEMA_reg_buffer_2011 ( .C (clk), .D (new_AGEMA_signal_3966), .Q (new_AGEMA_signal_3967) ) ;
    buf_clk new_AGEMA_reg_buffer_2015 ( .C (clk), .D (new_AGEMA_signal_3970), .Q (new_AGEMA_signal_3971) ) ;
    buf_clk new_AGEMA_reg_buffer_2019 ( .C (clk), .D (new_AGEMA_signal_3974), .Q (new_AGEMA_signal_3975) ) ;
    buf_clk new_AGEMA_reg_buffer_2023 ( .C (clk), .D (new_AGEMA_signal_3978), .Q (new_AGEMA_signal_3979) ) ;
    buf_clk new_AGEMA_reg_buffer_2027 ( .C (clk), .D (new_AGEMA_signal_3982), .Q (new_AGEMA_signal_3983) ) ;
    buf_clk new_AGEMA_reg_buffer_2031 ( .C (clk), .D (new_AGEMA_signal_3986), .Q (new_AGEMA_signal_3987) ) ;
    buf_clk new_AGEMA_reg_buffer_2035 ( .C (clk), .D (new_AGEMA_signal_3990), .Q (new_AGEMA_signal_3991) ) ;
    buf_clk new_AGEMA_reg_buffer_2039 ( .C (clk), .D (new_AGEMA_signal_3994), .Q (new_AGEMA_signal_3995) ) ;
    buf_clk new_AGEMA_reg_buffer_2043 ( .C (clk), .D (new_AGEMA_signal_3998), .Q (new_AGEMA_signal_3999) ) ;
    buf_clk new_AGEMA_reg_buffer_2047 ( .C (clk), .D (new_AGEMA_signal_4002), .Q (new_AGEMA_signal_4003) ) ;
    buf_clk new_AGEMA_reg_buffer_2051 ( .C (clk), .D (new_AGEMA_signal_4006), .Q (new_AGEMA_signal_4007) ) ;
    buf_clk new_AGEMA_reg_buffer_2055 ( .C (clk), .D (new_AGEMA_signal_4010), .Q (new_AGEMA_signal_4011) ) ;
    buf_clk new_AGEMA_reg_buffer_2059 ( .C (clk), .D (new_AGEMA_signal_4014), .Q (new_AGEMA_signal_4015) ) ;
    buf_clk new_AGEMA_reg_buffer_2063 ( .C (clk), .D (new_AGEMA_signal_4018), .Q (new_AGEMA_signal_4019) ) ;
    buf_clk new_AGEMA_reg_buffer_2067 ( .C (clk), .D (new_AGEMA_signal_4022), .Q (new_AGEMA_signal_4023) ) ;
    buf_clk new_AGEMA_reg_buffer_2071 ( .C (clk), .D (new_AGEMA_signal_4026), .Q (new_AGEMA_signal_4027) ) ;
    buf_clk new_AGEMA_reg_buffer_2075 ( .C (clk), .D (new_AGEMA_signal_4030), .Q (new_AGEMA_signal_4031) ) ;
    buf_clk new_AGEMA_reg_buffer_2079 ( .C (clk), .D (new_AGEMA_signal_4034), .Q (new_AGEMA_signal_4035) ) ;
    buf_clk new_AGEMA_reg_buffer_2083 ( .C (clk), .D (new_AGEMA_signal_4038), .Q (new_AGEMA_signal_4039) ) ;
    buf_clk new_AGEMA_reg_buffer_2087 ( .C (clk), .D (new_AGEMA_signal_4042), .Q (new_AGEMA_signal_4043) ) ;
    buf_clk new_AGEMA_reg_buffer_2091 ( .C (clk), .D (new_AGEMA_signal_4046), .Q (new_AGEMA_signal_4047) ) ;
    buf_clk new_AGEMA_reg_buffer_2095 ( .C (clk), .D (new_AGEMA_signal_4050), .Q (new_AGEMA_signal_4051) ) ;
    buf_clk new_AGEMA_reg_buffer_2099 ( .C (clk), .D (new_AGEMA_signal_4054), .Q (new_AGEMA_signal_4055) ) ;
    buf_clk new_AGEMA_reg_buffer_2103 ( .C (clk), .D (new_AGEMA_signal_4058), .Q (new_AGEMA_signal_4059) ) ;
    buf_clk new_AGEMA_reg_buffer_2107 ( .C (clk), .D (new_AGEMA_signal_4062), .Q (new_AGEMA_signal_4063) ) ;
    buf_clk new_AGEMA_reg_buffer_2111 ( .C (clk), .D (new_AGEMA_signal_4066), .Q (new_AGEMA_signal_4067) ) ;
    buf_clk new_AGEMA_reg_buffer_2115 ( .C (clk), .D (new_AGEMA_signal_4070), .Q (new_AGEMA_signal_4071) ) ;
    buf_clk new_AGEMA_reg_buffer_2119 ( .C (clk), .D (new_AGEMA_signal_4074), .Q (new_AGEMA_signal_4075) ) ;
    buf_clk new_AGEMA_reg_buffer_2123 ( .C (clk), .D (new_AGEMA_signal_4078), .Q (new_AGEMA_signal_4079) ) ;
    buf_clk new_AGEMA_reg_buffer_2127 ( .C (clk), .D (new_AGEMA_signal_4082), .Q (new_AGEMA_signal_4083) ) ;
    buf_clk new_AGEMA_reg_buffer_2131 ( .C (clk), .D (new_AGEMA_signal_4086), .Q (new_AGEMA_signal_4087) ) ;
    buf_clk new_AGEMA_reg_buffer_2135 ( .C (clk), .D (new_AGEMA_signal_4090), .Q (new_AGEMA_signal_4091) ) ;
    buf_clk new_AGEMA_reg_buffer_2139 ( .C (clk), .D (new_AGEMA_signal_4094), .Q (new_AGEMA_signal_4095) ) ;
    buf_clk new_AGEMA_reg_buffer_2143 ( .C (clk), .D (new_AGEMA_signal_4098), .Q (new_AGEMA_signal_4099) ) ;
    buf_clk new_AGEMA_reg_buffer_2147 ( .C (clk), .D (new_AGEMA_signal_4102), .Q (new_AGEMA_signal_4103) ) ;
    buf_clk new_AGEMA_reg_buffer_2151 ( .C (clk), .D (new_AGEMA_signal_4106), .Q (new_AGEMA_signal_4107) ) ;
    buf_clk new_AGEMA_reg_buffer_2155 ( .C (clk), .D (new_AGEMA_signal_4110), .Q (new_AGEMA_signal_4111) ) ;
    buf_clk new_AGEMA_reg_buffer_2159 ( .C (clk), .D (new_AGEMA_signal_4114), .Q (new_AGEMA_signal_4115) ) ;
    buf_clk new_AGEMA_reg_buffer_2163 ( .C (clk), .D (new_AGEMA_signal_4118), .Q (new_AGEMA_signal_4119) ) ;
    buf_clk new_AGEMA_reg_buffer_2167 ( .C (clk), .D (new_AGEMA_signal_4122), .Q (new_AGEMA_signal_4123) ) ;
    buf_clk new_AGEMA_reg_buffer_2171 ( .C (clk), .D (new_AGEMA_signal_4126), .Q (new_AGEMA_signal_4127) ) ;
    buf_clk new_AGEMA_reg_buffer_2175 ( .C (clk), .D (new_AGEMA_signal_4130), .Q (new_AGEMA_signal_4131) ) ;
    buf_clk new_AGEMA_reg_buffer_2179 ( .C (clk), .D (new_AGEMA_signal_4134), .Q (new_AGEMA_signal_4135) ) ;
    buf_clk new_AGEMA_reg_buffer_2183 ( .C (clk), .D (new_AGEMA_signal_4138), .Q (new_AGEMA_signal_4139) ) ;
    buf_clk new_AGEMA_reg_buffer_2187 ( .C (clk), .D (new_AGEMA_signal_4142), .Q (new_AGEMA_signal_4143) ) ;
    buf_clk new_AGEMA_reg_buffer_2191 ( .C (clk), .D (new_AGEMA_signal_4146), .Q (new_AGEMA_signal_4147) ) ;
    buf_clk new_AGEMA_reg_buffer_2195 ( .C (clk), .D (new_AGEMA_signal_4150), .Q (new_AGEMA_signal_4151) ) ;
    buf_clk new_AGEMA_reg_buffer_2199 ( .C (clk), .D (new_AGEMA_signal_4154), .Q (new_AGEMA_signal_4155) ) ;
    buf_clk new_AGEMA_reg_buffer_2203 ( .C (clk), .D (new_AGEMA_signal_4158), .Q (new_AGEMA_signal_4159) ) ;
    buf_clk new_AGEMA_reg_buffer_2207 ( .C (clk), .D (new_AGEMA_signal_4162), .Q (new_AGEMA_signal_4163) ) ;
    buf_clk new_AGEMA_reg_buffer_2211 ( .C (clk), .D (new_AGEMA_signal_4166), .Q (new_AGEMA_signal_4167) ) ;
    buf_clk new_AGEMA_reg_buffer_2215 ( .C (clk), .D (new_AGEMA_signal_4170), .Q (new_AGEMA_signal_4171) ) ;
    buf_clk new_AGEMA_reg_buffer_2219 ( .C (clk), .D (new_AGEMA_signal_4174), .Q (new_AGEMA_signal_4175) ) ;
    buf_clk new_AGEMA_reg_buffer_2223 ( .C (clk), .D (new_AGEMA_signal_4178), .Q (new_AGEMA_signal_4179) ) ;
    buf_clk new_AGEMA_reg_buffer_2227 ( .C (clk), .D (new_AGEMA_signal_4182), .Q (new_AGEMA_signal_4183) ) ;
    buf_clk new_AGEMA_reg_buffer_2231 ( .C (clk), .D (new_AGEMA_signal_4186), .Q (new_AGEMA_signal_4187) ) ;
    buf_clk new_AGEMA_reg_buffer_2235 ( .C (clk), .D (new_AGEMA_signal_4190), .Q (new_AGEMA_signal_4191) ) ;
    buf_clk new_AGEMA_reg_buffer_2239 ( .C (clk), .D (new_AGEMA_signal_4194), .Q (new_AGEMA_signal_4195) ) ;
    buf_clk new_AGEMA_reg_buffer_2243 ( .C (clk), .D (new_AGEMA_signal_4198), .Q (new_AGEMA_signal_4199) ) ;
    buf_clk new_AGEMA_reg_buffer_2246 ( .C (clk), .D (new_AGEMA_signal_4201), .Q (new_AGEMA_signal_4202) ) ;
    buf_clk new_AGEMA_reg_buffer_2249 ( .C (clk), .D (new_AGEMA_signal_4204), .Q (new_AGEMA_signal_4205) ) ;
    buf_clk new_AGEMA_reg_buffer_2252 ( .C (clk), .D (new_AGEMA_signal_4207), .Q (new_AGEMA_signal_4208) ) ;
    buf_clk new_AGEMA_reg_buffer_2255 ( .C (clk), .D (new_AGEMA_signal_4210), .Q (new_AGEMA_signal_4211) ) ;
    buf_clk new_AGEMA_reg_buffer_2258 ( .C (clk), .D (new_AGEMA_signal_4213), .Q (new_AGEMA_signal_4214) ) ;
    buf_clk new_AGEMA_reg_buffer_2261 ( .C (clk), .D (new_AGEMA_signal_4216), .Q (new_AGEMA_signal_4217) ) ;
    buf_clk new_AGEMA_reg_buffer_2264 ( .C (clk), .D (new_AGEMA_signal_4219), .Q (new_AGEMA_signal_4220) ) ;
    buf_clk new_AGEMA_reg_buffer_2267 ( .C (clk), .D (new_AGEMA_signal_4222), .Q (new_AGEMA_signal_4223) ) ;
    buf_clk new_AGEMA_reg_buffer_2270 ( .C (clk), .D (new_AGEMA_signal_4225), .Q (new_AGEMA_signal_4226) ) ;
    buf_clk new_AGEMA_reg_buffer_2273 ( .C (clk), .D (new_AGEMA_signal_4228), .Q (new_AGEMA_signal_4229) ) ;
    buf_clk new_AGEMA_reg_buffer_2276 ( .C (clk), .D (new_AGEMA_signal_4231), .Q (new_AGEMA_signal_4232) ) ;
    buf_clk new_AGEMA_reg_buffer_2279 ( .C (clk), .D (new_AGEMA_signal_4234), .Q (new_AGEMA_signal_4235) ) ;
    buf_clk new_AGEMA_reg_buffer_2282 ( .C (clk), .D (new_AGEMA_signal_4237), .Q (new_AGEMA_signal_4238) ) ;
    buf_clk new_AGEMA_reg_buffer_2285 ( .C (clk), .D (new_AGEMA_signal_4240), .Q (new_AGEMA_signal_4241) ) ;
    buf_clk new_AGEMA_reg_buffer_2288 ( .C (clk), .D (new_AGEMA_signal_4243), .Q (new_AGEMA_signal_4244) ) ;
    buf_clk new_AGEMA_reg_buffer_2291 ( .C (clk), .D (new_AGEMA_signal_4246), .Q (new_AGEMA_signal_4247) ) ;
    buf_clk new_AGEMA_reg_buffer_2294 ( .C (clk), .D (new_AGEMA_signal_4249), .Q (new_AGEMA_signal_4250) ) ;
    buf_clk new_AGEMA_reg_buffer_2297 ( .C (clk), .D (new_AGEMA_signal_4252), .Q (new_AGEMA_signal_4253) ) ;
    buf_clk new_AGEMA_reg_buffer_2300 ( .C (clk), .D (new_AGEMA_signal_4255), .Q (new_AGEMA_signal_4256) ) ;
    buf_clk new_AGEMA_reg_buffer_2303 ( .C (clk), .D (new_AGEMA_signal_4258), .Q (new_AGEMA_signal_4259) ) ;
    buf_clk new_AGEMA_reg_buffer_2306 ( .C (clk), .D (new_AGEMA_signal_4261), .Q (new_AGEMA_signal_4262) ) ;
    buf_clk new_AGEMA_reg_buffer_2309 ( .C (clk), .D (new_AGEMA_signal_4264), .Q (new_AGEMA_signal_4265) ) ;
    buf_clk new_AGEMA_reg_buffer_2312 ( .C (clk), .D (new_AGEMA_signal_4267), .Q (new_AGEMA_signal_4268) ) ;
    buf_clk new_AGEMA_reg_buffer_2315 ( .C (clk), .D (new_AGEMA_signal_4270), .Q (new_AGEMA_signal_4271) ) ;
    buf_clk new_AGEMA_reg_buffer_2318 ( .C (clk), .D (new_AGEMA_signal_4273), .Q (new_AGEMA_signal_4274) ) ;
    buf_clk new_AGEMA_reg_buffer_2321 ( .C (clk), .D (new_AGEMA_signal_4276), .Q (new_AGEMA_signal_4277) ) ;
    buf_clk new_AGEMA_reg_buffer_2324 ( .C (clk), .D (new_AGEMA_signal_4279), .Q (new_AGEMA_signal_4280) ) ;
    buf_clk new_AGEMA_reg_buffer_2327 ( .C (clk), .D (new_AGEMA_signal_4282), .Q (new_AGEMA_signal_4283) ) ;
    buf_clk new_AGEMA_reg_buffer_2330 ( .C (clk), .D (new_AGEMA_signal_4285), .Q (new_AGEMA_signal_4286) ) ;
    buf_clk new_AGEMA_reg_buffer_2333 ( .C (clk), .D (new_AGEMA_signal_4288), .Q (new_AGEMA_signal_4289) ) ;
    buf_clk new_AGEMA_reg_buffer_2336 ( .C (clk), .D (new_AGEMA_signal_4291), .Q (new_AGEMA_signal_4292) ) ;
    buf_clk new_AGEMA_reg_buffer_2339 ( .C (clk), .D (new_AGEMA_signal_4294), .Q (new_AGEMA_signal_4295) ) ;
    buf_clk new_AGEMA_reg_buffer_2342 ( .C (clk), .D (new_AGEMA_signal_4297), .Q (new_AGEMA_signal_4298) ) ;
    buf_clk new_AGEMA_reg_buffer_2345 ( .C (clk), .D (new_AGEMA_signal_4300), .Q (new_AGEMA_signal_4301) ) ;
    buf_clk new_AGEMA_reg_buffer_2348 ( .C (clk), .D (new_AGEMA_signal_4303), .Q (new_AGEMA_signal_4304) ) ;
    buf_clk new_AGEMA_reg_buffer_2351 ( .C (clk), .D (new_AGEMA_signal_4306), .Q (new_AGEMA_signal_4307) ) ;
    buf_clk new_AGEMA_reg_buffer_2355 ( .C (clk), .D (new_AGEMA_signal_4310), .Q (new_AGEMA_signal_4311) ) ;
    buf_clk new_AGEMA_reg_buffer_2359 ( .C (clk), .D (new_AGEMA_signal_4314), .Q (new_AGEMA_signal_4315) ) ;
    buf_clk new_AGEMA_reg_buffer_2363 ( .C (clk), .D (new_AGEMA_signal_4318), .Q (new_AGEMA_signal_4319) ) ;
    buf_clk new_AGEMA_reg_buffer_2367 ( .C (clk), .D (new_AGEMA_signal_4322), .Q (new_AGEMA_signal_4323) ) ;
    buf_clk new_AGEMA_reg_buffer_2371 ( .C (clk), .D (new_AGEMA_signal_4326), .Q (new_AGEMA_signal_4327) ) ;
    buf_clk new_AGEMA_reg_buffer_2375 ( .C (clk), .D (new_AGEMA_signal_4330), .Q (new_AGEMA_signal_4331) ) ;
    buf_clk new_AGEMA_reg_buffer_2379 ( .C (clk), .D (new_AGEMA_signal_4334), .Q (new_AGEMA_signal_4335) ) ;
    buf_clk new_AGEMA_reg_buffer_2383 ( .C (clk), .D (new_AGEMA_signal_4338), .Q (new_AGEMA_signal_4339) ) ;
    buf_clk new_AGEMA_reg_buffer_2387 ( .C (clk), .D (new_AGEMA_signal_4342), .Q (new_AGEMA_signal_4343) ) ;
    buf_clk new_AGEMA_reg_buffer_2391 ( .C (clk), .D (new_AGEMA_signal_4346), .Q (new_AGEMA_signal_4347) ) ;
    buf_clk new_AGEMA_reg_buffer_2395 ( .C (clk), .D (new_AGEMA_signal_4350), .Q (new_AGEMA_signal_4351) ) ;
    buf_clk new_AGEMA_reg_buffer_2399 ( .C (clk), .D (new_AGEMA_signal_4354), .Q (new_AGEMA_signal_4355) ) ;
    buf_clk new_AGEMA_reg_buffer_2403 ( .C (clk), .D (new_AGEMA_signal_4358), .Q (new_AGEMA_signal_4359) ) ;
    buf_clk new_AGEMA_reg_buffer_2407 ( .C (clk), .D (new_AGEMA_signal_4362), .Q (new_AGEMA_signal_4363) ) ;
    buf_clk new_AGEMA_reg_buffer_2411 ( .C (clk), .D (new_AGEMA_signal_4366), .Q (new_AGEMA_signal_4367) ) ;
    buf_clk new_AGEMA_reg_buffer_2415 ( .C (clk), .D (new_AGEMA_signal_4370), .Q (new_AGEMA_signal_4371) ) ;
    buf_clk new_AGEMA_reg_buffer_2419 ( .C (clk), .D (new_AGEMA_signal_4374), .Q (new_AGEMA_signal_4375) ) ;
    buf_clk new_AGEMA_reg_buffer_2423 ( .C (clk), .D (new_AGEMA_signal_4378), .Q (new_AGEMA_signal_4379) ) ;
    buf_clk new_AGEMA_reg_buffer_2427 ( .C (clk), .D (new_AGEMA_signal_4382), .Q (new_AGEMA_signal_4383) ) ;
    buf_clk new_AGEMA_reg_buffer_2431 ( .C (clk), .D (new_AGEMA_signal_4386), .Q (new_AGEMA_signal_4387) ) ;
    buf_clk new_AGEMA_reg_buffer_2435 ( .C (clk), .D (new_AGEMA_signal_4390), .Q (new_AGEMA_signal_4391) ) ;
    buf_clk new_AGEMA_reg_buffer_2439 ( .C (clk), .D (new_AGEMA_signal_4394), .Q (new_AGEMA_signal_4395) ) ;
    buf_clk new_AGEMA_reg_buffer_2443 ( .C (clk), .D (new_AGEMA_signal_4398), .Q (new_AGEMA_signal_4399) ) ;
    buf_clk new_AGEMA_reg_buffer_2447 ( .C (clk), .D (new_AGEMA_signal_4402), .Q (new_AGEMA_signal_4403) ) ;
    buf_clk new_AGEMA_reg_buffer_2451 ( .C (clk), .D (new_AGEMA_signal_4406), .Q (new_AGEMA_signal_4407) ) ;
    buf_clk new_AGEMA_reg_buffer_2455 ( .C (clk), .D (new_AGEMA_signal_4410), .Q (new_AGEMA_signal_4411) ) ;
    buf_clk new_AGEMA_reg_buffer_2459 ( .C (clk), .D (new_AGEMA_signal_4414), .Q (new_AGEMA_signal_4415) ) ;
    buf_clk new_AGEMA_reg_buffer_2463 ( .C (clk), .D (new_AGEMA_signal_4418), .Q (new_AGEMA_signal_4419) ) ;
    buf_clk new_AGEMA_reg_buffer_2467 ( .C (clk), .D (new_AGEMA_signal_4422), .Q (new_AGEMA_signal_4423) ) ;
    buf_clk new_AGEMA_reg_buffer_2471 ( .C (clk), .D (new_AGEMA_signal_4426), .Q (new_AGEMA_signal_4427) ) ;
    buf_clk new_AGEMA_reg_buffer_2475 ( .C (clk), .D (new_AGEMA_signal_4430), .Q (new_AGEMA_signal_4431) ) ;
    buf_clk new_AGEMA_reg_buffer_2479 ( .C (clk), .D (new_AGEMA_signal_4434), .Q (new_AGEMA_signal_4435) ) ;
    buf_clk new_AGEMA_reg_buffer_2483 ( .C (clk), .D (new_AGEMA_signal_4438), .Q (new_AGEMA_signal_4439) ) ;
    buf_clk new_AGEMA_reg_buffer_2487 ( .C (clk), .D (new_AGEMA_signal_4442), .Q (new_AGEMA_signal_4443) ) ;
    buf_clk new_AGEMA_reg_buffer_2491 ( .C (clk), .D (new_AGEMA_signal_4446), .Q (new_AGEMA_signal_4447) ) ;
    buf_clk new_AGEMA_reg_buffer_2495 ( .C (clk), .D (new_AGEMA_signal_4450), .Q (new_AGEMA_signal_4451) ) ;
    buf_clk new_AGEMA_reg_buffer_2499 ( .C (clk), .D (new_AGEMA_signal_4454), .Q (new_AGEMA_signal_4455) ) ;
    buf_clk new_AGEMA_reg_buffer_2503 ( .C (clk), .D (new_AGEMA_signal_4458), .Q (new_AGEMA_signal_4459) ) ;
    buf_clk new_AGEMA_reg_buffer_2507 ( .C (clk), .D (new_AGEMA_signal_4462), .Q (new_AGEMA_signal_4463) ) ;
    buf_clk new_AGEMA_reg_buffer_2511 ( .C (clk), .D (new_AGEMA_signal_4466), .Q (new_AGEMA_signal_4467) ) ;
    buf_clk new_AGEMA_reg_buffer_2515 ( .C (clk), .D (new_AGEMA_signal_4470), .Q (new_AGEMA_signal_4471) ) ;
    buf_clk new_AGEMA_reg_buffer_2519 ( .C (clk), .D (new_AGEMA_signal_4474), .Q (new_AGEMA_signal_4475) ) ;
    buf_clk new_AGEMA_reg_buffer_2523 ( .C (clk), .D (new_AGEMA_signal_4478), .Q (new_AGEMA_signal_4479) ) ;
    buf_clk new_AGEMA_reg_buffer_2527 ( .C (clk), .D (new_AGEMA_signal_4482), .Q (new_AGEMA_signal_4483) ) ;
    buf_clk new_AGEMA_reg_buffer_2531 ( .C (clk), .D (new_AGEMA_signal_4486), .Q (new_AGEMA_signal_4487) ) ;
    buf_clk new_AGEMA_reg_buffer_2535 ( .C (clk), .D (new_AGEMA_signal_4490), .Q (new_AGEMA_signal_4491) ) ;
    buf_clk new_AGEMA_reg_buffer_2539 ( .C (clk), .D (new_AGEMA_signal_4494), .Q (new_AGEMA_signal_4495) ) ;
    buf_clk new_AGEMA_reg_buffer_2543 ( .C (clk), .D (new_AGEMA_signal_4498), .Q (new_AGEMA_signal_4499) ) ;
    buf_clk new_AGEMA_reg_buffer_2547 ( .C (clk), .D (new_AGEMA_signal_4502), .Q (new_AGEMA_signal_4503) ) ;
    buf_clk new_AGEMA_reg_buffer_2551 ( .C (clk), .D (new_AGEMA_signal_4506), .Q (new_AGEMA_signal_4507) ) ;
    buf_clk new_AGEMA_reg_buffer_2555 ( .C (clk), .D (new_AGEMA_signal_4510), .Q (new_AGEMA_signal_4511) ) ;
    buf_clk new_AGEMA_reg_buffer_2559 ( .C (clk), .D (new_AGEMA_signal_4514), .Q (new_AGEMA_signal_4515) ) ;
    buf_clk new_AGEMA_reg_buffer_2563 ( .C (clk), .D (new_AGEMA_signal_4518), .Q (new_AGEMA_signal_4519) ) ;
    buf_clk new_AGEMA_reg_buffer_2567 ( .C (clk), .D (new_AGEMA_signal_4522), .Q (new_AGEMA_signal_4523) ) ;
    buf_clk new_AGEMA_reg_buffer_2571 ( .C (clk), .D (new_AGEMA_signal_4526), .Q (new_AGEMA_signal_4527) ) ;
    buf_clk new_AGEMA_reg_buffer_2575 ( .C (clk), .D (new_AGEMA_signal_4530), .Q (new_AGEMA_signal_4531) ) ;
    buf_clk new_AGEMA_reg_buffer_2579 ( .C (clk), .D (new_AGEMA_signal_4534), .Q (new_AGEMA_signal_4535) ) ;
    buf_clk new_AGEMA_reg_buffer_2583 ( .C (clk), .D (new_AGEMA_signal_4538), .Q (new_AGEMA_signal_4539) ) ;
    buf_clk new_AGEMA_reg_buffer_2587 ( .C (clk), .D (new_AGEMA_signal_4542), .Q (new_AGEMA_signal_4543) ) ;
    buf_clk new_AGEMA_reg_buffer_2591 ( .C (clk), .D (new_AGEMA_signal_4546), .Q (new_AGEMA_signal_4547) ) ;
    buf_clk new_AGEMA_reg_buffer_2595 ( .C (clk), .D (new_AGEMA_signal_4550), .Q (new_AGEMA_signal_4551) ) ;
    buf_clk new_AGEMA_reg_buffer_2599 ( .C (clk), .D (new_AGEMA_signal_4554), .Q (new_AGEMA_signal_4555) ) ;
    buf_clk new_AGEMA_reg_buffer_2603 ( .C (clk), .D (new_AGEMA_signal_4558), .Q (new_AGEMA_signal_4559) ) ;
    buf_clk new_AGEMA_reg_buffer_2607 ( .C (clk), .D (new_AGEMA_signal_4562), .Q (new_AGEMA_signal_4563) ) ;
    buf_clk new_AGEMA_reg_buffer_2611 ( .C (clk), .D (new_AGEMA_signal_4566), .Q (new_AGEMA_signal_4567) ) ;
    buf_clk new_AGEMA_reg_buffer_2615 ( .C (clk), .D (new_AGEMA_signal_4570), .Q (new_AGEMA_signal_4571) ) ;
    buf_clk new_AGEMA_reg_buffer_2619 ( .C (clk), .D (new_AGEMA_signal_4574), .Q (new_AGEMA_signal_4575) ) ;
    buf_clk new_AGEMA_reg_buffer_2623 ( .C (clk), .D (new_AGEMA_signal_4578), .Q (new_AGEMA_signal_4579) ) ;
    buf_clk new_AGEMA_reg_buffer_2627 ( .C (clk), .D (new_AGEMA_signal_4582), .Q (new_AGEMA_signal_4583) ) ;
    buf_clk new_AGEMA_reg_buffer_2631 ( .C (clk), .D (new_AGEMA_signal_4586), .Q (new_AGEMA_signal_4587) ) ;
    buf_clk new_AGEMA_reg_buffer_2635 ( .C (clk), .D (new_AGEMA_signal_4590), .Q (new_AGEMA_signal_4591) ) ;
    buf_clk new_AGEMA_reg_buffer_2639 ( .C (clk), .D (new_AGEMA_signal_4594), .Q (new_AGEMA_signal_4595) ) ;
    buf_clk new_AGEMA_reg_buffer_2643 ( .C (clk), .D (new_AGEMA_signal_4598), .Q (new_AGEMA_signal_4599) ) ;
    buf_clk new_AGEMA_reg_buffer_2647 ( .C (clk), .D (new_AGEMA_signal_4602), .Q (new_AGEMA_signal_4603) ) ;
    buf_clk new_AGEMA_reg_buffer_2651 ( .C (clk), .D (new_AGEMA_signal_4606), .Q (new_AGEMA_signal_4607) ) ;
    buf_clk new_AGEMA_reg_buffer_2655 ( .C (clk), .D (new_AGEMA_signal_4610), .Q (new_AGEMA_signal_4611) ) ;
    buf_clk new_AGEMA_reg_buffer_2659 ( .C (clk), .D (new_AGEMA_signal_4614), .Q (new_AGEMA_signal_4615) ) ;
    buf_clk new_AGEMA_reg_buffer_2663 ( .C (clk), .D (new_AGEMA_signal_4618), .Q (new_AGEMA_signal_4619) ) ;
    buf_clk new_AGEMA_reg_buffer_2667 ( .C (clk), .D (new_AGEMA_signal_4622), .Q (new_AGEMA_signal_4623) ) ;
    buf_clk new_AGEMA_reg_buffer_2671 ( .C (clk), .D (new_AGEMA_signal_4626), .Q (new_AGEMA_signal_4627) ) ;
    buf_clk new_AGEMA_reg_buffer_2675 ( .C (clk), .D (new_AGEMA_signal_4630), .Q (new_AGEMA_signal_4631) ) ;
    buf_clk new_AGEMA_reg_buffer_2679 ( .C (clk), .D (new_AGEMA_signal_4634), .Q (new_AGEMA_signal_4635) ) ;
    buf_clk new_AGEMA_reg_buffer_2683 ( .C (clk), .D (new_AGEMA_signal_4638), .Q (new_AGEMA_signal_4639) ) ;
    buf_clk new_AGEMA_reg_buffer_2687 ( .C (clk), .D (new_AGEMA_signal_4642), .Q (new_AGEMA_signal_4643) ) ;
    buf_clk new_AGEMA_reg_buffer_2691 ( .C (clk), .D (new_AGEMA_signal_4646), .Q (new_AGEMA_signal_4647) ) ;
    buf_clk new_AGEMA_reg_buffer_2695 ( .C (clk), .D (new_AGEMA_signal_4650), .Q (new_AGEMA_signal_4651) ) ;
    buf_clk new_AGEMA_reg_buffer_2699 ( .C (clk), .D (new_AGEMA_signal_4654), .Q (new_AGEMA_signal_4655) ) ;
    buf_clk new_AGEMA_reg_buffer_2703 ( .C (clk), .D (new_AGEMA_signal_4658), .Q (new_AGEMA_signal_4659) ) ;
    buf_clk new_AGEMA_reg_buffer_2707 ( .C (clk), .D (new_AGEMA_signal_4662), .Q (new_AGEMA_signal_4663) ) ;
    buf_clk new_AGEMA_reg_buffer_2711 ( .C (clk), .D (new_AGEMA_signal_4666), .Q (new_AGEMA_signal_4667) ) ;
    buf_clk new_AGEMA_reg_buffer_2715 ( .C (clk), .D (new_AGEMA_signal_4670), .Q (new_AGEMA_signal_4671) ) ;
    buf_clk new_AGEMA_reg_buffer_2719 ( .C (clk), .D (new_AGEMA_signal_4674), .Q (new_AGEMA_signal_4675) ) ;
    buf_clk new_AGEMA_reg_buffer_2723 ( .C (clk), .D (new_AGEMA_signal_4678), .Q (new_AGEMA_signal_4679) ) ;
    buf_clk new_AGEMA_reg_buffer_2727 ( .C (clk), .D (new_AGEMA_signal_4682), .Q (new_AGEMA_signal_4683) ) ;
    buf_clk new_AGEMA_reg_buffer_2731 ( .C (clk), .D (new_AGEMA_signal_4686), .Q (new_AGEMA_signal_4687) ) ;
    buf_clk new_AGEMA_reg_buffer_2735 ( .C (clk), .D (new_AGEMA_signal_4690), .Q (new_AGEMA_signal_4691) ) ;
    buf_clk new_AGEMA_reg_buffer_2739 ( .C (clk), .D (new_AGEMA_signal_4694), .Q (new_AGEMA_signal_4695) ) ;
    buf_clk new_AGEMA_reg_buffer_2743 ( .C (clk), .D (new_AGEMA_signal_4698), .Q (new_AGEMA_signal_4699) ) ;
    buf_clk new_AGEMA_reg_buffer_2747 ( .C (clk), .D (new_AGEMA_signal_4702), .Q (new_AGEMA_signal_4703) ) ;
    buf_clk new_AGEMA_reg_buffer_2751 ( .C (clk), .D (new_AGEMA_signal_4706), .Q (new_AGEMA_signal_4707) ) ;
    buf_clk new_AGEMA_reg_buffer_2755 ( .C (clk), .D (new_AGEMA_signal_4710), .Q (new_AGEMA_signal_4711) ) ;
    buf_clk new_AGEMA_reg_buffer_2759 ( .C (clk), .D (new_AGEMA_signal_4714), .Q (new_AGEMA_signal_4715) ) ;
    buf_clk new_AGEMA_reg_buffer_2763 ( .C (clk), .D (new_AGEMA_signal_4718), .Q (new_AGEMA_signal_4719) ) ;
    buf_clk new_AGEMA_reg_buffer_2767 ( .C (clk), .D (new_AGEMA_signal_4722), .Q (new_AGEMA_signal_4723) ) ;
    buf_clk new_AGEMA_reg_buffer_2771 ( .C (clk), .D (new_AGEMA_signal_4726), .Q (new_AGEMA_signal_4727) ) ;
    buf_clk new_AGEMA_reg_buffer_2775 ( .C (clk), .D (new_AGEMA_signal_4730), .Q (new_AGEMA_signal_4731) ) ;
    buf_clk new_AGEMA_reg_buffer_2779 ( .C (clk), .D (new_AGEMA_signal_4734), .Q (new_AGEMA_signal_4735) ) ;
    buf_clk new_AGEMA_reg_buffer_2783 ( .C (clk), .D (new_AGEMA_signal_4738), .Q (new_AGEMA_signal_4739) ) ;
    buf_clk new_AGEMA_reg_buffer_2787 ( .C (clk), .D (new_AGEMA_signal_4742), .Q (new_AGEMA_signal_4743) ) ;
    buf_clk new_AGEMA_reg_buffer_2791 ( .C (clk), .D (new_AGEMA_signal_4746), .Q (new_AGEMA_signal_4747) ) ;
    buf_clk new_AGEMA_reg_buffer_2795 ( .C (clk), .D (new_AGEMA_signal_4750), .Q (new_AGEMA_signal_4751) ) ;
    buf_clk new_AGEMA_reg_buffer_2799 ( .C (clk), .D (new_AGEMA_signal_4754), .Q (new_AGEMA_signal_4755) ) ;
    buf_clk new_AGEMA_reg_buffer_2803 ( .C (clk), .D (new_AGEMA_signal_4758), .Q (new_AGEMA_signal_4759) ) ;
    buf_clk new_AGEMA_reg_buffer_2807 ( .C (clk), .D (new_AGEMA_signal_4762), .Q (new_AGEMA_signal_4763) ) ;
    buf_clk new_AGEMA_reg_buffer_2811 ( .C (clk), .D (new_AGEMA_signal_4766), .Q (new_AGEMA_signal_4767) ) ;
    buf_clk new_AGEMA_reg_buffer_2815 ( .C (clk), .D (new_AGEMA_signal_4770), .Q (new_AGEMA_signal_4771) ) ;
    buf_clk new_AGEMA_reg_buffer_2819 ( .C (clk), .D (new_AGEMA_signal_4774), .Q (new_AGEMA_signal_4775) ) ;
    buf_clk new_AGEMA_reg_buffer_2823 ( .C (clk), .D (new_AGEMA_signal_4778), .Q (new_AGEMA_signal_4779) ) ;
    buf_clk new_AGEMA_reg_buffer_2827 ( .C (clk), .D (new_AGEMA_signal_4782), .Q (new_AGEMA_signal_4783) ) ;
    buf_clk new_AGEMA_reg_buffer_2831 ( .C (clk), .D (new_AGEMA_signal_4786), .Q (new_AGEMA_signal_4787) ) ;
    buf_clk new_AGEMA_reg_buffer_2835 ( .C (clk), .D (new_AGEMA_signal_4790), .Q (new_AGEMA_signal_4791) ) ;
    buf_clk new_AGEMA_reg_buffer_2839 ( .C (clk), .D (new_AGEMA_signal_4794), .Q (new_AGEMA_signal_4795) ) ;
    buf_clk new_AGEMA_reg_buffer_2843 ( .C (clk), .D (new_AGEMA_signal_4798), .Q (new_AGEMA_signal_4799) ) ;
    buf_clk new_AGEMA_reg_buffer_2847 ( .C (clk), .D (new_AGEMA_signal_4802), .Q (new_AGEMA_signal_4803) ) ;
    buf_clk new_AGEMA_reg_buffer_2851 ( .C (clk), .D (new_AGEMA_signal_4806), .Q (new_AGEMA_signal_4807) ) ;
    buf_clk new_AGEMA_reg_buffer_2855 ( .C (clk), .D (new_AGEMA_signal_4810), .Q (new_AGEMA_signal_4811) ) ;
    buf_clk new_AGEMA_reg_buffer_2859 ( .C (clk), .D (new_AGEMA_signal_4814), .Q (new_AGEMA_signal_4815) ) ;
    buf_clk new_AGEMA_reg_buffer_2863 ( .C (clk), .D (new_AGEMA_signal_4818), .Q (new_AGEMA_signal_4819) ) ;
    buf_clk new_AGEMA_reg_buffer_2867 ( .C (clk), .D (new_AGEMA_signal_4822), .Q (new_AGEMA_signal_4823) ) ;
    buf_clk new_AGEMA_reg_buffer_2871 ( .C (clk), .D (new_AGEMA_signal_4826), .Q (new_AGEMA_signal_4827) ) ;
    buf_clk new_AGEMA_reg_buffer_2875 ( .C (clk), .D (new_AGEMA_signal_4830), .Q (new_AGEMA_signal_4831) ) ;
    buf_clk new_AGEMA_reg_buffer_2879 ( .C (clk), .D (new_AGEMA_signal_4834), .Q (new_AGEMA_signal_4835) ) ;
    buf_clk new_AGEMA_reg_buffer_2883 ( .C (clk), .D (new_AGEMA_signal_4838), .Q (new_AGEMA_signal_4839) ) ;
    buf_clk new_AGEMA_reg_buffer_2887 ( .C (clk), .D (new_AGEMA_signal_4842), .Q (new_AGEMA_signal_4843) ) ;
    buf_clk new_AGEMA_reg_buffer_2891 ( .C (clk), .D (new_AGEMA_signal_4846), .Q (new_AGEMA_signal_4847) ) ;
    buf_clk new_AGEMA_reg_buffer_2895 ( .C (clk), .D (new_AGEMA_signal_4850), .Q (new_AGEMA_signal_4851) ) ;
    buf_clk new_AGEMA_reg_buffer_2899 ( .C (clk), .D (new_AGEMA_signal_4854), .Q (new_AGEMA_signal_4855) ) ;
    buf_clk new_AGEMA_reg_buffer_2903 ( .C (clk), .D (new_AGEMA_signal_4858), .Q (new_AGEMA_signal_4859) ) ;
    buf_clk new_AGEMA_reg_buffer_2907 ( .C (clk), .D (new_AGEMA_signal_4862), .Q (new_AGEMA_signal_4863) ) ;
    buf_clk new_AGEMA_reg_buffer_2911 ( .C (clk), .D (new_AGEMA_signal_4866), .Q (new_AGEMA_signal_4867) ) ;
    buf_clk new_AGEMA_reg_buffer_2915 ( .C (clk), .D (new_AGEMA_signal_4870), .Q (new_AGEMA_signal_4871) ) ;
    buf_clk new_AGEMA_reg_buffer_2919 ( .C (clk), .D (new_AGEMA_signal_4874), .Q (new_AGEMA_signal_4875) ) ;
    buf_clk new_AGEMA_reg_buffer_2923 ( .C (clk), .D (new_AGEMA_signal_4878), .Q (new_AGEMA_signal_4879) ) ;
    buf_clk new_AGEMA_reg_buffer_2927 ( .C (clk), .D (new_AGEMA_signal_4882), .Q (new_AGEMA_signal_4883) ) ;
    buf_clk new_AGEMA_reg_buffer_2931 ( .C (clk), .D (new_AGEMA_signal_4886), .Q (new_AGEMA_signal_4887) ) ;
    buf_clk new_AGEMA_reg_buffer_2935 ( .C (clk), .D (new_AGEMA_signal_4890), .Q (new_AGEMA_signal_4891) ) ;
    buf_clk new_AGEMA_reg_buffer_2939 ( .C (clk), .D (new_AGEMA_signal_4894), .Q (new_AGEMA_signal_4895) ) ;
    buf_clk new_AGEMA_reg_buffer_2943 ( .C (clk), .D (new_AGEMA_signal_4898), .Q (new_AGEMA_signal_4899) ) ;
    buf_clk new_AGEMA_reg_buffer_2947 ( .C (clk), .D (new_AGEMA_signal_4902), .Q (new_AGEMA_signal_4903) ) ;
    buf_clk new_AGEMA_reg_buffer_2951 ( .C (clk), .D (new_AGEMA_signal_4906), .Q (new_AGEMA_signal_4907) ) ;
    buf_clk new_AGEMA_reg_buffer_2955 ( .C (clk), .D (new_AGEMA_signal_4910), .Q (new_AGEMA_signal_4911) ) ;
    buf_clk new_AGEMA_reg_buffer_2959 ( .C (clk), .D (new_AGEMA_signal_4914), .Q (new_AGEMA_signal_4915) ) ;
    buf_clk new_AGEMA_reg_buffer_2963 ( .C (clk), .D (new_AGEMA_signal_4918), .Q (new_AGEMA_signal_4919) ) ;
    buf_clk new_AGEMA_reg_buffer_2967 ( .C (clk), .D (new_AGEMA_signal_4922), .Q (new_AGEMA_signal_4923) ) ;
    buf_clk new_AGEMA_reg_buffer_2971 ( .C (clk), .D (new_AGEMA_signal_4926), .Q (new_AGEMA_signal_4927) ) ;
    buf_clk new_AGEMA_reg_buffer_2975 ( .C (clk), .D (new_AGEMA_signal_4930), .Q (new_AGEMA_signal_4931) ) ;
    buf_clk new_AGEMA_reg_buffer_2979 ( .C (clk), .D (new_AGEMA_signal_4934), .Q (new_AGEMA_signal_4935) ) ;
    buf_clk new_AGEMA_reg_buffer_2983 ( .C (clk), .D (new_AGEMA_signal_4938), .Q (new_AGEMA_signal_4939) ) ;
    buf_clk new_AGEMA_reg_buffer_2987 ( .C (clk), .D (new_AGEMA_signal_4942), .Q (new_AGEMA_signal_4943) ) ;
    buf_clk new_AGEMA_reg_buffer_2991 ( .C (clk), .D (new_AGEMA_signal_4946), .Q (new_AGEMA_signal_4947) ) ;
    buf_clk new_AGEMA_reg_buffer_2995 ( .C (clk), .D (new_AGEMA_signal_4950), .Q (new_AGEMA_signal_4951) ) ;
    buf_clk new_AGEMA_reg_buffer_2999 ( .C (clk), .D (new_AGEMA_signal_4954), .Q (new_AGEMA_signal_4955) ) ;
    buf_clk new_AGEMA_reg_buffer_3003 ( .C (clk), .D (new_AGEMA_signal_4958), .Q (new_AGEMA_signal_4959) ) ;
    buf_clk new_AGEMA_reg_buffer_3007 ( .C (clk), .D (new_AGEMA_signal_4962), .Q (new_AGEMA_signal_4963) ) ;
    buf_clk new_AGEMA_reg_buffer_3011 ( .C (clk), .D (new_AGEMA_signal_4966), .Q (new_AGEMA_signal_4967) ) ;
    buf_clk new_AGEMA_reg_buffer_3015 ( .C (clk), .D (new_AGEMA_signal_4970), .Q (new_AGEMA_signal_4971) ) ;
    buf_clk new_AGEMA_reg_buffer_3019 ( .C (clk), .D (new_AGEMA_signal_4974), .Q (new_AGEMA_signal_4975) ) ;
    buf_clk new_AGEMA_reg_buffer_3023 ( .C (clk), .D (new_AGEMA_signal_4978), .Q (new_AGEMA_signal_4979) ) ;
    buf_clk new_AGEMA_reg_buffer_3027 ( .C (clk), .D (new_AGEMA_signal_4982), .Q (new_AGEMA_signal_4983) ) ;
    buf_clk new_AGEMA_reg_buffer_3031 ( .C (clk), .D (new_AGEMA_signal_4986), .Q (new_AGEMA_signal_4987) ) ;
    buf_clk new_AGEMA_reg_buffer_3035 ( .C (clk), .D (new_AGEMA_signal_4990), .Q (new_AGEMA_signal_4991) ) ;
    buf_clk new_AGEMA_reg_buffer_3039 ( .C (clk), .D (new_AGEMA_signal_4994), .Q (new_AGEMA_signal_4995) ) ;
    buf_clk new_AGEMA_reg_buffer_3043 ( .C (clk), .D (new_AGEMA_signal_4998), .Q (new_AGEMA_signal_4999) ) ;
    buf_clk new_AGEMA_reg_buffer_3047 ( .C (clk), .D (new_AGEMA_signal_5002), .Q (new_AGEMA_signal_5003) ) ;
    buf_clk new_AGEMA_reg_buffer_3051 ( .C (clk), .D (new_AGEMA_signal_5006), .Q (new_AGEMA_signal_5007) ) ;
    buf_clk new_AGEMA_reg_buffer_3055 ( .C (clk), .D (new_AGEMA_signal_5010), .Q (new_AGEMA_signal_5011) ) ;
    buf_clk new_AGEMA_reg_buffer_3059 ( .C (clk), .D (new_AGEMA_signal_5014), .Q (new_AGEMA_signal_5015) ) ;
    buf_clk new_AGEMA_reg_buffer_3063 ( .C (clk), .D (new_AGEMA_signal_5018), .Q (new_AGEMA_signal_5019) ) ;
    buf_clk new_AGEMA_reg_buffer_3067 ( .C (clk), .D (new_AGEMA_signal_5022), .Q (new_AGEMA_signal_5023) ) ;
    buf_clk new_AGEMA_reg_buffer_3071 ( .C (clk), .D (new_AGEMA_signal_5026), .Q (new_AGEMA_signal_5027) ) ;
    buf_clk new_AGEMA_reg_buffer_3075 ( .C (clk), .D (new_AGEMA_signal_5030), .Q (new_AGEMA_signal_5031) ) ;
    buf_clk new_AGEMA_reg_buffer_3079 ( .C (clk), .D (new_AGEMA_signal_5034), .Q (new_AGEMA_signal_5035) ) ;
    buf_clk new_AGEMA_reg_buffer_3083 ( .C (clk), .D (new_AGEMA_signal_5038), .Q (new_AGEMA_signal_5039) ) ;
    buf_clk new_AGEMA_reg_buffer_3087 ( .C (clk), .D (new_AGEMA_signal_5042), .Q (new_AGEMA_signal_5043) ) ;
    buf_clk new_AGEMA_reg_buffer_3091 ( .C (clk), .D (new_AGEMA_signal_5046), .Q (new_AGEMA_signal_5047) ) ;
    buf_clk new_AGEMA_reg_buffer_3095 ( .C (clk), .D (new_AGEMA_signal_5050), .Q (new_AGEMA_signal_5051) ) ;
    buf_clk new_AGEMA_reg_buffer_3099 ( .C (clk), .D (new_AGEMA_signal_5054), .Q (new_AGEMA_signal_5055) ) ;
    buf_clk new_AGEMA_reg_buffer_3103 ( .C (clk), .D (new_AGEMA_signal_5058), .Q (new_AGEMA_signal_5059) ) ;
    buf_clk new_AGEMA_reg_buffer_3107 ( .C (clk), .D (new_AGEMA_signal_5062), .Q (new_AGEMA_signal_5063) ) ;
    buf_clk new_AGEMA_reg_buffer_3111 ( .C (clk), .D (new_AGEMA_signal_5066), .Q (new_AGEMA_signal_5067) ) ;
    buf_clk new_AGEMA_reg_buffer_3115 ( .C (clk), .D (new_AGEMA_signal_5070), .Q (new_AGEMA_signal_5071) ) ;
    buf_clk new_AGEMA_reg_buffer_3119 ( .C (clk), .D (new_AGEMA_signal_5074), .Q (new_AGEMA_signal_5075) ) ;
    buf_clk new_AGEMA_reg_buffer_3123 ( .C (clk), .D (new_AGEMA_signal_5078), .Q (new_AGEMA_signal_5079) ) ;
    buf_clk new_AGEMA_reg_buffer_3127 ( .C (clk), .D (new_AGEMA_signal_5082), .Q (new_AGEMA_signal_5083) ) ;
    buf_clk new_AGEMA_reg_buffer_3131 ( .C (clk), .D (new_AGEMA_signal_5086), .Q (new_AGEMA_signal_5087) ) ;
    buf_clk new_AGEMA_reg_buffer_3135 ( .C (clk), .D (new_AGEMA_signal_5090), .Q (new_AGEMA_signal_5091) ) ;
    buf_clk new_AGEMA_reg_buffer_3139 ( .C (clk), .D (new_AGEMA_signal_5094), .Q (new_AGEMA_signal_5095) ) ;
    buf_clk new_AGEMA_reg_buffer_3143 ( .C (clk), .D (new_AGEMA_signal_5098), .Q (new_AGEMA_signal_5099) ) ;
    buf_clk new_AGEMA_reg_buffer_3147 ( .C (clk), .D (new_AGEMA_signal_5102), .Q (new_AGEMA_signal_5103) ) ;
    buf_clk new_AGEMA_reg_buffer_3151 ( .C (clk), .D (new_AGEMA_signal_5106), .Q (new_AGEMA_signal_5107) ) ;
    buf_clk new_AGEMA_reg_buffer_3155 ( .C (clk), .D (new_AGEMA_signal_5110), .Q (new_AGEMA_signal_5111) ) ;
    buf_clk new_AGEMA_reg_buffer_3159 ( .C (clk), .D (new_AGEMA_signal_5114), .Q (new_AGEMA_signal_5115) ) ;
    buf_clk new_AGEMA_reg_buffer_3163 ( .C (clk), .D (new_AGEMA_signal_5118), .Q (new_AGEMA_signal_5119) ) ;
    buf_clk new_AGEMA_reg_buffer_3167 ( .C (clk), .D (new_AGEMA_signal_5122), .Q (new_AGEMA_signal_5123) ) ;
    buf_clk new_AGEMA_reg_buffer_3171 ( .C (clk), .D (new_AGEMA_signal_5126), .Q (new_AGEMA_signal_5127) ) ;
    buf_clk new_AGEMA_reg_buffer_3175 ( .C (clk), .D (new_AGEMA_signal_5130), .Q (new_AGEMA_signal_5131) ) ;
    buf_clk new_AGEMA_reg_buffer_3179 ( .C (clk), .D (new_AGEMA_signal_5134), .Q (new_AGEMA_signal_5135) ) ;
    buf_clk new_AGEMA_reg_buffer_3183 ( .C (clk), .D (new_AGEMA_signal_5138), .Q (new_AGEMA_signal_5139) ) ;
    buf_clk new_AGEMA_reg_buffer_3187 ( .C (clk), .D (new_AGEMA_signal_5142), .Q (new_AGEMA_signal_5143) ) ;
    buf_clk new_AGEMA_reg_buffer_3191 ( .C (clk), .D (new_AGEMA_signal_5146), .Q (new_AGEMA_signal_5147) ) ;
    buf_clk new_AGEMA_reg_buffer_3195 ( .C (clk), .D (new_AGEMA_signal_5150), .Q (new_AGEMA_signal_5151) ) ;
    buf_clk new_AGEMA_reg_buffer_3199 ( .C (clk), .D (new_AGEMA_signal_5154), .Q (new_AGEMA_signal_5155) ) ;
    buf_clk new_AGEMA_reg_buffer_3203 ( .C (clk), .D (new_AGEMA_signal_5158), .Q (new_AGEMA_signal_5159) ) ;
    buf_clk new_AGEMA_reg_buffer_3207 ( .C (clk), .D (new_AGEMA_signal_5162), .Q (new_AGEMA_signal_5163) ) ;
    buf_clk new_AGEMA_reg_buffer_3211 ( .C (clk), .D (new_AGEMA_signal_5166), .Q (new_AGEMA_signal_5167) ) ;
    buf_clk new_AGEMA_reg_buffer_3215 ( .C (clk), .D (new_AGEMA_signal_5170), .Q (new_AGEMA_signal_5171) ) ;
    buf_clk new_AGEMA_reg_buffer_3219 ( .C (clk), .D (new_AGEMA_signal_5174), .Q (new_AGEMA_signal_5175) ) ;
    buf_clk new_AGEMA_reg_buffer_3223 ( .C (clk), .D (new_AGEMA_signal_5178), .Q (new_AGEMA_signal_5179) ) ;
    buf_clk new_AGEMA_reg_buffer_3227 ( .C (clk), .D (new_AGEMA_signal_5182), .Q (new_AGEMA_signal_5183) ) ;
    buf_clk new_AGEMA_reg_buffer_3231 ( .C (clk), .D (new_AGEMA_signal_5186), .Q (new_AGEMA_signal_5187) ) ;
    buf_clk new_AGEMA_reg_buffer_3235 ( .C (clk), .D (new_AGEMA_signal_5190), .Q (new_AGEMA_signal_5191) ) ;
    buf_clk new_AGEMA_reg_buffer_3239 ( .C (clk), .D (new_AGEMA_signal_5194), .Q (new_AGEMA_signal_5195) ) ;
    buf_clk new_AGEMA_reg_buffer_3243 ( .C (clk), .D (new_AGEMA_signal_5198), .Q (new_AGEMA_signal_5199) ) ;
    buf_clk new_AGEMA_reg_buffer_3247 ( .C (clk), .D (new_AGEMA_signal_5202), .Q (new_AGEMA_signal_5203) ) ;
    buf_clk new_AGEMA_reg_buffer_3251 ( .C (clk), .D (new_AGEMA_signal_5206), .Q (new_AGEMA_signal_5207) ) ;
    buf_clk new_AGEMA_reg_buffer_3255 ( .C (clk), .D (new_AGEMA_signal_5210), .Q (new_AGEMA_signal_5211) ) ;
    buf_clk new_AGEMA_reg_buffer_3259 ( .C (clk), .D (new_AGEMA_signal_5214), .Q (new_AGEMA_signal_5215) ) ;
    buf_clk new_AGEMA_reg_buffer_3263 ( .C (clk), .D (new_AGEMA_signal_5218), .Q (new_AGEMA_signal_5219) ) ;
    buf_clk new_AGEMA_reg_buffer_3267 ( .C (clk), .D (new_AGEMA_signal_5222), .Q (new_AGEMA_signal_5223) ) ;
    buf_clk new_AGEMA_reg_buffer_3271 ( .C (clk), .D (new_AGEMA_signal_5226), .Q (new_AGEMA_signal_5227) ) ;
    buf_clk new_AGEMA_reg_buffer_3275 ( .C (clk), .D (new_AGEMA_signal_5230), .Q (new_AGEMA_signal_5231) ) ;
    buf_clk new_AGEMA_reg_buffer_3279 ( .C (clk), .D (new_AGEMA_signal_5234), .Q (new_AGEMA_signal_5235) ) ;
    buf_clk new_AGEMA_reg_buffer_3283 ( .C (clk), .D (new_AGEMA_signal_5238), .Q (new_AGEMA_signal_5239) ) ;
    buf_clk new_AGEMA_reg_buffer_3287 ( .C (clk), .D (new_AGEMA_signal_5242), .Q (new_AGEMA_signal_5243) ) ;
    buf_clk new_AGEMA_reg_buffer_3291 ( .C (clk), .D (new_AGEMA_signal_5246), .Q (new_AGEMA_signal_5247) ) ;
    buf_clk new_AGEMA_reg_buffer_3295 ( .C (clk), .D (new_AGEMA_signal_5250), .Q (new_AGEMA_signal_5251) ) ;
    buf_clk new_AGEMA_reg_buffer_3299 ( .C (clk), .D (new_AGEMA_signal_5254), .Q (new_AGEMA_signal_5255) ) ;
    buf_clk new_AGEMA_reg_buffer_3303 ( .C (clk), .D (new_AGEMA_signal_5258), .Q (new_AGEMA_signal_5259) ) ;
    buf_clk new_AGEMA_reg_buffer_3307 ( .C (clk), .D (new_AGEMA_signal_5262), .Q (new_AGEMA_signal_5263) ) ;
    buf_clk new_AGEMA_reg_buffer_3311 ( .C (clk), .D (new_AGEMA_signal_5266), .Q (new_AGEMA_signal_5267) ) ;
    buf_clk new_AGEMA_reg_buffer_3315 ( .C (clk), .D (new_AGEMA_signal_5270), .Q (new_AGEMA_signal_5271) ) ;
    buf_clk new_AGEMA_reg_buffer_3319 ( .C (clk), .D (new_AGEMA_signal_5274), .Q (new_AGEMA_signal_5275) ) ;
    buf_clk new_AGEMA_reg_buffer_3323 ( .C (clk), .D (new_AGEMA_signal_5278), .Q (new_AGEMA_signal_5279) ) ;
    buf_clk new_AGEMA_reg_buffer_3327 ( .C (clk), .D (new_AGEMA_signal_5282), .Q (new_AGEMA_signal_5283) ) ;
    buf_clk new_AGEMA_reg_buffer_3331 ( .C (clk), .D (new_AGEMA_signal_5286), .Q (new_AGEMA_signal_5287) ) ;
    buf_clk new_AGEMA_reg_buffer_3335 ( .C (clk), .D (new_AGEMA_signal_5290), .Q (new_AGEMA_signal_5291) ) ;
    buf_clk new_AGEMA_reg_buffer_3339 ( .C (clk), .D (new_AGEMA_signal_5294), .Q (new_AGEMA_signal_5295) ) ;
    buf_clk new_AGEMA_reg_buffer_3343 ( .C (clk), .D (new_AGEMA_signal_5298), .Q (new_AGEMA_signal_5299) ) ;
    buf_clk new_AGEMA_reg_buffer_3347 ( .C (clk), .D (new_AGEMA_signal_5302), .Q (new_AGEMA_signal_5303) ) ;
    buf_clk new_AGEMA_reg_buffer_3351 ( .C (clk), .D (new_AGEMA_signal_5306), .Q (new_AGEMA_signal_5307) ) ;
    buf_clk new_AGEMA_reg_buffer_3355 ( .C (clk), .D (new_AGEMA_signal_5310), .Q (new_AGEMA_signal_5311) ) ;
    buf_clk new_AGEMA_reg_buffer_3359 ( .C (clk), .D (new_AGEMA_signal_5314), .Q (new_AGEMA_signal_5315) ) ;
    buf_clk new_AGEMA_reg_buffer_3363 ( .C (clk), .D (new_AGEMA_signal_5318), .Q (new_AGEMA_signal_5319) ) ;
    buf_clk new_AGEMA_reg_buffer_3367 ( .C (clk), .D (new_AGEMA_signal_5322), .Q (new_AGEMA_signal_5323) ) ;
    buf_clk new_AGEMA_reg_buffer_3371 ( .C (clk), .D (new_AGEMA_signal_5326), .Q (new_AGEMA_signal_5327) ) ;
    buf_clk new_AGEMA_reg_buffer_3375 ( .C (clk), .D (new_AGEMA_signal_5330), .Q (new_AGEMA_signal_5331) ) ;
    buf_clk new_AGEMA_reg_buffer_3379 ( .C (clk), .D (new_AGEMA_signal_5334), .Q (new_AGEMA_signal_5335) ) ;
    buf_clk new_AGEMA_reg_buffer_3383 ( .C (clk), .D (new_AGEMA_signal_5338), .Q (new_AGEMA_signal_5339) ) ;
    buf_clk new_AGEMA_reg_buffer_3387 ( .C (clk), .D (new_AGEMA_signal_5342), .Q (new_AGEMA_signal_5343) ) ;
    buf_clk new_AGEMA_reg_buffer_3391 ( .C (clk), .D (new_AGEMA_signal_5346), .Q (new_AGEMA_signal_5347) ) ;
    buf_clk new_AGEMA_reg_buffer_3395 ( .C (clk), .D (new_AGEMA_signal_5350), .Q (new_AGEMA_signal_5351) ) ;
    buf_clk new_AGEMA_reg_buffer_3399 ( .C (clk), .D (new_AGEMA_signal_5354), .Q (new_AGEMA_signal_5355) ) ;
    buf_clk new_AGEMA_reg_buffer_3403 ( .C (clk), .D (new_AGEMA_signal_5358), .Q (new_AGEMA_signal_5359) ) ;
    buf_clk new_AGEMA_reg_buffer_3407 ( .C (clk), .D (new_AGEMA_signal_5362), .Q (new_AGEMA_signal_5363) ) ;
    buf_clk new_AGEMA_reg_buffer_3411 ( .C (clk), .D (new_AGEMA_signal_5366), .Q (new_AGEMA_signal_5367) ) ;
    buf_clk new_AGEMA_reg_buffer_3415 ( .C (clk), .D (new_AGEMA_signal_5370), .Q (new_AGEMA_signal_5371) ) ;
    buf_clk new_AGEMA_reg_buffer_3419 ( .C (clk), .D (new_AGEMA_signal_5374), .Q (new_AGEMA_signal_5375) ) ;
    buf_clk new_AGEMA_reg_buffer_3423 ( .C (clk), .D (new_AGEMA_signal_5378), .Q (new_AGEMA_signal_5379) ) ;
    buf_clk new_AGEMA_reg_buffer_3427 ( .C (clk), .D (new_AGEMA_signal_5382), .Q (new_AGEMA_signal_5383) ) ;
    buf_clk new_AGEMA_reg_buffer_3431 ( .C (clk), .D (new_AGEMA_signal_5386), .Q (new_AGEMA_signal_5387) ) ;
    buf_clk new_AGEMA_reg_buffer_3435 ( .C (clk), .D (new_AGEMA_signal_5390), .Q (new_AGEMA_signal_5391) ) ;
    buf_clk new_AGEMA_reg_buffer_3439 ( .C (clk), .D (new_AGEMA_signal_5394), .Q (new_AGEMA_signal_5395) ) ;
    buf_clk new_AGEMA_reg_buffer_3443 ( .C (clk), .D (new_AGEMA_signal_5398), .Q (new_AGEMA_signal_5399) ) ;
    buf_clk new_AGEMA_reg_buffer_3447 ( .C (clk), .D (new_AGEMA_signal_5402), .Q (new_AGEMA_signal_5403) ) ;
    buf_clk new_AGEMA_reg_buffer_3451 ( .C (clk), .D (new_AGEMA_signal_5406), .Q (new_AGEMA_signal_5407) ) ;
    buf_clk new_AGEMA_reg_buffer_3455 ( .C (clk), .D (new_AGEMA_signal_5410), .Q (new_AGEMA_signal_5411) ) ;
    buf_clk new_AGEMA_reg_buffer_3459 ( .C (clk), .D (new_AGEMA_signal_5414), .Q (new_AGEMA_signal_5415) ) ;
    buf_clk new_AGEMA_reg_buffer_3463 ( .C (clk), .D (new_AGEMA_signal_5418), .Q (new_AGEMA_signal_5419) ) ;
    buf_clk new_AGEMA_reg_buffer_3467 ( .C (clk), .D (new_AGEMA_signal_5422), .Q (new_AGEMA_signal_5423) ) ;
    buf_clk new_AGEMA_reg_buffer_3471 ( .C (clk), .D (new_AGEMA_signal_5426), .Q (new_AGEMA_signal_5427) ) ;
    buf_clk new_AGEMA_reg_buffer_3475 ( .C (clk), .D (new_AGEMA_signal_5430), .Q (new_AGEMA_signal_5431) ) ;
    buf_clk new_AGEMA_reg_buffer_3479 ( .C (clk), .D (new_AGEMA_signal_5434), .Q (new_AGEMA_signal_5435) ) ;
    buf_clk new_AGEMA_reg_buffer_3483 ( .C (clk), .D (new_AGEMA_signal_5438), .Q (new_AGEMA_signal_5439) ) ;
    buf_clk new_AGEMA_reg_buffer_3487 ( .C (clk), .D (new_AGEMA_signal_5442), .Q (new_AGEMA_signal_5443) ) ;
    buf_clk new_AGEMA_reg_buffer_3491 ( .C (clk), .D (new_AGEMA_signal_5446), .Q (new_AGEMA_signal_5447) ) ;
    buf_clk new_AGEMA_reg_buffer_3495 ( .C (clk), .D (new_AGEMA_signal_5450), .Q (new_AGEMA_signal_5451) ) ;
    buf_clk new_AGEMA_reg_buffer_3499 ( .C (clk), .D (new_AGEMA_signal_5454), .Q (new_AGEMA_signal_5455) ) ;
    buf_clk new_AGEMA_reg_buffer_3503 ( .C (clk), .D (new_AGEMA_signal_5458), .Q (new_AGEMA_signal_5459) ) ;
    buf_clk new_AGEMA_reg_buffer_3507 ( .C (clk), .D (new_AGEMA_signal_5462), .Q (new_AGEMA_signal_5463) ) ;
    buf_clk new_AGEMA_reg_buffer_3511 ( .C (clk), .D (new_AGEMA_signal_5466), .Q (new_AGEMA_signal_5467) ) ;
    buf_clk new_AGEMA_reg_buffer_3515 ( .C (clk), .D (new_AGEMA_signal_5470), .Q (new_AGEMA_signal_5471) ) ;
    buf_clk new_AGEMA_reg_buffer_3519 ( .C (clk), .D (new_AGEMA_signal_5474), .Q (new_AGEMA_signal_5475) ) ;
    buf_clk new_AGEMA_reg_buffer_3523 ( .C (clk), .D (new_AGEMA_signal_5478), .Q (new_AGEMA_signal_5479) ) ;
    buf_clk new_AGEMA_reg_buffer_3527 ( .C (clk), .D (new_AGEMA_signal_5482), .Q (new_AGEMA_signal_5483) ) ;
    buf_clk new_AGEMA_reg_buffer_3531 ( .C (clk), .D (new_AGEMA_signal_5486), .Q (new_AGEMA_signal_5487) ) ;
    buf_clk new_AGEMA_reg_buffer_3535 ( .C (clk), .D (new_AGEMA_signal_5490), .Q (new_AGEMA_signal_5491) ) ;
    buf_clk new_AGEMA_reg_buffer_3539 ( .C (clk), .D (new_AGEMA_signal_5494), .Q (new_AGEMA_signal_5495) ) ;
    buf_clk new_AGEMA_reg_buffer_3543 ( .C (clk), .D (new_AGEMA_signal_5498), .Q (new_AGEMA_signal_5499) ) ;
    buf_clk new_AGEMA_reg_buffer_3547 ( .C (clk), .D (new_AGEMA_signal_5502), .Q (new_AGEMA_signal_5503) ) ;
    buf_clk new_AGEMA_reg_buffer_3551 ( .C (clk), .D (new_AGEMA_signal_5506), .Q (new_AGEMA_signal_5507) ) ;
    buf_clk new_AGEMA_reg_buffer_3555 ( .C (clk), .D (new_AGEMA_signal_5510), .Q (new_AGEMA_signal_5511) ) ;
    buf_clk new_AGEMA_reg_buffer_3559 ( .C (clk), .D (new_AGEMA_signal_5514), .Q (new_AGEMA_signal_5515) ) ;
    buf_clk new_AGEMA_reg_buffer_3563 ( .C (clk), .D (new_AGEMA_signal_5518), .Q (new_AGEMA_signal_5519) ) ;
    buf_clk new_AGEMA_reg_buffer_3567 ( .C (clk), .D (new_AGEMA_signal_5522), .Q (new_AGEMA_signal_5523) ) ;
    buf_clk new_AGEMA_reg_buffer_3571 ( .C (clk), .D (new_AGEMA_signal_5526), .Q (new_AGEMA_signal_5527) ) ;
    buf_clk new_AGEMA_reg_buffer_3575 ( .C (clk), .D (new_AGEMA_signal_5530), .Q (new_AGEMA_signal_5531) ) ;
    buf_clk new_AGEMA_reg_buffer_3579 ( .C (clk), .D (new_AGEMA_signal_5534), .Q (new_AGEMA_signal_5535) ) ;
    buf_clk new_AGEMA_reg_buffer_3583 ( .C (clk), .D (new_AGEMA_signal_5538), .Q (new_AGEMA_signal_5539) ) ;
    buf_clk new_AGEMA_reg_buffer_3587 ( .C (clk), .D (new_AGEMA_signal_5542), .Q (new_AGEMA_signal_5543) ) ;
    buf_clk new_AGEMA_reg_buffer_3591 ( .C (clk), .D (new_AGEMA_signal_5546), .Q (new_AGEMA_signal_5547) ) ;
    buf_clk new_AGEMA_reg_buffer_3595 ( .C (clk), .D (new_AGEMA_signal_5550), .Q (new_AGEMA_signal_5551) ) ;
    buf_clk new_AGEMA_reg_buffer_3599 ( .C (clk), .D (new_AGEMA_signal_5554), .Q (new_AGEMA_signal_5555) ) ;
    buf_clk new_AGEMA_reg_buffer_3603 ( .C (clk), .D (new_AGEMA_signal_5558), .Q (new_AGEMA_signal_5559) ) ;
    buf_clk new_AGEMA_reg_buffer_3607 ( .C (clk), .D (new_AGEMA_signal_5562), .Q (new_AGEMA_signal_5563) ) ;
    buf_clk new_AGEMA_reg_buffer_3611 ( .C (clk), .D (new_AGEMA_signal_5566), .Q (new_AGEMA_signal_5567) ) ;
    buf_clk new_AGEMA_reg_buffer_3615 ( .C (clk), .D (new_AGEMA_signal_5570), .Q (new_AGEMA_signal_5571) ) ;
    buf_clk new_AGEMA_reg_buffer_3619 ( .C (clk), .D (new_AGEMA_signal_5574), .Q (new_AGEMA_signal_5575) ) ;
    buf_clk new_AGEMA_reg_buffer_3623 ( .C (clk), .D (new_AGEMA_signal_5578), .Q (new_AGEMA_signal_5579) ) ;
    buf_clk new_AGEMA_reg_buffer_3627 ( .C (clk), .D (new_AGEMA_signal_5582), .Q (new_AGEMA_signal_5583) ) ;
    buf_clk new_AGEMA_reg_buffer_3631 ( .C (clk), .D (new_AGEMA_signal_5586), .Q (new_AGEMA_signal_5587) ) ;
    buf_clk new_AGEMA_reg_buffer_3635 ( .C (clk), .D (new_AGEMA_signal_5590), .Q (new_AGEMA_signal_5591) ) ;
    buf_clk new_AGEMA_reg_buffer_3639 ( .C (clk), .D (new_AGEMA_signal_5594), .Q (new_AGEMA_signal_5595) ) ;
    buf_clk new_AGEMA_reg_buffer_3643 ( .C (clk), .D (new_AGEMA_signal_5598), .Q (new_AGEMA_signal_5599) ) ;
    buf_clk new_AGEMA_reg_buffer_3647 ( .C (clk), .D (new_AGEMA_signal_5602), .Q (new_AGEMA_signal_5603) ) ;
    buf_clk new_AGEMA_reg_buffer_3651 ( .C (clk), .D (new_AGEMA_signal_5606), .Q (new_AGEMA_signal_5607) ) ;
    buf_clk new_AGEMA_reg_buffer_3655 ( .C (clk), .D (new_AGEMA_signal_5610), .Q (new_AGEMA_signal_5611) ) ;
    buf_clk new_AGEMA_reg_buffer_3659 ( .C (clk), .D (new_AGEMA_signal_5614), .Q (new_AGEMA_signal_5615) ) ;
    buf_clk new_AGEMA_reg_buffer_3663 ( .C (clk), .D (new_AGEMA_signal_5618), .Q (new_AGEMA_signal_5619) ) ;
    buf_clk new_AGEMA_reg_buffer_3667 ( .C (clk), .D (new_AGEMA_signal_5622), .Q (new_AGEMA_signal_5623) ) ;
    buf_clk new_AGEMA_reg_buffer_3671 ( .C (clk), .D (new_AGEMA_signal_5626), .Q (new_AGEMA_signal_5627) ) ;
    buf_clk new_AGEMA_reg_buffer_3675 ( .C (clk), .D (new_AGEMA_signal_5630), .Q (new_AGEMA_signal_5631) ) ;
    buf_clk new_AGEMA_reg_buffer_3679 ( .C (clk), .D (new_AGEMA_signal_5634), .Q (new_AGEMA_signal_5635) ) ;
    buf_clk new_AGEMA_reg_buffer_3683 ( .C (clk), .D (new_AGEMA_signal_5638), .Q (new_AGEMA_signal_5639) ) ;
    buf_clk new_AGEMA_reg_buffer_3687 ( .C (clk), .D (new_AGEMA_signal_5642), .Q (new_AGEMA_signal_5643) ) ;
    buf_clk new_AGEMA_reg_buffer_3691 ( .C (clk), .D (new_AGEMA_signal_5646), .Q (new_AGEMA_signal_5647) ) ;
    buf_clk new_AGEMA_reg_buffer_3695 ( .C (clk), .D (new_AGEMA_signal_5650), .Q (new_AGEMA_signal_5651) ) ;
    buf_clk new_AGEMA_reg_buffer_3699 ( .C (clk), .D (new_AGEMA_signal_5654), .Q (new_AGEMA_signal_5655) ) ;
    buf_clk new_AGEMA_reg_buffer_3703 ( .C (clk), .D (new_AGEMA_signal_5658), .Q (new_AGEMA_signal_5659) ) ;
    buf_clk new_AGEMA_reg_buffer_3707 ( .C (clk), .D (new_AGEMA_signal_5662), .Q (new_AGEMA_signal_5663) ) ;
    buf_clk new_AGEMA_reg_buffer_3711 ( .C (clk), .D (new_AGEMA_signal_5666), .Q (new_AGEMA_signal_5667) ) ;
    buf_clk new_AGEMA_reg_buffer_3715 ( .C (clk), .D (new_AGEMA_signal_5670), .Q (new_AGEMA_signal_5671) ) ;
    buf_clk new_AGEMA_reg_buffer_3719 ( .C (clk), .D (new_AGEMA_signal_5674), .Q (new_AGEMA_signal_5675) ) ;
    buf_clk new_AGEMA_reg_buffer_3723 ( .C (clk), .D (new_AGEMA_signal_5678), .Q (new_AGEMA_signal_5679) ) ;
    buf_clk new_AGEMA_reg_buffer_3727 ( .C (clk), .D (new_AGEMA_signal_5682), .Q (new_AGEMA_signal_5683) ) ;
    buf_clk new_AGEMA_reg_buffer_3731 ( .C (clk), .D (new_AGEMA_signal_5686), .Q (new_AGEMA_signal_5687) ) ;
    buf_clk new_AGEMA_reg_buffer_3735 ( .C (clk), .D (new_AGEMA_signal_5690), .Q (new_AGEMA_signal_5691) ) ;
    buf_clk new_AGEMA_reg_buffer_3739 ( .C (clk), .D (new_AGEMA_signal_5694), .Q (new_AGEMA_signal_5695) ) ;
    buf_clk new_AGEMA_reg_buffer_3743 ( .C (clk), .D (new_AGEMA_signal_5698), .Q (new_AGEMA_signal_5699) ) ;
    buf_clk new_AGEMA_reg_buffer_3747 ( .C (clk), .D (new_AGEMA_signal_5702), .Q (new_AGEMA_signal_5703) ) ;
    buf_clk new_AGEMA_reg_buffer_3751 ( .C (clk), .D (new_AGEMA_signal_5706), .Q (new_AGEMA_signal_5707) ) ;
    buf_clk new_AGEMA_reg_buffer_3755 ( .C (clk), .D (new_AGEMA_signal_5710), .Q (new_AGEMA_signal_5711) ) ;
    buf_clk new_AGEMA_reg_buffer_3759 ( .C (clk), .D (new_AGEMA_signal_5714), .Q (new_AGEMA_signal_5715) ) ;
    buf_clk new_AGEMA_reg_buffer_3763 ( .C (clk), .D (new_AGEMA_signal_5718), .Q (new_AGEMA_signal_5719) ) ;
    buf_clk new_AGEMA_reg_buffer_3767 ( .C (clk), .D (new_AGEMA_signal_5722), .Q (new_AGEMA_signal_5723) ) ;
    buf_clk new_AGEMA_reg_buffer_3771 ( .C (clk), .D (new_AGEMA_signal_5726), .Q (new_AGEMA_signal_5727) ) ;
    buf_clk new_AGEMA_reg_buffer_3775 ( .C (clk), .D (new_AGEMA_signal_5730), .Q (new_AGEMA_signal_5731) ) ;
    buf_clk new_AGEMA_reg_buffer_3779 ( .C (clk), .D (new_AGEMA_signal_5734), .Q (new_AGEMA_signal_5735) ) ;
    buf_clk new_AGEMA_reg_buffer_3783 ( .C (clk), .D (new_AGEMA_signal_5738), .Q (new_AGEMA_signal_5739) ) ;
    buf_clk new_AGEMA_reg_buffer_3787 ( .C (clk), .D (new_AGEMA_signal_5742), .Q (new_AGEMA_signal_5743) ) ;
    buf_clk new_AGEMA_reg_buffer_3791 ( .C (clk), .D (new_AGEMA_signal_5746), .Q (new_AGEMA_signal_5747) ) ;
    buf_clk new_AGEMA_reg_buffer_3795 ( .C (clk), .D (new_AGEMA_signal_5750), .Q (new_AGEMA_signal_5751) ) ;
    buf_clk new_AGEMA_reg_buffer_3799 ( .C (clk), .D (new_AGEMA_signal_5754), .Q (new_AGEMA_signal_5755) ) ;
    buf_clk new_AGEMA_reg_buffer_3803 ( .C (clk), .D (new_AGEMA_signal_5758), .Q (new_AGEMA_signal_5759) ) ;
    buf_clk new_AGEMA_reg_buffer_3807 ( .C (clk), .D (new_AGEMA_signal_5762), .Q (new_AGEMA_signal_5763) ) ;
    buf_clk new_AGEMA_reg_buffer_3811 ( .C (clk), .D (new_AGEMA_signal_5766), .Q (new_AGEMA_signal_5767) ) ;
    buf_clk new_AGEMA_reg_buffer_3815 ( .C (clk), .D (new_AGEMA_signal_5770), .Q (new_AGEMA_signal_5771) ) ;
    buf_clk new_AGEMA_reg_buffer_3819 ( .C (clk), .D (new_AGEMA_signal_5774), .Q (new_AGEMA_signal_5775) ) ;
    buf_clk new_AGEMA_reg_buffer_3823 ( .C (clk), .D (new_AGEMA_signal_5778), .Q (new_AGEMA_signal_5779) ) ;
    buf_clk new_AGEMA_reg_buffer_3827 ( .C (clk), .D (new_AGEMA_signal_5782), .Q (new_AGEMA_signal_5783) ) ;
    buf_clk new_AGEMA_reg_buffer_3831 ( .C (clk), .D (new_AGEMA_signal_5786), .Q (new_AGEMA_signal_5787) ) ;
    buf_clk new_AGEMA_reg_buffer_3835 ( .C (clk), .D (new_AGEMA_signal_5790), .Q (new_AGEMA_signal_5791) ) ;
    buf_clk new_AGEMA_reg_buffer_3839 ( .C (clk), .D (new_AGEMA_signal_5794), .Q (new_AGEMA_signal_5795) ) ;
    buf_clk new_AGEMA_reg_buffer_3843 ( .C (clk), .D (new_AGEMA_signal_5798), .Q (new_AGEMA_signal_5799) ) ;
    buf_clk new_AGEMA_reg_buffer_3847 ( .C (clk), .D (new_AGEMA_signal_5802), .Q (new_AGEMA_signal_5803) ) ;
    buf_clk new_AGEMA_reg_buffer_3851 ( .C (clk), .D (new_AGEMA_signal_5806), .Q (new_AGEMA_signal_5807) ) ;
    buf_clk new_AGEMA_reg_buffer_3855 ( .C (clk), .D (new_AGEMA_signal_5810), .Q (new_AGEMA_signal_5811) ) ;
    buf_clk new_AGEMA_reg_buffer_3859 ( .C (clk), .D (new_AGEMA_signal_5814), .Q (new_AGEMA_signal_5815) ) ;
    buf_clk new_AGEMA_reg_buffer_3863 ( .C (clk), .D (new_AGEMA_signal_5818), .Q (new_AGEMA_signal_5819) ) ;
    buf_clk new_AGEMA_reg_buffer_3867 ( .C (clk), .D (new_AGEMA_signal_5822), .Q (new_AGEMA_signal_5823) ) ;
    buf_clk new_AGEMA_reg_buffer_3871 ( .C (clk), .D (new_AGEMA_signal_5826), .Q (new_AGEMA_signal_5827) ) ;
    buf_clk new_AGEMA_reg_buffer_3875 ( .C (clk), .D (new_AGEMA_signal_5830), .Q (new_AGEMA_signal_5831) ) ;
    buf_clk new_AGEMA_reg_buffer_3879 ( .C (clk), .D (new_AGEMA_signal_5834), .Q (new_AGEMA_signal_5835) ) ;
    buf_clk new_AGEMA_reg_buffer_3883 ( .C (clk), .D (new_AGEMA_signal_5838), .Q (new_AGEMA_signal_5839) ) ;
    buf_clk new_AGEMA_reg_buffer_3887 ( .C (clk), .D (new_AGEMA_signal_5842), .Q (new_AGEMA_signal_5843) ) ;
    buf_clk new_AGEMA_reg_buffer_3891 ( .C (clk), .D (new_AGEMA_signal_5846), .Q (new_AGEMA_signal_5847) ) ;
    buf_clk new_AGEMA_reg_buffer_3895 ( .C (clk), .D (new_AGEMA_signal_5850), .Q (new_AGEMA_signal_5851) ) ;
    buf_clk new_AGEMA_reg_buffer_3899 ( .C (clk), .D (new_AGEMA_signal_5854), .Q (new_AGEMA_signal_5855) ) ;
    buf_clk new_AGEMA_reg_buffer_3903 ( .C (clk), .D (new_AGEMA_signal_5858), .Q (new_AGEMA_signal_5859) ) ;
    buf_clk new_AGEMA_reg_buffer_3907 ( .C (clk), .D (new_AGEMA_signal_5862), .Q (new_AGEMA_signal_5863) ) ;
    buf_clk new_AGEMA_reg_buffer_3911 ( .C (clk), .D (new_AGEMA_signal_5866), .Q (new_AGEMA_signal_5867) ) ;
    buf_clk new_AGEMA_reg_buffer_3915 ( .C (clk), .D (new_AGEMA_signal_5870), .Q (new_AGEMA_signal_5871) ) ;
    buf_clk new_AGEMA_reg_buffer_3919 ( .C (clk), .D (new_AGEMA_signal_5874), .Q (new_AGEMA_signal_5875) ) ;
    buf_clk new_AGEMA_reg_buffer_3923 ( .C (clk), .D (new_AGEMA_signal_5878), .Q (new_AGEMA_signal_5879) ) ;
    buf_clk new_AGEMA_reg_buffer_3927 ( .C (clk), .D (new_AGEMA_signal_5882), .Q (new_AGEMA_signal_5883) ) ;
    buf_clk new_AGEMA_reg_buffer_3931 ( .C (clk), .D (new_AGEMA_signal_5886), .Q (new_AGEMA_signal_5887) ) ;
    buf_clk new_AGEMA_reg_buffer_3935 ( .C (clk), .D (new_AGEMA_signal_5890), .Q (new_AGEMA_signal_5891) ) ;
    buf_clk new_AGEMA_reg_buffer_3939 ( .C (clk), .D (new_AGEMA_signal_5894), .Q (new_AGEMA_signal_5895) ) ;
    buf_clk new_AGEMA_reg_buffer_3943 ( .C (clk), .D (new_AGEMA_signal_5898), .Q (new_AGEMA_signal_5899) ) ;
    buf_clk new_AGEMA_reg_buffer_3947 ( .C (clk), .D (new_AGEMA_signal_5902), .Q (new_AGEMA_signal_5903) ) ;
    buf_clk new_AGEMA_reg_buffer_3951 ( .C (clk), .D (new_AGEMA_signal_5906), .Q (new_AGEMA_signal_5907) ) ;
    buf_clk new_AGEMA_reg_buffer_3955 ( .C (clk), .D (new_AGEMA_signal_5910), .Q (new_AGEMA_signal_5911) ) ;
    buf_clk new_AGEMA_reg_buffer_3959 ( .C (clk), .D (new_AGEMA_signal_5914), .Q (new_AGEMA_signal_5915) ) ;
    buf_clk new_AGEMA_reg_buffer_3963 ( .C (clk), .D (new_AGEMA_signal_5918), .Q (new_AGEMA_signal_5919) ) ;
    buf_clk new_AGEMA_reg_buffer_3967 ( .C (clk), .D (new_AGEMA_signal_5922), .Q (new_AGEMA_signal_5923) ) ;
    buf_clk new_AGEMA_reg_buffer_3971 ( .C (clk), .D (new_AGEMA_signal_5926), .Q (new_AGEMA_signal_5927) ) ;
    buf_clk new_AGEMA_reg_buffer_3975 ( .C (clk), .D (new_AGEMA_signal_5930), .Q (new_AGEMA_signal_5931) ) ;
    buf_clk new_AGEMA_reg_buffer_3979 ( .C (clk), .D (new_AGEMA_signal_5934), .Q (new_AGEMA_signal_5935) ) ;
    buf_clk new_AGEMA_reg_buffer_3983 ( .C (clk), .D (new_AGEMA_signal_5938), .Q (new_AGEMA_signal_5939) ) ;
    buf_clk new_AGEMA_reg_buffer_3987 ( .C (clk), .D (new_AGEMA_signal_5942), .Q (new_AGEMA_signal_5943) ) ;
    buf_clk new_AGEMA_reg_buffer_3991 ( .C (clk), .D (new_AGEMA_signal_5946), .Q (new_AGEMA_signal_5947) ) ;
    buf_clk new_AGEMA_reg_buffer_3995 ( .C (clk), .D (new_AGEMA_signal_5950), .Q (new_AGEMA_signal_5951) ) ;
    buf_clk new_AGEMA_reg_buffer_3999 ( .C (clk), .D (new_AGEMA_signal_5954), .Q (new_AGEMA_signal_5955) ) ;
    buf_clk new_AGEMA_reg_buffer_4003 ( .C (clk), .D (new_AGEMA_signal_5958), .Q (new_AGEMA_signal_5959) ) ;
    buf_clk new_AGEMA_reg_buffer_4007 ( .C (clk), .D (new_AGEMA_signal_5962), .Q (new_AGEMA_signal_5963) ) ;
    buf_clk new_AGEMA_reg_buffer_4011 ( .C (clk), .D (new_AGEMA_signal_5966), .Q (new_AGEMA_signal_5967) ) ;
    buf_clk new_AGEMA_reg_buffer_4015 ( .C (clk), .D (new_AGEMA_signal_5970), .Q (new_AGEMA_signal_5971) ) ;
    buf_clk new_AGEMA_reg_buffer_4019 ( .C (clk), .D (new_AGEMA_signal_5974), .Q (new_AGEMA_signal_5975) ) ;
    buf_clk new_AGEMA_reg_buffer_4023 ( .C (clk), .D (new_AGEMA_signal_5978), .Q (new_AGEMA_signal_5979) ) ;
    buf_clk new_AGEMA_reg_buffer_4027 ( .C (clk), .D (new_AGEMA_signal_5982), .Q (new_AGEMA_signal_5983) ) ;
    buf_clk new_AGEMA_reg_buffer_4031 ( .C (clk), .D (new_AGEMA_signal_5986), .Q (new_AGEMA_signal_5987) ) ;
    buf_clk new_AGEMA_reg_buffer_4035 ( .C (clk), .D (new_AGEMA_signal_5990), .Q (new_AGEMA_signal_5991) ) ;
    buf_clk new_AGEMA_reg_buffer_4039 ( .C (clk), .D (new_AGEMA_signal_5994), .Q (new_AGEMA_signal_5995) ) ;
    buf_clk new_AGEMA_reg_buffer_4043 ( .C (clk), .D (new_AGEMA_signal_5998), .Q (new_AGEMA_signal_5999) ) ;
    buf_clk new_AGEMA_reg_buffer_4047 ( .C (clk), .D (new_AGEMA_signal_6002), .Q (new_AGEMA_signal_6003) ) ;
    buf_clk new_AGEMA_reg_buffer_4051 ( .C (clk), .D (new_AGEMA_signal_6006), .Q (new_AGEMA_signal_6007) ) ;
    buf_clk new_AGEMA_reg_buffer_4055 ( .C (clk), .D (new_AGEMA_signal_6010), .Q (new_AGEMA_signal_6011) ) ;
    buf_clk new_AGEMA_reg_buffer_4059 ( .C (clk), .D (new_AGEMA_signal_6014), .Q (new_AGEMA_signal_6015) ) ;
    buf_clk new_AGEMA_reg_buffer_4063 ( .C (clk), .D (new_AGEMA_signal_6018), .Q (new_AGEMA_signal_6019) ) ;
    buf_clk new_AGEMA_reg_buffer_4067 ( .C (clk), .D (new_AGEMA_signal_6022), .Q (new_AGEMA_signal_6023) ) ;
    buf_clk new_AGEMA_reg_buffer_4071 ( .C (clk), .D (new_AGEMA_signal_6026), .Q (new_AGEMA_signal_6027) ) ;
    buf_clk new_AGEMA_reg_buffer_4075 ( .C (clk), .D (new_AGEMA_signal_6030), .Q (new_AGEMA_signal_6031) ) ;
    buf_clk new_AGEMA_reg_buffer_4079 ( .C (clk), .D (new_AGEMA_signal_6034), .Q (new_AGEMA_signal_6035) ) ;
    buf_clk new_AGEMA_reg_buffer_4083 ( .C (clk), .D (new_AGEMA_signal_6038), .Q (new_AGEMA_signal_6039) ) ;
    buf_clk new_AGEMA_reg_buffer_4087 ( .C (clk), .D (new_AGEMA_signal_6042), .Q (new_AGEMA_signal_6043) ) ;
    buf_clk new_AGEMA_reg_buffer_4091 ( .C (clk), .D (new_AGEMA_signal_6046), .Q (new_AGEMA_signal_6047) ) ;
    buf_clk new_AGEMA_reg_buffer_4095 ( .C (clk), .D (new_AGEMA_signal_6050), .Q (new_AGEMA_signal_6051) ) ;
    buf_clk new_AGEMA_reg_buffer_4099 ( .C (clk), .D (new_AGEMA_signal_6054), .Q (new_AGEMA_signal_6055) ) ;
    buf_clk new_AGEMA_reg_buffer_4103 ( .C (clk), .D (new_AGEMA_signal_6058), .Q (new_AGEMA_signal_6059) ) ;
    buf_clk new_AGEMA_reg_buffer_4107 ( .C (clk), .D (new_AGEMA_signal_6062), .Q (new_AGEMA_signal_6063) ) ;
    buf_clk new_AGEMA_reg_buffer_4111 ( .C (clk), .D (new_AGEMA_signal_6066), .Q (new_AGEMA_signal_6067) ) ;
    buf_clk new_AGEMA_reg_buffer_4115 ( .C (clk), .D (new_AGEMA_signal_6070), .Q (new_AGEMA_signal_6071) ) ;
    buf_clk new_AGEMA_reg_buffer_4119 ( .C (clk), .D (new_AGEMA_signal_6074), .Q (new_AGEMA_signal_6075) ) ;
    buf_clk new_AGEMA_reg_buffer_4123 ( .C (clk), .D (new_AGEMA_signal_6078), .Q (new_AGEMA_signal_6079) ) ;
    buf_clk new_AGEMA_reg_buffer_4127 ( .C (clk), .D (new_AGEMA_signal_6082), .Q (new_AGEMA_signal_6083) ) ;
    buf_clk new_AGEMA_reg_buffer_4131 ( .C (clk), .D (new_AGEMA_signal_6086), .Q (new_AGEMA_signal_6087) ) ;
    buf_clk new_AGEMA_reg_buffer_4135 ( .C (clk), .D (new_AGEMA_signal_6090), .Q (new_AGEMA_signal_6091) ) ;
    buf_clk new_AGEMA_reg_buffer_4139 ( .C (clk), .D (new_AGEMA_signal_6094), .Q (new_AGEMA_signal_6095) ) ;
    buf_clk new_AGEMA_reg_buffer_4143 ( .C (clk), .D (new_AGEMA_signal_6098), .Q (new_AGEMA_signal_6099) ) ;
    buf_clk new_AGEMA_reg_buffer_4147 ( .C (clk), .D (new_AGEMA_signal_6102), .Q (new_AGEMA_signal_6103) ) ;
    buf_clk new_AGEMA_reg_buffer_4151 ( .C (clk), .D (new_AGEMA_signal_6106), .Q (new_AGEMA_signal_6107) ) ;
    buf_clk new_AGEMA_reg_buffer_4155 ( .C (clk), .D (new_AGEMA_signal_6110), .Q (new_AGEMA_signal_6111) ) ;
    buf_clk new_AGEMA_reg_buffer_4159 ( .C (clk), .D (new_AGEMA_signal_6114), .Q (new_AGEMA_signal_6115) ) ;
    buf_clk new_AGEMA_reg_buffer_4163 ( .C (clk), .D (new_AGEMA_signal_6118), .Q (new_AGEMA_signal_6119) ) ;
    buf_clk new_AGEMA_reg_buffer_4167 ( .C (clk), .D (new_AGEMA_signal_6122), .Q (new_AGEMA_signal_6123) ) ;
    buf_clk new_AGEMA_reg_buffer_4171 ( .C (clk), .D (new_AGEMA_signal_6126), .Q (new_AGEMA_signal_6127) ) ;
    buf_clk new_AGEMA_reg_buffer_4175 ( .C (clk), .D (new_AGEMA_signal_6130), .Q (new_AGEMA_signal_6131) ) ;
    buf_clk new_AGEMA_reg_buffer_4179 ( .C (clk), .D (new_AGEMA_signal_6134), .Q (new_AGEMA_signal_6135) ) ;
    buf_clk new_AGEMA_reg_buffer_4183 ( .C (clk), .D (new_AGEMA_signal_6138), .Q (new_AGEMA_signal_6139) ) ;
    buf_clk new_AGEMA_reg_buffer_4187 ( .C (clk), .D (new_AGEMA_signal_6142), .Q (new_AGEMA_signal_6143) ) ;
    buf_clk new_AGEMA_reg_buffer_4191 ( .C (clk), .D (new_AGEMA_signal_6146), .Q (new_AGEMA_signal_6147) ) ;
    buf_clk new_AGEMA_reg_buffer_4195 ( .C (clk), .D (new_AGEMA_signal_6150), .Q (new_AGEMA_signal_6151) ) ;
    buf_clk new_AGEMA_reg_buffer_4199 ( .C (clk), .D (new_AGEMA_signal_6154), .Q (new_AGEMA_signal_6155) ) ;
    buf_clk new_AGEMA_reg_buffer_4203 ( .C (clk), .D (new_AGEMA_signal_6158), .Q (new_AGEMA_signal_6159) ) ;
    buf_clk new_AGEMA_reg_buffer_4207 ( .C (clk), .D (new_AGEMA_signal_6162), .Q (new_AGEMA_signal_6163) ) ;
    buf_clk new_AGEMA_reg_buffer_4211 ( .C (clk), .D (new_AGEMA_signal_6166), .Q (new_AGEMA_signal_6167) ) ;
    buf_clk new_AGEMA_reg_buffer_4215 ( .C (clk), .D (new_AGEMA_signal_6170), .Q (new_AGEMA_signal_6171) ) ;
    buf_clk new_AGEMA_reg_buffer_4219 ( .C (clk), .D (new_AGEMA_signal_6174), .Q (new_AGEMA_signal_6175) ) ;
    buf_clk new_AGEMA_reg_buffer_4223 ( .C (clk), .D (new_AGEMA_signal_6178), .Q (new_AGEMA_signal_6179) ) ;
    buf_clk new_AGEMA_reg_buffer_4227 ( .C (clk), .D (new_AGEMA_signal_6182), .Q (new_AGEMA_signal_6183) ) ;
    buf_clk new_AGEMA_reg_buffer_4231 ( .C (clk), .D (new_AGEMA_signal_6186), .Q (new_AGEMA_signal_6187) ) ;
    buf_clk new_AGEMA_reg_buffer_4235 ( .C (clk), .D (new_AGEMA_signal_6190), .Q (new_AGEMA_signal_6191) ) ;
    buf_clk new_AGEMA_reg_buffer_4239 ( .C (clk), .D (new_AGEMA_signal_6194), .Q (new_AGEMA_signal_6195) ) ;
    buf_clk new_AGEMA_reg_buffer_4243 ( .C (clk), .D (new_AGEMA_signal_6198), .Q (new_AGEMA_signal_6199) ) ;
    buf_clk new_AGEMA_reg_buffer_4247 ( .C (clk), .D (new_AGEMA_signal_6202), .Q (new_AGEMA_signal_6203) ) ;
    buf_clk new_AGEMA_reg_buffer_4251 ( .C (clk), .D (new_AGEMA_signal_6206), .Q (new_AGEMA_signal_6207) ) ;
    buf_clk new_AGEMA_reg_buffer_4255 ( .C (clk), .D (new_AGEMA_signal_6210), .Q (new_AGEMA_signal_6211) ) ;
    buf_clk new_AGEMA_reg_buffer_4259 ( .C (clk), .D (new_AGEMA_signal_6214), .Q (new_AGEMA_signal_6215) ) ;
    buf_clk new_AGEMA_reg_buffer_4263 ( .C (clk), .D (new_AGEMA_signal_6218), .Q (new_AGEMA_signal_6219) ) ;
    buf_clk new_AGEMA_reg_buffer_4267 ( .C (clk), .D (new_AGEMA_signal_6222), .Q (new_AGEMA_signal_6223) ) ;
    buf_clk new_AGEMA_reg_buffer_4271 ( .C (clk), .D (new_AGEMA_signal_6226), .Q (new_AGEMA_signal_6227) ) ;
    buf_clk new_AGEMA_reg_buffer_4275 ( .C (clk), .D (new_AGEMA_signal_6230), .Q (new_AGEMA_signal_6231) ) ;
    buf_clk new_AGEMA_reg_buffer_4279 ( .C (clk), .D (new_AGEMA_signal_6234), .Q (new_AGEMA_signal_6235) ) ;
    buf_clk new_AGEMA_reg_buffer_4283 ( .C (clk), .D (new_AGEMA_signal_6238), .Q (new_AGEMA_signal_6239) ) ;
    buf_clk new_AGEMA_reg_buffer_4287 ( .C (clk), .D (new_AGEMA_signal_6242), .Q (new_AGEMA_signal_6243) ) ;
    buf_clk new_AGEMA_reg_buffer_4291 ( .C (clk), .D (new_AGEMA_signal_6246), .Q (new_AGEMA_signal_6247) ) ;
    buf_clk new_AGEMA_reg_buffer_4295 ( .C (clk), .D (new_AGEMA_signal_6250), .Q (new_AGEMA_signal_6251) ) ;
    buf_clk new_AGEMA_reg_buffer_4299 ( .C (clk), .D (new_AGEMA_signal_6254), .Q (new_AGEMA_signal_6255) ) ;
    buf_clk new_AGEMA_reg_buffer_4303 ( .C (clk), .D (new_AGEMA_signal_6258), .Q (new_AGEMA_signal_6259) ) ;
    buf_clk new_AGEMA_reg_buffer_4307 ( .C (clk), .D (new_AGEMA_signal_6262), .Q (new_AGEMA_signal_6263) ) ;
    buf_clk new_AGEMA_reg_buffer_4311 ( .C (clk), .D (new_AGEMA_signal_6266), .Q (new_AGEMA_signal_6267) ) ;
    buf_clk new_AGEMA_reg_buffer_4315 ( .C (clk), .D (new_AGEMA_signal_6270), .Q (new_AGEMA_signal_6271) ) ;
    buf_clk new_AGEMA_reg_buffer_4319 ( .C (clk), .D (new_AGEMA_signal_6274), .Q (new_AGEMA_signal_6275) ) ;
    buf_clk new_AGEMA_reg_buffer_4323 ( .C (clk), .D (new_AGEMA_signal_6278), .Q (new_AGEMA_signal_6279) ) ;
    buf_clk new_AGEMA_reg_buffer_4327 ( .C (clk), .D (new_AGEMA_signal_6282), .Q (new_AGEMA_signal_6283) ) ;
    buf_clk new_AGEMA_reg_buffer_4331 ( .C (clk), .D (new_AGEMA_signal_6286), .Q (new_AGEMA_signal_6287) ) ;
    buf_clk new_AGEMA_reg_buffer_4335 ( .C (clk), .D (new_AGEMA_signal_6290), .Q (new_AGEMA_signal_6291) ) ;
    buf_clk new_AGEMA_reg_buffer_4339 ( .C (clk), .D (new_AGEMA_signal_6294), .Q (new_AGEMA_signal_6295) ) ;

    /* cells in depth 3 */
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M29_U1 ( .a ({new_AGEMA_signal_3389, Inst_bSbox_M28}), .b ({new_AGEMA_signal_3683, new_AGEMA_signal_3682}), .clk (clk), .r ({Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_3392, Inst_bSbox_M29}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M30_U1 ( .a ({new_AGEMA_signal_3388, Inst_bSbox_M26}), .b ({new_AGEMA_signal_3685, new_AGEMA_signal_3684}), .clk (clk), .r ({Fresh[55], Fresh[54], Fresh[53], Fresh[52]}), .c ({new_AGEMA_signal_3393, Inst_bSbox_M30}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M32_U1 ( .a ({new_AGEMA_signal_3683, new_AGEMA_signal_3682}), .b ({new_AGEMA_signal_3390, Inst_bSbox_M31}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56]}), .c ({new_AGEMA_signal_3394, Inst_bSbox_M32}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M35_U1 ( .a ({new_AGEMA_signal_3685, new_AGEMA_signal_3684}), .b ({new_AGEMA_signal_3386, Inst_bSbox_M34}), .clk (clk), .r ({Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_3395, Inst_bSbox_M35}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_M37_U1 ( .a ({new_AGEMA_signal_3687, new_AGEMA_signal_3686}), .b ({new_AGEMA_signal_3392, Inst_bSbox_M29}), .c ({new_AGEMA_signal_3397, Inst_bSbox_M37}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_M38_U1 ( .a ({new_AGEMA_signal_3394, Inst_bSbox_M32}), .b ({new_AGEMA_signal_3689, new_AGEMA_signal_3688}), .c ({new_AGEMA_signal_3398, Inst_bSbox_M38}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_M39_U1 ( .a ({new_AGEMA_signal_3691, new_AGEMA_signal_3690}), .b ({new_AGEMA_signal_3393, Inst_bSbox_M30}), .c ({new_AGEMA_signal_3399, Inst_bSbox_M39}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_M40_U1 ( .a ({new_AGEMA_signal_3395, Inst_bSbox_M35}), .b ({new_AGEMA_signal_3693, new_AGEMA_signal_3692}), .c ({new_AGEMA_signal_3400, Inst_bSbox_M40}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_M41_U1 ( .a ({new_AGEMA_signal_3398, Inst_bSbox_M38}), .b ({new_AGEMA_signal_3400, Inst_bSbox_M40}), .c ({new_AGEMA_signal_3401, Inst_bSbox_M41}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_M42_U1 ( .a ({new_AGEMA_signal_3397, Inst_bSbox_M37}), .b ({new_AGEMA_signal_3399, Inst_bSbox_M39}), .c ({new_AGEMA_signal_3402, Inst_bSbox_M42}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_M43_U1 ( .a ({new_AGEMA_signal_3397, Inst_bSbox_M37}), .b ({new_AGEMA_signal_3398, Inst_bSbox_M38}), .c ({new_AGEMA_signal_3403, Inst_bSbox_M43}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_M44_U1 ( .a ({new_AGEMA_signal_3399, Inst_bSbox_M39}), .b ({new_AGEMA_signal_3400, Inst_bSbox_M40}), .c ({new_AGEMA_signal_3404, Inst_bSbox_M44}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_M45_U1 ( .a ({new_AGEMA_signal_3402, Inst_bSbox_M42}), .b ({new_AGEMA_signal_3401, Inst_bSbox_M41}), .c ({new_AGEMA_signal_3413, Inst_bSbox_M45}) ) ;
    buf_clk new_AGEMA_reg_buffer_1730 ( .C (clk), .D (new_AGEMA_signal_3678), .Q (new_AGEMA_signal_3686) ) ;
    buf_clk new_AGEMA_reg_buffer_1731 ( .C (clk), .D (new_AGEMA_signal_3679), .Q (new_AGEMA_signal_3687) ) ;
    buf_clk new_AGEMA_reg_buffer_1732 ( .C (clk), .D (Inst_bSbox_M33), .Q (new_AGEMA_signal_3688) ) ;
    buf_clk new_AGEMA_reg_buffer_1733 ( .C (clk), .D (new_AGEMA_signal_3391), .Q (new_AGEMA_signal_3689) ) ;
    buf_clk new_AGEMA_reg_buffer_1734 ( .C (clk), .D (new_AGEMA_signal_3680), .Q (new_AGEMA_signal_3690) ) ;
    buf_clk new_AGEMA_reg_buffer_1735 ( .C (clk), .D (new_AGEMA_signal_3681), .Q (new_AGEMA_signal_3691) ) ;
    buf_clk new_AGEMA_reg_buffer_1736 ( .C (clk), .D (Inst_bSbox_M36), .Q (new_AGEMA_signal_3692) ) ;
    buf_clk new_AGEMA_reg_buffer_1737 ( .C (clk), .D (new_AGEMA_signal_3396), .Q (new_AGEMA_signal_3693) ) ;
    buf_clk new_AGEMA_reg_buffer_1740 ( .C (clk), .D (new_AGEMA_signal_3695), .Q (new_AGEMA_signal_3696) ) ;
    buf_clk new_AGEMA_reg_buffer_1744 ( .C (clk), .D (new_AGEMA_signal_3699), .Q (new_AGEMA_signal_3700) ) ;
    buf_clk new_AGEMA_reg_buffer_1748 ( .C (clk), .D (new_AGEMA_signal_3703), .Q (new_AGEMA_signal_3704) ) ;
    buf_clk new_AGEMA_reg_buffer_1752 ( .C (clk), .D (new_AGEMA_signal_3707), .Q (new_AGEMA_signal_3708) ) ;
    buf_clk new_AGEMA_reg_buffer_1756 ( .C (clk), .D (new_AGEMA_signal_3711), .Q (new_AGEMA_signal_3712) ) ;
    buf_clk new_AGEMA_reg_buffer_1760 ( .C (clk), .D (new_AGEMA_signal_3715), .Q (new_AGEMA_signal_3716) ) ;
    buf_clk new_AGEMA_reg_buffer_1764 ( .C (clk), .D (new_AGEMA_signal_3719), .Q (new_AGEMA_signal_3720) ) ;
    buf_clk new_AGEMA_reg_buffer_1768 ( .C (clk), .D (new_AGEMA_signal_3723), .Q (new_AGEMA_signal_3724) ) ;
    buf_clk new_AGEMA_reg_buffer_1772 ( .C (clk), .D (new_AGEMA_signal_3727), .Q (new_AGEMA_signal_3728) ) ;
    buf_clk new_AGEMA_reg_buffer_1776 ( .C (clk), .D (new_AGEMA_signal_3731), .Q (new_AGEMA_signal_3732) ) ;
    buf_clk new_AGEMA_reg_buffer_1780 ( .C (clk), .D (new_AGEMA_signal_3735), .Q (new_AGEMA_signal_3736) ) ;
    buf_clk new_AGEMA_reg_buffer_1784 ( .C (clk), .D (new_AGEMA_signal_3739), .Q (new_AGEMA_signal_3740) ) ;
    buf_clk new_AGEMA_reg_buffer_1788 ( .C (clk), .D (new_AGEMA_signal_3743), .Q (new_AGEMA_signal_3744) ) ;
    buf_clk new_AGEMA_reg_buffer_1792 ( .C (clk), .D (new_AGEMA_signal_3747), .Q (new_AGEMA_signal_3748) ) ;
    buf_clk new_AGEMA_reg_buffer_1796 ( .C (clk), .D (new_AGEMA_signal_3751), .Q (new_AGEMA_signal_3752) ) ;
    buf_clk new_AGEMA_reg_buffer_1800 ( .C (clk), .D (new_AGEMA_signal_3755), .Q (new_AGEMA_signal_3756) ) ;
    buf_clk new_AGEMA_reg_buffer_1804 ( .C (clk), .D (new_AGEMA_signal_3759), .Q (new_AGEMA_signal_3760) ) ;
    buf_clk new_AGEMA_reg_buffer_1808 ( .C (clk), .D (new_AGEMA_signal_3763), .Q (new_AGEMA_signal_3764) ) ;
    buf_clk new_AGEMA_reg_buffer_1812 ( .C (clk), .D (new_AGEMA_signal_3767), .Q (new_AGEMA_signal_3768) ) ;
    buf_clk new_AGEMA_reg_buffer_1816 ( .C (clk), .D (new_AGEMA_signal_3771), .Q (new_AGEMA_signal_3772) ) ;
    buf_clk new_AGEMA_reg_buffer_1820 ( .C (clk), .D (new_AGEMA_signal_3775), .Q (new_AGEMA_signal_3776) ) ;
    buf_clk new_AGEMA_reg_buffer_1824 ( .C (clk), .D (new_AGEMA_signal_3779), .Q (new_AGEMA_signal_3780) ) ;
    buf_clk new_AGEMA_reg_buffer_1828 ( .C (clk), .D (new_AGEMA_signal_3783), .Q (new_AGEMA_signal_3784) ) ;
    buf_clk new_AGEMA_reg_buffer_1832 ( .C (clk), .D (new_AGEMA_signal_3787), .Q (new_AGEMA_signal_3788) ) ;
    buf_clk new_AGEMA_reg_buffer_1836 ( .C (clk), .D (new_AGEMA_signal_3791), .Q (new_AGEMA_signal_3792) ) ;
    buf_clk new_AGEMA_reg_buffer_1840 ( .C (clk), .D (new_AGEMA_signal_3795), .Q (new_AGEMA_signal_3796) ) ;
    buf_clk new_AGEMA_reg_buffer_1844 ( .C (clk), .D (new_AGEMA_signal_3799), .Q (new_AGEMA_signal_3800) ) ;
    buf_clk new_AGEMA_reg_buffer_1848 ( .C (clk), .D (new_AGEMA_signal_3803), .Q (new_AGEMA_signal_3804) ) ;
    buf_clk new_AGEMA_reg_buffer_1852 ( .C (clk), .D (new_AGEMA_signal_3807), .Q (new_AGEMA_signal_3808) ) ;
    buf_clk new_AGEMA_reg_buffer_1856 ( .C (clk), .D (new_AGEMA_signal_3811), .Q (new_AGEMA_signal_3812) ) ;
    buf_clk new_AGEMA_reg_buffer_1860 ( .C (clk), .D (new_AGEMA_signal_3815), .Q (new_AGEMA_signal_3816) ) ;
    buf_clk new_AGEMA_reg_buffer_1864 ( .C (clk), .D (new_AGEMA_signal_3819), .Q (new_AGEMA_signal_3820) ) ;
    buf_clk new_AGEMA_reg_buffer_1868 ( .C (clk), .D (new_AGEMA_signal_3823), .Q (new_AGEMA_signal_3824) ) ;
    buf_clk new_AGEMA_reg_buffer_1872 ( .C (clk), .D (new_AGEMA_signal_3827), .Q (new_AGEMA_signal_3828) ) ;
    buf_clk new_AGEMA_reg_buffer_1876 ( .C (clk), .D (new_AGEMA_signal_3831), .Q (new_AGEMA_signal_3832) ) ;
    buf_clk new_AGEMA_reg_buffer_1880 ( .C (clk), .D (new_AGEMA_signal_3835), .Q (new_AGEMA_signal_3836) ) ;
    buf_clk new_AGEMA_reg_buffer_1884 ( .C (clk), .D (new_AGEMA_signal_3839), .Q (new_AGEMA_signal_3840) ) ;
    buf_clk new_AGEMA_reg_buffer_1888 ( .C (clk), .D (new_AGEMA_signal_3843), .Q (new_AGEMA_signal_3844) ) ;
    buf_clk new_AGEMA_reg_buffer_1892 ( .C (clk), .D (new_AGEMA_signal_3847), .Q (new_AGEMA_signal_3848) ) ;
    buf_clk new_AGEMA_reg_buffer_1896 ( .C (clk), .D (new_AGEMA_signal_3851), .Q (new_AGEMA_signal_3852) ) ;
    buf_clk new_AGEMA_reg_buffer_1900 ( .C (clk), .D (new_AGEMA_signal_3855), .Q (new_AGEMA_signal_3856) ) ;
    buf_clk new_AGEMA_reg_buffer_1904 ( .C (clk), .D (new_AGEMA_signal_3859), .Q (new_AGEMA_signal_3860) ) ;
    buf_clk new_AGEMA_reg_buffer_1908 ( .C (clk), .D (new_AGEMA_signal_3863), .Q (new_AGEMA_signal_3864) ) ;
    buf_clk new_AGEMA_reg_buffer_1912 ( .C (clk), .D (new_AGEMA_signal_3867), .Q (new_AGEMA_signal_3868) ) ;
    buf_clk new_AGEMA_reg_buffer_1916 ( .C (clk), .D (new_AGEMA_signal_3871), .Q (new_AGEMA_signal_3872) ) ;
    buf_clk new_AGEMA_reg_buffer_1920 ( .C (clk), .D (new_AGEMA_signal_3875), .Q (new_AGEMA_signal_3876) ) ;
    buf_clk new_AGEMA_reg_buffer_1924 ( .C (clk), .D (new_AGEMA_signal_3879), .Q (new_AGEMA_signal_3880) ) ;
    buf_clk new_AGEMA_reg_buffer_1928 ( .C (clk), .D (new_AGEMA_signal_3883), .Q (new_AGEMA_signal_3884) ) ;
    buf_clk new_AGEMA_reg_buffer_1932 ( .C (clk), .D (new_AGEMA_signal_3887), .Q (new_AGEMA_signal_3888) ) ;
    buf_clk new_AGEMA_reg_buffer_1936 ( .C (clk), .D (new_AGEMA_signal_3891), .Q (new_AGEMA_signal_3892) ) ;
    buf_clk new_AGEMA_reg_buffer_1940 ( .C (clk), .D (new_AGEMA_signal_3895), .Q (new_AGEMA_signal_3896) ) ;
    buf_clk new_AGEMA_reg_buffer_1944 ( .C (clk), .D (new_AGEMA_signal_3899), .Q (new_AGEMA_signal_3900) ) ;
    buf_clk new_AGEMA_reg_buffer_1948 ( .C (clk), .D (new_AGEMA_signal_3903), .Q (new_AGEMA_signal_3904) ) ;
    buf_clk new_AGEMA_reg_buffer_1952 ( .C (clk), .D (new_AGEMA_signal_3907), .Q (new_AGEMA_signal_3908) ) ;
    buf_clk new_AGEMA_reg_buffer_1956 ( .C (clk), .D (new_AGEMA_signal_3911), .Q (new_AGEMA_signal_3912) ) ;
    buf_clk new_AGEMA_reg_buffer_1960 ( .C (clk), .D (new_AGEMA_signal_3915), .Q (new_AGEMA_signal_3916) ) ;
    buf_clk new_AGEMA_reg_buffer_1964 ( .C (clk), .D (new_AGEMA_signal_3919), .Q (new_AGEMA_signal_3920) ) ;
    buf_clk new_AGEMA_reg_buffer_1968 ( .C (clk), .D (new_AGEMA_signal_3923), .Q (new_AGEMA_signal_3924) ) ;
    buf_clk new_AGEMA_reg_buffer_1972 ( .C (clk), .D (new_AGEMA_signal_3927), .Q (new_AGEMA_signal_3928) ) ;
    buf_clk new_AGEMA_reg_buffer_1976 ( .C (clk), .D (new_AGEMA_signal_3931), .Q (new_AGEMA_signal_3932) ) ;
    buf_clk new_AGEMA_reg_buffer_1980 ( .C (clk), .D (new_AGEMA_signal_3935), .Q (new_AGEMA_signal_3936) ) ;
    buf_clk new_AGEMA_reg_buffer_1984 ( .C (clk), .D (new_AGEMA_signal_3939), .Q (new_AGEMA_signal_3940) ) ;
    buf_clk new_AGEMA_reg_buffer_1988 ( .C (clk), .D (new_AGEMA_signal_3943), .Q (new_AGEMA_signal_3944) ) ;
    buf_clk new_AGEMA_reg_buffer_1992 ( .C (clk), .D (new_AGEMA_signal_3947), .Q (new_AGEMA_signal_3948) ) ;
    buf_clk new_AGEMA_reg_buffer_1996 ( .C (clk), .D (new_AGEMA_signal_3951), .Q (new_AGEMA_signal_3952) ) ;
    buf_clk new_AGEMA_reg_buffer_2000 ( .C (clk), .D (new_AGEMA_signal_3955), .Q (new_AGEMA_signal_3956) ) ;
    buf_clk new_AGEMA_reg_buffer_2004 ( .C (clk), .D (new_AGEMA_signal_3959), .Q (new_AGEMA_signal_3960) ) ;
    buf_clk new_AGEMA_reg_buffer_2008 ( .C (clk), .D (new_AGEMA_signal_3963), .Q (new_AGEMA_signal_3964) ) ;
    buf_clk new_AGEMA_reg_buffer_2012 ( .C (clk), .D (new_AGEMA_signal_3967), .Q (new_AGEMA_signal_3968) ) ;
    buf_clk new_AGEMA_reg_buffer_2016 ( .C (clk), .D (new_AGEMA_signal_3971), .Q (new_AGEMA_signal_3972) ) ;
    buf_clk new_AGEMA_reg_buffer_2020 ( .C (clk), .D (new_AGEMA_signal_3975), .Q (new_AGEMA_signal_3976) ) ;
    buf_clk new_AGEMA_reg_buffer_2024 ( .C (clk), .D (new_AGEMA_signal_3979), .Q (new_AGEMA_signal_3980) ) ;
    buf_clk new_AGEMA_reg_buffer_2028 ( .C (clk), .D (new_AGEMA_signal_3983), .Q (new_AGEMA_signal_3984) ) ;
    buf_clk new_AGEMA_reg_buffer_2032 ( .C (clk), .D (new_AGEMA_signal_3987), .Q (new_AGEMA_signal_3988) ) ;
    buf_clk new_AGEMA_reg_buffer_2036 ( .C (clk), .D (new_AGEMA_signal_3991), .Q (new_AGEMA_signal_3992) ) ;
    buf_clk new_AGEMA_reg_buffer_2040 ( .C (clk), .D (new_AGEMA_signal_3995), .Q (new_AGEMA_signal_3996) ) ;
    buf_clk new_AGEMA_reg_buffer_2044 ( .C (clk), .D (new_AGEMA_signal_3999), .Q (new_AGEMA_signal_4000) ) ;
    buf_clk new_AGEMA_reg_buffer_2048 ( .C (clk), .D (new_AGEMA_signal_4003), .Q (new_AGEMA_signal_4004) ) ;
    buf_clk new_AGEMA_reg_buffer_2052 ( .C (clk), .D (new_AGEMA_signal_4007), .Q (new_AGEMA_signal_4008) ) ;
    buf_clk new_AGEMA_reg_buffer_2056 ( .C (clk), .D (new_AGEMA_signal_4011), .Q (new_AGEMA_signal_4012) ) ;
    buf_clk new_AGEMA_reg_buffer_2060 ( .C (clk), .D (new_AGEMA_signal_4015), .Q (new_AGEMA_signal_4016) ) ;
    buf_clk new_AGEMA_reg_buffer_2064 ( .C (clk), .D (new_AGEMA_signal_4019), .Q (new_AGEMA_signal_4020) ) ;
    buf_clk new_AGEMA_reg_buffer_2068 ( .C (clk), .D (new_AGEMA_signal_4023), .Q (new_AGEMA_signal_4024) ) ;
    buf_clk new_AGEMA_reg_buffer_2072 ( .C (clk), .D (new_AGEMA_signal_4027), .Q (new_AGEMA_signal_4028) ) ;
    buf_clk new_AGEMA_reg_buffer_2076 ( .C (clk), .D (new_AGEMA_signal_4031), .Q (new_AGEMA_signal_4032) ) ;
    buf_clk new_AGEMA_reg_buffer_2080 ( .C (clk), .D (new_AGEMA_signal_4035), .Q (new_AGEMA_signal_4036) ) ;
    buf_clk new_AGEMA_reg_buffer_2084 ( .C (clk), .D (new_AGEMA_signal_4039), .Q (new_AGEMA_signal_4040) ) ;
    buf_clk new_AGEMA_reg_buffer_2088 ( .C (clk), .D (new_AGEMA_signal_4043), .Q (new_AGEMA_signal_4044) ) ;
    buf_clk new_AGEMA_reg_buffer_2092 ( .C (clk), .D (new_AGEMA_signal_4047), .Q (new_AGEMA_signal_4048) ) ;
    buf_clk new_AGEMA_reg_buffer_2096 ( .C (clk), .D (new_AGEMA_signal_4051), .Q (new_AGEMA_signal_4052) ) ;
    buf_clk new_AGEMA_reg_buffer_2100 ( .C (clk), .D (new_AGEMA_signal_4055), .Q (new_AGEMA_signal_4056) ) ;
    buf_clk new_AGEMA_reg_buffer_2104 ( .C (clk), .D (new_AGEMA_signal_4059), .Q (new_AGEMA_signal_4060) ) ;
    buf_clk new_AGEMA_reg_buffer_2108 ( .C (clk), .D (new_AGEMA_signal_4063), .Q (new_AGEMA_signal_4064) ) ;
    buf_clk new_AGEMA_reg_buffer_2112 ( .C (clk), .D (new_AGEMA_signal_4067), .Q (new_AGEMA_signal_4068) ) ;
    buf_clk new_AGEMA_reg_buffer_2116 ( .C (clk), .D (new_AGEMA_signal_4071), .Q (new_AGEMA_signal_4072) ) ;
    buf_clk new_AGEMA_reg_buffer_2120 ( .C (clk), .D (new_AGEMA_signal_4075), .Q (new_AGEMA_signal_4076) ) ;
    buf_clk new_AGEMA_reg_buffer_2124 ( .C (clk), .D (new_AGEMA_signal_4079), .Q (new_AGEMA_signal_4080) ) ;
    buf_clk new_AGEMA_reg_buffer_2128 ( .C (clk), .D (new_AGEMA_signal_4083), .Q (new_AGEMA_signal_4084) ) ;
    buf_clk new_AGEMA_reg_buffer_2132 ( .C (clk), .D (new_AGEMA_signal_4087), .Q (new_AGEMA_signal_4088) ) ;
    buf_clk new_AGEMA_reg_buffer_2136 ( .C (clk), .D (new_AGEMA_signal_4091), .Q (new_AGEMA_signal_4092) ) ;
    buf_clk new_AGEMA_reg_buffer_2140 ( .C (clk), .D (new_AGEMA_signal_4095), .Q (new_AGEMA_signal_4096) ) ;
    buf_clk new_AGEMA_reg_buffer_2144 ( .C (clk), .D (new_AGEMA_signal_4099), .Q (new_AGEMA_signal_4100) ) ;
    buf_clk new_AGEMA_reg_buffer_2148 ( .C (clk), .D (new_AGEMA_signal_4103), .Q (new_AGEMA_signal_4104) ) ;
    buf_clk new_AGEMA_reg_buffer_2152 ( .C (clk), .D (new_AGEMA_signal_4107), .Q (new_AGEMA_signal_4108) ) ;
    buf_clk new_AGEMA_reg_buffer_2156 ( .C (clk), .D (new_AGEMA_signal_4111), .Q (new_AGEMA_signal_4112) ) ;
    buf_clk new_AGEMA_reg_buffer_2160 ( .C (clk), .D (new_AGEMA_signal_4115), .Q (new_AGEMA_signal_4116) ) ;
    buf_clk new_AGEMA_reg_buffer_2164 ( .C (clk), .D (new_AGEMA_signal_4119), .Q (new_AGEMA_signal_4120) ) ;
    buf_clk new_AGEMA_reg_buffer_2168 ( .C (clk), .D (new_AGEMA_signal_4123), .Q (new_AGEMA_signal_4124) ) ;
    buf_clk new_AGEMA_reg_buffer_2172 ( .C (clk), .D (new_AGEMA_signal_4127), .Q (new_AGEMA_signal_4128) ) ;
    buf_clk new_AGEMA_reg_buffer_2176 ( .C (clk), .D (new_AGEMA_signal_4131), .Q (new_AGEMA_signal_4132) ) ;
    buf_clk new_AGEMA_reg_buffer_2180 ( .C (clk), .D (new_AGEMA_signal_4135), .Q (new_AGEMA_signal_4136) ) ;
    buf_clk new_AGEMA_reg_buffer_2184 ( .C (clk), .D (new_AGEMA_signal_4139), .Q (new_AGEMA_signal_4140) ) ;
    buf_clk new_AGEMA_reg_buffer_2188 ( .C (clk), .D (new_AGEMA_signal_4143), .Q (new_AGEMA_signal_4144) ) ;
    buf_clk new_AGEMA_reg_buffer_2192 ( .C (clk), .D (new_AGEMA_signal_4147), .Q (new_AGEMA_signal_4148) ) ;
    buf_clk new_AGEMA_reg_buffer_2196 ( .C (clk), .D (new_AGEMA_signal_4151), .Q (new_AGEMA_signal_4152) ) ;
    buf_clk new_AGEMA_reg_buffer_2200 ( .C (clk), .D (new_AGEMA_signal_4155), .Q (new_AGEMA_signal_4156) ) ;
    buf_clk new_AGEMA_reg_buffer_2204 ( .C (clk), .D (new_AGEMA_signal_4159), .Q (new_AGEMA_signal_4160) ) ;
    buf_clk new_AGEMA_reg_buffer_2208 ( .C (clk), .D (new_AGEMA_signal_4163), .Q (new_AGEMA_signal_4164) ) ;
    buf_clk new_AGEMA_reg_buffer_2212 ( .C (clk), .D (new_AGEMA_signal_4167), .Q (new_AGEMA_signal_4168) ) ;
    buf_clk new_AGEMA_reg_buffer_2216 ( .C (clk), .D (new_AGEMA_signal_4171), .Q (new_AGEMA_signal_4172) ) ;
    buf_clk new_AGEMA_reg_buffer_2220 ( .C (clk), .D (new_AGEMA_signal_4175), .Q (new_AGEMA_signal_4176) ) ;
    buf_clk new_AGEMA_reg_buffer_2224 ( .C (clk), .D (new_AGEMA_signal_4179), .Q (new_AGEMA_signal_4180) ) ;
    buf_clk new_AGEMA_reg_buffer_2228 ( .C (clk), .D (new_AGEMA_signal_4183), .Q (new_AGEMA_signal_4184) ) ;
    buf_clk new_AGEMA_reg_buffer_2232 ( .C (clk), .D (new_AGEMA_signal_4187), .Q (new_AGEMA_signal_4188) ) ;
    buf_clk new_AGEMA_reg_buffer_2236 ( .C (clk), .D (new_AGEMA_signal_4191), .Q (new_AGEMA_signal_4192) ) ;
    buf_clk new_AGEMA_reg_buffer_2240 ( .C (clk), .D (new_AGEMA_signal_4195), .Q (new_AGEMA_signal_4196) ) ;
    buf_clk new_AGEMA_reg_buffer_2244 ( .C (clk), .D (new_AGEMA_signal_4199), .Q (new_AGEMA_signal_4200) ) ;
    buf_clk new_AGEMA_reg_buffer_2247 ( .C (clk), .D (new_AGEMA_signal_4202), .Q (new_AGEMA_signal_4203) ) ;
    buf_clk new_AGEMA_reg_buffer_2250 ( .C (clk), .D (new_AGEMA_signal_4205), .Q (new_AGEMA_signal_4206) ) ;
    buf_clk new_AGEMA_reg_buffer_2253 ( .C (clk), .D (new_AGEMA_signal_4208), .Q (new_AGEMA_signal_4209) ) ;
    buf_clk new_AGEMA_reg_buffer_2256 ( .C (clk), .D (new_AGEMA_signal_4211), .Q (new_AGEMA_signal_4212) ) ;
    buf_clk new_AGEMA_reg_buffer_2259 ( .C (clk), .D (new_AGEMA_signal_4214), .Q (new_AGEMA_signal_4215) ) ;
    buf_clk new_AGEMA_reg_buffer_2262 ( .C (clk), .D (new_AGEMA_signal_4217), .Q (new_AGEMA_signal_4218) ) ;
    buf_clk new_AGEMA_reg_buffer_2265 ( .C (clk), .D (new_AGEMA_signal_4220), .Q (new_AGEMA_signal_4221) ) ;
    buf_clk new_AGEMA_reg_buffer_2268 ( .C (clk), .D (new_AGEMA_signal_4223), .Q (new_AGEMA_signal_4224) ) ;
    buf_clk new_AGEMA_reg_buffer_2271 ( .C (clk), .D (new_AGEMA_signal_4226), .Q (new_AGEMA_signal_4227) ) ;
    buf_clk new_AGEMA_reg_buffer_2274 ( .C (clk), .D (new_AGEMA_signal_4229), .Q (new_AGEMA_signal_4230) ) ;
    buf_clk new_AGEMA_reg_buffer_2277 ( .C (clk), .D (new_AGEMA_signal_4232), .Q (new_AGEMA_signal_4233) ) ;
    buf_clk new_AGEMA_reg_buffer_2280 ( .C (clk), .D (new_AGEMA_signal_4235), .Q (new_AGEMA_signal_4236) ) ;
    buf_clk new_AGEMA_reg_buffer_2283 ( .C (clk), .D (new_AGEMA_signal_4238), .Q (new_AGEMA_signal_4239) ) ;
    buf_clk new_AGEMA_reg_buffer_2286 ( .C (clk), .D (new_AGEMA_signal_4241), .Q (new_AGEMA_signal_4242) ) ;
    buf_clk new_AGEMA_reg_buffer_2289 ( .C (clk), .D (new_AGEMA_signal_4244), .Q (new_AGEMA_signal_4245) ) ;
    buf_clk new_AGEMA_reg_buffer_2292 ( .C (clk), .D (new_AGEMA_signal_4247), .Q (new_AGEMA_signal_4248) ) ;
    buf_clk new_AGEMA_reg_buffer_2295 ( .C (clk), .D (new_AGEMA_signal_4250), .Q (new_AGEMA_signal_4251) ) ;
    buf_clk new_AGEMA_reg_buffer_2298 ( .C (clk), .D (new_AGEMA_signal_4253), .Q (new_AGEMA_signal_4254) ) ;
    buf_clk new_AGEMA_reg_buffer_2301 ( .C (clk), .D (new_AGEMA_signal_4256), .Q (new_AGEMA_signal_4257) ) ;
    buf_clk new_AGEMA_reg_buffer_2304 ( .C (clk), .D (new_AGEMA_signal_4259), .Q (new_AGEMA_signal_4260) ) ;
    buf_clk new_AGEMA_reg_buffer_2307 ( .C (clk), .D (new_AGEMA_signal_4262), .Q (new_AGEMA_signal_4263) ) ;
    buf_clk new_AGEMA_reg_buffer_2310 ( .C (clk), .D (new_AGEMA_signal_4265), .Q (new_AGEMA_signal_4266) ) ;
    buf_clk new_AGEMA_reg_buffer_2313 ( .C (clk), .D (new_AGEMA_signal_4268), .Q (new_AGEMA_signal_4269) ) ;
    buf_clk new_AGEMA_reg_buffer_2316 ( .C (clk), .D (new_AGEMA_signal_4271), .Q (new_AGEMA_signal_4272) ) ;
    buf_clk new_AGEMA_reg_buffer_2319 ( .C (clk), .D (new_AGEMA_signal_4274), .Q (new_AGEMA_signal_4275) ) ;
    buf_clk new_AGEMA_reg_buffer_2322 ( .C (clk), .D (new_AGEMA_signal_4277), .Q (new_AGEMA_signal_4278) ) ;
    buf_clk new_AGEMA_reg_buffer_2325 ( .C (clk), .D (new_AGEMA_signal_4280), .Q (new_AGEMA_signal_4281) ) ;
    buf_clk new_AGEMA_reg_buffer_2328 ( .C (clk), .D (new_AGEMA_signal_4283), .Q (new_AGEMA_signal_4284) ) ;
    buf_clk new_AGEMA_reg_buffer_2331 ( .C (clk), .D (new_AGEMA_signal_4286), .Q (new_AGEMA_signal_4287) ) ;
    buf_clk new_AGEMA_reg_buffer_2334 ( .C (clk), .D (new_AGEMA_signal_4289), .Q (new_AGEMA_signal_4290) ) ;
    buf_clk new_AGEMA_reg_buffer_2337 ( .C (clk), .D (new_AGEMA_signal_4292), .Q (new_AGEMA_signal_4293) ) ;
    buf_clk new_AGEMA_reg_buffer_2340 ( .C (clk), .D (new_AGEMA_signal_4295), .Q (new_AGEMA_signal_4296) ) ;
    buf_clk new_AGEMA_reg_buffer_2343 ( .C (clk), .D (new_AGEMA_signal_4298), .Q (new_AGEMA_signal_4299) ) ;
    buf_clk new_AGEMA_reg_buffer_2346 ( .C (clk), .D (new_AGEMA_signal_4301), .Q (new_AGEMA_signal_4302) ) ;
    buf_clk new_AGEMA_reg_buffer_2349 ( .C (clk), .D (new_AGEMA_signal_4304), .Q (new_AGEMA_signal_4305) ) ;
    buf_clk new_AGEMA_reg_buffer_2352 ( .C (clk), .D (new_AGEMA_signal_4307), .Q (new_AGEMA_signal_4308) ) ;
    buf_clk new_AGEMA_reg_buffer_2356 ( .C (clk), .D (new_AGEMA_signal_4311), .Q (new_AGEMA_signal_4312) ) ;
    buf_clk new_AGEMA_reg_buffer_2360 ( .C (clk), .D (new_AGEMA_signal_4315), .Q (new_AGEMA_signal_4316) ) ;
    buf_clk new_AGEMA_reg_buffer_2364 ( .C (clk), .D (new_AGEMA_signal_4319), .Q (new_AGEMA_signal_4320) ) ;
    buf_clk new_AGEMA_reg_buffer_2368 ( .C (clk), .D (new_AGEMA_signal_4323), .Q (new_AGEMA_signal_4324) ) ;
    buf_clk new_AGEMA_reg_buffer_2372 ( .C (clk), .D (new_AGEMA_signal_4327), .Q (new_AGEMA_signal_4328) ) ;
    buf_clk new_AGEMA_reg_buffer_2376 ( .C (clk), .D (new_AGEMA_signal_4331), .Q (new_AGEMA_signal_4332) ) ;
    buf_clk new_AGEMA_reg_buffer_2380 ( .C (clk), .D (new_AGEMA_signal_4335), .Q (new_AGEMA_signal_4336) ) ;
    buf_clk new_AGEMA_reg_buffer_2384 ( .C (clk), .D (new_AGEMA_signal_4339), .Q (new_AGEMA_signal_4340) ) ;
    buf_clk new_AGEMA_reg_buffer_2388 ( .C (clk), .D (new_AGEMA_signal_4343), .Q (new_AGEMA_signal_4344) ) ;
    buf_clk new_AGEMA_reg_buffer_2392 ( .C (clk), .D (new_AGEMA_signal_4347), .Q (new_AGEMA_signal_4348) ) ;
    buf_clk new_AGEMA_reg_buffer_2396 ( .C (clk), .D (new_AGEMA_signal_4351), .Q (new_AGEMA_signal_4352) ) ;
    buf_clk new_AGEMA_reg_buffer_2400 ( .C (clk), .D (new_AGEMA_signal_4355), .Q (new_AGEMA_signal_4356) ) ;
    buf_clk new_AGEMA_reg_buffer_2404 ( .C (clk), .D (new_AGEMA_signal_4359), .Q (new_AGEMA_signal_4360) ) ;
    buf_clk new_AGEMA_reg_buffer_2408 ( .C (clk), .D (new_AGEMA_signal_4363), .Q (new_AGEMA_signal_4364) ) ;
    buf_clk new_AGEMA_reg_buffer_2412 ( .C (clk), .D (new_AGEMA_signal_4367), .Q (new_AGEMA_signal_4368) ) ;
    buf_clk new_AGEMA_reg_buffer_2416 ( .C (clk), .D (new_AGEMA_signal_4371), .Q (new_AGEMA_signal_4372) ) ;
    buf_clk new_AGEMA_reg_buffer_2420 ( .C (clk), .D (new_AGEMA_signal_4375), .Q (new_AGEMA_signal_4376) ) ;
    buf_clk new_AGEMA_reg_buffer_2424 ( .C (clk), .D (new_AGEMA_signal_4379), .Q (new_AGEMA_signal_4380) ) ;
    buf_clk new_AGEMA_reg_buffer_2428 ( .C (clk), .D (new_AGEMA_signal_4383), .Q (new_AGEMA_signal_4384) ) ;
    buf_clk new_AGEMA_reg_buffer_2432 ( .C (clk), .D (new_AGEMA_signal_4387), .Q (new_AGEMA_signal_4388) ) ;
    buf_clk new_AGEMA_reg_buffer_2436 ( .C (clk), .D (new_AGEMA_signal_4391), .Q (new_AGEMA_signal_4392) ) ;
    buf_clk new_AGEMA_reg_buffer_2440 ( .C (clk), .D (new_AGEMA_signal_4395), .Q (new_AGEMA_signal_4396) ) ;
    buf_clk new_AGEMA_reg_buffer_2444 ( .C (clk), .D (new_AGEMA_signal_4399), .Q (new_AGEMA_signal_4400) ) ;
    buf_clk new_AGEMA_reg_buffer_2448 ( .C (clk), .D (new_AGEMA_signal_4403), .Q (new_AGEMA_signal_4404) ) ;
    buf_clk new_AGEMA_reg_buffer_2452 ( .C (clk), .D (new_AGEMA_signal_4407), .Q (new_AGEMA_signal_4408) ) ;
    buf_clk new_AGEMA_reg_buffer_2456 ( .C (clk), .D (new_AGEMA_signal_4411), .Q (new_AGEMA_signal_4412) ) ;
    buf_clk new_AGEMA_reg_buffer_2460 ( .C (clk), .D (new_AGEMA_signal_4415), .Q (new_AGEMA_signal_4416) ) ;
    buf_clk new_AGEMA_reg_buffer_2464 ( .C (clk), .D (new_AGEMA_signal_4419), .Q (new_AGEMA_signal_4420) ) ;
    buf_clk new_AGEMA_reg_buffer_2468 ( .C (clk), .D (new_AGEMA_signal_4423), .Q (new_AGEMA_signal_4424) ) ;
    buf_clk new_AGEMA_reg_buffer_2472 ( .C (clk), .D (new_AGEMA_signal_4427), .Q (new_AGEMA_signal_4428) ) ;
    buf_clk new_AGEMA_reg_buffer_2476 ( .C (clk), .D (new_AGEMA_signal_4431), .Q (new_AGEMA_signal_4432) ) ;
    buf_clk new_AGEMA_reg_buffer_2480 ( .C (clk), .D (new_AGEMA_signal_4435), .Q (new_AGEMA_signal_4436) ) ;
    buf_clk new_AGEMA_reg_buffer_2484 ( .C (clk), .D (new_AGEMA_signal_4439), .Q (new_AGEMA_signal_4440) ) ;
    buf_clk new_AGEMA_reg_buffer_2488 ( .C (clk), .D (new_AGEMA_signal_4443), .Q (new_AGEMA_signal_4444) ) ;
    buf_clk new_AGEMA_reg_buffer_2492 ( .C (clk), .D (new_AGEMA_signal_4447), .Q (new_AGEMA_signal_4448) ) ;
    buf_clk new_AGEMA_reg_buffer_2496 ( .C (clk), .D (new_AGEMA_signal_4451), .Q (new_AGEMA_signal_4452) ) ;
    buf_clk new_AGEMA_reg_buffer_2500 ( .C (clk), .D (new_AGEMA_signal_4455), .Q (new_AGEMA_signal_4456) ) ;
    buf_clk new_AGEMA_reg_buffer_2504 ( .C (clk), .D (new_AGEMA_signal_4459), .Q (new_AGEMA_signal_4460) ) ;
    buf_clk new_AGEMA_reg_buffer_2508 ( .C (clk), .D (new_AGEMA_signal_4463), .Q (new_AGEMA_signal_4464) ) ;
    buf_clk new_AGEMA_reg_buffer_2512 ( .C (clk), .D (new_AGEMA_signal_4467), .Q (new_AGEMA_signal_4468) ) ;
    buf_clk new_AGEMA_reg_buffer_2516 ( .C (clk), .D (new_AGEMA_signal_4471), .Q (new_AGEMA_signal_4472) ) ;
    buf_clk new_AGEMA_reg_buffer_2520 ( .C (clk), .D (new_AGEMA_signal_4475), .Q (new_AGEMA_signal_4476) ) ;
    buf_clk new_AGEMA_reg_buffer_2524 ( .C (clk), .D (new_AGEMA_signal_4479), .Q (new_AGEMA_signal_4480) ) ;
    buf_clk new_AGEMA_reg_buffer_2528 ( .C (clk), .D (new_AGEMA_signal_4483), .Q (new_AGEMA_signal_4484) ) ;
    buf_clk new_AGEMA_reg_buffer_2532 ( .C (clk), .D (new_AGEMA_signal_4487), .Q (new_AGEMA_signal_4488) ) ;
    buf_clk new_AGEMA_reg_buffer_2536 ( .C (clk), .D (new_AGEMA_signal_4491), .Q (new_AGEMA_signal_4492) ) ;
    buf_clk new_AGEMA_reg_buffer_2540 ( .C (clk), .D (new_AGEMA_signal_4495), .Q (new_AGEMA_signal_4496) ) ;
    buf_clk new_AGEMA_reg_buffer_2544 ( .C (clk), .D (new_AGEMA_signal_4499), .Q (new_AGEMA_signal_4500) ) ;
    buf_clk new_AGEMA_reg_buffer_2548 ( .C (clk), .D (new_AGEMA_signal_4503), .Q (new_AGEMA_signal_4504) ) ;
    buf_clk new_AGEMA_reg_buffer_2552 ( .C (clk), .D (new_AGEMA_signal_4507), .Q (new_AGEMA_signal_4508) ) ;
    buf_clk new_AGEMA_reg_buffer_2556 ( .C (clk), .D (new_AGEMA_signal_4511), .Q (new_AGEMA_signal_4512) ) ;
    buf_clk new_AGEMA_reg_buffer_2560 ( .C (clk), .D (new_AGEMA_signal_4515), .Q (new_AGEMA_signal_4516) ) ;
    buf_clk new_AGEMA_reg_buffer_2564 ( .C (clk), .D (new_AGEMA_signal_4519), .Q (new_AGEMA_signal_4520) ) ;
    buf_clk new_AGEMA_reg_buffer_2568 ( .C (clk), .D (new_AGEMA_signal_4523), .Q (new_AGEMA_signal_4524) ) ;
    buf_clk new_AGEMA_reg_buffer_2572 ( .C (clk), .D (new_AGEMA_signal_4527), .Q (new_AGEMA_signal_4528) ) ;
    buf_clk new_AGEMA_reg_buffer_2576 ( .C (clk), .D (new_AGEMA_signal_4531), .Q (new_AGEMA_signal_4532) ) ;
    buf_clk new_AGEMA_reg_buffer_2580 ( .C (clk), .D (new_AGEMA_signal_4535), .Q (new_AGEMA_signal_4536) ) ;
    buf_clk new_AGEMA_reg_buffer_2584 ( .C (clk), .D (new_AGEMA_signal_4539), .Q (new_AGEMA_signal_4540) ) ;
    buf_clk new_AGEMA_reg_buffer_2588 ( .C (clk), .D (new_AGEMA_signal_4543), .Q (new_AGEMA_signal_4544) ) ;
    buf_clk new_AGEMA_reg_buffer_2592 ( .C (clk), .D (new_AGEMA_signal_4547), .Q (new_AGEMA_signal_4548) ) ;
    buf_clk new_AGEMA_reg_buffer_2596 ( .C (clk), .D (new_AGEMA_signal_4551), .Q (new_AGEMA_signal_4552) ) ;
    buf_clk new_AGEMA_reg_buffer_2600 ( .C (clk), .D (new_AGEMA_signal_4555), .Q (new_AGEMA_signal_4556) ) ;
    buf_clk new_AGEMA_reg_buffer_2604 ( .C (clk), .D (new_AGEMA_signal_4559), .Q (new_AGEMA_signal_4560) ) ;
    buf_clk new_AGEMA_reg_buffer_2608 ( .C (clk), .D (new_AGEMA_signal_4563), .Q (new_AGEMA_signal_4564) ) ;
    buf_clk new_AGEMA_reg_buffer_2612 ( .C (clk), .D (new_AGEMA_signal_4567), .Q (new_AGEMA_signal_4568) ) ;
    buf_clk new_AGEMA_reg_buffer_2616 ( .C (clk), .D (new_AGEMA_signal_4571), .Q (new_AGEMA_signal_4572) ) ;
    buf_clk new_AGEMA_reg_buffer_2620 ( .C (clk), .D (new_AGEMA_signal_4575), .Q (new_AGEMA_signal_4576) ) ;
    buf_clk new_AGEMA_reg_buffer_2624 ( .C (clk), .D (new_AGEMA_signal_4579), .Q (new_AGEMA_signal_4580) ) ;
    buf_clk new_AGEMA_reg_buffer_2628 ( .C (clk), .D (new_AGEMA_signal_4583), .Q (new_AGEMA_signal_4584) ) ;
    buf_clk new_AGEMA_reg_buffer_2632 ( .C (clk), .D (new_AGEMA_signal_4587), .Q (new_AGEMA_signal_4588) ) ;
    buf_clk new_AGEMA_reg_buffer_2636 ( .C (clk), .D (new_AGEMA_signal_4591), .Q (new_AGEMA_signal_4592) ) ;
    buf_clk new_AGEMA_reg_buffer_2640 ( .C (clk), .D (new_AGEMA_signal_4595), .Q (new_AGEMA_signal_4596) ) ;
    buf_clk new_AGEMA_reg_buffer_2644 ( .C (clk), .D (new_AGEMA_signal_4599), .Q (new_AGEMA_signal_4600) ) ;
    buf_clk new_AGEMA_reg_buffer_2648 ( .C (clk), .D (new_AGEMA_signal_4603), .Q (new_AGEMA_signal_4604) ) ;
    buf_clk new_AGEMA_reg_buffer_2652 ( .C (clk), .D (new_AGEMA_signal_4607), .Q (new_AGEMA_signal_4608) ) ;
    buf_clk new_AGEMA_reg_buffer_2656 ( .C (clk), .D (new_AGEMA_signal_4611), .Q (new_AGEMA_signal_4612) ) ;
    buf_clk new_AGEMA_reg_buffer_2660 ( .C (clk), .D (new_AGEMA_signal_4615), .Q (new_AGEMA_signal_4616) ) ;
    buf_clk new_AGEMA_reg_buffer_2664 ( .C (clk), .D (new_AGEMA_signal_4619), .Q (new_AGEMA_signal_4620) ) ;
    buf_clk new_AGEMA_reg_buffer_2668 ( .C (clk), .D (new_AGEMA_signal_4623), .Q (new_AGEMA_signal_4624) ) ;
    buf_clk new_AGEMA_reg_buffer_2672 ( .C (clk), .D (new_AGEMA_signal_4627), .Q (new_AGEMA_signal_4628) ) ;
    buf_clk new_AGEMA_reg_buffer_2676 ( .C (clk), .D (new_AGEMA_signal_4631), .Q (new_AGEMA_signal_4632) ) ;
    buf_clk new_AGEMA_reg_buffer_2680 ( .C (clk), .D (new_AGEMA_signal_4635), .Q (new_AGEMA_signal_4636) ) ;
    buf_clk new_AGEMA_reg_buffer_2684 ( .C (clk), .D (new_AGEMA_signal_4639), .Q (new_AGEMA_signal_4640) ) ;
    buf_clk new_AGEMA_reg_buffer_2688 ( .C (clk), .D (new_AGEMA_signal_4643), .Q (new_AGEMA_signal_4644) ) ;
    buf_clk new_AGEMA_reg_buffer_2692 ( .C (clk), .D (new_AGEMA_signal_4647), .Q (new_AGEMA_signal_4648) ) ;
    buf_clk new_AGEMA_reg_buffer_2696 ( .C (clk), .D (new_AGEMA_signal_4651), .Q (new_AGEMA_signal_4652) ) ;
    buf_clk new_AGEMA_reg_buffer_2700 ( .C (clk), .D (new_AGEMA_signal_4655), .Q (new_AGEMA_signal_4656) ) ;
    buf_clk new_AGEMA_reg_buffer_2704 ( .C (clk), .D (new_AGEMA_signal_4659), .Q (new_AGEMA_signal_4660) ) ;
    buf_clk new_AGEMA_reg_buffer_2708 ( .C (clk), .D (new_AGEMA_signal_4663), .Q (new_AGEMA_signal_4664) ) ;
    buf_clk new_AGEMA_reg_buffer_2712 ( .C (clk), .D (new_AGEMA_signal_4667), .Q (new_AGEMA_signal_4668) ) ;
    buf_clk new_AGEMA_reg_buffer_2716 ( .C (clk), .D (new_AGEMA_signal_4671), .Q (new_AGEMA_signal_4672) ) ;
    buf_clk new_AGEMA_reg_buffer_2720 ( .C (clk), .D (new_AGEMA_signal_4675), .Q (new_AGEMA_signal_4676) ) ;
    buf_clk new_AGEMA_reg_buffer_2724 ( .C (clk), .D (new_AGEMA_signal_4679), .Q (new_AGEMA_signal_4680) ) ;
    buf_clk new_AGEMA_reg_buffer_2728 ( .C (clk), .D (new_AGEMA_signal_4683), .Q (new_AGEMA_signal_4684) ) ;
    buf_clk new_AGEMA_reg_buffer_2732 ( .C (clk), .D (new_AGEMA_signal_4687), .Q (new_AGEMA_signal_4688) ) ;
    buf_clk new_AGEMA_reg_buffer_2736 ( .C (clk), .D (new_AGEMA_signal_4691), .Q (new_AGEMA_signal_4692) ) ;
    buf_clk new_AGEMA_reg_buffer_2740 ( .C (clk), .D (new_AGEMA_signal_4695), .Q (new_AGEMA_signal_4696) ) ;
    buf_clk new_AGEMA_reg_buffer_2744 ( .C (clk), .D (new_AGEMA_signal_4699), .Q (new_AGEMA_signal_4700) ) ;
    buf_clk new_AGEMA_reg_buffer_2748 ( .C (clk), .D (new_AGEMA_signal_4703), .Q (new_AGEMA_signal_4704) ) ;
    buf_clk new_AGEMA_reg_buffer_2752 ( .C (clk), .D (new_AGEMA_signal_4707), .Q (new_AGEMA_signal_4708) ) ;
    buf_clk new_AGEMA_reg_buffer_2756 ( .C (clk), .D (new_AGEMA_signal_4711), .Q (new_AGEMA_signal_4712) ) ;
    buf_clk new_AGEMA_reg_buffer_2760 ( .C (clk), .D (new_AGEMA_signal_4715), .Q (new_AGEMA_signal_4716) ) ;
    buf_clk new_AGEMA_reg_buffer_2764 ( .C (clk), .D (new_AGEMA_signal_4719), .Q (new_AGEMA_signal_4720) ) ;
    buf_clk new_AGEMA_reg_buffer_2768 ( .C (clk), .D (new_AGEMA_signal_4723), .Q (new_AGEMA_signal_4724) ) ;
    buf_clk new_AGEMA_reg_buffer_2772 ( .C (clk), .D (new_AGEMA_signal_4727), .Q (new_AGEMA_signal_4728) ) ;
    buf_clk new_AGEMA_reg_buffer_2776 ( .C (clk), .D (new_AGEMA_signal_4731), .Q (new_AGEMA_signal_4732) ) ;
    buf_clk new_AGEMA_reg_buffer_2780 ( .C (clk), .D (new_AGEMA_signal_4735), .Q (new_AGEMA_signal_4736) ) ;
    buf_clk new_AGEMA_reg_buffer_2784 ( .C (clk), .D (new_AGEMA_signal_4739), .Q (new_AGEMA_signal_4740) ) ;
    buf_clk new_AGEMA_reg_buffer_2788 ( .C (clk), .D (new_AGEMA_signal_4743), .Q (new_AGEMA_signal_4744) ) ;
    buf_clk new_AGEMA_reg_buffer_2792 ( .C (clk), .D (new_AGEMA_signal_4747), .Q (new_AGEMA_signal_4748) ) ;
    buf_clk new_AGEMA_reg_buffer_2796 ( .C (clk), .D (new_AGEMA_signal_4751), .Q (new_AGEMA_signal_4752) ) ;
    buf_clk new_AGEMA_reg_buffer_2800 ( .C (clk), .D (new_AGEMA_signal_4755), .Q (new_AGEMA_signal_4756) ) ;
    buf_clk new_AGEMA_reg_buffer_2804 ( .C (clk), .D (new_AGEMA_signal_4759), .Q (new_AGEMA_signal_4760) ) ;
    buf_clk new_AGEMA_reg_buffer_2808 ( .C (clk), .D (new_AGEMA_signal_4763), .Q (new_AGEMA_signal_4764) ) ;
    buf_clk new_AGEMA_reg_buffer_2812 ( .C (clk), .D (new_AGEMA_signal_4767), .Q (new_AGEMA_signal_4768) ) ;
    buf_clk new_AGEMA_reg_buffer_2816 ( .C (clk), .D (new_AGEMA_signal_4771), .Q (new_AGEMA_signal_4772) ) ;
    buf_clk new_AGEMA_reg_buffer_2820 ( .C (clk), .D (new_AGEMA_signal_4775), .Q (new_AGEMA_signal_4776) ) ;
    buf_clk new_AGEMA_reg_buffer_2824 ( .C (clk), .D (new_AGEMA_signal_4779), .Q (new_AGEMA_signal_4780) ) ;
    buf_clk new_AGEMA_reg_buffer_2828 ( .C (clk), .D (new_AGEMA_signal_4783), .Q (new_AGEMA_signal_4784) ) ;
    buf_clk new_AGEMA_reg_buffer_2832 ( .C (clk), .D (new_AGEMA_signal_4787), .Q (new_AGEMA_signal_4788) ) ;
    buf_clk new_AGEMA_reg_buffer_2836 ( .C (clk), .D (new_AGEMA_signal_4791), .Q (new_AGEMA_signal_4792) ) ;
    buf_clk new_AGEMA_reg_buffer_2840 ( .C (clk), .D (new_AGEMA_signal_4795), .Q (new_AGEMA_signal_4796) ) ;
    buf_clk new_AGEMA_reg_buffer_2844 ( .C (clk), .D (new_AGEMA_signal_4799), .Q (new_AGEMA_signal_4800) ) ;
    buf_clk new_AGEMA_reg_buffer_2848 ( .C (clk), .D (new_AGEMA_signal_4803), .Q (new_AGEMA_signal_4804) ) ;
    buf_clk new_AGEMA_reg_buffer_2852 ( .C (clk), .D (new_AGEMA_signal_4807), .Q (new_AGEMA_signal_4808) ) ;
    buf_clk new_AGEMA_reg_buffer_2856 ( .C (clk), .D (new_AGEMA_signal_4811), .Q (new_AGEMA_signal_4812) ) ;
    buf_clk new_AGEMA_reg_buffer_2860 ( .C (clk), .D (new_AGEMA_signal_4815), .Q (new_AGEMA_signal_4816) ) ;
    buf_clk new_AGEMA_reg_buffer_2864 ( .C (clk), .D (new_AGEMA_signal_4819), .Q (new_AGEMA_signal_4820) ) ;
    buf_clk new_AGEMA_reg_buffer_2868 ( .C (clk), .D (new_AGEMA_signal_4823), .Q (new_AGEMA_signal_4824) ) ;
    buf_clk new_AGEMA_reg_buffer_2872 ( .C (clk), .D (new_AGEMA_signal_4827), .Q (new_AGEMA_signal_4828) ) ;
    buf_clk new_AGEMA_reg_buffer_2876 ( .C (clk), .D (new_AGEMA_signal_4831), .Q (new_AGEMA_signal_4832) ) ;
    buf_clk new_AGEMA_reg_buffer_2880 ( .C (clk), .D (new_AGEMA_signal_4835), .Q (new_AGEMA_signal_4836) ) ;
    buf_clk new_AGEMA_reg_buffer_2884 ( .C (clk), .D (new_AGEMA_signal_4839), .Q (new_AGEMA_signal_4840) ) ;
    buf_clk new_AGEMA_reg_buffer_2888 ( .C (clk), .D (new_AGEMA_signal_4843), .Q (new_AGEMA_signal_4844) ) ;
    buf_clk new_AGEMA_reg_buffer_2892 ( .C (clk), .D (new_AGEMA_signal_4847), .Q (new_AGEMA_signal_4848) ) ;
    buf_clk new_AGEMA_reg_buffer_2896 ( .C (clk), .D (new_AGEMA_signal_4851), .Q (new_AGEMA_signal_4852) ) ;
    buf_clk new_AGEMA_reg_buffer_2900 ( .C (clk), .D (new_AGEMA_signal_4855), .Q (new_AGEMA_signal_4856) ) ;
    buf_clk new_AGEMA_reg_buffer_2904 ( .C (clk), .D (new_AGEMA_signal_4859), .Q (new_AGEMA_signal_4860) ) ;
    buf_clk new_AGEMA_reg_buffer_2908 ( .C (clk), .D (new_AGEMA_signal_4863), .Q (new_AGEMA_signal_4864) ) ;
    buf_clk new_AGEMA_reg_buffer_2912 ( .C (clk), .D (new_AGEMA_signal_4867), .Q (new_AGEMA_signal_4868) ) ;
    buf_clk new_AGEMA_reg_buffer_2916 ( .C (clk), .D (new_AGEMA_signal_4871), .Q (new_AGEMA_signal_4872) ) ;
    buf_clk new_AGEMA_reg_buffer_2920 ( .C (clk), .D (new_AGEMA_signal_4875), .Q (new_AGEMA_signal_4876) ) ;
    buf_clk new_AGEMA_reg_buffer_2924 ( .C (clk), .D (new_AGEMA_signal_4879), .Q (new_AGEMA_signal_4880) ) ;
    buf_clk new_AGEMA_reg_buffer_2928 ( .C (clk), .D (new_AGEMA_signal_4883), .Q (new_AGEMA_signal_4884) ) ;
    buf_clk new_AGEMA_reg_buffer_2932 ( .C (clk), .D (new_AGEMA_signal_4887), .Q (new_AGEMA_signal_4888) ) ;
    buf_clk new_AGEMA_reg_buffer_2936 ( .C (clk), .D (new_AGEMA_signal_4891), .Q (new_AGEMA_signal_4892) ) ;
    buf_clk new_AGEMA_reg_buffer_2940 ( .C (clk), .D (new_AGEMA_signal_4895), .Q (new_AGEMA_signal_4896) ) ;
    buf_clk new_AGEMA_reg_buffer_2944 ( .C (clk), .D (new_AGEMA_signal_4899), .Q (new_AGEMA_signal_4900) ) ;
    buf_clk new_AGEMA_reg_buffer_2948 ( .C (clk), .D (new_AGEMA_signal_4903), .Q (new_AGEMA_signal_4904) ) ;
    buf_clk new_AGEMA_reg_buffer_2952 ( .C (clk), .D (new_AGEMA_signal_4907), .Q (new_AGEMA_signal_4908) ) ;
    buf_clk new_AGEMA_reg_buffer_2956 ( .C (clk), .D (new_AGEMA_signal_4911), .Q (new_AGEMA_signal_4912) ) ;
    buf_clk new_AGEMA_reg_buffer_2960 ( .C (clk), .D (new_AGEMA_signal_4915), .Q (new_AGEMA_signal_4916) ) ;
    buf_clk new_AGEMA_reg_buffer_2964 ( .C (clk), .D (new_AGEMA_signal_4919), .Q (new_AGEMA_signal_4920) ) ;
    buf_clk new_AGEMA_reg_buffer_2968 ( .C (clk), .D (new_AGEMA_signal_4923), .Q (new_AGEMA_signal_4924) ) ;
    buf_clk new_AGEMA_reg_buffer_2972 ( .C (clk), .D (new_AGEMA_signal_4927), .Q (new_AGEMA_signal_4928) ) ;
    buf_clk new_AGEMA_reg_buffer_2976 ( .C (clk), .D (new_AGEMA_signal_4931), .Q (new_AGEMA_signal_4932) ) ;
    buf_clk new_AGEMA_reg_buffer_2980 ( .C (clk), .D (new_AGEMA_signal_4935), .Q (new_AGEMA_signal_4936) ) ;
    buf_clk new_AGEMA_reg_buffer_2984 ( .C (clk), .D (new_AGEMA_signal_4939), .Q (new_AGEMA_signal_4940) ) ;
    buf_clk new_AGEMA_reg_buffer_2988 ( .C (clk), .D (new_AGEMA_signal_4943), .Q (new_AGEMA_signal_4944) ) ;
    buf_clk new_AGEMA_reg_buffer_2992 ( .C (clk), .D (new_AGEMA_signal_4947), .Q (new_AGEMA_signal_4948) ) ;
    buf_clk new_AGEMA_reg_buffer_2996 ( .C (clk), .D (new_AGEMA_signal_4951), .Q (new_AGEMA_signal_4952) ) ;
    buf_clk new_AGEMA_reg_buffer_3000 ( .C (clk), .D (new_AGEMA_signal_4955), .Q (new_AGEMA_signal_4956) ) ;
    buf_clk new_AGEMA_reg_buffer_3004 ( .C (clk), .D (new_AGEMA_signal_4959), .Q (new_AGEMA_signal_4960) ) ;
    buf_clk new_AGEMA_reg_buffer_3008 ( .C (clk), .D (new_AGEMA_signal_4963), .Q (new_AGEMA_signal_4964) ) ;
    buf_clk new_AGEMA_reg_buffer_3012 ( .C (clk), .D (new_AGEMA_signal_4967), .Q (new_AGEMA_signal_4968) ) ;
    buf_clk new_AGEMA_reg_buffer_3016 ( .C (clk), .D (new_AGEMA_signal_4971), .Q (new_AGEMA_signal_4972) ) ;
    buf_clk new_AGEMA_reg_buffer_3020 ( .C (clk), .D (new_AGEMA_signal_4975), .Q (new_AGEMA_signal_4976) ) ;
    buf_clk new_AGEMA_reg_buffer_3024 ( .C (clk), .D (new_AGEMA_signal_4979), .Q (new_AGEMA_signal_4980) ) ;
    buf_clk new_AGEMA_reg_buffer_3028 ( .C (clk), .D (new_AGEMA_signal_4983), .Q (new_AGEMA_signal_4984) ) ;
    buf_clk new_AGEMA_reg_buffer_3032 ( .C (clk), .D (new_AGEMA_signal_4987), .Q (new_AGEMA_signal_4988) ) ;
    buf_clk new_AGEMA_reg_buffer_3036 ( .C (clk), .D (new_AGEMA_signal_4991), .Q (new_AGEMA_signal_4992) ) ;
    buf_clk new_AGEMA_reg_buffer_3040 ( .C (clk), .D (new_AGEMA_signal_4995), .Q (new_AGEMA_signal_4996) ) ;
    buf_clk new_AGEMA_reg_buffer_3044 ( .C (clk), .D (new_AGEMA_signal_4999), .Q (new_AGEMA_signal_5000) ) ;
    buf_clk new_AGEMA_reg_buffer_3048 ( .C (clk), .D (new_AGEMA_signal_5003), .Q (new_AGEMA_signal_5004) ) ;
    buf_clk new_AGEMA_reg_buffer_3052 ( .C (clk), .D (new_AGEMA_signal_5007), .Q (new_AGEMA_signal_5008) ) ;
    buf_clk new_AGEMA_reg_buffer_3056 ( .C (clk), .D (new_AGEMA_signal_5011), .Q (new_AGEMA_signal_5012) ) ;
    buf_clk new_AGEMA_reg_buffer_3060 ( .C (clk), .D (new_AGEMA_signal_5015), .Q (new_AGEMA_signal_5016) ) ;
    buf_clk new_AGEMA_reg_buffer_3064 ( .C (clk), .D (new_AGEMA_signal_5019), .Q (new_AGEMA_signal_5020) ) ;
    buf_clk new_AGEMA_reg_buffer_3068 ( .C (clk), .D (new_AGEMA_signal_5023), .Q (new_AGEMA_signal_5024) ) ;
    buf_clk new_AGEMA_reg_buffer_3072 ( .C (clk), .D (new_AGEMA_signal_5027), .Q (new_AGEMA_signal_5028) ) ;
    buf_clk new_AGEMA_reg_buffer_3076 ( .C (clk), .D (new_AGEMA_signal_5031), .Q (new_AGEMA_signal_5032) ) ;
    buf_clk new_AGEMA_reg_buffer_3080 ( .C (clk), .D (new_AGEMA_signal_5035), .Q (new_AGEMA_signal_5036) ) ;
    buf_clk new_AGEMA_reg_buffer_3084 ( .C (clk), .D (new_AGEMA_signal_5039), .Q (new_AGEMA_signal_5040) ) ;
    buf_clk new_AGEMA_reg_buffer_3088 ( .C (clk), .D (new_AGEMA_signal_5043), .Q (new_AGEMA_signal_5044) ) ;
    buf_clk new_AGEMA_reg_buffer_3092 ( .C (clk), .D (new_AGEMA_signal_5047), .Q (new_AGEMA_signal_5048) ) ;
    buf_clk new_AGEMA_reg_buffer_3096 ( .C (clk), .D (new_AGEMA_signal_5051), .Q (new_AGEMA_signal_5052) ) ;
    buf_clk new_AGEMA_reg_buffer_3100 ( .C (clk), .D (new_AGEMA_signal_5055), .Q (new_AGEMA_signal_5056) ) ;
    buf_clk new_AGEMA_reg_buffer_3104 ( .C (clk), .D (new_AGEMA_signal_5059), .Q (new_AGEMA_signal_5060) ) ;
    buf_clk new_AGEMA_reg_buffer_3108 ( .C (clk), .D (new_AGEMA_signal_5063), .Q (new_AGEMA_signal_5064) ) ;
    buf_clk new_AGEMA_reg_buffer_3112 ( .C (clk), .D (new_AGEMA_signal_5067), .Q (new_AGEMA_signal_5068) ) ;
    buf_clk new_AGEMA_reg_buffer_3116 ( .C (clk), .D (new_AGEMA_signal_5071), .Q (new_AGEMA_signal_5072) ) ;
    buf_clk new_AGEMA_reg_buffer_3120 ( .C (clk), .D (new_AGEMA_signal_5075), .Q (new_AGEMA_signal_5076) ) ;
    buf_clk new_AGEMA_reg_buffer_3124 ( .C (clk), .D (new_AGEMA_signal_5079), .Q (new_AGEMA_signal_5080) ) ;
    buf_clk new_AGEMA_reg_buffer_3128 ( .C (clk), .D (new_AGEMA_signal_5083), .Q (new_AGEMA_signal_5084) ) ;
    buf_clk new_AGEMA_reg_buffer_3132 ( .C (clk), .D (new_AGEMA_signal_5087), .Q (new_AGEMA_signal_5088) ) ;
    buf_clk new_AGEMA_reg_buffer_3136 ( .C (clk), .D (new_AGEMA_signal_5091), .Q (new_AGEMA_signal_5092) ) ;
    buf_clk new_AGEMA_reg_buffer_3140 ( .C (clk), .D (new_AGEMA_signal_5095), .Q (new_AGEMA_signal_5096) ) ;
    buf_clk new_AGEMA_reg_buffer_3144 ( .C (clk), .D (new_AGEMA_signal_5099), .Q (new_AGEMA_signal_5100) ) ;
    buf_clk new_AGEMA_reg_buffer_3148 ( .C (clk), .D (new_AGEMA_signal_5103), .Q (new_AGEMA_signal_5104) ) ;
    buf_clk new_AGEMA_reg_buffer_3152 ( .C (clk), .D (new_AGEMA_signal_5107), .Q (new_AGEMA_signal_5108) ) ;
    buf_clk new_AGEMA_reg_buffer_3156 ( .C (clk), .D (new_AGEMA_signal_5111), .Q (new_AGEMA_signal_5112) ) ;
    buf_clk new_AGEMA_reg_buffer_3160 ( .C (clk), .D (new_AGEMA_signal_5115), .Q (new_AGEMA_signal_5116) ) ;
    buf_clk new_AGEMA_reg_buffer_3164 ( .C (clk), .D (new_AGEMA_signal_5119), .Q (new_AGEMA_signal_5120) ) ;
    buf_clk new_AGEMA_reg_buffer_3168 ( .C (clk), .D (new_AGEMA_signal_5123), .Q (new_AGEMA_signal_5124) ) ;
    buf_clk new_AGEMA_reg_buffer_3172 ( .C (clk), .D (new_AGEMA_signal_5127), .Q (new_AGEMA_signal_5128) ) ;
    buf_clk new_AGEMA_reg_buffer_3176 ( .C (clk), .D (new_AGEMA_signal_5131), .Q (new_AGEMA_signal_5132) ) ;
    buf_clk new_AGEMA_reg_buffer_3180 ( .C (clk), .D (new_AGEMA_signal_5135), .Q (new_AGEMA_signal_5136) ) ;
    buf_clk new_AGEMA_reg_buffer_3184 ( .C (clk), .D (new_AGEMA_signal_5139), .Q (new_AGEMA_signal_5140) ) ;
    buf_clk new_AGEMA_reg_buffer_3188 ( .C (clk), .D (new_AGEMA_signal_5143), .Q (new_AGEMA_signal_5144) ) ;
    buf_clk new_AGEMA_reg_buffer_3192 ( .C (clk), .D (new_AGEMA_signal_5147), .Q (new_AGEMA_signal_5148) ) ;
    buf_clk new_AGEMA_reg_buffer_3196 ( .C (clk), .D (new_AGEMA_signal_5151), .Q (new_AGEMA_signal_5152) ) ;
    buf_clk new_AGEMA_reg_buffer_3200 ( .C (clk), .D (new_AGEMA_signal_5155), .Q (new_AGEMA_signal_5156) ) ;
    buf_clk new_AGEMA_reg_buffer_3204 ( .C (clk), .D (new_AGEMA_signal_5159), .Q (new_AGEMA_signal_5160) ) ;
    buf_clk new_AGEMA_reg_buffer_3208 ( .C (clk), .D (new_AGEMA_signal_5163), .Q (new_AGEMA_signal_5164) ) ;
    buf_clk new_AGEMA_reg_buffer_3212 ( .C (clk), .D (new_AGEMA_signal_5167), .Q (new_AGEMA_signal_5168) ) ;
    buf_clk new_AGEMA_reg_buffer_3216 ( .C (clk), .D (new_AGEMA_signal_5171), .Q (new_AGEMA_signal_5172) ) ;
    buf_clk new_AGEMA_reg_buffer_3220 ( .C (clk), .D (new_AGEMA_signal_5175), .Q (new_AGEMA_signal_5176) ) ;
    buf_clk new_AGEMA_reg_buffer_3224 ( .C (clk), .D (new_AGEMA_signal_5179), .Q (new_AGEMA_signal_5180) ) ;
    buf_clk new_AGEMA_reg_buffer_3228 ( .C (clk), .D (new_AGEMA_signal_5183), .Q (new_AGEMA_signal_5184) ) ;
    buf_clk new_AGEMA_reg_buffer_3232 ( .C (clk), .D (new_AGEMA_signal_5187), .Q (new_AGEMA_signal_5188) ) ;
    buf_clk new_AGEMA_reg_buffer_3236 ( .C (clk), .D (new_AGEMA_signal_5191), .Q (new_AGEMA_signal_5192) ) ;
    buf_clk new_AGEMA_reg_buffer_3240 ( .C (clk), .D (new_AGEMA_signal_5195), .Q (new_AGEMA_signal_5196) ) ;
    buf_clk new_AGEMA_reg_buffer_3244 ( .C (clk), .D (new_AGEMA_signal_5199), .Q (new_AGEMA_signal_5200) ) ;
    buf_clk new_AGEMA_reg_buffer_3248 ( .C (clk), .D (new_AGEMA_signal_5203), .Q (new_AGEMA_signal_5204) ) ;
    buf_clk new_AGEMA_reg_buffer_3252 ( .C (clk), .D (new_AGEMA_signal_5207), .Q (new_AGEMA_signal_5208) ) ;
    buf_clk new_AGEMA_reg_buffer_3256 ( .C (clk), .D (new_AGEMA_signal_5211), .Q (new_AGEMA_signal_5212) ) ;
    buf_clk new_AGEMA_reg_buffer_3260 ( .C (clk), .D (new_AGEMA_signal_5215), .Q (new_AGEMA_signal_5216) ) ;
    buf_clk new_AGEMA_reg_buffer_3264 ( .C (clk), .D (new_AGEMA_signal_5219), .Q (new_AGEMA_signal_5220) ) ;
    buf_clk new_AGEMA_reg_buffer_3268 ( .C (clk), .D (new_AGEMA_signal_5223), .Q (new_AGEMA_signal_5224) ) ;
    buf_clk new_AGEMA_reg_buffer_3272 ( .C (clk), .D (new_AGEMA_signal_5227), .Q (new_AGEMA_signal_5228) ) ;
    buf_clk new_AGEMA_reg_buffer_3276 ( .C (clk), .D (new_AGEMA_signal_5231), .Q (new_AGEMA_signal_5232) ) ;
    buf_clk new_AGEMA_reg_buffer_3280 ( .C (clk), .D (new_AGEMA_signal_5235), .Q (new_AGEMA_signal_5236) ) ;
    buf_clk new_AGEMA_reg_buffer_3284 ( .C (clk), .D (new_AGEMA_signal_5239), .Q (new_AGEMA_signal_5240) ) ;
    buf_clk new_AGEMA_reg_buffer_3288 ( .C (clk), .D (new_AGEMA_signal_5243), .Q (new_AGEMA_signal_5244) ) ;
    buf_clk new_AGEMA_reg_buffer_3292 ( .C (clk), .D (new_AGEMA_signal_5247), .Q (new_AGEMA_signal_5248) ) ;
    buf_clk new_AGEMA_reg_buffer_3296 ( .C (clk), .D (new_AGEMA_signal_5251), .Q (new_AGEMA_signal_5252) ) ;
    buf_clk new_AGEMA_reg_buffer_3300 ( .C (clk), .D (new_AGEMA_signal_5255), .Q (new_AGEMA_signal_5256) ) ;
    buf_clk new_AGEMA_reg_buffer_3304 ( .C (clk), .D (new_AGEMA_signal_5259), .Q (new_AGEMA_signal_5260) ) ;
    buf_clk new_AGEMA_reg_buffer_3308 ( .C (clk), .D (new_AGEMA_signal_5263), .Q (new_AGEMA_signal_5264) ) ;
    buf_clk new_AGEMA_reg_buffer_3312 ( .C (clk), .D (new_AGEMA_signal_5267), .Q (new_AGEMA_signal_5268) ) ;
    buf_clk new_AGEMA_reg_buffer_3316 ( .C (clk), .D (new_AGEMA_signal_5271), .Q (new_AGEMA_signal_5272) ) ;
    buf_clk new_AGEMA_reg_buffer_3320 ( .C (clk), .D (new_AGEMA_signal_5275), .Q (new_AGEMA_signal_5276) ) ;
    buf_clk new_AGEMA_reg_buffer_3324 ( .C (clk), .D (new_AGEMA_signal_5279), .Q (new_AGEMA_signal_5280) ) ;
    buf_clk new_AGEMA_reg_buffer_3328 ( .C (clk), .D (new_AGEMA_signal_5283), .Q (new_AGEMA_signal_5284) ) ;
    buf_clk new_AGEMA_reg_buffer_3332 ( .C (clk), .D (new_AGEMA_signal_5287), .Q (new_AGEMA_signal_5288) ) ;
    buf_clk new_AGEMA_reg_buffer_3336 ( .C (clk), .D (new_AGEMA_signal_5291), .Q (new_AGEMA_signal_5292) ) ;
    buf_clk new_AGEMA_reg_buffer_3340 ( .C (clk), .D (new_AGEMA_signal_5295), .Q (new_AGEMA_signal_5296) ) ;
    buf_clk new_AGEMA_reg_buffer_3344 ( .C (clk), .D (new_AGEMA_signal_5299), .Q (new_AGEMA_signal_5300) ) ;
    buf_clk new_AGEMA_reg_buffer_3348 ( .C (clk), .D (new_AGEMA_signal_5303), .Q (new_AGEMA_signal_5304) ) ;
    buf_clk new_AGEMA_reg_buffer_3352 ( .C (clk), .D (new_AGEMA_signal_5307), .Q (new_AGEMA_signal_5308) ) ;
    buf_clk new_AGEMA_reg_buffer_3356 ( .C (clk), .D (new_AGEMA_signal_5311), .Q (new_AGEMA_signal_5312) ) ;
    buf_clk new_AGEMA_reg_buffer_3360 ( .C (clk), .D (new_AGEMA_signal_5315), .Q (new_AGEMA_signal_5316) ) ;
    buf_clk new_AGEMA_reg_buffer_3364 ( .C (clk), .D (new_AGEMA_signal_5319), .Q (new_AGEMA_signal_5320) ) ;
    buf_clk new_AGEMA_reg_buffer_3368 ( .C (clk), .D (new_AGEMA_signal_5323), .Q (new_AGEMA_signal_5324) ) ;
    buf_clk new_AGEMA_reg_buffer_3372 ( .C (clk), .D (new_AGEMA_signal_5327), .Q (new_AGEMA_signal_5328) ) ;
    buf_clk new_AGEMA_reg_buffer_3376 ( .C (clk), .D (new_AGEMA_signal_5331), .Q (new_AGEMA_signal_5332) ) ;
    buf_clk new_AGEMA_reg_buffer_3380 ( .C (clk), .D (new_AGEMA_signal_5335), .Q (new_AGEMA_signal_5336) ) ;
    buf_clk new_AGEMA_reg_buffer_3384 ( .C (clk), .D (new_AGEMA_signal_5339), .Q (new_AGEMA_signal_5340) ) ;
    buf_clk new_AGEMA_reg_buffer_3388 ( .C (clk), .D (new_AGEMA_signal_5343), .Q (new_AGEMA_signal_5344) ) ;
    buf_clk new_AGEMA_reg_buffer_3392 ( .C (clk), .D (new_AGEMA_signal_5347), .Q (new_AGEMA_signal_5348) ) ;
    buf_clk new_AGEMA_reg_buffer_3396 ( .C (clk), .D (new_AGEMA_signal_5351), .Q (new_AGEMA_signal_5352) ) ;
    buf_clk new_AGEMA_reg_buffer_3400 ( .C (clk), .D (new_AGEMA_signal_5355), .Q (new_AGEMA_signal_5356) ) ;
    buf_clk new_AGEMA_reg_buffer_3404 ( .C (clk), .D (new_AGEMA_signal_5359), .Q (new_AGEMA_signal_5360) ) ;
    buf_clk new_AGEMA_reg_buffer_3408 ( .C (clk), .D (new_AGEMA_signal_5363), .Q (new_AGEMA_signal_5364) ) ;
    buf_clk new_AGEMA_reg_buffer_3412 ( .C (clk), .D (new_AGEMA_signal_5367), .Q (new_AGEMA_signal_5368) ) ;
    buf_clk new_AGEMA_reg_buffer_3416 ( .C (clk), .D (new_AGEMA_signal_5371), .Q (new_AGEMA_signal_5372) ) ;
    buf_clk new_AGEMA_reg_buffer_3420 ( .C (clk), .D (new_AGEMA_signal_5375), .Q (new_AGEMA_signal_5376) ) ;
    buf_clk new_AGEMA_reg_buffer_3424 ( .C (clk), .D (new_AGEMA_signal_5379), .Q (new_AGEMA_signal_5380) ) ;
    buf_clk new_AGEMA_reg_buffer_3428 ( .C (clk), .D (new_AGEMA_signal_5383), .Q (new_AGEMA_signal_5384) ) ;
    buf_clk new_AGEMA_reg_buffer_3432 ( .C (clk), .D (new_AGEMA_signal_5387), .Q (new_AGEMA_signal_5388) ) ;
    buf_clk new_AGEMA_reg_buffer_3436 ( .C (clk), .D (new_AGEMA_signal_5391), .Q (new_AGEMA_signal_5392) ) ;
    buf_clk new_AGEMA_reg_buffer_3440 ( .C (clk), .D (new_AGEMA_signal_5395), .Q (new_AGEMA_signal_5396) ) ;
    buf_clk new_AGEMA_reg_buffer_3444 ( .C (clk), .D (new_AGEMA_signal_5399), .Q (new_AGEMA_signal_5400) ) ;
    buf_clk new_AGEMA_reg_buffer_3448 ( .C (clk), .D (new_AGEMA_signal_5403), .Q (new_AGEMA_signal_5404) ) ;
    buf_clk new_AGEMA_reg_buffer_3452 ( .C (clk), .D (new_AGEMA_signal_5407), .Q (new_AGEMA_signal_5408) ) ;
    buf_clk new_AGEMA_reg_buffer_3456 ( .C (clk), .D (new_AGEMA_signal_5411), .Q (new_AGEMA_signal_5412) ) ;
    buf_clk new_AGEMA_reg_buffer_3460 ( .C (clk), .D (new_AGEMA_signal_5415), .Q (new_AGEMA_signal_5416) ) ;
    buf_clk new_AGEMA_reg_buffer_3464 ( .C (clk), .D (new_AGEMA_signal_5419), .Q (new_AGEMA_signal_5420) ) ;
    buf_clk new_AGEMA_reg_buffer_3468 ( .C (clk), .D (new_AGEMA_signal_5423), .Q (new_AGEMA_signal_5424) ) ;
    buf_clk new_AGEMA_reg_buffer_3472 ( .C (clk), .D (new_AGEMA_signal_5427), .Q (new_AGEMA_signal_5428) ) ;
    buf_clk new_AGEMA_reg_buffer_3476 ( .C (clk), .D (new_AGEMA_signal_5431), .Q (new_AGEMA_signal_5432) ) ;
    buf_clk new_AGEMA_reg_buffer_3480 ( .C (clk), .D (new_AGEMA_signal_5435), .Q (new_AGEMA_signal_5436) ) ;
    buf_clk new_AGEMA_reg_buffer_3484 ( .C (clk), .D (new_AGEMA_signal_5439), .Q (new_AGEMA_signal_5440) ) ;
    buf_clk new_AGEMA_reg_buffer_3488 ( .C (clk), .D (new_AGEMA_signal_5443), .Q (new_AGEMA_signal_5444) ) ;
    buf_clk new_AGEMA_reg_buffer_3492 ( .C (clk), .D (new_AGEMA_signal_5447), .Q (new_AGEMA_signal_5448) ) ;
    buf_clk new_AGEMA_reg_buffer_3496 ( .C (clk), .D (new_AGEMA_signal_5451), .Q (new_AGEMA_signal_5452) ) ;
    buf_clk new_AGEMA_reg_buffer_3500 ( .C (clk), .D (new_AGEMA_signal_5455), .Q (new_AGEMA_signal_5456) ) ;
    buf_clk new_AGEMA_reg_buffer_3504 ( .C (clk), .D (new_AGEMA_signal_5459), .Q (new_AGEMA_signal_5460) ) ;
    buf_clk new_AGEMA_reg_buffer_3508 ( .C (clk), .D (new_AGEMA_signal_5463), .Q (new_AGEMA_signal_5464) ) ;
    buf_clk new_AGEMA_reg_buffer_3512 ( .C (clk), .D (new_AGEMA_signal_5467), .Q (new_AGEMA_signal_5468) ) ;
    buf_clk new_AGEMA_reg_buffer_3516 ( .C (clk), .D (new_AGEMA_signal_5471), .Q (new_AGEMA_signal_5472) ) ;
    buf_clk new_AGEMA_reg_buffer_3520 ( .C (clk), .D (new_AGEMA_signal_5475), .Q (new_AGEMA_signal_5476) ) ;
    buf_clk new_AGEMA_reg_buffer_3524 ( .C (clk), .D (new_AGEMA_signal_5479), .Q (new_AGEMA_signal_5480) ) ;
    buf_clk new_AGEMA_reg_buffer_3528 ( .C (clk), .D (new_AGEMA_signal_5483), .Q (new_AGEMA_signal_5484) ) ;
    buf_clk new_AGEMA_reg_buffer_3532 ( .C (clk), .D (new_AGEMA_signal_5487), .Q (new_AGEMA_signal_5488) ) ;
    buf_clk new_AGEMA_reg_buffer_3536 ( .C (clk), .D (new_AGEMA_signal_5491), .Q (new_AGEMA_signal_5492) ) ;
    buf_clk new_AGEMA_reg_buffer_3540 ( .C (clk), .D (new_AGEMA_signal_5495), .Q (new_AGEMA_signal_5496) ) ;
    buf_clk new_AGEMA_reg_buffer_3544 ( .C (clk), .D (new_AGEMA_signal_5499), .Q (new_AGEMA_signal_5500) ) ;
    buf_clk new_AGEMA_reg_buffer_3548 ( .C (clk), .D (new_AGEMA_signal_5503), .Q (new_AGEMA_signal_5504) ) ;
    buf_clk new_AGEMA_reg_buffer_3552 ( .C (clk), .D (new_AGEMA_signal_5507), .Q (new_AGEMA_signal_5508) ) ;
    buf_clk new_AGEMA_reg_buffer_3556 ( .C (clk), .D (new_AGEMA_signal_5511), .Q (new_AGEMA_signal_5512) ) ;
    buf_clk new_AGEMA_reg_buffer_3560 ( .C (clk), .D (new_AGEMA_signal_5515), .Q (new_AGEMA_signal_5516) ) ;
    buf_clk new_AGEMA_reg_buffer_3564 ( .C (clk), .D (new_AGEMA_signal_5519), .Q (new_AGEMA_signal_5520) ) ;
    buf_clk new_AGEMA_reg_buffer_3568 ( .C (clk), .D (new_AGEMA_signal_5523), .Q (new_AGEMA_signal_5524) ) ;
    buf_clk new_AGEMA_reg_buffer_3572 ( .C (clk), .D (new_AGEMA_signal_5527), .Q (new_AGEMA_signal_5528) ) ;
    buf_clk new_AGEMA_reg_buffer_3576 ( .C (clk), .D (new_AGEMA_signal_5531), .Q (new_AGEMA_signal_5532) ) ;
    buf_clk new_AGEMA_reg_buffer_3580 ( .C (clk), .D (new_AGEMA_signal_5535), .Q (new_AGEMA_signal_5536) ) ;
    buf_clk new_AGEMA_reg_buffer_3584 ( .C (clk), .D (new_AGEMA_signal_5539), .Q (new_AGEMA_signal_5540) ) ;
    buf_clk new_AGEMA_reg_buffer_3588 ( .C (clk), .D (new_AGEMA_signal_5543), .Q (new_AGEMA_signal_5544) ) ;
    buf_clk new_AGEMA_reg_buffer_3592 ( .C (clk), .D (new_AGEMA_signal_5547), .Q (new_AGEMA_signal_5548) ) ;
    buf_clk new_AGEMA_reg_buffer_3596 ( .C (clk), .D (new_AGEMA_signal_5551), .Q (new_AGEMA_signal_5552) ) ;
    buf_clk new_AGEMA_reg_buffer_3600 ( .C (clk), .D (new_AGEMA_signal_5555), .Q (new_AGEMA_signal_5556) ) ;
    buf_clk new_AGEMA_reg_buffer_3604 ( .C (clk), .D (new_AGEMA_signal_5559), .Q (new_AGEMA_signal_5560) ) ;
    buf_clk new_AGEMA_reg_buffer_3608 ( .C (clk), .D (new_AGEMA_signal_5563), .Q (new_AGEMA_signal_5564) ) ;
    buf_clk new_AGEMA_reg_buffer_3612 ( .C (clk), .D (new_AGEMA_signal_5567), .Q (new_AGEMA_signal_5568) ) ;
    buf_clk new_AGEMA_reg_buffer_3616 ( .C (clk), .D (new_AGEMA_signal_5571), .Q (new_AGEMA_signal_5572) ) ;
    buf_clk new_AGEMA_reg_buffer_3620 ( .C (clk), .D (new_AGEMA_signal_5575), .Q (new_AGEMA_signal_5576) ) ;
    buf_clk new_AGEMA_reg_buffer_3624 ( .C (clk), .D (new_AGEMA_signal_5579), .Q (new_AGEMA_signal_5580) ) ;
    buf_clk new_AGEMA_reg_buffer_3628 ( .C (clk), .D (new_AGEMA_signal_5583), .Q (new_AGEMA_signal_5584) ) ;
    buf_clk new_AGEMA_reg_buffer_3632 ( .C (clk), .D (new_AGEMA_signal_5587), .Q (new_AGEMA_signal_5588) ) ;
    buf_clk new_AGEMA_reg_buffer_3636 ( .C (clk), .D (new_AGEMA_signal_5591), .Q (new_AGEMA_signal_5592) ) ;
    buf_clk new_AGEMA_reg_buffer_3640 ( .C (clk), .D (new_AGEMA_signal_5595), .Q (new_AGEMA_signal_5596) ) ;
    buf_clk new_AGEMA_reg_buffer_3644 ( .C (clk), .D (new_AGEMA_signal_5599), .Q (new_AGEMA_signal_5600) ) ;
    buf_clk new_AGEMA_reg_buffer_3648 ( .C (clk), .D (new_AGEMA_signal_5603), .Q (new_AGEMA_signal_5604) ) ;
    buf_clk new_AGEMA_reg_buffer_3652 ( .C (clk), .D (new_AGEMA_signal_5607), .Q (new_AGEMA_signal_5608) ) ;
    buf_clk new_AGEMA_reg_buffer_3656 ( .C (clk), .D (new_AGEMA_signal_5611), .Q (new_AGEMA_signal_5612) ) ;
    buf_clk new_AGEMA_reg_buffer_3660 ( .C (clk), .D (new_AGEMA_signal_5615), .Q (new_AGEMA_signal_5616) ) ;
    buf_clk new_AGEMA_reg_buffer_3664 ( .C (clk), .D (new_AGEMA_signal_5619), .Q (new_AGEMA_signal_5620) ) ;
    buf_clk new_AGEMA_reg_buffer_3668 ( .C (clk), .D (new_AGEMA_signal_5623), .Q (new_AGEMA_signal_5624) ) ;
    buf_clk new_AGEMA_reg_buffer_3672 ( .C (clk), .D (new_AGEMA_signal_5627), .Q (new_AGEMA_signal_5628) ) ;
    buf_clk new_AGEMA_reg_buffer_3676 ( .C (clk), .D (new_AGEMA_signal_5631), .Q (new_AGEMA_signal_5632) ) ;
    buf_clk new_AGEMA_reg_buffer_3680 ( .C (clk), .D (new_AGEMA_signal_5635), .Q (new_AGEMA_signal_5636) ) ;
    buf_clk new_AGEMA_reg_buffer_3684 ( .C (clk), .D (new_AGEMA_signal_5639), .Q (new_AGEMA_signal_5640) ) ;
    buf_clk new_AGEMA_reg_buffer_3688 ( .C (clk), .D (new_AGEMA_signal_5643), .Q (new_AGEMA_signal_5644) ) ;
    buf_clk new_AGEMA_reg_buffer_3692 ( .C (clk), .D (new_AGEMA_signal_5647), .Q (new_AGEMA_signal_5648) ) ;
    buf_clk new_AGEMA_reg_buffer_3696 ( .C (clk), .D (new_AGEMA_signal_5651), .Q (new_AGEMA_signal_5652) ) ;
    buf_clk new_AGEMA_reg_buffer_3700 ( .C (clk), .D (new_AGEMA_signal_5655), .Q (new_AGEMA_signal_5656) ) ;
    buf_clk new_AGEMA_reg_buffer_3704 ( .C (clk), .D (new_AGEMA_signal_5659), .Q (new_AGEMA_signal_5660) ) ;
    buf_clk new_AGEMA_reg_buffer_3708 ( .C (clk), .D (new_AGEMA_signal_5663), .Q (new_AGEMA_signal_5664) ) ;
    buf_clk new_AGEMA_reg_buffer_3712 ( .C (clk), .D (new_AGEMA_signal_5667), .Q (new_AGEMA_signal_5668) ) ;
    buf_clk new_AGEMA_reg_buffer_3716 ( .C (clk), .D (new_AGEMA_signal_5671), .Q (new_AGEMA_signal_5672) ) ;
    buf_clk new_AGEMA_reg_buffer_3720 ( .C (clk), .D (new_AGEMA_signal_5675), .Q (new_AGEMA_signal_5676) ) ;
    buf_clk new_AGEMA_reg_buffer_3724 ( .C (clk), .D (new_AGEMA_signal_5679), .Q (new_AGEMA_signal_5680) ) ;
    buf_clk new_AGEMA_reg_buffer_3728 ( .C (clk), .D (new_AGEMA_signal_5683), .Q (new_AGEMA_signal_5684) ) ;
    buf_clk new_AGEMA_reg_buffer_3732 ( .C (clk), .D (new_AGEMA_signal_5687), .Q (new_AGEMA_signal_5688) ) ;
    buf_clk new_AGEMA_reg_buffer_3736 ( .C (clk), .D (new_AGEMA_signal_5691), .Q (new_AGEMA_signal_5692) ) ;
    buf_clk new_AGEMA_reg_buffer_3740 ( .C (clk), .D (new_AGEMA_signal_5695), .Q (new_AGEMA_signal_5696) ) ;
    buf_clk new_AGEMA_reg_buffer_3744 ( .C (clk), .D (new_AGEMA_signal_5699), .Q (new_AGEMA_signal_5700) ) ;
    buf_clk new_AGEMA_reg_buffer_3748 ( .C (clk), .D (new_AGEMA_signal_5703), .Q (new_AGEMA_signal_5704) ) ;
    buf_clk new_AGEMA_reg_buffer_3752 ( .C (clk), .D (new_AGEMA_signal_5707), .Q (new_AGEMA_signal_5708) ) ;
    buf_clk new_AGEMA_reg_buffer_3756 ( .C (clk), .D (new_AGEMA_signal_5711), .Q (new_AGEMA_signal_5712) ) ;
    buf_clk new_AGEMA_reg_buffer_3760 ( .C (clk), .D (new_AGEMA_signal_5715), .Q (new_AGEMA_signal_5716) ) ;
    buf_clk new_AGEMA_reg_buffer_3764 ( .C (clk), .D (new_AGEMA_signal_5719), .Q (new_AGEMA_signal_5720) ) ;
    buf_clk new_AGEMA_reg_buffer_3768 ( .C (clk), .D (new_AGEMA_signal_5723), .Q (new_AGEMA_signal_5724) ) ;
    buf_clk new_AGEMA_reg_buffer_3772 ( .C (clk), .D (new_AGEMA_signal_5727), .Q (new_AGEMA_signal_5728) ) ;
    buf_clk new_AGEMA_reg_buffer_3776 ( .C (clk), .D (new_AGEMA_signal_5731), .Q (new_AGEMA_signal_5732) ) ;
    buf_clk new_AGEMA_reg_buffer_3780 ( .C (clk), .D (new_AGEMA_signal_5735), .Q (new_AGEMA_signal_5736) ) ;
    buf_clk new_AGEMA_reg_buffer_3784 ( .C (clk), .D (new_AGEMA_signal_5739), .Q (new_AGEMA_signal_5740) ) ;
    buf_clk new_AGEMA_reg_buffer_3788 ( .C (clk), .D (new_AGEMA_signal_5743), .Q (new_AGEMA_signal_5744) ) ;
    buf_clk new_AGEMA_reg_buffer_3792 ( .C (clk), .D (new_AGEMA_signal_5747), .Q (new_AGEMA_signal_5748) ) ;
    buf_clk new_AGEMA_reg_buffer_3796 ( .C (clk), .D (new_AGEMA_signal_5751), .Q (new_AGEMA_signal_5752) ) ;
    buf_clk new_AGEMA_reg_buffer_3800 ( .C (clk), .D (new_AGEMA_signal_5755), .Q (new_AGEMA_signal_5756) ) ;
    buf_clk new_AGEMA_reg_buffer_3804 ( .C (clk), .D (new_AGEMA_signal_5759), .Q (new_AGEMA_signal_5760) ) ;
    buf_clk new_AGEMA_reg_buffer_3808 ( .C (clk), .D (new_AGEMA_signal_5763), .Q (new_AGEMA_signal_5764) ) ;
    buf_clk new_AGEMA_reg_buffer_3812 ( .C (clk), .D (new_AGEMA_signal_5767), .Q (new_AGEMA_signal_5768) ) ;
    buf_clk new_AGEMA_reg_buffer_3816 ( .C (clk), .D (new_AGEMA_signal_5771), .Q (new_AGEMA_signal_5772) ) ;
    buf_clk new_AGEMA_reg_buffer_3820 ( .C (clk), .D (new_AGEMA_signal_5775), .Q (new_AGEMA_signal_5776) ) ;
    buf_clk new_AGEMA_reg_buffer_3824 ( .C (clk), .D (new_AGEMA_signal_5779), .Q (new_AGEMA_signal_5780) ) ;
    buf_clk new_AGEMA_reg_buffer_3828 ( .C (clk), .D (new_AGEMA_signal_5783), .Q (new_AGEMA_signal_5784) ) ;
    buf_clk new_AGEMA_reg_buffer_3832 ( .C (clk), .D (new_AGEMA_signal_5787), .Q (new_AGEMA_signal_5788) ) ;
    buf_clk new_AGEMA_reg_buffer_3836 ( .C (clk), .D (new_AGEMA_signal_5791), .Q (new_AGEMA_signal_5792) ) ;
    buf_clk new_AGEMA_reg_buffer_3840 ( .C (clk), .D (new_AGEMA_signal_5795), .Q (new_AGEMA_signal_5796) ) ;
    buf_clk new_AGEMA_reg_buffer_3844 ( .C (clk), .D (new_AGEMA_signal_5799), .Q (new_AGEMA_signal_5800) ) ;
    buf_clk new_AGEMA_reg_buffer_3848 ( .C (clk), .D (new_AGEMA_signal_5803), .Q (new_AGEMA_signal_5804) ) ;
    buf_clk new_AGEMA_reg_buffer_3852 ( .C (clk), .D (new_AGEMA_signal_5807), .Q (new_AGEMA_signal_5808) ) ;
    buf_clk new_AGEMA_reg_buffer_3856 ( .C (clk), .D (new_AGEMA_signal_5811), .Q (new_AGEMA_signal_5812) ) ;
    buf_clk new_AGEMA_reg_buffer_3860 ( .C (clk), .D (new_AGEMA_signal_5815), .Q (new_AGEMA_signal_5816) ) ;
    buf_clk new_AGEMA_reg_buffer_3864 ( .C (clk), .D (new_AGEMA_signal_5819), .Q (new_AGEMA_signal_5820) ) ;
    buf_clk new_AGEMA_reg_buffer_3868 ( .C (clk), .D (new_AGEMA_signal_5823), .Q (new_AGEMA_signal_5824) ) ;
    buf_clk new_AGEMA_reg_buffer_3872 ( .C (clk), .D (new_AGEMA_signal_5827), .Q (new_AGEMA_signal_5828) ) ;
    buf_clk new_AGEMA_reg_buffer_3876 ( .C (clk), .D (new_AGEMA_signal_5831), .Q (new_AGEMA_signal_5832) ) ;
    buf_clk new_AGEMA_reg_buffer_3880 ( .C (clk), .D (new_AGEMA_signal_5835), .Q (new_AGEMA_signal_5836) ) ;
    buf_clk new_AGEMA_reg_buffer_3884 ( .C (clk), .D (new_AGEMA_signal_5839), .Q (new_AGEMA_signal_5840) ) ;
    buf_clk new_AGEMA_reg_buffer_3888 ( .C (clk), .D (new_AGEMA_signal_5843), .Q (new_AGEMA_signal_5844) ) ;
    buf_clk new_AGEMA_reg_buffer_3892 ( .C (clk), .D (new_AGEMA_signal_5847), .Q (new_AGEMA_signal_5848) ) ;
    buf_clk new_AGEMA_reg_buffer_3896 ( .C (clk), .D (new_AGEMA_signal_5851), .Q (new_AGEMA_signal_5852) ) ;
    buf_clk new_AGEMA_reg_buffer_3900 ( .C (clk), .D (new_AGEMA_signal_5855), .Q (new_AGEMA_signal_5856) ) ;
    buf_clk new_AGEMA_reg_buffer_3904 ( .C (clk), .D (new_AGEMA_signal_5859), .Q (new_AGEMA_signal_5860) ) ;
    buf_clk new_AGEMA_reg_buffer_3908 ( .C (clk), .D (new_AGEMA_signal_5863), .Q (new_AGEMA_signal_5864) ) ;
    buf_clk new_AGEMA_reg_buffer_3912 ( .C (clk), .D (new_AGEMA_signal_5867), .Q (new_AGEMA_signal_5868) ) ;
    buf_clk new_AGEMA_reg_buffer_3916 ( .C (clk), .D (new_AGEMA_signal_5871), .Q (new_AGEMA_signal_5872) ) ;
    buf_clk new_AGEMA_reg_buffer_3920 ( .C (clk), .D (new_AGEMA_signal_5875), .Q (new_AGEMA_signal_5876) ) ;
    buf_clk new_AGEMA_reg_buffer_3924 ( .C (clk), .D (new_AGEMA_signal_5879), .Q (new_AGEMA_signal_5880) ) ;
    buf_clk new_AGEMA_reg_buffer_3928 ( .C (clk), .D (new_AGEMA_signal_5883), .Q (new_AGEMA_signal_5884) ) ;
    buf_clk new_AGEMA_reg_buffer_3932 ( .C (clk), .D (new_AGEMA_signal_5887), .Q (new_AGEMA_signal_5888) ) ;
    buf_clk new_AGEMA_reg_buffer_3936 ( .C (clk), .D (new_AGEMA_signal_5891), .Q (new_AGEMA_signal_5892) ) ;
    buf_clk new_AGEMA_reg_buffer_3940 ( .C (clk), .D (new_AGEMA_signal_5895), .Q (new_AGEMA_signal_5896) ) ;
    buf_clk new_AGEMA_reg_buffer_3944 ( .C (clk), .D (new_AGEMA_signal_5899), .Q (new_AGEMA_signal_5900) ) ;
    buf_clk new_AGEMA_reg_buffer_3948 ( .C (clk), .D (new_AGEMA_signal_5903), .Q (new_AGEMA_signal_5904) ) ;
    buf_clk new_AGEMA_reg_buffer_3952 ( .C (clk), .D (new_AGEMA_signal_5907), .Q (new_AGEMA_signal_5908) ) ;
    buf_clk new_AGEMA_reg_buffer_3956 ( .C (clk), .D (new_AGEMA_signal_5911), .Q (new_AGEMA_signal_5912) ) ;
    buf_clk new_AGEMA_reg_buffer_3960 ( .C (clk), .D (new_AGEMA_signal_5915), .Q (new_AGEMA_signal_5916) ) ;
    buf_clk new_AGEMA_reg_buffer_3964 ( .C (clk), .D (new_AGEMA_signal_5919), .Q (new_AGEMA_signal_5920) ) ;
    buf_clk new_AGEMA_reg_buffer_3968 ( .C (clk), .D (new_AGEMA_signal_5923), .Q (new_AGEMA_signal_5924) ) ;
    buf_clk new_AGEMA_reg_buffer_3972 ( .C (clk), .D (new_AGEMA_signal_5927), .Q (new_AGEMA_signal_5928) ) ;
    buf_clk new_AGEMA_reg_buffer_3976 ( .C (clk), .D (new_AGEMA_signal_5931), .Q (new_AGEMA_signal_5932) ) ;
    buf_clk new_AGEMA_reg_buffer_3980 ( .C (clk), .D (new_AGEMA_signal_5935), .Q (new_AGEMA_signal_5936) ) ;
    buf_clk new_AGEMA_reg_buffer_3984 ( .C (clk), .D (new_AGEMA_signal_5939), .Q (new_AGEMA_signal_5940) ) ;
    buf_clk new_AGEMA_reg_buffer_3988 ( .C (clk), .D (new_AGEMA_signal_5943), .Q (new_AGEMA_signal_5944) ) ;
    buf_clk new_AGEMA_reg_buffer_3992 ( .C (clk), .D (new_AGEMA_signal_5947), .Q (new_AGEMA_signal_5948) ) ;
    buf_clk new_AGEMA_reg_buffer_3996 ( .C (clk), .D (new_AGEMA_signal_5951), .Q (new_AGEMA_signal_5952) ) ;
    buf_clk new_AGEMA_reg_buffer_4000 ( .C (clk), .D (new_AGEMA_signal_5955), .Q (new_AGEMA_signal_5956) ) ;
    buf_clk new_AGEMA_reg_buffer_4004 ( .C (clk), .D (new_AGEMA_signal_5959), .Q (new_AGEMA_signal_5960) ) ;
    buf_clk new_AGEMA_reg_buffer_4008 ( .C (clk), .D (new_AGEMA_signal_5963), .Q (new_AGEMA_signal_5964) ) ;
    buf_clk new_AGEMA_reg_buffer_4012 ( .C (clk), .D (new_AGEMA_signal_5967), .Q (new_AGEMA_signal_5968) ) ;
    buf_clk new_AGEMA_reg_buffer_4016 ( .C (clk), .D (new_AGEMA_signal_5971), .Q (new_AGEMA_signal_5972) ) ;
    buf_clk new_AGEMA_reg_buffer_4020 ( .C (clk), .D (new_AGEMA_signal_5975), .Q (new_AGEMA_signal_5976) ) ;
    buf_clk new_AGEMA_reg_buffer_4024 ( .C (clk), .D (new_AGEMA_signal_5979), .Q (new_AGEMA_signal_5980) ) ;
    buf_clk new_AGEMA_reg_buffer_4028 ( .C (clk), .D (new_AGEMA_signal_5983), .Q (new_AGEMA_signal_5984) ) ;
    buf_clk new_AGEMA_reg_buffer_4032 ( .C (clk), .D (new_AGEMA_signal_5987), .Q (new_AGEMA_signal_5988) ) ;
    buf_clk new_AGEMA_reg_buffer_4036 ( .C (clk), .D (new_AGEMA_signal_5991), .Q (new_AGEMA_signal_5992) ) ;
    buf_clk new_AGEMA_reg_buffer_4040 ( .C (clk), .D (new_AGEMA_signal_5995), .Q (new_AGEMA_signal_5996) ) ;
    buf_clk new_AGEMA_reg_buffer_4044 ( .C (clk), .D (new_AGEMA_signal_5999), .Q (new_AGEMA_signal_6000) ) ;
    buf_clk new_AGEMA_reg_buffer_4048 ( .C (clk), .D (new_AGEMA_signal_6003), .Q (new_AGEMA_signal_6004) ) ;
    buf_clk new_AGEMA_reg_buffer_4052 ( .C (clk), .D (new_AGEMA_signal_6007), .Q (new_AGEMA_signal_6008) ) ;
    buf_clk new_AGEMA_reg_buffer_4056 ( .C (clk), .D (new_AGEMA_signal_6011), .Q (new_AGEMA_signal_6012) ) ;
    buf_clk new_AGEMA_reg_buffer_4060 ( .C (clk), .D (new_AGEMA_signal_6015), .Q (new_AGEMA_signal_6016) ) ;
    buf_clk new_AGEMA_reg_buffer_4064 ( .C (clk), .D (new_AGEMA_signal_6019), .Q (new_AGEMA_signal_6020) ) ;
    buf_clk new_AGEMA_reg_buffer_4068 ( .C (clk), .D (new_AGEMA_signal_6023), .Q (new_AGEMA_signal_6024) ) ;
    buf_clk new_AGEMA_reg_buffer_4072 ( .C (clk), .D (new_AGEMA_signal_6027), .Q (new_AGEMA_signal_6028) ) ;
    buf_clk new_AGEMA_reg_buffer_4076 ( .C (clk), .D (new_AGEMA_signal_6031), .Q (new_AGEMA_signal_6032) ) ;
    buf_clk new_AGEMA_reg_buffer_4080 ( .C (clk), .D (new_AGEMA_signal_6035), .Q (new_AGEMA_signal_6036) ) ;
    buf_clk new_AGEMA_reg_buffer_4084 ( .C (clk), .D (new_AGEMA_signal_6039), .Q (new_AGEMA_signal_6040) ) ;
    buf_clk new_AGEMA_reg_buffer_4088 ( .C (clk), .D (new_AGEMA_signal_6043), .Q (new_AGEMA_signal_6044) ) ;
    buf_clk new_AGEMA_reg_buffer_4092 ( .C (clk), .D (new_AGEMA_signal_6047), .Q (new_AGEMA_signal_6048) ) ;
    buf_clk new_AGEMA_reg_buffer_4096 ( .C (clk), .D (new_AGEMA_signal_6051), .Q (new_AGEMA_signal_6052) ) ;
    buf_clk new_AGEMA_reg_buffer_4100 ( .C (clk), .D (new_AGEMA_signal_6055), .Q (new_AGEMA_signal_6056) ) ;
    buf_clk new_AGEMA_reg_buffer_4104 ( .C (clk), .D (new_AGEMA_signal_6059), .Q (new_AGEMA_signal_6060) ) ;
    buf_clk new_AGEMA_reg_buffer_4108 ( .C (clk), .D (new_AGEMA_signal_6063), .Q (new_AGEMA_signal_6064) ) ;
    buf_clk new_AGEMA_reg_buffer_4112 ( .C (clk), .D (new_AGEMA_signal_6067), .Q (new_AGEMA_signal_6068) ) ;
    buf_clk new_AGEMA_reg_buffer_4116 ( .C (clk), .D (new_AGEMA_signal_6071), .Q (new_AGEMA_signal_6072) ) ;
    buf_clk new_AGEMA_reg_buffer_4120 ( .C (clk), .D (new_AGEMA_signal_6075), .Q (new_AGEMA_signal_6076) ) ;
    buf_clk new_AGEMA_reg_buffer_4124 ( .C (clk), .D (new_AGEMA_signal_6079), .Q (new_AGEMA_signal_6080) ) ;
    buf_clk new_AGEMA_reg_buffer_4128 ( .C (clk), .D (new_AGEMA_signal_6083), .Q (new_AGEMA_signal_6084) ) ;
    buf_clk new_AGEMA_reg_buffer_4132 ( .C (clk), .D (new_AGEMA_signal_6087), .Q (new_AGEMA_signal_6088) ) ;
    buf_clk new_AGEMA_reg_buffer_4136 ( .C (clk), .D (new_AGEMA_signal_6091), .Q (new_AGEMA_signal_6092) ) ;
    buf_clk new_AGEMA_reg_buffer_4140 ( .C (clk), .D (new_AGEMA_signal_6095), .Q (new_AGEMA_signal_6096) ) ;
    buf_clk new_AGEMA_reg_buffer_4144 ( .C (clk), .D (new_AGEMA_signal_6099), .Q (new_AGEMA_signal_6100) ) ;
    buf_clk new_AGEMA_reg_buffer_4148 ( .C (clk), .D (new_AGEMA_signal_6103), .Q (new_AGEMA_signal_6104) ) ;
    buf_clk new_AGEMA_reg_buffer_4152 ( .C (clk), .D (new_AGEMA_signal_6107), .Q (new_AGEMA_signal_6108) ) ;
    buf_clk new_AGEMA_reg_buffer_4156 ( .C (clk), .D (new_AGEMA_signal_6111), .Q (new_AGEMA_signal_6112) ) ;
    buf_clk new_AGEMA_reg_buffer_4160 ( .C (clk), .D (new_AGEMA_signal_6115), .Q (new_AGEMA_signal_6116) ) ;
    buf_clk new_AGEMA_reg_buffer_4164 ( .C (clk), .D (new_AGEMA_signal_6119), .Q (new_AGEMA_signal_6120) ) ;
    buf_clk new_AGEMA_reg_buffer_4168 ( .C (clk), .D (new_AGEMA_signal_6123), .Q (new_AGEMA_signal_6124) ) ;
    buf_clk new_AGEMA_reg_buffer_4172 ( .C (clk), .D (new_AGEMA_signal_6127), .Q (new_AGEMA_signal_6128) ) ;
    buf_clk new_AGEMA_reg_buffer_4176 ( .C (clk), .D (new_AGEMA_signal_6131), .Q (new_AGEMA_signal_6132) ) ;
    buf_clk new_AGEMA_reg_buffer_4180 ( .C (clk), .D (new_AGEMA_signal_6135), .Q (new_AGEMA_signal_6136) ) ;
    buf_clk new_AGEMA_reg_buffer_4184 ( .C (clk), .D (new_AGEMA_signal_6139), .Q (new_AGEMA_signal_6140) ) ;
    buf_clk new_AGEMA_reg_buffer_4188 ( .C (clk), .D (new_AGEMA_signal_6143), .Q (new_AGEMA_signal_6144) ) ;
    buf_clk new_AGEMA_reg_buffer_4192 ( .C (clk), .D (new_AGEMA_signal_6147), .Q (new_AGEMA_signal_6148) ) ;
    buf_clk new_AGEMA_reg_buffer_4196 ( .C (clk), .D (new_AGEMA_signal_6151), .Q (new_AGEMA_signal_6152) ) ;
    buf_clk new_AGEMA_reg_buffer_4200 ( .C (clk), .D (new_AGEMA_signal_6155), .Q (new_AGEMA_signal_6156) ) ;
    buf_clk new_AGEMA_reg_buffer_4204 ( .C (clk), .D (new_AGEMA_signal_6159), .Q (new_AGEMA_signal_6160) ) ;
    buf_clk new_AGEMA_reg_buffer_4208 ( .C (clk), .D (new_AGEMA_signal_6163), .Q (new_AGEMA_signal_6164) ) ;
    buf_clk new_AGEMA_reg_buffer_4212 ( .C (clk), .D (new_AGEMA_signal_6167), .Q (new_AGEMA_signal_6168) ) ;
    buf_clk new_AGEMA_reg_buffer_4216 ( .C (clk), .D (new_AGEMA_signal_6171), .Q (new_AGEMA_signal_6172) ) ;
    buf_clk new_AGEMA_reg_buffer_4220 ( .C (clk), .D (new_AGEMA_signal_6175), .Q (new_AGEMA_signal_6176) ) ;
    buf_clk new_AGEMA_reg_buffer_4224 ( .C (clk), .D (new_AGEMA_signal_6179), .Q (new_AGEMA_signal_6180) ) ;
    buf_clk new_AGEMA_reg_buffer_4228 ( .C (clk), .D (new_AGEMA_signal_6183), .Q (new_AGEMA_signal_6184) ) ;
    buf_clk new_AGEMA_reg_buffer_4232 ( .C (clk), .D (new_AGEMA_signal_6187), .Q (new_AGEMA_signal_6188) ) ;
    buf_clk new_AGEMA_reg_buffer_4236 ( .C (clk), .D (new_AGEMA_signal_6191), .Q (new_AGEMA_signal_6192) ) ;
    buf_clk new_AGEMA_reg_buffer_4240 ( .C (clk), .D (new_AGEMA_signal_6195), .Q (new_AGEMA_signal_6196) ) ;
    buf_clk new_AGEMA_reg_buffer_4244 ( .C (clk), .D (new_AGEMA_signal_6199), .Q (new_AGEMA_signal_6200) ) ;
    buf_clk new_AGEMA_reg_buffer_4248 ( .C (clk), .D (new_AGEMA_signal_6203), .Q (new_AGEMA_signal_6204) ) ;
    buf_clk new_AGEMA_reg_buffer_4252 ( .C (clk), .D (new_AGEMA_signal_6207), .Q (new_AGEMA_signal_6208) ) ;
    buf_clk new_AGEMA_reg_buffer_4256 ( .C (clk), .D (new_AGEMA_signal_6211), .Q (new_AGEMA_signal_6212) ) ;
    buf_clk new_AGEMA_reg_buffer_4260 ( .C (clk), .D (new_AGEMA_signal_6215), .Q (new_AGEMA_signal_6216) ) ;
    buf_clk new_AGEMA_reg_buffer_4264 ( .C (clk), .D (new_AGEMA_signal_6219), .Q (new_AGEMA_signal_6220) ) ;
    buf_clk new_AGEMA_reg_buffer_4268 ( .C (clk), .D (new_AGEMA_signal_6223), .Q (new_AGEMA_signal_6224) ) ;
    buf_clk new_AGEMA_reg_buffer_4272 ( .C (clk), .D (new_AGEMA_signal_6227), .Q (new_AGEMA_signal_6228) ) ;
    buf_clk new_AGEMA_reg_buffer_4276 ( .C (clk), .D (new_AGEMA_signal_6231), .Q (new_AGEMA_signal_6232) ) ;
    buf_clk new_AGEMA_reg_buffer_4280 ( .C (clk), .D (new_AGEMA_signal_6235), .Q (new_AGEMA_signal_6236) ) ;
    buf_clk new_AGEMA_reg_buffer_4284 ( .C (clk), .D (new_AGEMA_signal_6239), .Q (new_AGEMA_signal_6240) ) ;
    buf_clk new_AGEMA_reg_buffer_4288 ( .C (clk), .D (new_AGEMA_signal_6243), .Q (new_AGEMA_signal_6244) ) ;
    buf_clk new_AGEMA_reg_buffer_4292 ( .C (clk), .D (new_AGEMA_signal_6247), .Q (new_AGEMA_signal_6248) ) ;
    buf_clk new_AGEMA_reg_buffer_4296 ( .C (clk), .D (new_AGEMA_signal_6251), .Q (new_AGEMA_signal_6252) ) ;
    buf_clk new_AGEMA_reg_buffer_4300 ( .C (clk), .D (new_AGEMA_signal_6255), .Q (new_AGEMA_signal_6256) ) ;
    buf_clk new_AGEMA_reg_buffer_4304 ( .C (clk), .D (new_AGEMA_signal_6259), .Q (new_AGEMA_signal_6260) ) ;
    buf_clk new_AGEMA_reg_buffer_4308 ( .C (clk), .D (new_AGEMA_signal_6263), .Q (new_AGEMA_signal_6264) ) ;
    buf_clk new_AGEMA_reg_buffer_4312 ( .C (clk), .D (new_AGEMA_signal_6267), .Q (new_AGEMA_signal_6268) ) ;
    buf_clk new_AGEMA_reg_buffer_4316 ( .C (clk), .D (new_AGEMA_signal_6271), .Q (new_AGEMA_signal_6272) ) ;
    buf_clk new_AGEMA_reg_buffer_4320 ( .C (clk), .D (new_AGEMA_signal_6275), .Q (new_AGEMA_signal_6276) ) ;
    buf_clk new_AGEMA_reg_buffer_4324 ( .C (clk), .D (new_AGEMA_signal_6279), .Q (new_AGEMA_signal_6280) ) ;
    buf_clk new_AGEMA_reg_buffer_4328 ( .C (clk), .D (new_AGEMA_signal_6283), .Q (new_AGEMA_signal_6284) ) ;
    buf_clk new_AGEMA_reg_buffer_4332 ( .C (clk), .D (new_AGEMA_signal_6287), .Q (new_AGEMA_signal_6288) ) ;
    buf_clk new_AGEMA_reg_buffer_4336 ( .C (clk), .D (new_AGEMA_signal_6291), .Q (new_AGEMA_signal_6292) ) ;
    buf_clk new_AGEMA_reg_buffer_4340 ( .C (clk), .D (new_AGEMA_signal_6295), .Q (new_AGEMA_signal_6296) ) ;

    /* cells in depth 4 */
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateIn_mux_inst_0_U1 ( .s (new_AGEMA_signal_3697), .b ({new_AGEMA_signal_3454, SboxOut[0]}), .a ({new_AGEMA_signal_3705, new_AGEMA_signal_3701}), .c ({new_AGEMA_signal_3455, StateIn[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateIn_mux_inst_1_U1 ( .s (new_AGEMA_signal_3697), .b ({new_AGEMA_signal_3463, SboxOut[1]}), .a ({new_AGEMA_signal_3713, new_AGEMA_signal_3709}), .c ({new_AGEMA_signal_3464, StateIn[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateIn_mux_inst_2_U1 ( .s (new_AGEMA_signal_3697), .b ({new_AGEMA_signal_3462, SboxOut[2]}), .a ({new_AGEMA_signal_3721, new_AGEMA_signal_3717}), .c ({new_AGEMA_signal_3465, StateIn[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateIn_mux_inst_3_U1 ( .s (new_AGEMA_signal_3697), .b ({new_AGEMA_signal_3461, SboxOut[3]}), .a ({new_AGEMA_signal_3729, new_AGEMA_signal_3725}), .c ({new_AGEMA_signal_3466, StateIn[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateIn_mux_inst_4_U1 ( .s (new_AGEMA_signal_3697), .b ({new_AGEMA_signal_3460, SboxOut[4]}), .a ({new_AGEMA_signal_3737, new_AGEMA_signal_3733}), .c ({new_AGEMA_signal_3467, StateIn[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateIn_mux_inst_5_U1 ( .s (new_AGEMA_signal_3697), .b ({new_AGEMA_signal_3459, SboxOut[5]}), .a ({new_AGEMA_signal_3745, new_AGEMA_signal_3741}), .c ({new_AGEMA_signal_3468, StateIn[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateIn_mux_inst_6_U1 ( .s (new_AGEMA_signal_3697), .b ({new_AGEMA_signal_3458, SboxOut[6]}), .a ({new_AGEMA_signal_3753, new_AGEMA_signal_3749}), .c ({new_AGEMA_signal_3469, StateIn[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) MUX_StateIn_mux_inst_7_U1 ( .s (new_AGEMA_signal_3697), .b ({new_AGEMA_signal_3457, SboxOut[7]}), .a ({new_AGEMA_signal_3761, new_AGEMA_signal_3757}), .c ({new_AGEMA_signal_3470, StateIn[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S33reg_gff_1_SFF_0_MUXInst_U1 ( .s (new_AGEMA_signal_3765), .b ({new_AGEMA_signal_3488, stateArray_inS33ser[0]}), .a ({new_AGEMA_signal_3773, new_AGEMA_signal_3769}), .c ({new_AGEMA_signal_3497, stateArray_S33reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S33reg_gff_1_SFF_1_MUXInst_U1 ( .s (new_AGEMA_signal_3765), .b ({new_AGEMA_signal_3499, stateArray_inS33ser[1]}), .a ({new_AGEMA_signal_3781, new_AGEMA_signal_3777}), .c ({new_AGEMA_signal_3520, stateArray_S33reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S33reg_gff_1_SFF_2_MUXInst_U1 ( .s (new_AGEMA_signal_3765), .b ({new_AGEMA_signal_3501, stateArray_inS33ser[2]}), .a ({new_AGEMA_signal_3789, new_AGEMA_signal_3785}), .c ({new_AGEMA_signal_3521, stateArray_S33reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S33reg_gff_1_SFF_3_MUXInst_U1 ( .s (new_AGEMA_signal_3765), .b ({new_AGEMA_signal_3503, stateArray_inS33ser[3]}), .a ({new_AGEMA_signal_3797, new_AGEMA_signal_3793}), .c ({new_AGEMA_signal_3522, stateArray_S33reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S33reg_gff_1_SFF_4_MUXInst_U1 ( .s (new_AGEMA_signal_3765), .b ({new_AGEMA_signal_3505, stateArray_inS33ser[4]}), .a ({new_AGEMA_signal_3805, new_AGEMA_signal_3801}), .c ({new_AGEMA_signal_3523, stateArray_S33reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S33reg_gff_1_SFF_5_MUXInst_U1 ( .s (new_AGEMA_signal_3765), .b ({new_AGEMA_signal_3507, stateArray_inS33ser[5]}), .a ({new_AGEMA_signal_3813, new_AGEMA_signal_3809}), .c ({new_AGEMA_signal_3524, stateArray_S33reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S33reg_gff_1_SFF_6_MUXInst_U1 ( .s (new_AGEMA_signal_3765), .b ({new_AGEMA_signal_3509, stateArray_inS33ser[6]}), .a ({new_AGEMA_signal_3821, new_AGEMA_signal_3817}), .c ({new_AGEMA_signal_3525, stateArray_S33reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_S33reg_gff_1_SFF_7_MUXInst_U1 ( .s (new_AGEMA_signal_3765), .b ({new_AGEMA_signal_3511, stateArray_inS33ser[7]}), .a ({new_AGEMA_signal_3829, new_AGEMA_signal_3825}), .c ({new_AGEMA_signal_3526, stateArray_S33reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_input_MC_mux_inst_0_U1 ( .s (new_AGEMA_signal_3833), .b ({new_AGEMA_signal_3455, StateIn[0]}), .a ({new_AGEMA_signal_3841, new_AGEMA_signal_3837}), .c ({new_AGEMA_signal_3471, stateArray_input_MC[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_input_MC_mux_inst_1_U1 ( .s (new_AGEMA_signal_3833), .b ({new_AGEMA_signal_3464, StateIn[1]}), .a ({new_AGEMA_signal_3849, new_AGEMA_signal_3845}), .c ({new_AGEMA_signal_3480, stateArray_input_MC[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_input_MC_mux_inst_2_U1 ( .s (new_AGEMA_signal_3833), .b ({new_AGEMA_signal_3465, StateIn[2]}), .a ({new_AGEMA_signal_3857, new_AGEMA_signal_3853}), .c ({new_AGEMA_signal_3481, stateArray_input_MC[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_input_MC_mux_inst_3_U1 ( .s (new_AGEMA_signal_3833), .b ({new_AGEMA_signal_3466, StateIn[3]}), .a ({new_AGEMA_signal_3865, new_AGEMA_signal_3861}), .c ({new_AGEMA_signal_3482, stateArray_input_MC[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_input_MC_mux_inst_4_U1 ( .s (new_AGEMA_signal_3833), .b ({new_AGEMA_signal_3467, StateIn[4]}), .a ({new_AGEMA_signal_3873, new_AGEMA_signal_3869}), .c ({new_AGEMA_signal_3483, stateArray_input_MC[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_input_MC_mux_inst_5_U1 ( .s (new_AGEMA_signal_3833), .b ({new_AGEMA_signal_3468, StateIn[5]}), .a ({new_AGEMA_signal_3881, new_AGEMA_signal_3877}), .c ({new_AGEMA_signal_3484, stateArray_input_MC[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_input_MC_mux_inst_6_U1 ( .s (new_AGEMA_signal_3833), .b ({new_AGEMA_signal_3469, StateIn[6]}), .a ({new_AGEMA_signal_3889, new_AGEMA_signal_3885}), .c ({new_AGEMA_signal_3485, stateArray_input_MC[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_input_MC_mux_inst_7_U1 ( .s (new_AGEMA_signal_3833), .b ({new_AGEMA_signal_3470, StateIn[7]}), .a ({new_AGEMA_signal_3897, new_AGEMA_signal_3893}), .c ({new_AGEMA_signal_3486, stateArray_input_MC[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS33ser_mux_inst_0_U1 ( .s (new_AGEMA_signal_3901), .b ({new_AGEMA_signal_3909, new_AGEMA_signal_3905}), .a ({new_AGEMA_signal_3471, stateArray_input_MC[0]}), .c ({new_AGEMA_signal_3488, stateArray_inS33ser[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS33ser_mux_inst_1_U1 ( .s (new_AGEMA_signal_3901), .b ({new_AGEMA_signal_3917, new_AGEMA_signal_3913}), .a ({new_AGEMA_signal_3480, stateArray_input_MC[1]}), .c ({new_AGEMA_signal_3499, stateArray_inS33ser[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS33ser_mux_inst_2_U1 ( .s (new_AGEMA_signal_3901), .b ({new_AGEMA_signal_3925, new_AGEMA_signal_3921}), .a ({new_AGEMA_signal_3481, stateArray_input_MC[2]}), .c ({new_AGEMA_signal_3501, stateArray_inS33ser[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS33ser_mux_inst_3_U1 ( .s (new_AGEMA_signal_3901), .b ({new_AGEMA_signal_3933, new_AGEMA_signal_3929}), .a ({new_AGEMA_signal_3482, stateArray_input_MC[3]}), .c ({new_AGEMA_signal_3503, stateArray_inS33ser[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS33ser_mux_inst_4_U1 ( .s (new_AGEMA_signal_3901), .b ({new_AGEMA_signal_3941, new_AGEMA_signal_3937}), .a ({new_AGEMA_signal_3483, stateArray_input_MC[4]}), .c ({new_AGEMA_signal_3505, stateArray_inS33ser[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS33ser_mux_inst_5_U1 ( .s (new_AGEMA_signal_3901), .b ({new_AGEMA_signal_3949, new_AGEMA_signal_3945}), .a ({new_AGEMA_signal_3484, stateArray_input_MC[5]}), .c ({new_AGEMA_signal_3507, stateArray_inS33ser[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS33ser_mux_inst_6_U1 ( .s (new_AGEMA_signal_3901), .b ({new_AGEMA_signal_3957, new_AGEMA_signal_3953}), .a ({new_AGEMA_signal_3485, stateArray_input_MC[6]}), .c ({new_AGEMA_signal_3509, stateArray_inS33ser[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) stateArray_MUX_inS33ser_mux_inst_7_U1 ( .s (new_AGEMA_signal_3901), .b ({new_AGEMA_signal_3965, new_AGEMA_signal_3961}), .a ({new_AGEMA_signal_3486, stateArray_input_MC[7]}), .c ({new_AGEMA_signal_3511, stateArray_inS33ser[7]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) KeyArray_U42 ( .a ({new_AGEMA_signal_3472, KeyArray_n55}), .b ({new_AGEMA_signal_3973, new_AGEMA_signal_3969}), .c ({new_AGEMA_signal_3489, KeyArray_inS30par[7]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) KeyArray_U41 ( .a ({1'b0, new_AGEMA_signal_3977}), .b ({new_AGEMA_signal_3457, SboxOut[7]}), .c ({new_AGEMA_signal_3472, KeyArray_n55}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) KeyArray_U40 ( .a ({new_AGEMA_signal_3473, KeyArray_n54}), .b ({new_AGEMA_signal_3985, new_AGEMA_signal_3981}), .c ({new_AGEMA_signal_3490, KeyArray_inS30par[6]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) KeyArray_U39 ( .a ({1'b0, new_AGEMA_signal_3989}), .b ({new_AGEMA_signal_3458, SboxOut[6]}), .c ({new_AGEMA_signal_3473, KeyArray_n54}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) KeyArray_U38 ( .a ({new_AGEMA_signal_3474, KeyArray_n53}), .b ({new_AGEMA_signal_3997, new_AGEMA_signal_3993}), .c ({new_AGEMA_signal_3491, KeyArray_inS30par[5]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) KeyArray_U37 ( .a ({1'b0, new_AGEMA_signal_4001}), .b ({new_AGEMA_signal_3459, SboxOut[5]}), .c ({new_AGEMA_signal_3474, KeyArray_n53}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) KeyArray_U36 ( .a ({new_AGEMA_signal_3475, KeyArray_n52}), .b ({new_AGEMA_signal_4009, new_AGEMA_signal_4005}), .c ({new_AGEMA_signal_3492, KeyArray_inS30par[4]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) KeyArray_U35 ( .a ({1'b0, new_AGEMA_signal_4013}), .b ({new_AGEMA_signal_3460, SboxOut[4]}), .c ({new_AGEMA_signal_3475, KeyArray_n52}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) KeyArray_U34 ( .a ({new_AGEMA_signal_3476, KeyArray_n51}), .b ({new_AGEMA_signal_4021, new_AGEMA_signal_4017}), .c ({new_AGEMA_signal_3493, KeyArray_inS30par[3]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) KeyArray_U33 ( .a ({1'b0, new_AGEMA_signal_4025}), .b ({new_AGEMA_signal_3461, SboxOut[3]}), .c ({new_AGEMA_signal_3476, KeyArray_n51}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) KeyArray_U32 ( .a ({new_AGEMA_signal_3477, KeyArray_n50}), .b ({new_AGEMA_signal_4033, new_AGEMA_signal_4029}), .c ({new_AGEMA_signal_3494, KeyArray_inS30par[2]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) KeyArray_U31 ( .a ({1'b0, new_AGEMA_signal_4037}), .b ({new_AGEMA_signal_3462, SboxOut[2]}), .c ({new_AGEMA_signal_3477, KeyArray_n50}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) KeyArray_U30 ( .a ({new_AGEMA_signal_3478, KeyArray_n49}), .b ({new_AGEMA_signal_4045, new_AGEMA_signal_4041}), .c ({new_AGEMA_signal_3495, KeyArray_inS30par[1]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) KeyArray_U29 ( .a ({1'b0, new_AGEMA_signal_4049}), .b ({new_AGEMA_signal_3463, SboxOut[1]}), .c ({new_AGEMA_signal_3478, KeyArray_n49}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) KeyArray_U28 ( .a ({new_AGEMA_signal_3456, KeyArray_n48}), .b ({new_AGEMA_signal_4057, new_AGEMA_signal_4053}), .c ({new_AGEMA_signal_3479, KeyArray_inS30par[0]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) KeyArray_U27 ( .a ({1'b0, new_AGEMA_signal_4061}), .b ({new_AGEMA_signal_3454, SboxOut[0]}), .c ({new_AGEMA_signal_3456, KeyArray_n48}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S30reg_gff_1_SFF_0_U1 ( .s (new_AGEMA_signal_4065), .b ({new_AGEMA_signal_4073, new_AGEMA_signal_4069}), .a ({new_AGEMA_signal_3496, KeyArray_S30reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_3512, KeyArray_S30reg_gff_1_SFF_0_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1 ( .s (new_AGEMA_signal_4077), .b ({new_AGEMA_signal_4085, new_AGEMA_signal_4081}), .a ({new_AGEMA_signal_3479, KeyArray_inS30par[0]}), .c ({new_AGEMA_signal_3496, KeyArray_S30reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S30reg_gff_1_SFF_1_U1 ( .s (new_AGEMA_signal_4065), .b ({new_AGEMA_signal_4093, new_AGEMA_signal_4089}), .a ({new_AGEMA_signal_3513, KeyArray_S30reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_3527, KeyArray_S30reg_gff_1_SFF_1_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1 ( .s (new_AGEMA_signal_4077), .b ({new_AGEMA_signal_4101, new_AGEMA_signal_4097}), .a ({new_AGEMA_signal_3495, KeyArray_inS30par[1]}), .c ({new_AGEMA_signal_3513, KeyArray_S30reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S30reg_gff_1_SFF_2_U1 ( .s (new_AGEMA_signal_4065), .b ({new_AGEMA_signal_4109, new_AGEMA_signal_4105}), .a ({new_AGEMA_signal_3514, KeyArray_S30reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_3528, KeyArray_S30reg_gff_1_SFF_2_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1 ( .s (new_AGEMA_signal_4077), .b ({new_AGEMA_signal_4117, new_AGEMA_signal_4113}), .a ({new_AGEMA_signal_3494, KeyArray_inS30par[2]}), .c ({new_AGEMA_signal_3514, KeyArray_S30reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S30reg_gff_1_SFF_3_U1 ( .s (new_AGEMA_signal_4065), .b ({new_AGEMA_signal_4125, new_AGEMA_signal_4121}), .a ({new_AGEMA_signal_3515, KeyArray_S30reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_3529, KeyArray_S30reg_gff_1_SFF_3_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1 ( .s (new_AGEMA_signal_4077), .b ({new_AGEMA_signal_4133, new_AGEMA_signal_4129}), .a ({new_AGEMA_signal_3493, KeyArray_inS30par[3]}), .c ({new_AGEMA_signal_3515, KeyArray_S30reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S30reg_gff_1_SFF_4_U1 ( .s (new_AGEMA_signal_4065), .b ({new_AGEMA_signal_4141, new_AGEMA_signal_4137}), .a ({new_AGEMA_signal_3516, KeyArray_S30reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_3530, KeyArray_S30reg_gff_1_SFF_4_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1 ( .s (new_AGEMA_signal_4077), .b ({new_AGEMA_signal_4149, new_AGEMA_signal_4145}), .a ({new_AGEMA_signal_3492, KeyArray_inS30par[4]}), .c ({new_AGEMA_signal_3516, KeyArray_S30reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S30reg_gff_1_SFF_5_U1 ( .s (new_AGEMA_signal_4065), .b ({new_AGEMA_signal_4157, new_AGEMA_signal_4153}), .a ({new_AGEMA_signal_3517, KeyArray_S30reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_3531, KeyArray_S30reg_gff_1_SFF_5_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1 ( .s (new_AGEMA_signal_4077), .b ({new_AGEMA_signal_4165, new_AGEMA_signal_4161}), .a ({new_AGEMA_signal_3491, KeyArray_inS30par[5]}), .c ({new_AGEMA_signal_3517, KeyArray_S30reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S30reg_gff_1_SFF_6_U1 ( .s (new_AGEMA_signal_4065), .b ({new_AGEMA_signal_4173, new_AGEMA_signal_4169}), .a ({new_AGEMA_signal_3518, KeyArray_S30reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_3532, KeyArray_S30reg_gff_1_SFF_6_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1 ( .s (new_AGEMA_signal_4077), .b ({new_AGEMA_signal_4181, new_AGEMA_signal_4177}), .a ({new_AGEMA_signal_3490, KeyArray_inS30par[6]}), .c ({new_AGEMA_signal_3518, KeyArray_S30reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S30reg_gff_1_SFF_7_U1 ( .s (new_AGEMA_signal_4065), .b ({new_AGEMA_signal_4189, new_AGEMA_signal_4185}), .a ({new_AGEMA_signal_3519, KeyArray_S30reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_3533, KeyArray_S30reg_gff_1_SFF_7_n5}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1 ( .s (new_AGEMA_signal_4077), .b ({new_AGEMA_signal_4197, new_AGEMA_signal_4193}), .a ({new_AGEMA_signal_3489, KeyArray_inS30par[7]}), .c ({new_AGEMA_signal_3519, KeyArray_S30reg_gff_1_SFF_7_QD}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M46_U1 ( .a ({new_AGEMA_signal_3404, Inst_bSbox_M44}), .b ({new_AGEMA_signal_4203, new_AGEMA_signal_4200}), .clk (clk), .r ({Fresh[67], Fresh[66], Fresh[65], Fresh[64]}), .c ({new_AGEMA_signal_3414, Inst_bSbox_M46}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M47_U1 ( .a ({new_AGEMA_signal_3400, Inst_bSbox_M40}), .b ({new_AGEMA_signal_4209, new_AGEMA_signal_4206}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69], Fresh[68]}), .c ({new_AGEMA_signal_3405, Inst_bSbox_M47}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M48_U1 ( .a ({new_AGEMA_signal_3399, Inst_bSbox_M39}), .b ({new_AGEMA_signal_4215, new_AGEMA_signal_4212}), .clk (clk), .r ({Fresh[75], Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_3406, Inst_bSbox_M48}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M49_U1 ( .a ({new_AGEMA_signal_3403, Inst_bSbox_M43}), .b ({new_AGEMA_signal_4221, new_AGEMA_signal_4218}), .clk (clk), .r ({Fresh[79], Fresh[78], Fresh[77], Fresh[76]}), .c ({new_AGEMA_signal_3415, Inst_bSbox_M49}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M50_U1 ( .a ({new_AGEMA_signal_3398, Inst_bSbox_M38}), .b ({new_AGEMA_signal_4227, new_AGEMA_signal_4224}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81], Fresh[80]}), .c ({new_AGEMA_signal_3407, Inst_bSbox_M50}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M51_U1 ( .a ({new_AGEMA_signal_3397, Inst_bSbox_M37}), .b ({new_AGEMA_signal_4233, new_AGEMA_signal_4230}), .clk (clk), .r ({Fresh[87], Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_3408, Inst_bSbox_M51}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M52_U1 ( .a ({new_AGEMA_signal_3402, Inst_bSbox_M42}), .b ({new_AGEMA_signal_4239, new_AGEMA_signal_4236}), .clk (clk), .r ({Fresh[91], Fresh[90], Fresh[89], Fresh[88]}), .c ({new_AGEMA_signal_3416, Inst_bSbox_M52}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M53_U1 ( .a ({new_AGEMA_signal_3413, Inst_bSbox_M45}), .b ({new_AGEMA_signal_4245, new_AGEMA_signal_4242}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92]}), .c ({new_AGEMA_signal_3425, Inst_bSbox_M53}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M54_U1 ( .a ({new_AGEMA_signal_3401, Inst_bSbox_M41}), .b ({new_AGEMA_signal_4251, new_AGEMA_signal_4248}), .clk (clk), .r ({Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_3417, Inst_bSbox_M54}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M55_U1 ( .a ({new_AGEMA_signal_3404, Inst_bSbox_M44}), .b ({new_AGEMA_signal_4257, new_AGEMA_signal_4254}), .clk (clk), .r ({Fresh[103], Fresh[102], Fresh[101], Fresh[100]}), .c ({new_AGEMA_signal_3418, Inst_bSbox_M55}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M56_U1 ( .a ({new_AGEMA_signal_3400, Inst_bSbox_M40}), .b ({new_AGEMA_signal_4263, new_AGEMA_signal_4260}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105], Fresh[104]}), .c ({new_AGEMA_signal_3409, Inst_bSbox_M56}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M57_U1 ( .a ({new_AGEMA_signal_3399, Inst_bSbox_M39}), .b ({new_AGEMA_signal_4269, new_AGEMA_signal_4266}), .clk (clk), .r ({Fresh[111], Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_3410, Inst_bSbox_M57}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M58_U1 ( .a ({new_AGEMA_signal_3403, Inst_bSbox_M43}), .b ({new_AGEMA_signal_4275, new_AGEMA_signal_4272}), .clk (clk), .r ({Fresh[115], Fresh[114], Fresh[113], Fresh[112]}), .c ({new_AGEMA_signal_3419, Inst_bSbox_M58}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M59_U1 ( .a ({new_AGEMA_signal_3398, Inst_bSbox_M38}), .b ({new_AGEMA_signal_4281, new_AGEMA_signal_4278}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116]}), .c ({new_AGEMA_signal_3411, Inst_bSbox_M59}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M60_U1 ( .a ({new_AGEMA_signal_3397, Inst_bSbox_M37}), .b ({new_AGEMA_signal_4287, new_AGEMA_signal_4284}), .clk (clk), .r ({Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_3412, Inst_bSbox_M60}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M61_U1 ( .a ({new_AGEMA_signal_3402, Inst_bSbox_M42}), .b ({new_AGEMA_signal_4293, new_AGEMA_signal_4290}), .clk (clk), .r ({Fresh[127], Fresh[126], Fresh[125], Fresh[124]}), .c ({new_AGEMA_signal_3420, Inst_bSbox_M61}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M62_U1 ( .a ({new_AGEMA_signal_3413, Inst_bSbox_M45}), .b ({new_AGEMA_signal_4299, new_AGEMA_signal_4296}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129], Fresh[128]}), .c ({new_AGEMA_signal_3426, Inst_bSbox_M62}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_AND_M63_U1 ( .a ({new_AGEMA_signal_3401, Inst_bSbox_M41}), .b ({new_AGEMA_signal_4305, new_AGEMA_signal_4302}), .clk (clk), .r ({Fresh[135], Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_3421, Inst_bSbox_M63}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_L0_U1 ( .a ({new_AGEMA_signal_3420, Inst_bSbox_M61}), .b ({new_AGEMA_signal_3426, Inst_bSbox_M62}), .c ({new_AGEMA_signal_3435, Inst_bSbox_L0}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_L1_U1 ( .a ({new_AGEMA_signal_3407, Inst_bSbox_M50}), .b ({new_AGEMA_signal_3409, Inst_bSbox_M56}), .c ({new_AGEMA_signal_3422, Inst_bSbox_L1}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_L2_U1 ( .a ({new_AGEMA_signal_3414, Inst_bSbox_M46}), .b ({new_AGEMA_signal_3406, Inst_bSbox_M48}), .c ({new_AGEMA_signal_3427, Inst_bSbox_L2}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_L3_U1 ( .a ({new_AGEMA_signal_3405, Inst_bSbox_M47}), .b ({new_AGEMA_signal_3418, Inst_bSbox_M55}), .c ({new_AGEMA_signal_3428, Inst_bSbox_L3}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_L4_U1 ( .a ({new_AGEMA_signal_3417, Inst_bSbox_M54}), .b ({new_AGEMA_signal_3419, Inst_bSbox_M58}), .c ({new_AGEMA_signal_3429, Inst_bSbox_L4}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_L5_U1 ( .a ({new_AGEMA_signal_3415, Inst_bSbox_M49}), .b ({new_AGEMA_signal_3420, Inst_bSbox_M61}), .c ({new_AGEMA_signal_3430, Inst_bSbox_L5}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_L6_U1 ( .a ({new_AGEMA_signal_3426, Inst_bSbox_M62}), .b ({new_AGEMA_signal_3430, Inst_bSbox_L5}), .c ({new_AGEMA_signal_3436, Inst_bSbox_L6}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_L7_U1 ( .a ({new_AGEMA_signal_3414, Inst_bSbox_M46}), .b ({new_AGEMA_signal_3428, Inst_bSbox_L3}), .c ({new_AGEMA_signal_3437, Inst_bSbox_L7}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_L8_U1 ( .a ({new_AGEMA_signal_3408, Inst_bSbox_M51}), .b ({new_AGEMA_signal_3411, Inst_bSbox_M59}), .c ({new_AGEMA_signal_3423, Inst_bSbox_L8}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_L9_U1 ( .a ({new_AGEMA_signal_3416, Inst_bSbox_M52}), .b ({new_AGEMA_signal_3425, Inst_bSbox_M53}), .c ({new_AGEMA_signal_3438, Inst_bSbox_L9}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_L10_U1 ( .a ({new_AGEMA_signal_3425, Inst_bSbox_M53}), .b ({new_AGEMA_signal_3429, Inst_bSbox_L4}), .c ({new_AGEMA_signal_3439, Inst_bSbox_L10}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_L11_U1 ( .a ({new_AGEMA_signal_3412, Inst_bSbox_M60}), .b ({new_AGEMA_signal_3427, Inst_bSbox_L2}), .c ({new_AGEMA_signal_3440, Inst_bSbox_L11}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_L12_U1 ( .a ({new_AGEMA_signal_3406, Inst_bSbox_M48}), .b ({new_AGEMA_signal_3408, Inst_bSbox_M51}), .c ({new_AGEMA_signal_3424, Inst_bSbox_L12}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_L13_U1 ( .a ({new_AGEMA_signal_3407, Inst_bSbox_M50}), .b ({new_AGEMA_signal_3435, Inst_bSbox_L0}), .c ({new_AGEMA_signal_3444, Inst_bSbox_L13}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_L14_U1 ( .a ({new_AGEMA_signal_3416, Inst_bSbox_M52}), .b ({new_AGEMA_signal_3420, Inst_bSbox_M61}), .c ({new_AGEMA_signal_3431, Inst_bSbox_L14}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_L15_U1 ( .a ({new_AGEMA_signal_3418, Inst_bSbox_M55}), .b ({new_AGEMA_signal_3422, Inst_bSbox_L1}), .c ({new_AGEMA_signal_3432, Inst_bSbox_L15}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_L16_U1 ( .a ({new_AGEMA_signal_3409, Inst_bSbox_M56}), .b ({new_AGEMA_signal_3435, Inst_bSbox_L0}), .c ({new_AGEMA_signal_3445, Inst_bSbox_L16}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_L17_U1 ( .a ({new_AGEMA_signal_3410, Inst_bSbox_M57}), .b ({new_AGEMA_signal_3422, Inst_bSbox_L1}), .c ({new_AGEMA_signal_3433, Inst_bSbox_L17}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_L18_U1 ( .a ({new_AGEMA_signal_3419, Inst_bSbox_M58}), .b ({new_AGEMA_signal_3423, Inst_bSbox_L8}), .c ({new_AGEMA_signal_3434, Inst_bSbox_L18}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_L19_U1 ( .a ({new_AGEMA_signal_3421, Inst_bSbox_M63}), .b ({new_AGEMA_signal_3429, Inst_bSbox_L4}), .c ({new_AGEMA_signal_3441, Inst_bSbox_L19}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_L20_U1 ( .a ({new_AGEMA_signal_3435, Inst_bSbox_L0}), .b ({new_AGEMA_signal_3422, Inst_bSbox_L1}), .c ({new_AGEMA_signal_3446, Inst_bSbox_L20}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_L21_U1 ( .a ({new_AGEMA_signal_3422, Inst_bSbox_L1}), .b ({new_AGEMA_signal_3437, Inst_bSbox_L7}), .c ({new_AGEMA_signal_3447, Inst_bSbox_L21}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_L22_U1 ( .a ({new_AGEMA_signal_3428, Inst_bSbox_L3}), .b ({new_AGEMA_signal_3424, Inst_bSbox_L12}), .c ({new_AGEMA_signal_3442, Inst_bSbox_L22}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_L23_U1 ( .a ({new_AGEMA_signal_3434, Inst_bSbox_L18}), .b ({new_AGEMA_signal_3427, Inst_bSbox_L2}), .c ({new_AGEMA_signal_3443, Inst_bSbox_L23}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_L24_U1 ( .a ({new_AGEMA_signal_3432, Inst_bSbox_L15}), .b ({new_AGEMA_signal_3438, Inst_bSbox_L9}), .c ({new_AGEMA_signal_3448, Inst_bSbox_L24}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_L25_U1 ( .a ({new_AGEMA_signal_3436, Inst_bSbox_L6}), .b ({new_AGEMA_signal_3439, Inst_bSbox_L10}), .c ({new_AGEMA_signal_3449, Inst_bSbox_L25}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_L26_U1 ( .a ({new_AGEMA_signal_3437, Inst_bSbox_L7}), .b ({new_AGEMA_signal_3438, Inst_bSbox_L9}), .c ({new_AGEMA_signal_3450, Inst_bSbox_L26}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_L27_U1 ( .a ({new_AGEMA_signal_3423, Inst_bSbox_L8}), .b ({new_AGEMA_signal_3439, Inst_bSbox_L10}), .c ({new_AGEMA_signal_3451, Inst_bSbox_L27}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_L28_U1 ( .a ({new_AGEMA_signal_3440, Inst_bSbox_L11}), .b ({new_AGEMA_signal_3431, Inst_bSbox_L14}), .c ({new_AGEMA_signal_3452, Inst_bSbox_L28}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_L29_U1 ( .a ({new_AGEMA_signal_3440, Inst_bSbox_L11}), .b ({new_AGEMA_signal_3433, Inst_bSbox_L17}), .c ({new_AGEMA_signal_3453, Inst_bSbox_L29}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_S0_U1 ( .a ({new_AGEMA_signal_3436, Inst_bSbox_L6}), .b ({new_AGEMA_signal_3448, Inst_bSbox_L24}), .c ({new_AGEMA_signal_3457, SboxOut[7]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_S1_U1 ( .a ({new_AGEMA_signal_3445, Inst_bSbox_L16}), .b ({new_AGEMA_signal_3450, Inst_bSbox_L26}), .c ({new_AGEMA_signal_3458, SboxOut[6]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_S2_U1 ( .a ({new_AGEMA_signal_3441, Inst_bSbox_L19}), .b ({new_AGEMA_signal_3452, Inst_bSbox_L28}), .c ({new_AGEMA_signal_3459, SboxOut[5]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_S3_U1 ( .a ({new_AGEMA_signal_3436, Inst_bSbox_L6}), .b ({new_AGEMA_signal_3447, Inst_bSbox_L21}), .c ({new_AGEMA_signal_3460, SboxOut[4]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_S4_U1 ( .a ({new_AGEMA_signal_3446, Inst_bSbox_L20}), .b ({new_AGEMA_signal_3442, Inst_bSbox_L22}), .c ({new_AGEMA_signal_3461, SboxOut[3]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_S5_U1 ( .a ({new_AGEMA_signal_3449, Inst_bSbox_L25}), .b ({new_AGEMA_signal_3453, Inst_bSbox_L29}), .c ({new_AGEMA_signal_3462, SboxOut[2]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_S6_U1 ( .a ({new_AGEMA_signal_3444, Inst_bSbox_L13}), .b ({new_AGEMA_signal_3451, Inst_bSbox_L27}), .c ({new_AGEMA_signal_3463, SboxOut[1]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) Inst_bSbox_XOR_S7_U1 ( .a ({new_AGEMA_signal_3436, Inst_bSbox_L6}), .b ({new_AGEMA_signal_3443, Inst_bSbox_L23}), .c ({new_AGEMA_signal_3454, SboxOut[0]}) ) ;
    buf_clk new_AGEMA_reg_buffer_1741 ( .C (clk), .D (new_AGEMA_signal_3696), .Q (new_AGEMA_signal_3697) ) ;
    buf_clk new_AGEMA_reg_buffer_1745 ( .C (clk), .D (new_AGEMA_signal_3700), .Q (new_AGEMA_signal_3701) ) ;
    buf_clk new_AGEMA_reg_buffer_1749 ( .C (clk), .D (new_AGEMA_signal_3704), .Q (new_AGEMA_signal_3705) ) ;
    buf_clk new_AGEMA_reg_buffer_1753 ( .C (clk), .D (new_AGEMA_signal_3708), .Q (new_AGEMA_signal_3709) ) ;
    buf_clk new_AGEMA_reg_buffer_1757 ( .C (clk), .D (new_AGEMA_signal_3712), .Q (new_AGEMA_signal_3713) ) ;
    buf_clk new_AGEMA_reg_buffer_1761 ( .C (clk), .D (new_AGEMA_signal_3716), .Q (new_AGEMA_signal_3717) ) ;
    buf_clk new_AGEMA_reg_buffer_1765 ( .C (clk), .D (new_AGEMA_signal_3720), .Q (new_AGEMA_signal_3721) ) ;
    buf_clk new_AGEMA_reg_buffer_1769 ( .C (clk), .D (new_AGEMA_signal_3724), .Q (new_AGEMA_signal_3725) ) ;
    buf_clk new_AGEMA_reg_buffer_1773 ( .C (clk), .D (new_AGEMA_signal_3728), .Q (new_AGEMA_signal_3729) ) ;
    buf_clk new_AGEMA_reg_buffer_1777 ( .C (clk), .D (new_AGEMA_signal_3732), .Q (new_AGEMA_signal_3733) ) ;
    buf_clk new_AGEMA_reg_buffer_1781 ( .C (clk), .D (new_AGEMA_signal_3736), .Q (new_AGEMA_signal_3737) ) ;
    buf_clk new_AGEMA_reg_buffer_1785 ( .C (clk), .D (new_AGEMA_signal_3740), .Q (new_AGEMA_signal_3741) ) ;
    buf_clk new_AGEMA_reg_buffer_1789 ( .C (clk), .D (new_AGEMA_signal_3744), .Q (new_AGEMA_signal_3745) ) ;
    buf_clk new_AGEMA_reg_buffer_1793 ( .C (clk), .D (new_AGEMA_signal_3748), .Q (new_AGEMA_signal_3749) ) ;
    buf_clk new_AGEMA_reg_buffer_1797 ( .C (clk), .D (new_AGEMA_signal_3752), .Q (new_AGEMA_signal_3753) ) ;
    buf_clk new_AGEMA_reg_buffer_1801 ( .C (clk), .D (new_AGEMA_signal_3756), .Q (new_AGEMA_signal_3757) ) ;
    buf_clk new_AGEMA_reg_buffer_1805 ( .C (clk), .D (new_AGEMA_signal_3760), .Q (new_AGEMA_signal_3761) ) ;
    buf_clk new_AGEMA_reg_buffer_1809 ( .C (clk), .D (new_AGEMA_signal_3764), .Q (new_AGEMA_signal_3765) ) ;
    buf_clk new_AGEMA_reg_buffer_1813 ( .C (clk), .D (new_AGEMA_signal_3768), .Q (new_AGEMA_signal_3769) ) ;
    buf_clk new_AGEMA_reg_buffer_1817 ( .C (clk), .D (new_AGEMA_signal_3772), .Q (new_AGEMA_signal_3773) ) ;
    buf_clk new_AGEMA_reg_buffer_1821 ( .C (clk), .D (new_AGEMA_signal_3776), .Q (new_AGEMA_signal_3777) ) ;
    buf_clk new_AGEMA_reg_buffer_1825 ( .C (clk), .D (new_AGEMA_signal_3780), .Q (new_AGEMA_signal_3781) ) ;
    buf_clk new_AGEMA_reg_buffer_1829 ( .C (clk), .D (new_AGEMA_signal_3784), .Q (new_AGEMA_signal_3785) ) ;
    buf_clk new_AGEMA_reg_buffer_1833 ( .C (clk), .D (new_AGEMA_signal_3788), .Q (new_AGEMA_signal_3789) ) ;
    buf_clk new_AGEMA_reg_buffer_1837 ( .C (clk), .D (new_AGEMA_signal_3792), .Q (new_AGEMA_signal_3793) ) ;
    buf_clk new_AGEMA_reg_buffer_1841 ( .C (clk), .D (new_AGEMA_signal_3796), .Q (new_AGEMA_signal_3797) ) ;
    buf_clk new_AGEMA_reg_buffer_1845 ( .C (clk), .D (new_AGEMA_signal_3800), .Q (new_AGEMA_signal_3801) ) ;
    buf_clk new_AGEMA_reg_buffer_1849 ( .C (clk), .D (new_AGEMA_signal_3804), .Q (new_AGEMA_signal_3805) ) ;
    buf_clk new_AGEMA_reg_buffer_1853 ( .C (clk), .D (new_AGEMA_signal_3808), .Q (new_AGEMA_signal_3809) ) ;
    buf_clk new_AGEMA_reg_buffer_1857 ( .C (clk), .D (new_AGEMA_signal_3812), .Q (new_AGEMA_signal_3813) ) ;
    buf_clk new_AGEMA_reg_buffer_1861 ( .C (clk), .D (new_AGEMA_signal_3816), .Q (new_AGEMA_signal_3817) ) ;
    buf_clk new_AGEMA_reg_buffer_1865 ( .C (clk), .D (new_AGEMA_signal_3820), .Q (new_AGEMA_signal_3821) ) ;
    buf_clk new_AGEMA_reg_buffer_1869 ( .C (clk), .D (new_AGEMA_signal_3824), .Q (new_AGEMA_signal_3825) ) ;
    buf_clk new_AGEMA_reg_buffer_1873 ( .C (clk), .D (new_AGEMA_signal_3828), .Q (new_AGEMA_signal_3829) ) ;
    buf_clk new_AGEMA_reg_buffer_1877 ( .C (clk), .D (new_AGEMA_signal_3832), .Q (new_AGEMA_signal_3833) ) ;
    buf_clk new_AGEMA_reg_buffer_1881 ( .C (clk), .D (new_AGEMA_signal_3836), .Q (new_AGEMA_signal_3837) ) ;
    buf_clk new_AGEMA_reg_buffer_1885 ( .C (clk), .D (new_AGEMA_signal_3840), .Q (new_AGEMA_signal_3841) ) ;
    buf_clk new_AGEMA_reg_buffer_1889 ( .C (clk), .D (new_AGEMA_signal_3844), .Q (new_AGEMA_signal_3845) ) ;
    buf_clk new_AGEMA_reg_buffer_1893 ( .C (clk), .D (new_AGEMA_signal_3848), .Q (new_AGEMA_signal_3849) ) ;
    buf_clk new_AGEMA_reg_buffer_1897 ( .C (clk), .D (new_AGEMA_signal_3852), .Q (new_AGEMA_signal_3853) ) ;
    buf_clk new_AGEMA_reg_buffer_1901 ( .C (clk), .D (new_AGEMA_signal_3856), .Q (new_AGEMA_signal_3857) ) ;
    buf_clk new_AGEMA_reg_buffer_1905 ( .C (clk), .D (new_AGEMA_signal_3860), .Q (new_AGEMA_signal_3861) ) ;
    buf_clk new_AGEMA_reg_buffer_1909 ( .C (clk), .D (new_AGEMA_signal_3864), .Q (new_AGEMA_signal_3865) ) ;
    buf_clk new_AGEMA_reg_buffer_1913 ( .C (clk), .D (new_AGEMA_signal_3868), .Q (new_AGEMA_signal_3869) ) ;
    buf_clk new_AGEMA_reg_buffer_1917 ( .C (clk), .D (new_AGEMA_signal_3872), .Q (new_AGEMA_signal_3873) ) ;
    buf_clk new_AGEMA_reg_buffer_1921 ( .C (clk), .D (new_AGEMA_signal_3876), .Q (new_AGEMA_signal_3877) ) ;
    buf_clk new_AGEMA_reg_buffer_1925 ( .C (clk), .D (new_AGEMA_signal_3880), .Q (new_AGEMA_signal_3881) ) ;
    buf_clk new_AGEMA_reg_buffer_1929 ( .C (clk), .D (new_AGEMA_signal_3884), .Q (new_AGEMA_signal_3885) ) ;
    buf_clk new_AGEMA_reg_buffer_1933 ( .C (clk), .D (new_AGEMA_signal_3888), .Q (new_AGEMA_signal_3889) ) ;
    buf_clk new_AGEMA_reg_buffer_1937 ( .C (clk), .D (new_AGEMA_signal_3892), .Q (new_AGEMA_signal_3893) ) ;
    buf_clk new_AGEMA_reg_buffer_1941 ( .C (clk), .D (new_AGEMA_signal_3896), .Q (new_AGEMA_signal_3897) ) ;
    buf_clk new_AGEMA_reg_buffer_1945 ( .C (clk), .D (new_AGEMA_signal_3900), .Q (new_AGEMA_signal_3901) ) ;
    buf_clk new_AGEMA_reg_buffer_1949 ( .C (clk), .D (new_AGEMA_signal_3904), .Q (new_AGEMA_signal_3905) ) ;
    buf_clk new_AGEMA_reg_buffer_1953 ( .C (clk), .D (new_AGEMA_signal_3908), .Q (new_AGEMA_signal_3909) ) ;
    buf_clk new_AGEMA_reg_buffer_1957 ( .C (clk), .D (new_AGEMA_signal_3912), .Q (new_AGEMA_signal_3913) ) ;
    buf_clk new_AGEMA_reg_buffer_1961 ( .C (clk), .D (new_AGEMA_signal_3916), .Q (new_AGEMA_signal_3917) ) ;
    buf_clk new_AGEMA_reg_buffer_1965 ( .C (clk), .D (new_AGEMA_signal_3920), .Q (new_AGEMA_signal_3921) ) ;
    buf_clk new_AGEMA_reg_buffer_1969 ( .C (clk), .D (new_AGEMA_signal_3924), .Q (new_AGEMA_signal_3925) ) ;
    buf_clk new_AGEMA_reg_buffer_1973 ( .C (clk), .D (new_AGEMA_signal_3928), .Q (new_AGEMA_signal_3929) ) ;
    buf_clk new_AGEMA_reg_buffer_1977 ( .C (clk), .D (new_AGEMA_signal_3932), .Q (new_AGEMA_signal_3933) ) ;
    buf_clk new_AGEMA_reg_buffer_1981 ( .C (clk), .D (new_AGEMA_signal_3936), .Q (new_AGEMA_signal_3937) ) ;
    buf_clk new_AGEMA_reg_buffer_1985 ( .C (clk), .D (new_AGEMA_signal_3940), .Q (new_AGEMA_signal_3941) ) ;
    buf_clk new_AGEMA_reg_buffer_1989 ( .C (clk), .D (new_AGEMA_signal_3944), .Q (new_AGEMA_signal_3945) ) ;
    buf_clk new_AGEMA_reg_buffer_1993 ( .C (clk), .D (new_AGEMA_signal_3948), .Q (new_AGEMA_signal_3949) ) ;
    buf_clk new_AGEMA_reg_buffer_1997 ( .C (clk), .D (new_AGEMA_signal_3952), .Q (new_AGEMA_signal_3953) ) ;
    buf_clk new_AGEMA_reg_buffer_2001 ( .C (clk), .D (new_AGEMA_signal_3956), .Q (new_AGEMA_signal_3957) ) ;
    buf_clk new_AGEMA_reg_buffer_2005 ( .C (clk), .D (new_AGEMA_signal_3960), .Q (new_AGEMA_signal_3961) ) ;
    buf_clk new_AGEMA_reg_buffer_2009 ( .C (clk), .D (new_AGEMA_signal_3964), .Q (new_AGEMA_signal_3965) ) ;
    buf_clk new_AGEMA_reg_buffer_2013 ( .C (clk), .D (new_AGEMA_signal_3968), .Q (new_AGEMA_signal_3969) ) ;
    buf_clk new_AGEMA_reg_buffer_2017 ( .C (clk), .D (new_AGEMA_signal_3972), .Q (new_AGEMA_signal_3973) ) ;
    buf_clk new_AGEMA_reg_buffer_2021 ( .C (clk), .D (new_AGEMA_signal_3976), .Q (new_AGEMA_signal_3977) ) ;
    buf_clk new_AGEMA_reg_buffer_2025 ( .C (clk), .D (new_AGEMA_signal_3980), .Q (new_AGEMA_signal_3981) ) ;
    buf_clk new_AGEMA_reg_buffer_2029 ( .C (clk), .D (new_AGEMA_signal_3984), .Q (new_AGEMA_signal_3985) ) ;
    buf_clk new_AGEMA_reg_buffer_2033 ( .C (clk), .D (new_AGEMA_signal_3988), .Q (new_AGEMA_signal_3989) ) ;
    buf_clk new_AGEMA_reg_buffer_2037 ( .C (clk), .D (new_AGEMA_signal_3992), .Q (new_AGEMA_signal_3993) ) ;
    buf_clk new_AGEMA_reg_buffer_2041 ( .C (clk), .D (new_AGEMA_signal_3996), .Q (new_AGEMA_signal_3997) ) ;
    buf_clk new_AGEMA_reg_buffer_2045 ( .C (clk), .D (new_AGEMA_signal_4000), .Q (new_AGEMA_signal_4001) ) ;
    buf_clk new_AGEMA_reg_buffer_2049 ( .C (clk), .D (new_AGEMA_signal_4004), .Q (new_AGEMA_signal_4005) ) ;
    buf_clk new_AGEMA_reg_buffer_2053 ( .C (clk), .D (new_AGEMA_signal_4008), .Q (new_AGEMA_signal_4009) ) ;
    buf_clk new_AGEMA_reg_buffer_2057 ( .C (clk), .D (new_AGEMA_signal_4012), .Q (new_AGEMA_signal_4013) ) ;
    buf_clk new_AGEMA_reg_buffer_2061 ( .C (clk), .D (new_AGEMA_signal_4016), .Q (new_AGEMA_signal_4017) ) ;
    buf_clk new_AGEMA_reg_buffer_2065 ( .C (clk), .D (new_AGEMA_signal_4020), .Q (new_AGEMA_signal_4021) ) ;
    buf_clk new_AGEMA_reg_buffer_2069 ( .C (clk), .D (new_AGEMA_signal_4024), .Q (new_AGEMA_signal_4025) ) ;
    buf_clk new_AGEMA_reg_buffer_2073 ( .C (clk), .D (new_AGEMA_signal_4028), .Q (new_AGEMA_signal_4029) ) ;
    buf_clk new_AGEMA_reg_buffer_2077 ( .C (clk), .D (new_AGEMA_signal_4032), .Q (new_AGEMA_signal_4033) ) ;
    buf_clk new_AGEMA_reg_buffer_2081 ( .C (clk), .D (new_AGEMA_signal_4036), .Q (new_AGEMA_signal_4037) ) ;
    buf_clk new_AGEMA_reg_buffer_2085 ( .C (clk), .D (new_AGEMA_signal_4040), .Q (new_AGEMA_signal_4041) ) ;
    buf_clk new_AGEMA_reg_buffer_2089 ( .C (clk), .D (new_AGEMA_signal_4044), .Q (new_AGEMA_signal_4045) ) ;
    buf_clk new_AGEMA_reg_buffer_2093 ( .C (clk), .D (new_AGEMA_signal_4048), .Q (new_AGEMA_signal_4049) ) ;
    buf_clk new_AGEMA_reg_buffer_2097 ( .C (clk), .D (new_AGEMA_signal_4052), .Q (new_AGEMA_signal_4053) ) ;
    buf_clk new_AGEMA_reg_buffer_2101 ( .C (clk), .D (new_AGEMA_signal_4056), .Q (new_AGEMA_signal_4057) ) ;
    buf_clk new_AGEMA_reg_buffer_2105 ( .C (clk), .D (new_AGEMA_signal_4060), .Q (new_AGEMA_signal_4061) ) ;
    buf_clk new_AGEMA_reg_buffer_2109 ( .C (clk), .D (new_AGEMA_signal_4064), .Q (new_AGEMA_signal_4065) ) ;
    buf_clk new_AGEMA_reg_buffer_2113 ( .C (clk), .D (new_AGEMA_signal_4068), .Q (new_AGEMA_signal_4069) ) ;
    buf_clk new_AGEMA_reg_buffer_2117 ( .C (clk), .D (new_AGEMA_signal_4072), .Q (new_AGEMA_signal_4073) ) ;
    buf_clk new_AGEMA_reg_buffer_2121 ( .C (clk), .D (new_AGEMA_signal_4076), .Q (new_AGEMA_signal_4077) ) ;
    buf_clk new_AGEMA_reg_buffer_2125 ( .C (clk), .D (new_AGEMA_signal_4080), .Q (new_AGEMA_signal_4081) ) ;
    buf_clk new_AGEMA_reg_buffer_2129 ( .C (clk), .D (new_AGEMA_signal_4084), .Q (new_AGEMA_signal_4085) ) ;
    buf_clk new_AGEMA_reg_buffer_2133 ( .C (clk), .D (new_AGEMA_signal_4088), .Q (new_AGEMA_signal_4089) ) ;
    buf_clk new_AGEMA_reg_buffer_2137 ( .C (clk), .D (new_AGEMA_signal_4092), .Q (new_AGEMA_signal_4093) ) ;
    buf_clk new_AGEMA_reg_buffer_2141 ( .C (clk), .D (new_AGEMA_signal_4096), .Q (new_AGEMA_signal_4097) ) ;
    buf_clk new_AGEMA_reg_buffer_2145 ( .C (clk), .D (new_AGEMA_signal_4100), .Q (new_AGEMA_signal_4101) ) ;
    buf_clk new_AGEMA_reg_buffer_2149 ( .C (clk), .D (new_AGEMA_signal_4104), .Q (new_AGEMA_signal_4105) ) ;
    buf_clk new_AGEMA_reg_buffer_2153 ( .C (clk), .D (new_AGEMA_signal_4108), .Q (new_AGEMA_signal_4109) ) ;
    buf_clk new_AGEMA_reg_buffer_2157 ( .C (clk), .D (new_AGEMA_signal_4112), .Q (new_AGEMA_signal_4113) ) ;
    buf_clk new_AGEMA_reg_buffer_2161 ( .C (clk), .D (new_AGEMA_signal_4116), .Q (new_AGEMA_signal_4117) ) ;
    buf_clk new_AGEMA_reg_buffer_2165 ( .C (clk), .D (new_AGEMA_signal_4120), .Q (new_AGEMA_signal_4121) ) ;
    buf_clk new_AGEMA_reg_buffer_2169 ( .C (clk), .D (new_AGEMA_signal_4124), .Q (new_AGEMA_signal_4125) ) ;
    buf_clk new_AGEMA_reg_buffer_2173 ( .C (clk), .D (new_AGEMA_signal_4128), .Q (new_AGEMA_signal_4129) ) ;
    buf_clk new_AGEMA_reg_buffer_2177 ( .C (clk), .D (new_AGEMA_signal_4132), .Q (new_AGEMA_signal_4133) ) ;
    buf_clk new_AGEMA_reg_buffer_2181 ( .C (clk), .D (new_AGEMA_signal_4136), .Q (new_AGEMA_signal_4137) ) ;
    buf_clk new_AGEMA_reg_buffer_2185 ( .C (clk), .D (new_AGEMA_signal_4140), .Q (new_AGEMA_signal_4141) ) ;
    buf_clk new_AGEMA_reg_buffer_2189 ( .C (clk), .D (new_AGEMA_signal_4144), .Q (new_AGEMA_signal_4145) ) ;
    buf_clk new_AGEMA_reg_buffer_2193 ( .C (clk), .D (new_AGEMA_signal_4148), .Q (new_AGEMA_signal_4149) ) ;
    buf_clk new_AGEMA_reg_buffer_2197 ( .C (clk), .D (new_AGEMA_signal_4152), .Q (new_AGEMA_signal_4153) ) ;
    buf_clk new_AGEMA_reg_buffer_2201 ( .C (clk), .D (new_AGEMA_signal_4156), .Q (new_AGEMA_signal_4157) ) ;
    buf_clk new_AGEMA_reg_buffer_2205 ( .C (clk), .D (new_AGEMA_signal_4160), .Q (new_AGEMA_signal_4161) ) ;
    buf_clk new_AGEMA_reg_buffer_2209 ( .C (clk), .D (new_AGEMA_signal_4164), .Q (new_AGEMA_signal_4165) ) ;
    buf_clk new_AGEMA_reg_buffer_2213 ( .C (clk), .D (new_AGEMA_signal_4168), .Q (new_AGEMA_signal_4169) ) ;
    buf_clk new_AGEMA_reg_buffer_2217 ( .C (clk), .D (new_AGEMA_signal_4172), .Q (new_AGEMA_signal_4173) ) ;
    buf_clk new_AGEMA_reg_buffer_2221 ( .C (clk), .D (new_AGEMA_signal_4176), .Q (new_AGEMA_signal_4177) ) ;
    buf_clk new_AGEMA_reg_buffer_2225 ( .C (clk), .D (new_AGEMA_signal_4180), .Q (new_AGEMA_signal_4181) ) ;
    buf_clk new_AGEMA_reg_buffer_2229 ( .C (clk), .D (new_AGEMA_signal_4184), .Q (new_AGEMA_signal_4185) ) ;
    buf_clk new_AGEMA_reg_buffer_2233 ( .C (clk), .D (new_AGEMA_signal_4188), .Q (new_AGEMA_signal_4189) ) ;
    buf_clk new_AGEMA_reg_buffer_2237 ( .C (clk), .D (new_AGEMA_signal_4192), .Q (new_AGEMA_signal_4193) ) ;
    buf_clk new_AGEMA_reg_buffer_2241 ( .C (clk), .D (new_AGEMA_signal_4196), .Q (new_AGEMA_signal_4197) ) ;
    buf_clk new_AGEMA_reg_buffer_2353 ( .C (clk), .D (new_AGEMA_signal_4308), .Q (new_AGEMA_signal_4309) ) ;
    buf_clk new_AGEMA_reg_buffer_2357 ( .C (clk), .D (new_AGEMA_signal_4312), .Q (new_AGEMA_signal_4313) ) ;
    buf_clk new_AGEMA_reg_buffer_2361 ( .C (clk), .D (new_AGEMA_signal_4316), .Q (new_AGEMA_signal_4317) ) ;
    buf_clk new_AGEMA_reg_buffer_2365 ( .C (clk), .D (new_AGEMA_signal_4320), .Q (new_AGEMA_signal_4321) ) ;
    buf_clk new_AGEMA_reg_buffer_2369 ( .C (clk), .D (new_AGEMA_signal_4324), .Q (new_AGEMA_signal_4325) ) ;
    buf_clk new_AGEMA_reg_buffer_2373 ( .C (clk), .D (new_AGEMA_signal_4328), .Q (new_AGEMA_signal_4329) ) ;
    buf_clk new_AGEMA_reg_buffer_2377 ( .C (clk), .D (new_AGEMA_signal_4332), .Q (new_AGEMA_signal_4333) ) ;
    buf_clk new_AGEMA_reg_buffer_2381 ( .C (clk), .D (new_AGEMA_signal_4336), .Q (new_AGEMA_signal_4337) ) ;
    buf_clk new_AGEMA_reg_buffer_2385 ( .C (clk), .D (new_AGEMA_signal_4340), .Q (new_AGEMA_signal_4341) ) ;
    buf_clk new_AGEMA_reg_buffer_2389 ( .C (clk), .D (new_AGEMA_signal_4344), .Q (new_AGEMA_signal_4345) ) ;
    buf_clk new_AGEMA_reg_buffer_2393 ( .C (clk), .D (new_AGEMA_signal_4348), .Q (new_AGEMA_signal_4349) ) ;
    buf_clk new_AGEMA_reg_buffer_2397 ( .C (clk), .D (new_AGEMA_signal_4352), .Q (new_AGEMA_signal_4353) ) ;
    buf_clk new_AGEMA_reg_buffer_2401 ( .C (clk), .D (new_AGEMA_signal_4356), .Q (new_AGEMA_signal_4357) ) ;
    buf_clk new_AGEMA_reg_buffer_2405 ( .C (clk), .D (new_AGEMA_signal_4360), .Q (new_AGEMA_signal_4361) ) ;
    buf_clk new_AGEMA_reg_buffer_2409 ( .C (clk), .D (new_AGEMA_signal_4364), .Q (new_AGEMA_signal_4365) ) ;
    buf_clk new_AGEMA_reg_buffer_2413 ( .C (clk), .D (new_AGEMA_signal_4368), .Q (new_AGEMA_signal_4369) ) ;
    buf_clk new_AGEMA_reg_buffer_2417 ( .C (clk), .D (new_AGEMA_signal_4372), .Q (new_AGEMA_signal_4373) ) ;
    buf_clk new_AGEMA_reg_buffer_2421 ( .C (clk), .D (new_AGEMA_signal_4376), .Q (new_AGEMA_signal_4377) ) ;
    buf_clk new_AGEMA_reg_buffer_2425 ( .C (clk), .D (new_AGEMA_signal_4380), .Q (new_AGEMA_signal_4381) ) ;
    buf_clk new_AGEMA_reg_buffer_2429 ( .C (clk), .D (new_AGEMA_signal_4384), .Q (new_AGEMA_signal_4385) ) ;
    buf_clk new_AGEMA_reg_buffer_2433 ( .C (clk), .D (new_AGEMA_signal_4388), .Q (new_AGEMA_signal_4389) ) ;
    buf_clk new_AGEMA_reg_buffer_2437 ( .C (clk), .D (new_AGEMA_signal_4392), .Q (new_AGEMA_signal_4393) ) ;
    buf_clk new_AGEMA_reg_buffer_2441 ( .C (clk), .D (new_AGEMA_signal_4396), .Q (new_AGEMA_signal_4397) ) ;
    buf_clk new_AGEMA_reg_buffer_2445 ( .C (clk), .D (new_AGEMA_signal_4400), .Q (new_AGEMA_signal_4401) ) ;
    buf_clk new_AGEMA_reg_buffer_2449 ( .C (clk), .D (new_AGEMA_signal_4404), .Q (new_AGEMA_signal_4405) ) ;
    buf_clk new_AGEMA_reg_buffer_2453 ( .C (clk), .D (new_AGEMA_signal_4408), .Q (new_AGEMA_signal_4409) ) ;
    buf_clk new_AGEMA_reg_buffer_2457 ( .C (clk), .D (new_AGEMA_signal_4412), .Q (new_AGEMA_signal_4413) ) ;
    buf_clk new_AGEMA_reg_buffer_2461 ( .C (clk), .D (new_AGEMA_signal_4416), .Q (new_AGEMA_signal_4417) ) ;
    buf_clk new_AGEMA_reg_buffer_2465 ( .C (clk), .D (new_AGEMA_signal_4420), .Q (new_AGEMA_signal_4421) ) ;
    buf_clk new_AGEMA_reg_buffer_2469 ( .C (clk), .D (new_AGEMA_signal_4424), .Q (new_AGEMA_signal_4425) ) ;
    buf_clk new_AGEMA_reg_buffer_2473 ( .C (clk), .D (new_AGEMA_signal_4428), .Q (new_AGEMA_signal_4429) ) ;
    buf_clk new_AGEMA_reg_buffer_2477 ( .C (clk), .D (new_AGEMA_signal_4432), .Q (new_AGEMA_signal_4433) ) ;
    buf_clk new_AGEMA_reg_buffer_2481 ( .C (clk), .D (new_AGEMA_signal_4436), .Q (new_AGEMA_signal_4437) ) ;
    buf_clk new_AGEMA_reg_buffer_2485 ( .C (clk), .D (new_AGEMA_signal_4440), .Q (new_AGEMA_signal_4441) ) ;
    buf_clk new_AGEMA_reg_buffer_2489 ( .C (clk), .D (new_AGEMA_signal_4444), .Q (new_AGEMA_signal_4445) ) ;
    buf_clk new_AGEMA_reg_buffer_2493 ( .C (clk), .D (new_AGEMA_signal_4448), .Q (new_AGEMA_signal_4449) ) ;
    buf_clk new_AGEMA_reg_buffer_2497 ( .C (clk), .D (new_AGEMA_signal_4452), .Q (new_AGEMA_signal_4453) ) ;
    buf_clk new_AGEMA_reg_buffer_2501 ( .C (clk), .D (new_AGEMA_signal_4456), .Q (new_AGEMA_signal_4457) ) ;
    buf_clk new_AGEMA_reg_buffer_2505 ( .C (clk), .D (new_AGEMA_signal_4460), .Q (new_AGEMA_signal_4461) ) ;
    buf_clk new_AGEMA_reg_buffer_2509 ( .C (clk), .D (new_AGEMA_signal_4464), .Q (new_AGEMA_signal_4465) ) ;
    buf_clk new_AGEMA_reg_buffer_2513 ( .C (clk), .D (new_AGEMA_signal_4468), .Q (new_AGEMA_signal_4469) ) ;
    buf_clk new_AGEMA_reg_buffer_2517 ( .C (clk), .D (new_AGEMA_signal_4472), .Q (new_AGEMA_signal_4473) ) ;
    buf_clk new_AGEMA_reg_buffer_2521 ( .C (clk), .D (new_AGEMA_signal_4476), .Q (new_AGEMA_signal_4477) ) ;
    buf_clk new_AGEMA_reg_buffer_2525 ( .C (clk), .D (new_AGEMA_signal_4480), .Q (new_AGEMA_signal_4481) ) ;
    buf_clk new_AGEMA_reg_buffer_2529 ( .C (clk), .D (new_AGEMA_signal_4484), .Q (new_AGEMA_signal_4485) ) ;
    buf_clk new_AGEMA_reg_buffer_2533 ( .C (clk), .D (new_AGEMA_signal_4488), .Q (new_AGEMA_signal_4489) ) ;
    buf_clk new_AGEMA_reg_buffer_2537 ( .C (clk), .D (new_AGEMA_signal_4492), .Q (new_AGEMA_signal_4493) ) ;
    buf_clk new_AGEMA_reg_buffer_2541 ( .C (clk), .D (new_AGEMA_signal_4496), .Q (new_AGEMA_signal_4497) ) ;
    buf_clk new_AGEMA_reg_buffer_2545 ( .C (clk), .D (new_AGEMA_signal_4500), .Q (new_AGEMA_signal_4501) ) ;
    buf_clk new_AGEMA_reg_buffer_2549 ( .C (clk), .D (new_AGEMA_signal_4504), .Q (new_AGEMA_signal_4505) ) ;
    buf_clk new_AGEMA_reg_buffer_2553 ( .C (clk), .D (new_AGEMA_signal_4508), .Q (new_AGEMA_signal_4509) ) ;
    buf_clk new_AGEMA_reg_buffer_2557 ( .C (clk), .D (new_AGEMA_signal_4512), .Q (new_AGEMA_signal_4513) ) ;
    buf_clk new_AGEMA_reg_buffer_2561 ( .C (clk), .D (new_AGEMA_signal_4516), .Q (new_AGEMA_signal_4517) ) ;
    buf_clk new_AGEMA_reg_buffer_2565 ( .C (clk), .D (new_AGEMA_signal_4520), .Q (new_AGEMA_signal_4521) ) ;
    buf_clk new_AGEMA_reg_buffer_2569 ( .C (clk), .D (new_AGEMA_signal_4524), .Q (new_AGEMA_signal_4525) ) ;
    buf_clk new_AGEMA_reg_buffer_2573 ( .C (clk), .D (new_AGEMA_signal_4528), .Q (new_AGEMA_signal_4529) ) ;
    buf_clk new_AGEMA_reg_buffer_2577 ( .C (clk), .D (new_AGEMA_signal_4532), .Q (new_AGEMA_signal_4533) ) ;
    buf_clk new_AGEMA_reg_buffer_2581 ( .C (clk), .D (new_AGEMA_signal_4536), .Q (new_AGEMA_signal_4537) ) ;
    buf_clk new_AGEMA_reg_buffer_2585 ( .C (clk), .D (new_AGEMA_signal_4540), .Q (new_AGEMA_signal_4541) ) ;
    buf_clk new_AGEMA_reg_buffer_2589 ( .C (clk), .D (new_AGEMA_signal_4544), .Q (new_AGEMA_signal_4545) ) ;
    buf_clk new_AGEMA_reg_buffer_2593 ( .C (clk), .D (new_AGEMA_signal_4548), .Q (new_AGEMA_signal_4549) ) ;
    buf_clk new_AGEMA_reg_buffer_2597 ( .C (clk), .D (new_AGEMA_signal_4552), .Q (new_AGEMA_signal_4553) ) ;
    buf_clk new_AGEMA_reg_buffer_2601 ( .C (clk), .D (new_AGEMA_signal_4556), .Q (new_AGEMA_signal_4557) ) ;
    buf_clk new_AGEMA_reg_buffer_2605 ( .C (clk), .D (new_AGEMA_signal_4560), .Q (new_AGEMA_signal_4561) ) ;
    buf_clk new_AGEMA_reg_buffer_2609 ( .C (clk), .D (new_AGEMA_signal_4564), .Q (new_AGEMA_signal_4565) ) ;
    buf_clk new_AGEMA_reg_buffer_2613 ( .C (clk), .D (new_AGEMA_signal_4568), .Q (new_AGEMA_signal_4569) ) ;
    buf_clk new_AGEMA_reg_buffer_2617 ( .C (clk), .D (new_AGEMA_signal_4572), .Q (new_AGEMA_signal_4573) ) ;
    buf_clk new_AGEMA_reg_buffer_2621 ( .C (clk), .D (new_AGEMA_signal_4576), .Q (new_AGEMA_signal_4577) ) ;
    buf_clk new_AGEMA_reg_buffer_2625 ( .C (clk), .D (new_AGEMA_signal_4580), .Q (new_AGEMA_signal_4581) ) ;
    buf_clk new_AGEMA_reg_buffer_2629 ( .C (clk), .D (new_AGEMA_signal_4584), .Q (new_AGEMA_signal_4585) ) ;
    buf_clk new_AGEMA_reg_buffer_2633 ( .C (clk), .D (new_AGEMA_signal_4588), .Q (new_AGEMA_signal_4589) ) ;
    buf_clk new_AGEMA_reg_buffer_2637 ( .C (clk), .D (new_AGEMA_signal_4592), .Q (new_AGEMA_signal_4593) ) ;
    buf_clk new_AGEMA_reg_buffer_2641 ( .C (clk), .D (new_AGEMA_signal_4596), .Q (new_AGEMA_signal_4597) ) ;
    buf_clk new_AGEMA_reg_buffer_2645 ( .C (clk), .D (new_AGEMA_signal_4600), .Q (new_AGEMA_signal_4601) ) ;
    buf_clk new_AGEMA_reg_buffer_2649 ( .C (clk), .D (new_AGEMA_signal_4604), .Q (new_AGEMA_signal_4605) ) ;
    buf_clk new_AGEMA_reg_buffer_2653 ( .C (clk), .D (new_AGEMA_signal_4608), .Q (new_AGEMA_signal_4609) ) ;
    buf_clk new_AGEMA_reg_buffer_2657 ( .C (clk), .D (new_AGEMA_signal_4612), .Q (new_AGEMA_signal_4613) ) ;
    buf_clk new_AGEMA_reg_buffer_2661 ( .C (clk), .D (new_AGEMA_signal_4616), .Q (new_AGEMA_signal_4617) ) ;
    buf_clk new_AGEMA_reg_buffer_2665 ( .C (clk), .D (new_AGEMA_signal_4620), .Q (new_AGEMA_signal_4621) ) ;
    buf_clk new_AGEMA_reg_buffer_2669 ( .C (clk), .D (new_AGEMA_signal_4624), .Q (new_AGEMA_signal_4625) ) ;
    buf_clk new_AGEMA_reg_buffer_2673 ( .C (clk), .D (new_AGEMA_signal_4628), .Q (new_AGEMA_signal_4629) ) ;
    buf_clk new_AGEMA_reg_buffer_2677 ( .C (clk), .D (new_AGEMA_signal_4632), .Q (new_AGEMA_signal_4633) ) ;
    buf_clk new_AGEMA_reg_buffer_2681 ( .C (clk), .D (new_AGEMA_signal_4636), .Q (new_AGEMA_signal_4637) ) ;
    buf_clk new_AGEMA_reg_buffer_2685 ( .C (clk), .D (new_AGEMA_signal_4640), .Q (new_AGEMA_signal_4641) ) ;
    buf_clk new_AGEMA_reg_buffer_2689 ( .C (clk), .D (new_AGEMA_signal_4644), .Q (new_AGEMA_signal_4645) ) ;
    buf_clk new_AGEMA_reg_buffer_2693 ( .C (clk), .D (new_AGEMA_signal_4648), .Q (new_AGEMA_signal_4649) ) ;
    buf_clk new_AGEMA_reg_buffer_2697 ( .C (clk), .D (new_AGEMA_signal_4652), .Q (new_AGEMA_signal_4653) ) ;
    buf_clk new_AGEMA_reg_buffer_2701 ( .C (clk), .D (new_AGEMA_signal_4656), .Q (new_AGEMA_signal_4657) ) ;
    buf_clk new_AGEMA_reg_buffer_2705 ( .C (clk), .D (new_AGEMA_signal_4660), .Q (new_AGEMA_signal_4661) ) ;
    buf_clk new_AGEMA_reg_buffer_2709 ( .C (clk), .D (new_AGEMA_signal_4664), .Q (new_AGEMA_signal_4665) ) ;
    buf_clk new_AGEMA_reg_buffer_2713 ( .C (clk), .D (new_AGEMA_signal_4668), .Q (new_AGEMA_signal_4669) ) ;
    buf_clk new_AGEMA_reg_buffer_2717 ( .C (clk), .D (new_AGEMA_signal_4672), .Q (new_AGEMA_signal_4673) ) ;
    buf_clk new_AGEMA_reg_buffer_2721 ( .C (clk), .D (new_AGEMA_signal_4676), .Q (new_AGEMA_signal_4677) ) ;
    buf_clk new_AGEMA_reg_buffer_2725 ( .C (clk), .D (new_AGEMA_signal_4680), .Q (new_AGEMA_signal_4681) ) ;
    buf_clk new_AGEMA_reg_buffer_2729 ( .C (clk), .D (new_AGEMA_signal_4684), .Q (new_AGEMA_signal_4685) ) ;
    buf_clk new_AGEMA_reg_buffer_2733 ( .C (clk), .D (new_AGEMA_signal_4688), .Q (new_AGEMA_signal_4689) ) ;
    buf_clk new_AGEMA_reg_buffer_2737 ( .C (clk), .D (new_AGEMA_signal_4692), .Q (new_AGEMA_signal_4693) ) ;
    buf_clk new_AGEMA_reg_buffer_2741 ( .C (clk), .D (new_AGEMA_signal_4696), .Q (new_AGEMA_signal_4697) ) ;
    buf_clk new_AGEMA_reg_buffer_2745 ( .C (clk), .D (new_AGEMA_signal_4700), .Q (new_AGEMA_signal_4701) ) ;
    buf_clk new_AGEMA_reg_buffer_2749 ( .C (clk), .D (new_AGEMA_signal_4704), .Q (new_AGEMA_signal_4705) ) ;
    buf_clk new_AGEMA_reg_buffer_2753 ( .C (clk), .D (new_AGEMA_signal_4708), .Q (new_AGEMA_signal_4709) ) ;
    buf_clk new_AGEMA_reg_buffer_2757 ( .C (clk), .D (new_AGEMA_signal_4712), .Q (new_AGEMA_signal_4713) ) ;
    buf_clk new_AGEMA_reg_buffer_2761 ( .C (clk), .D (new_AGEMA_signal_4716), .Q (new_AGEMA_signal_4717) ) ;
    buf_clk new_AGEMA_reg_buffer_2765 ( .C (clk), .D (new_AGEMA_signal_4720), .Q (new_AGEMA_signal_4721) ) ;
    buf_clk new_AGEMA_reg_buffer_2769 ( .C (clk), .D (new_AGEMA_signal_4724), .Q (new_AGEMA_signal_4725) ) ;
    buf_clk new_AGEMA_reg_buffer_2773 ( .C (clk), .D (new_AGEMA_signal_4728), .Q (new_AGEMA_signal_4729) ) ;
    buf_clk new_AGEMA_reg_buffer_2777 ( .C (clk), .D (new_AGEMA_signal_4732), .Q (new_AGEMA_signal_4733) ) ;
    buf_clk new_AGEMA_reg_buffer_2781 ( .C (clk), .D (new_AGEMA_signal_4736), .Q (new_AGEMA_signal_4737) ) ;
    buf_clk new_AGEMA_reg_buffer_2785 ( .C (clk), .D (new_AGEMA_signal_4740), .Q (new_AGEMA_signal_4741) ) ;
    buf_clk new_AGEMA_reg_buffer_2789 ( .C (clk), .D (new_AGEMA_signal_4744), .Q (new_AGEMA_signal_4745) ) ;
    buf_clk new_AGEMA_reg_buffer_2793 ( .C (clk), .D (new_AGEMA_signal_4748), .Q (new_AGEMA_signal_4749) ) ;
    buf_clk new_AGEMA_reg_buffer_2797 ( .C (clk), .D (new_AGEMA_signal_4752), .Q (new_AGEMA_signal_4753) ) ;
    buf_clk new_AGEMA_reg_buffer_2801 ( .C (clk), .D (new_AGEMA_signal_4756), .Q (new_AGEMA_signal_4757) ) ;
    buf_clk new_AGEMA_reg_buffer_2805 ( .C (clk), .D (new_AGEMA_signal_4760), .Q (new_AGEMA_signal_4761) ) ;
    buf_clk new_AGEMA_reg_buffer_2809 ( .C (clk), .D (new_AGEMA_signal_4764), .Q (new_AGEMA_signal_4765) ) ;
    buf_clk new_AGEMA_reg_buffer_2813 ( .C (clk), .D (new_AGEMA_signal_4768), .Q (new_AGEMA_signal_4769) ) ;
    buf_clk new_AGEMA_reg_buffer_2817 ( .C (clk), .D (new_AGEMA_signal_4772), .Q (new_AGEMA_signal_4773) ) ;
    buf_clk new_AGEMA_reg_buffer_2821 ( .C (clk), .D (new_AGEMA_signal_4776), .Q (new_AGEMA_signal_4777) ) ;
    buf_clk new_AGEMA_reg_buffer_2825 ( .C (clk), .D (new_AGEMA_signal_4780), .Q (new_AGEMA_signal_4781) ) ;
    buf_clk new_AGEMA_reg_buffer_2829 ( .C (clk), .D (new_AGEMA_signal_4784), .Q (new_AGEMA_signal_4785) ) ;
    buf_clk new_AGEMA_reg_buffer_2833 ( .C (clk), .D (new_AGEMA_signal_4788), .Q (new_AGEMA_signal_4789) ) ;
    buf_clk new_AGEMA_reg_buffer_2837 ( .C (clk), .D (new_AGEMA_signal_4792), .Q (new_AGEMA_signal_4793) ) ;
    buf_clk new_AGEMA_reg_buffer_2841 ( .C (clk), .D (new_AGEMA_signal_4796), .Q (new_AGEMA_signal_4797) ) ;
    buf_clk new_AGEMA_reg_buffer_2845 ( .C (clk), .D (new_AGEMA_signal_4800), .Q (new_AGEMA_signal_4801) ) ;
    buf_clk new_AGEMA_reg_buffer_2849 ( .C (clk), .D (new_AGEMA_signal_4804), .Q (new_AGEMA_signal_4805) ) ;
    buf_clk new_AGEMA_reg_buffer_2853 ( .C (clk), .D (new_AGEMA_signal_4808), .Q (new_AGEMA_signal_4809) ) ;
    buf_clk new_AGEMA_reg_buffer_2857 ( .C (clk), .D (new_AGEMA_signal_4812), .Q (new_AGEMA_signal_4813) ) ;
    buf_clk new_AGEMA_reg_buffer_2861 ( .C (clk), .D (new_AGEMA_signal_4816), .Q (new_AGEMA_signal_4817) ) ;
    buf_clk new_AGEMA_reg_buffer_2865 ( .C (clk), .D (new_AGEMA_signal_4820), .Q (new_AGEMA_signal_4821) ) ;
    buf_clk new_AGEMA_reg_buffer_2869 ( .C (clk), .D (new_AGEMA_signal_4824), .Q (new_AGEMA_signal_4825) ) ;
    buf_clk new_AGEMA_reg_buffer_2873 ( .C (clk), .D (new_AGEMA_signal_4828), .Q (new_AGEMA_signal_4829) ) ;
    buf_clk new_AGEMA_reg_buffer_2877 ( .C (clk), .D (new_AGEMA_signal_4832), .Q (new_AGEMA_signal_4833) ) ;
    buf_clk new_AGEMA_reg_buffer_2881 ( .C (clk), .D (new_AGEMA_signal_4836), .Q (new_AGEMA_signal_4837) ) ;
    buf_clk new_AGEMA_reg_buffer_2885 ( .C (clk), .D (new_AGEMA_signal_4840), .Q (new_AGEMA_signal_4841) ) ;
    buf_clk new_AGEMA_reg_buffer_2889 ( .C (clk), .D (new_AGEMA_signal_4844), .Q (new_AGEMA_signal_4845) ) ;
    buf_clk new_AGEMA_reg_buffer_2893 ( .C (clk), .D (new_AGEMA_signal_4848), .Q (new_AGEMA_signal_4849) ) ;
    buf_clk new_AGEMA_reg_buffer_2897 ( .C (clk), .D (new_AGEMA_signal_4852), .Q (new_AGEMA_signal_4853) ) ;
    buf_clk new_AGEMA_reg_buffer_2901 ( .C (clk), .D (new_AGEMA_signal_4856), .Q (new_AGEMA_signal_4857) ) ;
    buf_clk new_AGEMA_reg_buffer_2905 ( .C (clk), .D (new_AGEMA_signal_4860), .Q (new_AGEMA_signal_4861) ) ;
    buf_clk new_AGEMA_reg_buffer_2909 ( .C (clk), .D (new_AGEMA_signal_4864), .Q (new_AGEMA_signal_4865) ) ;
    buf_clk new_AGEMA_reg_buffer_2913 ( .C (clk), .D (new_AGEMA_signal_4868), .Q (new_AGEMA_signal_4869) ) ;
    buf_clk new_AGEMA_reg_buffer_2917 ( .C (clk), .D (new_AGEMA_signal_4872), .Q (new_AGEMA_signal_4873) ) ;
    buf_clk new_AGEMA_reg_buffer_2921 ( .C (clk), .D (new_AGEMA_signal_4876), .Q (new_AGEMA_signal_4877) ) ;
    buf_clk new_AGEMA_reg_buffer_2925 ( .C (clk), .D (new_AGEMA_signal_4880), .Q (new_AGEMA_signal_4881) ) ;
    buf_clk new_AGEMA_reg_buffer_2929 ( .C (clk), .D (new_AGEMA_signal_4884), .Q (new_AGEMA_signal_4885) ) ;
    buf_clk new_AGEMA_reg_buffer_2933 ( .C (clk), .D (new_AGEMA_signal_4888), .Q (new_AGEMA_signal_4889) ) ;
    buf_clk new_AGEMA_reg_buffer_2937 ( .C (clk), .D (new_AGEMA_signal_4892), .Q (new_AGEMA_signal_4893) ) ;
    buf_clk new_AGEMA_reg_buffer_2941 ( .C (clk), .D (new_AGEMA_signal_4896), .Q (new_AGEMA_signal_4897) ) ;
    buf_clk new_AGEMA_reg_buffer_2945 ( .C (clk), .D (new_AGEMA_signal_4900), .Q (new_AGEMA_signal_4901) ) ;
    buf_clk new_AGEMA_reg_buffer_2949 ( .C (clk), .D (new_AGEMA_signal_4904), .Q (new_AGEMA_signal_4905) ) ;
    buf_clk new_AGEMA_reg_buffer_2953 ( .C (clk), .D (new_AGEMA_signal_4908), .Q (new_AGEMA_signal_4909) ) ;
    buf_clk new_AGEMA_reg_buffer_2957 ( .C (clk), .D (new_AGEMA_signal_4912), .Q (new_AGEMA_signal_4913) ) ;
    buf_clk new_AGEMA_reg_buffer_2961 ( .C (clk), .D (new_AGEMA_signal_4916), .Q (new_AGEMA_signal_4917) ) ;
    buf_clk new_AGEMA_reg_buffer_2965 ( .C (clk), .D (new_AGEMA_signal_4920), .Q (new_AGEMA_signal_4921) ) ;
    buf_clk new_AGEMA_reg_buffer_2969 ( .C (clk), .D (new_AGEMA_signal_4924), .Q (new_AGEMA_signal_4925) ) ;
    buf_clk new_AGEMA_reg_buffer_2973 ( .C (clk), .D (new_AGEMA_signal_4928), .Q (new_AGEMA_signal_4929) ) ;
    buf_clk new_AGEMA_reg_buffer_2977 ( .C (clk), .D (new_AGEMA_signal_4932), .Q (new_AGEMA_signal_4933) ) ;
    buf_clk new_AGEMA_reg_buffer_2981 ( .C (clk), .D (new_AGEMA_signal_4936), .Q (new_AGEMA_signal_4937) ) ;
    buf_clk new_AGEMA_reg_buffer_2985 ( .C (clk), .D (new_AGEMA_signal_4940), .Q (new_AGEMA_signal_4941) ) ;
    buf_clk new_AGEMA_reg_buffer_2989 ( .C (clk), .D (new_AGEMA_signal_4944), .Q (new_AGEMA_signal_4945) ) ;
    buf_clk new_AGEMA_reg_buffer_2993 ( .C (clk), .D (new_AGEMA_signal_4948), .Q (new_AGEMA_signal_4949) ) ;
    buf_clk new_AGEMA_reg_buffer_2997 ( .C (clk), .D (new_AGEMA_signal_4952), .Q (new_AGEMA_signal_4953) ) ;
    buf_clk new_AGEMA_reg_buffer_3001 ( .C (clk), .D (new_AGEMA_signal_4956), .Q (new_AGEMA_signal_4957) ) ;
    buf_clk new_AGEMA_reg_buffer_3005 ( .C (clk), .D (new_AGEMA_signal_4960), .Q (new_AGEMA_signal_4961) ) ;
    buf_clk new_AGEMA_reg_buffer_3009 ( .C (clk), .D (new_AGEMA_signal_4964), .Q (new_AGEMA_signal_4965) ) ;
    buf_clk new_AGEMA_reg_buffer_3013 ( .C (clk), .D (new_AGEMA_signal_4968), .Q (new_AGEMA_signal_4969) ) ;
    buf_clk new_AGEMA_reg_buffer_3017 ( .C (clk), .D (new_AGEMA_signal_4972), .Q (new_AGEMA_signal_4973) ) ;
    buf_clk new_AGEMA_reg_buffer_3021 ( .C (clk), .D (new_AGEMA_signal_4976), .Q (new_AGEMA_signal_4977) ) ;
    buf_clk new_AGEMA_reg_buffer_3025 ( .C (clk), .D (new_AGEMA_signal_4980), .Q (new_AGEMA_signal_4981) ) ;
    buf_clk new_AGEMA_reg_buffer_3029 ( .C (clk), .D (new_AGEMA_signal_4984), .Q (new_AGEMA_signal_4985) ) ;
    buf_clk new_AGEMA_reg_buffer_3033 ( .C (clk), .D (new_AGEMA_signal_4988), .Q (new_AGEMA_signal_4989) ) ;
    buf_clk new_AGEMA_reg_buffer_3037 ( .C (clk), .D (new_AGEMA_signal_4992), .Q (new_AGEMA_signal_4993) ) ;
    buf_clk new_AGEMA_reg_buffer_3041 ( .C (clk), .D (new_AGEMA_signal_4996), .Q (new_AGEMA_signal_4997) ) ;
    buf_clk new_AGEMA_reg_buffer_3045 ( .C (clk), .D (new_AGEMA_signal_5000), .Q (new_AGEMA_signal_5001) ) ;
    buf_clk new_AGEMA_reg_buffer_3049 ( .C (clk), .D (new_AGEMA_signal_5004), .Q (new_AGEMA_signal_5005) ) ;
    buf_clk new_AGEMA_reg_buffer_3053 ( .C (clk), .D (new_AGEMA_signal_5008), .Q (new_AGEMA_signal_5009) ) ;
    buf_clk new_AGEMA_reg_buffer_3057 ( .C (clk), .D (new_AGEMA_signal_5012), .Q (new_AGEMA_signal_5013) ) ;
    buf_clk new_AGEMA_reg_buffer_3061 ( .C (clk), .D (new_AGEMA_signal_5016), .Q (new_AGEMA_signal_5017) ) ;
    buf_clk new_AGEMA_reg_buffer_3065 ( .C (clk), .D (new_AGEMA_signal_5020), .Q (new_AGEMA_signal_5021) ) ;
    buf_clk new_AGEMA_reg_buffer_3069 ( .C (clk), .D (new_AGEMA_signal_5024), .Q (new_AGEMA_signal_5025) ) ;
    buf_clk new_AGEMA_reg_buffer_3073 ( .C (clk), .D (new_AGEMA_signal_5028), .Q (new_AGEMA_signal_5029) ) ;
    buf_clk new_AGEMA_reg_buffer_3077 ( .C (clk), .D (new_AGEMA_signal_5032), .Q (new_AGEMA_signal_5033) ) ;
    buf_clk new_AGEMA_reg_buffer_3081 ( .C (clk), .D (new_AGEMA_signal_5036), .Q (new_AGEMA_signal_5037) ) ;
    buf_clk new_AGEMA_reg_buffer_3085 ( .C (clk), .D (new_AGEMA_signal_5040), .Q (new_AGEMA_signal_5041) ) ;
    buf_clk new_AGEMA_reg_buffer_3089 ( .C (clk), .D (new_AGEMA_signal_5044), .Q (new_AGEMA_signal_5045) ) ;
    buf_clk new_AGEMA_reg_buffer_3093 ( .C (clk), .D (new_AGEMA_signal_5048), .Q (new_AGEMA_signal_5049) ) ;
    buf_clk new_AGEMA_reg_buffer_3097 ( .C (clk), .D (new_AGEMA_signal_5052), .Q (new_AGEMA_signal_5053) ) ;
    buf_clk new_AGEMA_reg_buffer_3101 ( .C (clk), .D (new_AGEMA_signal_5056), .Q (new_AGEMA_signal_5057) ) ;
    buf_clk new_AGEMA_reg_buffer_3105 ( .C (clk), .D (new_AGEMA_signal_5060), .Q (new_AGEMA_signal_5061) ) ;
    buf_clk new_AGEMA_reg_buffer_3109 ( .C (clk), .D (new_AGEMA_signal_5064), .Q (new_AGEMA_signal_5065) ) ;
    buf_clk new_AGEMA_reg_buffer_3113 ( .C (clk), .D (new_AGEMA_signal_5068), .Q (new_AGEMA_signal_5069) ) ;
    buf_clk new_AGEMA_reg_buffer_3117 ( .C (clk), .D (new_AGEMA_signal_5072), .Q (new_AGEMA_signal_5073) ) ;
    buf_clk new_AGEMA_reg_buffer_3121 ( .C (clk), .D (new_AGEMA_signal_5076), .Q (new_AGEMA_signal_5077) ) ;
    buf_clk new_AGEMA_reg_buffer_3125 ( .C (clk), .D (new_AGEMA_signal_5080), .Q (new_AGEMA_signal_5081) ) ;
    buf_clk new_AGEMA_reg_buffer_3129 ( .C (clk), .D (new_AGEMA_signal_5084), .Q (new_AGEMA_signal_5085) ) ;
    buf_clk new_AGEMA_reg_buffer_3133 ( .C (clk), .D (new_AGEMA_signal_5088), .Q (new_AGEMA_signal_5089) ) ;
    buf_clk new_AGEMA_reg_buffer_3137 ( .C (clk), .D (new_AGEMA_signal_5092), .Q (new_AGEMA_signal_5093) ) ;
    buf_clk new_AGEMA_reg_buffer_3141 ( .C (clk), .D (new_AGEMA_signal_5096), .Q (new_AGEMA_signal_5097) ) ;
    buf_clk new_AGEMA_reg_buffer_3145 ( .C (clk), .D (new_AGEMA_signal_5100), .Q (new_AGEMA_signal_5101) ) ;
    buf_clk new_AGEMA_reg_buffer_3149 ( .C (clk), .D (new_AGEMA_signal_5104), .Q (new_AGEMA_signal_5105) ) ;
    buf_clk new_AGEMA_reg_buffer_3153 ( .C (clk), .D (new_AGEMA_signal_5108), .Q (new_AGEMA_signal_5109) ) ;
    buf_clk new_AGEMA_reg_buffer_3157 ( .C (clk), .D (new_AGEMA_signal_5112), .Q (new_AGEMA_signal_5113) ) ;
    buf_clk new_AGEMA_reg_buffer_3161 ( .C (clk), .D (new_AGEMA_signal_5116), .Q (new_AGEMA_signal_5117) ) ;
    buf_clk new_AGEMA_reg_buffer_3165 ( .C (clk), .D (new_AGEMA_signal_5120), .Q (new_AGEMA_signal_5121) ) ;
    buf_clk new_AGEMA_reg_buffer_3169 ( .C (clk), .D (new_AGEMA_signal_5124), .Q (new_AGEMA_signal_5125) ) ;
    buf_clk new_AGEMA_reg_buffer_3173 ( .C (clk), .D (new_AGEMA_signal_5128), .Q (new_AGEMA_signal_5129) ) ;
    buf_clk new_AGEMA_reg_buffer_3177 ( .C (clk), .D (new_AGEMA_signal_5132), .Q (new_AGEMA_signal_5133) ) ;
    buf_clk new_AGEMA_reg_buffer_3181 ( .C (clk), .D (new_AGEMA_signal_5136), .Q (new_AGEMA_signal_5137) ) ;
    buf_clk new_AGEMA_reg_buffer_3185 ( .C (clk), .D (new_AGEMA_signal_5140), .Q (new_AGEMA_signal_5141) ) ;
    buf_clk new_AGEMA_reg_buffer_3189 ( .C (clk), .D (new_AGEMA_signal_5144), .Q (new_AGEMA_signal_5145) ) ;
    buf_clk new_AGEMA_reg_buffer_3193 ( .C (clk), .D (new_AGEMA_signal_5148), .Q (new_AGEMA_signal_5149) ) ;
    buf_clk new_AGEMA_reg_buffer_3197 ( .C (clk), .D (new_AGEMA_signal_5152), .Q (new_AGEMA_signal_5153) ) ;
    buf_clk new_AGEMA_reg_buffer_3201 ( .C (clk), .D (new_AGEMA_signal_5156), .Q (new_AGEMA_signal_5157) ) ;
    buf_clk new_AGEMA_reg_buffer_3205 ( .C (clk), .D (new_AGEMA_signal_5160), .Q (new_AGEMA_signal_5161) ) ;
    buf_clk new_AGEMA_reg_buffer_3209 ( .C (clk), .D (new_AGEMA_signal_5164), .Q (new_AGEMA_signal_5165) ) ;
    buf_clk new_AGEMA_reg_buffer_3213 ( .C (clk), .D (new_AGEMA_signal_5168), .Q (new_AGEMA_signal_5169) ) ;
    buf_clk new_AGEMA_reg_buffer_3217 ( .C (clk), .D (new_AGEMA_signal_5172), .Q (new_AGEMA_signal_5173) ) ;
    buf_clk new_AGEMA_reg_buffer_3221 ( .C (clk), .D (new_AGEMA_signal_5176), .Q (new_AGEMA_signal_5177) ) ;
    buf_clk new_AGEMA_reg_buffer_3225 ( .C (clk), .D (new_AGEMA_signal_5180), .Q (new_AGEMA_signal_5181) ) ;
    buf_clk new_AGEMA_reg_buffer_3229 ( .C (clk), .D (new_AGEMA_signal_5184), .Q (new_AGEMA_signal_5185) ) ;
    buf_clk new_AGEMA_reg_buffer_3233 ( .C (clk), .D (new_AGEMA_signal_5188), .Q (new_AGEMA_signal_5189) ) ;
    buf_clk new_AGEMA_reg_buffer_3237 ( .C (clk), .D (new_AGEMA_signal_5192), .Q (new_AGEMA_signal_5193) ) ;
    buf_clk new_AGEMA_reg_buffer_3241 ( .C (clk), .D (new_AGEMA_signal_5196), .Q (new_AGEMA_signal_5197) ) ;
    buf_clk new_AGEMA_reg_buffer_3245 ( .C (clk), .D (new_AGEMA_signal_5200), .Q (new_AGEMA_signal_5201) ) ;
    buf_clk new_AGEMA_reg_buffer_3249 ( .C (clk), .D (new_AGEMA_signal_5204), .Q (new_AGEMA_signal_5205) ) ;
    buf_clk new_AGEMA_reg_buffer_3253 ( .C (clk), .D (new_AGEMA_signal_5208), .Q (new_AGEMA_signal_5209) ) ;
    buf_clk new_AGEMA_reg_buffer_3257 ( .C (clk), .D (new_AGEMA_signal_5212), .Q (new_AGEMA_signal_5213) ) ;
    buf_clk new_AGEMA_reg_buffer_3261 ( .C (clk), .D (new_AGEMA_signal_5216), .Q (new_AGEMA_signal_5217) ) ;
    buf_clk new_AGEMA_reg_buffer_3265 ( .C (clk), .D (new_AGEMA_signal_5220), .Q (new_AGEMA_signal_5221) ) ;
    buf_clk new_AGEMA_reg_buffer_3269 ( .C (clk), .D (new_AGEMA_signal_5224), .Q (new_AGEMA_signal_5225) ) ;
    buf_clk new_AGEMA_reg_buffer_3273 ( .C (clk), .D (new_AGEMA_signal_5228), .Q (new_AGEMA_signal_5229) ) ;
    buf_clk new_AGEMA_reg_buffer_3277 ( .C (clk), .D (new_AGEMA_signal_5232), .Q (new_AGEMA_signal_5233) ) ;
    buf_clk new_AGEMA_reg_buffer_3281 ( .C (clk), .D (new_AGEMA_signal_5236), .Q (new_AGEMA_signal_5237) ) ;
    buf_clk new_AGEMA_reg_buffer_3285 ( .C (clk), .D (new_AGEMA_signal_5240), .Q (new_AGEMA_signal_5241) ) ;
    buf_clk new_AGEMA_reg_buffer_3289 ( .C (clk), .D (new_AGEMA_signal_5244), .Q (new_AGEMA_signal_5245) ) ;
    buf_clk new_AGEMA_reg_buffer_3293 ( .C (clk), .D (new_AGEMA_signal_5248), .Q (new_AGEMA_signal_5249) ) ;
    buf_clk new_AGEMA_reg_buffer_3297 ( .C (clk), .D (new_AGEMA_signal_5252), .Q (new_AGEMA_signal_5253) ) ;
    buf_clk new_AGEMA_reg_buffer_3301 ( .C (clk), .D (new_AGEMA_signal_5256), .Q (new_AGEMA_signal_5257) ) ;
    buf_clk new_AGEMA_reg_buffer_3305 ( .C (clk), .D (new_AGEMA_signal_5260), .Q (new_AGEMA_signal_5261) ) ;
    buf_clk new_AGEMA_reg_buffer_3309 ( .C (clk), .D (new_AGEMA_signal_5264), .Q (new_AGEMA_signal_5265) ) ;
    buf_clk new_AGEMA_reg_buffer_3313 ( .C (clk), .D (new_AGEMA_signal_5268), .Q (new_AGEMA_signal_5269) ) ;
    buf_clk new_AGEMA_reg_buffer_3317 ( .C (clk), .D (new_AGEMA_signal_5272), .Q (new_AGEMA_signal_5273) ) ;
    buf_clk new_AGEMA_reg_buffer_3321 ( .C (clk), .D (new_AGEMA_signal_5276), .Q (new_AGEMA_signal_5277) ) ;
    buf_clk new_AGEMA_reg_buffer_3325 ( .C (clk), .D (new_AGEMA_signal_5280), .Q (new_AGEMA_signal_5281) ) ;
    buf_clk new_AGEMA_reg_buffer_3329 ( .C (clk), .D (new_AGEMA_signal_5284), .Q (new_AGEMA_signal_5285) ) ;
    buf_clk new_AGEMA_reg_buffer_3333 ( .C (clk), .D (new_AGEMA_signal_5288), .Q (new_AGEMA_signal_5289) ) ;
    buf_clk new_AGEMA_reg_buffer_3337 ( .C (clk), .D (new_AGEMA_signal_5292), .Q (new_AGEMA_signal_5293) ) ;
    buf_clk new_AGEMA_reg_buffer_3341 ( .C (clk), .D (new_AGEMA_signal_5296), .Q (new_AGEMA_signal_5297) ) ;
    buf_clk new_AGEMA_reg_buffer_3345 ( .C (clk), .D (new_AGEMA_signal_5300), .Q (new_AGEMA_signal_5301) ) ;
    buf_clk new_AGEMA_reg_buffer_3349 ( .C (clk), .D (new_AGEMA_signal_5304), .Q (new_AGEMA_signal_5305) ) ;
    buf_clk new_AGEMA_reg_buffer_3353 ( .C (clk), .D (new_AGEMA_signal_5308), .Q (new_AGEMA_signal_5309) ) ;
    buf_clk new_AGEMA_reg_buffer_3357 ( .C (clk), .D (new_AGEMA_signal_5312), .Q (new_AGEMA_signal_5313) ) ;
    buf_clk new_AGEMA_reg_buffer_3361 ( .C (clk), .D (new_AGEMA_signal_5316), .Q (new_AGEMA_signal_5317) ) ;
    buf_clk new_AGEMA_reg_buffer_3365 ( .C (clk), .D (new_AGEMA_signal_5320), .Q (new_AGEMA_signal_5321) ) ;
    buf_clk new_AGEMA_reg_buffer_3369 ( .C (clk), .D (new_AGEMA_signal_5324), .Q (new_AGEMA_signal_5325) ) ;
    buf_clk new_AGEMA_reg_buffer_3373 ( .C (clk), .D (new_AGEMA_signal_5328), .Q (new_AGEMA_signal_5329) ) ;
    buf_clk new_AGEMA_reg_buffer_3377 ( .C (clk), .D (new_AGEMA_signal_5332), .Q (new_AGEMA_signal_5333) ) ;
    buf_clk new_AGEMA_reg_buffer_3381 ( .C (clk), .D (new_AGEMA_signal_5336), .Q (new_AGEMA_signal_5337) ) ;
    buf_clk new_AGEMA_reg_buffer_3385 ( .C (clk), .D (new_AGEMA_signal_5340), .Q (new_AGEMA_signal_5341) ) ;
    buf_clk new_AGEMA_reg_buffer_3389 ( .C (clk), .D (new_AGEMA_signal_5344), .Q (new_AGEMA_signal_5345) ) ;
    buf_clk new_AGEMA_reg_buffer_3393 ( .C (clk), .D (new_AGEMA_signal_5348), .Q (new_AGEMA_signal_5349) ) ;
    buf_clk new_AGEMA_reg_buffer_3397 ( .C (clk), .D (new_AGEMA_signal_5352), .Q (new_AGEMA_signal_5353) ) ;
    buf_clk new_AGEMA_reg_buffer_3401 ( .C (clk), .D (new_AGEMA_signal_5356), .Q (new_AGEMA_signal_5357) ) ;
    buf_clk new_AGEMA_reg_buffer_3405 ( .C (clk), .D (new_AGEMA_signal_5360), .Q (new_AGEMA_signal_5361) ) ;
    buf_clk new_AGEMA_reg_buffer_3409 ( .C (clk), .D (new_AGEMA_signal_5364), .Q (new_AGEMA_signal_5365) ) ;
    buf_clk new_AGEMA_reg_buffer_3413 ( .C (clk), .D (new_AGEMA_signal_5368), .Q (new_AGEMA_signal_5369) ) ;
    buf_clk new_AGEMA_reg_buffer_3417 ( .C (clk), .D (new_AGEMA_signal_5372), .Q (new_AGEMA_signal_5373) ) ;
    buf_clk new_AGEMA_reg_buffer_3421 ( .C (clk), .D (new_AGEMA_signal_5376), .Q (new_AGEMA_signal_5377) ) ;
    buf_clk new_AGEMA_reg_buffer_3425 ( .C (clk), .D (new_AGEMA_signal_5380), .Q (new_AGEMA_signal_5381) ) ;
    buf_clk new_AGEMA_reg_buffer_3429 ( .C (clk), .D (new_AGEMA_signal_5384), .Q (new_AGEMA_signal_5385) ) ;
    buf_clk new_AGEMA_reg_buffer_3433 ( .C (clk), .D (new_AGEMA_signal_5388), .Q (new_AGEMA_signal_5389) ) ;
    buf_clk new_AGEMA_reg_buffer_3437 ( .C (clk), .D (new_AGEMA_signal_5392), .Q (new_AGEMA_signal_5393) ) ;
    buf_clk new_AGEMA_reg_buffer_3441 ( .C (clk), .D (new_AGEMA_signal_5396), .Q (new_AGEMA_signal_5397) ) ;
    buf_clk new_AGEMA_reg_buffer_3445 ( .C (clk), .D (new_AGEMA_signal_5400), .Q (new_AGEMA_signal_5401) ) ;
    buf_clk new_AGEMA_reg_buffer_3449 ( .C (clk), .D (new_AGEMA_signal_5404), .Q (new_AGEMA_signal_5405) ) ;
    buf_clk new_AGEMA_reg_buffer_3453 ( .C (clk), .D (new_AGEMA_signal_5408), .Q (new_AGEMA_signal_5409) ) ;
    buf_clk new_AGEMA_reg_buffer_3457 ( .C (clk), .D (new_AGEMA_signal_5412), .Q (new_AGEMA_signal_5413) ) ;
    buf_clk new_AGEMA_reg_buffer_3461 ( .C (clk), .D (new_AGEMA_signal_5416), .Q (new_AGEMA_signal_5417) ) ;
    buf_clk new_AGEMA_reg_buffer_3465 ( .C (clk), .D (new_AGEMA_signal_5420), .Q (new_AGEMA_signal_5421) ) ;
    buf_clk new_AGEMA_reg_buffer_3469 ( .C (clk), .D (new_AGEMA_signal_5424), .Q (new_AGEMA_signal_5425) ) ;
    buf_clk new_AGEMA_reg_buffer_3473 ( .C (clk), .D (new_AGEMA_signal_5428), .Q (new_AGEMA_signal_5429) ) ;
    buf_clk new_AGEMA_reg_buffer_3477 ( .C (clk), .D (new_AGEMA_signal_5432), .Q (new_AGEMA_signal_5433) ) ;
    buf_clk new_AGEMA_reg_buffer_3481 ( .C (clk), .D (new_AGEMA_signal_5436), .Q (new_AGEMA_signal_5437) ) ;
    buf_clk new_AGEMA_reg_buffer_3485 ( .C (clk), .D (new_AGEMA_signal_5440), .Q (new_AGEMA_signal_5441) ) ;
    buf_clk new_AGEMA_reg_buffer_3489 ( .C (clk), .D (new_AGEMA_signal_5444), .Q (new_AGEMA_signal_5445) ) ;
    buf_clk new_AGEMA_reg_buffer_3493 ( .C (clk), .D (new_AGEMA_signal_5448), .Q (new_AGEMA_signal_5449) ) ;
    buf_clk new_AGEMA_reg_buffer_3497 ( .C (clk), .D (new_AGEMA_signal_5452), .Q (new_AGEMA_signal_5453) ) ;
    buf_clk new_AGEMA_reg_buffer_3501 ( .C (clk), .D (new_AGEMA_signal_5456), .Q (new_AGEMA_signal_5457) ) ;
    buf_clk new_AGEMA_reg_buffer_3505 ( .C (clk), .D (new_AGEMA_signal_5460), .Q (new_AGEMA_signal_5461) ) ;
    buf_clk new_AGEMA_reg_buffer_3509 ( .C (clk), .D (new_AGEMA_signal_5464), .Q (new_AGEMA_signal_5465) ) ;
    buf_clk new_AGEMA_reg_buffer_3513 ( .C (clk), .D (new_AGEMA_signal_5468), .Q (new_AGEMA_signal_5469) ) ;
    buf_clk new_AGEMA_reg_buffer_3517 ( .C (clk), .D (new_AGEMA_signal_5472), .Q (new_AGEMA_signal_5473) ) ;
    buf_clk new_AGEMA_reg_buffer_3521 ( .C (clk), .D (new_AGEMA_signal_5476), .Q (new_AGEMA_signal_5477) ) ;
    buf_clk new_AGEMA_reg_buffer_3525 ( .C (clk), .D (new_AGEMA_signal_5480), .Q (new_AGEMA_signal_5481) ) ;
    buf_clk new_AGEMA_reg_buffer_3529 ( .C (clk), .D (new_AGEMA_signal_5484), .Q (new_AGEMA_signal_5485) ) ;
    buf_clk new_AGEMA_reg_buffer_3533 ( .C (clk), .D (new_AGEMA_signal_5488), .Q (new_AGEMA_signal_5489) ) ;
    buf_clk new_AGEMA_reg_buffer_3537 ( .C (clk), .D (new_AGEMA_signal_5492), .Q (new_AGEMA_signal_5493) ) ;
    buf_clk new_AGEMA_reg_buffer_3541 ( .C (clk), .D (new_AGEMA_signal_5496), .Q (new_AGEMA_signal_5497) ) ;
    buf_clk new_AGEMA_reg_buffer_3545 ( .C (clk), .D (new_AGEMA_signal_5500), .Q (new_AGEMA_signal_5501) ) ;
    buf_clk new_AGEMA_reg_buffer_3549 ( .C (clk), .D (new_AGEMA_signal_5504), .Q (new_AGEMA_signal_5505) ) ;
    buf_clk new_AGEMA_reg_buffer_3553 ( .C (clk), .D (new_AGEMA_signal_5508), .Q (new_AGEMA_signal_5509) ) ;
    buf_clk new_AGEMA_reg_buffer_3557 ( .C (clk), .D (new_AGEMA_signal_5512), .Q (new_AGEMA_signal_5513) ) ;
    buf_clk new_AGEMA_reg_buffer_3561 ( .C (clk), .D (new_AGEMA_signal_5516), .Q (new_AGEMA_signal_5517) ) ;
    buf_clk new_AGEMA_reg_buffer_3565 ( .C (clk), .D (new_AGEMA_signal_5520), .Q (new_AGEMA_signal_5521) ) ;
    buf_clk new_AGEMA_reg_buffer_3569 ( .C (clk), .D (new_AGEMA_signal_5524), .Q (new_AGEMA_signal_5525) ) ;
    buf_clk new_AGEMA_reg_buffer_3573 ( .C (clk), .D (new_AGEMA_signal_5528), .Q (new_AGEMA_signal_5529) ) ;
    buf_clk new_AGEMA_reg_buffer_3577 ( .C (clk), .D (new_AGEMA_signal_5532), .Q (new_AGEMA_signal_5533) ) ;
    buf_clk new_AGEMA_reg_buffer_3581 ( .C (clk), .D (new_AGEMA_signal_5536), .Q (new_AGEMA_signal_5537) ) ;
    buf_clk new_AGEMA_reg_buffer_3585 ( .C (clk), .D (new_AGEMA_signal_5540), .Q (new_AGEMA_signal_5541) ) ;
    buf_clk new_AGEMA_reg_buffer_3589 ( .C (clk), .D (new_AGEMA_signal_5544), .Q (new_AGEMA_signal_5545) ) ;
    buf_clk new_AGEMA_reg_buffer_3593 ( .C (clk), .D (new_AGEMA_signal_5548), .Q (new_AGEMA_signal_5549) ) ;
    buf_clk new_AGEMA_reg_buffer_3597 ( .C (clk), .D (new_AGEMA_signal_5552), .Q (new_AGEMA_signal_5553) ) ;
    buf_clk new_AGEMA_reg_buffer_3601 ( .C (clk), .D (new_AGEMA_signal_5556), .Q (new_AGEMA_signal_5557) ) ;
    buf_clk new_AGEMA_reg_buffer_3605 ( .C (clk), .D (new_AGEMA_signal_5560), .Q (new_AGEMA_signal_5561) ) ;
    buf_clk new_AGEMA_reg_buffer_3609 ( .C (clk), .D (new_AGEMA_signal_5564), .Q (new_AGEMA_signal_5565) ) ;
    buf_clk new_AGEMA_reg_buffer_3613 ( .C (clk), .D (new_AGEMA_signal_5568), .Q (new_AGEMA_signal_5569) ) ;
    buf_clk new_AGEMA_reg_buffer_3617 ( .C (clk), .D (new_AGEMA_signal_5572), .Q (new_AGEMA_signal_5573) ) ;
    buf_clk new_AGEMA_reg_buffer_3621 ( .C (clk), .D (new_AGEMA_signal_5576), .Q (new_AGEMA_signal_5577) ) ;
    buf_clk new_AGEMA_reg_buffer_3625 ( .C (clk), .D (new_AGEMA_signal_5580), .Q (new_AGEMA_signal_5581) ) ;
    buf_clk new_AGEMA_reg_buffer_3629 ( .C (clk), .D (new_AGEMA_signal_5584), .Q (new_AGEMA_signal_5585) ) ;
    buf_clk new_AGEMA_reg_buffer_3633 ( .C (clk), .D (new_AGEMA_signal_5588), .Q (new_AGEMA_signal_5589) ) ;
    buf_clk new_AGEMA_reg_buffer_3637 ( .C (clk), .D (new_AGEMA_signal_5592), .Q (new_AGEMA_signal_5593) ) ;
    buf_clk new_AGEMA_reg_buffer_3641 ( .C (clk), .D (new_AGEMA_signal_5596), .Q (new_AGEMA_signal_5597) ) ;
    buf_clk new_AGEMA_reg_buffer_3645 ( .C (clk), .D (new_AGEMA_signal_5600), .Q (new_AGEMA_signal_5601) ) ;
    buf_clk new_AGEMA_reg_buffer_3649 ( .C (clk), .D (new_AGEMA_signal_5604), .Q (new_AGEMA_signal_5605) ) ;
    buf_clk new_AGEMA_reg_buffer_3653 ( .C (clk), .D (new_AGEMA_signal_5608), .Q (new_AGEMA_signal_5609) ) ;
    buf_clk new_AGEMA_reg_buffer_3657 ( .C (clk), .D (new_AGEMA_signal_5612), .Q (new_AGEMA_signal_5613) ) ;
    buf_clk new_AGEMA_reg_buffer_3661 ( .C (clk), .D (new_AGEMA_signal_5616), .Q (new_AGEMA_signal_5617) ) ;
    buf_clk new_AGEMA_reg_buffer_3665 ( .C (clk), .D (new_AGEMA_signal_5620), .Q (new_AGEMA_signal_5621) ) ;
    buf_clk new_AGEMA_reg_buffer_3669 ( .C (clk), .D (new_AGEMA_signal_5624), .Q (new_AGEMA_signal_5625) ) ;
    buf_clk new_AGEMA_reg_buffer_3673 ( .C (clk), .D (new_AGEMA_signal_5628), .Q (new_AGEMA_signal_5629) ) ;
    buf_clk new_AGEMA_reg_buffer_3677 ( .C (clk), .D (new_AGEMA_signal_5632), .Q (new_AGEMA_signal_5633) ) ;
    buf_clk new_AGEMA_reg_buffer_3681 ( .C (clk), .D (new_AGEMA_signal_5636), .Q (new_AGEMA_signal_5637) ) ;
    buf_clk new_AGEMA_reg_buffer_3685 ( .C (clk), .D (new_AGEMA_signal_5640), .Q (new_AGEMA_signal_5641) ) ;
    buf_clk new_AGEMA_reg_buffer_3689 ( .C (clk), .D (new_AGEMA_signal_5644), .Q (new_AGEMA_signal_5645) ) ;
    buf_clk new_AGEMA_reg_buffer_3693 ( .C (clk), .D (new_AGEMA_signal_5648), .Q (new_AGEMA_signal_5649) ) ;
    buf_clk new_AGEMA_reg_buffer_3697 ( .C (clk), .D (new_AGEMA_signal_5652), .Q (new_AGEMA_signal_5653) ) ;
    buf_clk new_AGEMA_reg_buffer_3701 ( .C (clk), .D (new_AGEMA_signal_5656), .Q (new_AGEMA_signal_5657) ) ;
    buf_clk new_AGEMA_reg_buffer_3705 ( .C (clk), .D (new_AGEMA_signal_5660), .Q (new_AGEMA_signal_5661) ) ;
    buf_clk new_AGEMA_reg_buffer_3709 ( .C (clk), .D (new_AGEMA_signal_5664), .Q (new_AGEMA_signal_5665) ) ;
    buf_clk new_AGEMA_reg_buffer_3713 ( .C (clk), .D (new_AGEMA_signal_5668), .Q (new_AGEMA_signal_5669) ) ;
    buf_clk new_AGEMA_reg_buffer_3717 ( .C (clk), .D (new_AGEMA_signal_5672), .Q (new_AGEMA_signal_5673) ) ;
    buf_clk new_AGEMA_reg_buffer_3721 ( .C (clk), .D (new_AGEMA_signal_5676), .Q (new_AGEMA_signal_5677) ) ;
    buf_clk new_AGEMA_reg_buffer_3725 ( .C (clk), .D (new_AGEMA_signal_5680), .Q (new_AGEMA_signal_5681) ) ;
    buf_clk new_AGEMA_reg_buffer_3729 ( .C (clk), .D (new_AGEMA_signal_5684), .Q (new_AGEMA_signal_5685) ) ;
    buf_clk new_AGEMA_reg_buffer_3733 ( .C (clk), .D (new_AGEMA_signal_5688), .Q (new_AGEMA_signal_5689) ) ;
    buf_clk new_AGEMA_reg_buffer_3737 ( .C (clk), .D (new_AGEMA_signal_5692), .Q (new_AGEMA_signal_5693) ) ;
    buf_clk new_AGEMA_reg_buffer_3741 ( .C (clk), .D (new_AGEMA_signal_5696), .Q (new_AGEMA_signal_5697) ) ;
    buf_clk new_AGEMA_reg_buffer_3745 ( .C (clk), .D (new_AGEMA_signal_5700), .Q (new_AGEMA_signal_5701) ) ;
    buf_clk new_AGEMA_reg_buffer_3749 ( .C (clk), .D (new_AGEMA_signal_5704), .Q (new_AGEMA_signal_5705) ) ;
    buf_clk new_AGEMA_reg_buffer_3753 ( .C (clk), .D (new_AGEMA_signal_5708), .Q (new_AGEMA_signal_5709) ) ;
    buf_clk new_AGEMA_reg_buffer_3757 ( .C (clk), .D (new_AGEMA_signal_5712), .Q (new_AGEMA_signal_5713) ) ;
    buf_clk new_AGEMA_reg_buffer_3761 ( .C (clk), .D (new_AGEMA_signal_5716), .Q (new_AGEMA_signal_5717) ) ;
    buf_clk new_AGEMA_reg_buffer_3765 ( .C (clk), .D (new_AGEMA_signal_5720), .Q (new_AGEMA_signal_5721) ) ;
    buf_clk new_AGEMA_reg_buffer_3769 ( .C (clk), .D (new_AGEMA_signal_5724), .Q (new_AGEMA_signal_5725) ) ;
    buf_clk new_AGEMA_reg_buffer_3773 ( .C (clk), .D (new_AGEMA_signal_5728), .Q (new_AGEMA_signal_5729) ) ;
    buf_clk new_AGEMA_reg_buffer_3777 ( .C (clk), .D (new_AGEMA_signal_5732), .Q (new_AGEMA_signal_5733) ) ;
    buf_clk new_AGEMA_reg_buffer_3781 ( .C (clk), .D (new_AGEMA_signal_5736), .Q (new_AGEMA_signal_5737) ) ;
    buf_clk new_AGEMA_reg_buffer_3785 ( .C (clk), .D (new_AGEMA_signal_5740), .Q (new_AGEMA_signal_5741) ) ;
    buf_clk new_AGEMA_reg_buffer_3789 ( .C (clk), .D (new_AGEMA_signal_5744), .Q (new_AGEMA_signal_5745) ) ;
    buf_clk new_AGEMA_reg_buffer_3793 ( .C (clk), .D (new_AGEMA_signal_5748), .Q (new_AGEMA_signal_5749) ) ;
    buf_clk new_AGEMA_reg_buffer_3797 ( .C (clk), .D (new_AGEMA_signal_5752), .Q (new_AGEMA_signal_5753) ) ;
    buf_clk new_AGEMA_reg_buffer_3801 ( .C (clk), .D (new_AGEMA_signal_5756), .Q (new_AGEMA_signal_5757) ) ;
    buf_clk new_AGEMA_reg_buffer_3805 ( .C (clk), .D (new_AGEMA_signal_5760), .Q (new_AGEMA_signal_5761) ) ;
    buf_clk new_AGEMA_reg_buffer_3809 ( .C (clk), .D (new_AGEMA_signal_5764), .Q (new_AGEMA_signal_5765) ) ;
    buf_clk new_AGEMA_reg_buffer_3813 ( .C (clk), .D (new_AGEMA_signal_5768), .Q (new_AGEMA_signal_5769) ) ;
    buf_clk new_AGEMA_reg_buffer_3817 ( .C (clk), .D (new_AGEMA_signal_5772), .Q (new_AGEMA_signal_5773) ) ;
    buf_clk new_AGEMA_reg_buffer_3821 ( .C (clk), .D (new_AGEMA_signal_5776), .Q (new_AGEMA_signal_5777) ) ;
    buf_clk new_AGEMA_reg_buffer_3825 ( .C (clk), .D (new_AGEMA_signal_5780), .Q (new_AGEMA_signal_5781) ) ;
    buf_clk new_AGEMA_reg_buffer_3829 ( .C (clk), .D (new_AGEMA_signal_5784), .Q (new_AGEMA_signal_5785) ) ;
    buf_clk new_AGEMA_reg_buffer_3833 ( .C (clk), .D (new_AGEMA_signal_5788), .Q (new_AGEMA_signal_5789) ) ;
    buf_clk new_AGEMA_reg_buffer_3837 ( .C (clk), .D (new_AGEMA_signal_5792), .Q (new_AGEMA_signal_5793) ) ;
    buf_clk new_AGEMA_reg_buffer_3841 ( .C (clk), .D (new_AGEMA_signal_5796), .Q (new_AGEMA_signal_5797) ) ;
    buf_clk new_AGEMA_reg_buffer_3845 ( .C (clk), .D (new_AGEMA_signal_5800), .Q (new_AGEMA_signal_5801) ) ;
    buf_clk new_AGEMA_reg_buffer_3849 ( .C (clk), .D (new_AGEMA_signal_5804), .Q (new_AGEMA_signal_5805) ) ;
    buf_clk new_AGEMA_reg_buffer_3853 ( .C (clk), .D (new_AGEMA_signal_5808), .Q (new_AGEMA_signal_5809) ) ;
    buf_clk new_AGEMA_reg_buffer_3857 ( .C (clk), .D (new_AGEMA_signal_5812), .Q (new_AGEMA_signal_5813) ) ;
    buf_clk new_AGEMA_reg_buffer_3861 ( .C (clk), .D (new_AGEMA_signal_5816), .Q (new_AGEMA_signal_5817) ) ;
    buf_clk new_AGEMA_reg_buffer_3865 ( .C (clk), .D (new_AGEMA_signal_5820), .Q (new_AGEMA_signal_5821) ) ;
    buf_clk new_AGEMA_reg_buffer_3869 ( .C (clk), .D (new_AGEMA_signal_5824), .Q (new_AGEMA_signal_5825) ) ;
    buf_clk new_AGEMA_reg_buffer_3873 ( .C (clk), .D (new_AGEMA_signal_5828), .Q (new_AGEMA_signal_5829) ) ;
    buf_clk new_AGEMA_reg_buffer_3877 ( .C (clk), .D (new_AGEMA_signal_5832), .Q (new_AGEMA_signal_5833) ) ;
    buf_clk new_AGEMA_reg_buffer_3881 ( .C (clk), .D (new_AGEMA_signal_5836), .Q (new_AGEMA_signal_5837) ) ;
    buf_clk new_AGEMA_reg_buffer_3885 ( .C (clk), .D (new_AGEMA_signal_5840), .Q (new_AGEMA_signal_5841) ) ;
    buf_clk new_AGEMA_reg_buffer_3889 ( .C (clk), .D (new_AGEMA_signal_5844), .Q (new_AGEMA_signal_5845) ) ;
    buf_clk new_AGEMA_reg_buffer_3893 ( .C (clk), .D (new_AGEMA_signal_5848), .Q (new_AGEMA_signal_5849) ) ;
    buf_clk new_AGEMA_reg_buffer_3897 ( .C (clk), .D (new_AGEMA_signal_5852), .Q (new_AGEMA_signal_5853) ) ;
    buf_clk new_AGEMA_reg_buffer_3901 ( .C (clk), .D (new_AGEMA_signal_5856), .Q (new_AGEMA_signal_5857) ) ;
    buf_clk new_AGEMA_reg_buffer_3905 ( .C (clk), .D (new_AGEMA_signal_5860), .Q (new_AGEMA_signal_5861) ) ;
    buf_clk new_AGEMA_reg_buffer_3909 ( .C (clk), .D (new_AGEMA_signal_5864), .Q (new_AGEMA_signal_5865) ) ;
    buf_clk new_AGEMA_reg_buffer_3913 ( .C (clk), .D (new_AGEMA_signal_5868), .Q (new_AGEMA_signal_5869) ) ;
    buf_clk new_AGEMA_reg_buffer_3917 ( .C (clk), .D (new_AGEMA_signal_5872), .Q (new_AGEMA_signal_5873) ) ;
    buf_clk new_AGEMA_reg_buffer_3921 ( .C (clk), .D (new_AGEMA_signal_5876), .Q (new_AGEMA_signal_5877) ) ;
    buf_clk new_AGEMA_reg_buffer_3925 ( .C (clk), .D (new_AGEMA_signal_5880), .Q (new_AGEMA_signal_5881) ) ;
    buf_clk new_AGEMA_reg_buffer_3929 ( .C (clk), .D (new_AGEMA_signal_5884), .Q (new_AGEMA_signal_5885) ) ;
    buf_clk new_AGEMA_reg_buffer_3933 ( .C (clk), .D (new_AGEMA_signal_5888), .Q (new_AGEMA_signal_5889) ) ;
    buf_clk new_AGEMA_reg_buffer_3937 ( .C (clk), .D (new_AGEMA_signal_5892), .Q (new_AGEMA_signal_5893) ) ;
    buf_clk new_AGEMA_reg_buffer_3941 ( .C (clk), .D (new_AGEMA_signal_5896), .Q (new_AGEMA_signal_5897) ) ;
    buf_clk new_AGEMA_reg_buffer_3945 ( .C (clk), .D (new_AGEMA_signal_5900), .Q (new_AGEMA_signal_5901) ) ;
    buf_clk new_AGEMA_reg_buffer_3949 ( .C (clk), .D (new_AGEMA_signal_5904), .Q (new_AGEMA_signal_5905) ) ;
    buf_clk new_AGEMA_reg_buffer_3953 ( .C (clk), .D (new_AGEMA_signal_5908), .Q (new_AGEMA_signal_5909) ) ;
    buf_clk new_AGEMA_reg_buffer_3957 ( .C (clk), .D (new_AGEMA_signal_5912), .Q (new_AGEMA_signal_5913) ) ;
    buf_clk new_AGEMA_reg_buffer_3961 ( .C (clk), .D (new_AGEMA_signal_5916), .Q (new_AGEMA_signal_5917) ) ;
    buf_clk new_AGEMA_reg_buffer_3965 ( .C (clk), .D (new_AGEMA_signal_5920), .Q (new_AGEMA_signal_5921) ) ;
    buf_clk new_AGEMA_reg_buffer_3969 ( .C (clk), .D (new_AGEMA_signal_5924), .Q (new_AGEMA_signal_5925) ) ;
    buf_clk new_AGEMA_reg_buffer_3973 ( .C (clk), .D (new_AGEMA_signal_5928), .Q (new_AGEMA_signal_5929) ) ;
    buf_clk new_AGEMA_reg_buffer_3977 ( .C (clk), .D (new_AGEMA_signal_5932), .Q (new_AGEMA_signal_5933) ) ;
    buf_clk new_AGEMA_reg_buffer_3981 ( .C (clk), .D (new_AGEMA_signal_5936), .Q (new_AGEMA_signal_5937) ) ;
    buf_clk new_AGEMA_reg_buffer_3985 ( .C (clk), .D (new_AGEMA_signal_5940), .Q (new_AGEMA_signal_5941) ) ;
    buf_clk new_AGEMA_reg_buffer_3989 ( .C (clk), .D (new_AGEMA_signal_5944), .Q (new_AGEMA_signal_5945) ) ;
    buf_clk new_AGEMA_reg_buffer_3993 ( .C (clk), .D (new_AGEMA_signal_5948), .Q (new_AGEMA_signal_5949) ) ;
    buf_clk new_AGEMA_reg_buffer_3997 ( .C (clk), .D (new_AGEMA_signal_5952), .Q (new_AGEMA_signal_5953) ) ;
    buf_clk new_AGEMA_reg_buffer_4001 ( .C (clk), .D (new_AGEMA_signal_5956), .Q (new_AGEMA_signal_5957) ) ;
    buf_clk new_AGEMA_reg_buffer_4005 ( .C (clk), .D (new_AGEMA_signal_5960), .Q (new_AGEMA_signal_5961) ) ;
    buf_clk new_AGEMA_reg_buffer_4009 ( .C (clk), .D (new_AGEMA_signal_5964), .Q (new_AGEMA_signal_5965) ) ;
    buf_clk new_AGEMA_reg_buffer_4013 ( .C (clk), .D (new_AGEMA_signal_5968), .Q (new_AGEMA_signal_5969) ) ;
    buf_clk new_AGEMA_reg_buffer_4017 ( .C (clk), .D (new_AGEMA_signal_5972), .Q (new_AGEMA_signal_5973) ) ;
    buf_clk new_AGEMA_reg_buffer_4021 ( .C (clk), .D (new_AGEMA_signal_5976), .Q (new_AGEMA_signal_5977) ) ;
    buf_clk new_AGEMA_reg_buffer_4025 ( .C (clk), .D (new_AGEMA_signal_5980), .Q (new_AGEMA_signal_5981) ) ;
    buf_clk new_AGEMA_reg_buffer_4029 ( .C (clk), .D (new_AGEMA_signal_5984), .Q (new_AGEMA_signal_5985) ) ;
    buf_clk new_AGEMA_reg_buffer_4033 ( .C (clk), .D (new_AGEMA_signal_5988), .Q (new_AGEMA_signal_5989) ) ;
    buf_clk new_AGEMA_reg_buffer_4037 ( .C (clk), .D (new_AGEMA_signal_5992), .Q (new_AGEMA_signal_5993) ) ;
    buf_clk new_AGEMA_reg_buffer_4041 ( .C (clk), .D (new_AGEMA_signal_5996), .Q (new_AGEMA_signal_5997) ) ;
    buf_clk new_AGEMA_reg_buffer_4045 ( .C (clk), .D (new_AGEMA_signal_6000), .Q (new_AGEMA_signal_6001) ) ;
    buf_clk new_AGEMA_reg_buffer_4049 ( .C (clk), .D (new_AGEMA_signal_6004), .Q (new_AGEMA_signal_6005) ) ;
    buf_clk new_AGEMA_reg_buffer_4053 ( .C (clk), .D (new_AGEMA_signal_6008), .Q (new_AGEMA_signal_6009) ) ;
    buf_clk new_AGEMA_reg_buffer_4057 ( .C (clk), .D (new_AGEMA_signal_6012), .Q (new_AGEMA_signal_6013) ) ;
    buf_clk new_AGEMA_reg_buffer_4061 ( .C (clk), .D (new_AGEMA_signal_6016), .Q (new_AGEMA_signal_6017) ) ;
    buf_clk new_AGEMA_reg_buffer_4065 ( .C (clk), .D (new_AGEMA_signal_6020), .Q (new_AGEMA_signal_6021) ) ;
    buf_clk new_AGEMA_reg_buffer_4069 ( .C (clk), .D (new_AGEMA_signal_6024), .Q (new_AGEMA_signal_6025) ) ;
    buf_clk new_AGEMA_reg_buffer_4073 ( .C (clk), .D (new_AGEMA_signal_6028), .Q (new_AGEMA_signal_6029) ) ;
    buf_clk new_AGEMA_reg_buffer_4077 ( .C (clk), .D (new_AGEMA_signal_6032), .Q (new_AGEMA_signal_6033) ) ;
    buf_clk new_AGEMA_reg_buffer_4081 ( .C (clk), .D (new_AGEMA_signal_6036), .Q (new_AGEMA_signal_6037) ) ;
    buf_clk new_AGEMA_reg_buffer_4085 ( .C (clk), .D (new_AGEMA_signal_6040), .Q (new_AGEMA_signal_6041) ) ;
    buf_clk new_AGEMA_reg_buffer_4089 ( .C (clk), .D (new_AGEMA_signal_6044), .Q (new_AGEMA_signal_6045) ) ;
    buf_clk new_AGEMA_reg_buffer_4093 ( .C (clk), .D (new_AGEMA_signal_6048), .Q (new_AGEMA_signal_6049) ) ;
    buf_clk new_AGEMA_reg_buffer_4097 ( .C (clk), .D (new_AGEMA_signal_6052), .Q (new_AGEMA_signal_6053) ) ;
    buf_clk new_AGEMA_reg_buffer_4101 ( .C (clk), .D (new_AGEMA_signal_6056), .Q (new_AGEMA_signal_6057) ) ;
    buf_clk new_AGEMA_reg_buffer_4105 ( .C (clk), .D (new_AGEMA_signal_6060), .Q (new_AGEMA_signal_6061) ) ;
    buf_clk new_AGEMA_reg_buffer_4109 ( .C (clk), .D (new_AGEMA_signal_6064), .Q (new_AGEMA_signal_6065) ) ;
    buf_clk new_AGEMA_reg_buffer_4113 ( .C (clk), .D (new_AGEMA_signal_6068), .Q (new_AGEMA_signal_6069) ) ;
    buf_clk new_AGEMA_reg_buffer_4117 ( .C (clk), .D (new_AGEMA_signal_6072), .Q (new_AGEMA_signal_6073) ) ;
    buf_clk new_AGEMA_reg_buffer_4121 ( .C (clk), .D (new_AGEMA_signal_6076), .Q (new_AGEMA_signal_6077) ) ;
    buf_clk new_AGEMA_reg_buffer_4125 ( .C (clk), .D (new_AGEMA_signal_6080), .Q (new_AGEMA_signal_6081) ) ;
    buf_clk new_AGEMA_reg_buffer_4129 ( .C (clk), .D (new_AGEMA_signal_6084), .Q (new_AGEMA_signal_6085) ) ;
    buf_clk new_AGEMA_reg_buffer_4133 ( .C (clk), .D (new_AGEMA_signal_6088), .Q (new_AGEMA_signal_6089) ) ;
    buf_clk new_AGEMA_reg_buffer_4137 ( .C (clk), .D (new_AGEMA_signal_6092), .Q (new_AGEMA_signal_6093) ) ;
    buf_clk new_AGEMA_reg_buffer_4141 ( .C (clk), .D (new_AGEMA_signal_6096), .Q (new_AGEMA_signal_6097) ) ;
    buf_clk new_AGEMA_reg_buffer_4145 ( .C (clk), .D (new_AGEMA_signal_6100), .Q (new_AGEMA_signal_6101) ) ;
    buf_clk new_AGEMA_reg_buffer_4149 ( .C (clk), .D (new_AGEMA_signal_6104), .Q (new_AGEMA_signal_6105) ) ;
    buf_clk new_AGEMA_reg_buffer_4153 ( .C (clk), .D (new_AGEMA_signal_6108), .Q (new_AGEMA_signal_6109) ) ;
    buf_clk new_AGEMA_reg_buffer_4157 ( .C (clk), .D (new_AGEMA_signal_6112), .Q (new_AGEMA_signal_6113) ) ;
    buf_clk new_AGEMA_reg_buffer_4161 ( .C (clk), .D (new_AGEMA_signal_6116), .Q (new_AGEMA_signal_6117) ) ;
    buf_clk new_AGEMA_reg_buffer_4165 ( .C (clk), .D (new_AGEMA_signal_6120), .Q (new_AGEMA_signal_6121) ) ;
    buf_clk new_AGEMA_reg_buffer_4169 ( .C (clk), .D (new_AGEMA_signal_6124), .Q (new_AGEMA_signal_6125) ) ;
    buf_clk new_AGEMA_reg_buffer_4173 ( .C (clk), .D (new_AGEMA_signal_6128), .Q (new_AGEMA_signal_6129) ) ;
    buf_clk new_AGEMA_reg_buffer_4177 ( .C (clk), .D (new_AGEMA_signal_6132), .Q (new_AGEMA_signal_6133) ) ;
    buf_clk new_AGEMA_reg_buffer_4181 ( .C (clk), .D (new_AGEMA_signal_6136), .Q (new_AGEMA_signal_6137) ) ;
    buf_clk new_AGEMA_reg_buffer_4185 ( .C (clk), .D (new_AGEMA_signal_6140), .Q (new_AGEMA_signal_6141) ) ;
    buf_clk new_AGEMA_reg_buffer_4189 ( .C (clk), .D (new_AGEMA_signal_6144), .Q (new_AGEMA_signal_6145) ) ;
    buf_clk new_AGEMA_reg_buffer_4193 ( .C (clk), .D (new_AGEMA_signal_6148), .Q (new_AGEMA_signal_6149) ) ;
    buf_clk new_AGEMA_reg_buffer_4197 ( .C (clk), .D (new_AGEMA_signal_6152), .Q (new_AGEMA_signal_6153) ) ;
    buf_clk new_AGEMA_reg_buffer_4201 ( .C (clk), .D (new_AGEMA_signal_6156), .Q (new_AGEMA_signal_6157) ) ;
    buf_clk new_AGEMA_reg_buffer_4205 ( .C (clk), .D (new_AGEMA_signal_6160), .Q (new_AGEMA_signal_6161) ) ;
    buf_clk new_AGEMA_reg_buffer_4209 ( .C (clk), .D (new_AGEMA_signal_6164), .Q (new_AGEMA_signal_6165) ) ;
    buf_clk new_AGEMA_reg_buffer_4213 ( .C (clk), .D (new_AGEMA_signal_6168), .Q (new_AGEMA_signal_6169) ) ;
    buf_clk new_AGEMA_reg_buffer_4217 ( .C (clk), .D (new_AGEMA_signal_6172), .Q (new_AGEMA_signal_6173) ) ;
    buf_clk new_AGEMA_reg_buffer_4221 ( .C (clk), .D (new_AGEMA_signal_6176), .Q (new_AGEMA_signal_6177) ) ;
    buf_clk new_AGEMA_reg_buffer_4225 ( .C (clk), .D (new_AGEMA_signal_6180), .Q (new_AGEMA_signal_6181) ) ;
    buf_clk new_AGEMA_reg_buffer_4229 ( .C (clk), .D (new_AGEMA_signal_6184), .Q (new_AGEMA_signal_6185) ) ;
    buf_clk new_AGEMA_reg_buffer_4233 ( .C (clk), .D (new_AGEMA_signal_6188), .Q (new_AGEMA_signal_6189) ) ;
    buf_clk new_AGEMA_reg_buffer_4237 ( .C (clk), .D (new_AGEMA_signal_6192), .Q (new_AGEMA_signal_6193) ) ;
    buf_clk new_AGEMA_reg_buffer_4241 ( .C (clk), .D (new_AGEMA_signal_6196), .Q (new_AGEMA_signal_6197) ) ;
    buf_clk new_AGEMA_reg_buffer_4245 ( .C (clk), .D (new_AGEMA_signal_6200), .Q (new_AGEMA_signal_6201) ) ;
    buf_clk new_AGEMA_reg_buffer_4249 ( .C (clk), .D (new_AGEMA_signal_6204), .Q (new_AGEMA_signal_6205) ) ;
    buf_clk new_AGEMA_reg_buffer_4253 ( .C (clk), .D (new_AGEMA_signal_6208), .Q (new_AGEMA_signal_6209) ) ;
    buf_clk new_AGEMA_reg_buffer_4257 ( .C (clk), .D (new_AGEMA_signal_6212), .Q (new_AGEMA_signal_6213) ) ;
    buf_clk new_AGEMA_reg_buffer_4261 ( .C (clk), .D (new_AGEMA_signal_6216), .Q (new_AGEMA_signal_6217) ) ;
    buf_clk new_AGEMA_reg_buffer_4265 ( .C (clk), .D (new_AGEMA_signal_6220), .Q (new_AGEMA_signal_6221) ) ;
    buf_clk new_AGEMA_reg_buffer_4269 ( .C (clk), .D (new_AGEMA_signal_6224), .Q (new_AGEMA_signal_6225) ) ;
    buf_clk new_AGEMA_reg_buffer_4273 ( .C (clk), .D (new_AGEMA_signal_6228), .Q (new_AGEMA_signal_6229) ) ;
    buf_clk new_AGEMA_reg_buffer_4277 ( .C (clk), .D (new_AGEMA_signal_6232), .Q (new_AGEMA_signal_6233) ) ;
    buf_clk new_AGEMA_reg_buffer_4281 ( .C (clk), .D (new_AGEMA_signal_6236), .Q (new_AGEMA_signal_6237) ) ;
    buf_clk new_AGEMA_reg_buffer_4285 ( .C (clk), .D (new_AGEMA_signal_6240), .Q (new_AGEMA_signal_6241) ) ;
    buf_clk new_AGEMA_reg_buffer_4289 ( .C (clk), .D (new_AGEMA_signal_6244), .Q (new_AGEMA_signal_6245) ) ;
    buf_clk new_AGEMA_reg_buffer_4293 ( .C (clk), .D (new_AGEMA_signal_6248), .Q (new_AGEMA_signal_6249) ) ;
    buf_clk new_AGEMA_reg_buffer_4297 ( .C (clk), .D (new_AGEMA_signal_6252), .Q (new_AGEMA_signal_6253) ) ;
    buf_clk new_AGEMA_reg_buffer_4301 ( .C (clk), .D (new_AGEMA_signal_6256), .Q (new_AGEMA_signal_6257) ) ;
    buf_clk new_AGEMA_reg_buffer_4305 ( .C (clk), .D (new_AGEMA_signal_6260), .Q (new_AGEMA_signal_6261) ) ;
    buf_clk new_AGEMA_reg_buffer_4309 ( .C (clk), .D (new_AGEMA_signal_6264), .Q (new_AGEMA_signal_6265) ) ;
    buf_clk new_AGEMA_reg_buffer_4313 ( .C (clk), .D (new_AGEMA_signal_6268), .Q (new_AGEMA_signal_6269) ) ;
    buf_clk new_AGEMA_reg_buffer_4317 ( .C (clk), .D (new_AGEMA_signal_6272), .Q (new_AGEMA_signal_6273) ) ;
    buf_clk new_AGEMA_reg_buffer_4321 ( .C (clk), .D (new_AGEMA_signal_6276), .Q (new_AGEMA_signal_6277) ) ;
    buf_clk new_AGEMA_reg_buffer_4325 ( .C (clk), .D (new_AGEMA_signal_6280), .Q (new_AGEMA_signal_6281) ) ;
    buf_clk new_AGEMA_reg_buffer_4329 ( .C (clk), .D (new_AGEMA_signal_6284), .Q (new_AGEMA_signal_6285) ) ;
    buf_clk new_AGEMA_reg_buffer_4333 ( .C (clk), .D (new_AGEMA_signal_6288), .Q (new_AGEMA_signal_6289) ) ;
    buf_clk new_AGEMA_reg_buffer_4337 ( .C (clk), .D (new_AGEMA_signal_6292), .Q (new_AGEMA_signal_6293) ) ;
    buf_clk new_AGEMA_reg_buffer_4341 ( .C (clk), .D (new_AGEMA_signal_6296), .Q (new_AGEMA_signal_6297) ) ;

    /* register cells */
    DFF_X1 ctrl_seq6_SFF_0_Q_reg_FF_FF ( .CK (clk), .D (new_AGEMA_signal_4309), .Q (ctrl_seq6In_1_), .QN () ) ;
    DFF_X1 ctrl_seq6_SFF_1_Q_reg_FF_FF ( .CK (clk), .D (new_AGEMA_signal_4313), .Q (ctrl_seq6In_2_), .QN () ) ;
    DFF_X1 ctrl_seq6_SFF_2_Q_reg_FF_FF ( .CK (clk), .D (new_AGEMA_signal_4317), .Q (ctrl_seq6In_3_), .QN () ) ;
    DFF_X1 ctrl_seq6_SFF_3_Q_reg_FF_FF ( .CK (clk), .D (new_AGEMA_signal_4321), .Q (ctrl_seq6In_4_), .QN () ) ;
    DFF_X1 ctrl_seq6_SFF_4_Q_reg_FF_FF ( .CK (clk), .D (new_AGEMA_signal_4325), .Q (ctrl_seq6Out_4_), .QN () ) ;
    DFF_X1 ctrl_seq4_SFF_0_Q_reg_FF_FF ( .CK (clk), .D (new_AGEMA_signal_4329), .Q (ctrl_seq4In_1_), .QN () ) ;
    DFF_X1 ctrl_seq4_SFF_1_Q_reg_FF_FF ( .CK (clk), .D (new_AGEMA_signal_4333), .Q (ctrl_seq4Out_1_), .QN () ) ;
    DFF_X1 ctrl_CSselMC_reg_FF_FF ( .CK (clk), .D (new_AGEMA_signal_4337), .Q (ctrl_n6), .QN () ) ;
    DFF_X1 ctrl_CSenRC_reg_FF_FF ( .CK (clk), .D (new_AGEMA_signal_4341), .Q (enRCon), .QN () ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S00reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4349, new_AGEMA_signal_4345}), .Q ({ciphertext_s1[120], ciphertext_s0[120]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S00reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4357, new_AGEMA_signal_4353}), .Q ({ciphertext_s1[121], ciphertext_s0[121]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S00reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4365, new_AGEMA_signal_4361}), .Q ({ciphertext_s1[122], ciphertext_s0[122]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S00reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4373, new_AGEMA_signal_4369}), .Q ({ciphertext_s1[123], ciphertext_s0[123]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S00reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4381, new_AGEMA_signal_4377}), .Q ({ciphertext_s1[124], ciphertext_s0[124]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S00reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4389, new_AGEMA_signal_4385}), .Q ({ciphertext_s1[125], ciphertext_s0[125]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S00reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4397, new_AGEMA_signal_4393}), .Q ({ciphertext_s1[126], ciphertext_s0[126]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S00reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4405, new_AGEMA_signal_4401}), .Q ({ciphertext_s1[127], ciphertext_s0[127]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S01reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4413, new_AGEMA_signal_4409}), .Q ({ciphertext_s1[112], ciphertext_s0[112]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S01reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4421, new_AGEMA_signal_4417}), .Q ({ciphertext_s1[113], ciphertext_s0[113]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S01reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4429, new_AGEMA_signal_4425}), .Q ({ciphertext_s1[114], ciphertext_s0[114]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S01reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4437, new_AGEMA_signal_4433}), .Q ({ciphertext_s1[115], ciphertext_s0[115]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S01reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4445, new_AGEMA_signal_4441}), .Q ({ciphertext_s1[116], ciphertext_s0[116]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S01reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4453, new_AGEMA_signal_4449}), .Q ({ciphertext_s1[117], ciphertext_s0[117]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S01reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4461, new_AGEMA_signal_4457}), .Q ({ciphertext_s1[118], ciphertext_s0[118]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S01reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4469, new_AGEMA_signal_4465}), .Q ({ciphertext_s1[119], ciphertext_s0[119]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S02reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4477, new_AGEMA_signal_4473}), .Q ({ciphertext_s1[104], ciphertext_s0[104]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S02reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4485, new_AGEMA_signal_4481}), .Q ({ciphertext_s1[105], ciphertext_s0[105]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S02reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4493, new_AGEMA_signal_4489}), .Q ({ciphertext_s1[106], ciphertext_s0[106]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S02reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4501, new_AGEMA_signal_4497}), .Q ({ciphertext_s1[107], ciphertext_s0[107]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S02reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4509, new_AGEMA_signal_4505}), .Q ({ciphertext_s1[108], ciphertext_s0[108]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S02reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4517, new_AGEMA_signal_4513}), .Q ({ciphertext_s1[109], ciphertext_s0[109]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S02reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4525, new_AGEMA_signal_4521}), .Q ({ciphertext_s1[110], ciphertext_s0[110]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S02reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4533, new_AGEMA_signal_4529}), .Q ({ciphertext_s1[111], ciphertext_s0[111]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S03reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4541, new_AGEMA_signal_4537}), .Q ({ciphertext_s1[96], ciphertext_s0[96]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S03reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4549, new_AGEMA_signal_4545}), .Q ({ciphertext_s1[97], ciphertext_s0[97]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S03reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4557, new_AGEMA_signal_4553}), .Q ({ciphertext_s1[98], ciphertext_s0[98]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S03reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4565, new_AGEMA_signal_4561}), .Q ({ciphertext_s1[99], ciphertext_s0[99]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S03reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4573, new_AGEMA_signal_4569}), .Q ({ciphertext_s1[100], ciphertext_s0[100]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S03reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4581, new_AGEMA_signal_4577}), .Q ({ciphertext_s1[101], ciphertext_s0[101]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S03reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4589, new_AGEMA_signal_4585}), .Q ({ciphertext_s1[102], ciphertext_s0[102]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S03reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4597, new_AGEMA_signal_4593}), .Q ({ciphertext_s1[103], ciphertext_s0[103]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S10reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4605, new_AGEMA_signal_4601}), .Q ({ciphertext_s1[88], ciphertext_s0[88]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S10reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4613, new_AGEMA_signal_4609}), .Q ({ciphertext_s1[89], ciphertext_s0[89]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S10reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4621, new_AGEMA_signal_4617}), .Q ({ciphertext_s1[90], ciphertext_s0[90]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S10reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4629, new_AGEMA_signal_4625}), .Q ({ciphertext_s1[91], ciphertext_s0[91]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S10reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4637, new_AGEMA_signal_4633}), .Q ({ciphertext_s1[92], ciphertext_s0[92]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S10reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4645, new_AGEMA_signal_4641}), .Q ({ciphertext_s1[93], ciphertext_s0[93]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S10reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4653, new_AGEMA_signal_4649}), .Q ({ciphertext_s1[94], ciphertext_s0[94]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S10reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4661, new_AGEMA_signal_4657}), .Q ({ciphertext_s1[95], ciphertext_s0[95]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S11reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4669, new_AGEMA_signal_4665}), .Q ({ciphertext_s1[80], ciphertext_s0[80]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S11reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4677, new_AGEMA_signal_4673}), .Q ({ciphertext_s1[81], ciphertext_s0[81]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S11reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4685, new_AGEMA_signal_4681}), .Q ({ciphertext_s1[82], ciphertext_s0[82]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S11reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4693, new_AGEMA_signal_4689}), .Q ({ciphertext_s1[83], ciphertext_s0[83]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S11reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4701, new_AGEMA_signal_4697}), .Q ({ciphertext_s1[84], ciphertext_s0[84]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S11reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4709, new_AGEMA_signal_4705}), .Q ({ciphertext_s1[85], ciphertext_s0[85]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S11reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4717, new_AGEMA_signal_4713}), .Q ({ciphertext_s1[86], ciphertext_s0[86]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S11reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4725, new_AGEMA_signal_4721}), .Q ({ciphertext_s1[87], ciphertext_s0[87]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S12reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4733, new_AGEMA_signal_4729}), .Q ({ciphertext_s1[72], ciphertext_s0[72]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S12reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4741, new_AGEMA_signal_4737}), .Q ({ciphertext_s1[73], ciphertext_s0[73]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S12reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4749, new_AGEMA_signal_4745}), .Q ({ciphertext_s1[74], ciphertext_s0[74]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S12reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4757, new_AGEMA_signal_4753}), .Q ({ciphertext_s1[75], ciphertext_s0[75]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S12reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4765, new_AGEMA_signal_4761}), .Q ({ciphertext_s1[76], ciphertext_s0[76]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S12reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4773, new_AGEMA_signal_4769}), .Q ({ciphertext_s1[77], ciphertext_s0[77]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S12reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4781, new_AGEMA_signal_4777}), .Q ({ciphertext_s1[78], ciphertext_s0[78]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S12reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4789, new_AGEMA_signal_4785}), .Q ({ciphertext_s1[79], ciphertext_s0[79]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S13reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4797, new_AGEMA_signal_4793}), .Q ({ciphertext_s1[64], ciphertext_s0[64]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S13reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4805, new_AGEMA_signal_4801}), .Q ({ciphertext_s1[65], ciphertext_s0[65]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S13reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4813, new_AGEMA_signal_4809}), .Q ({ciphertext_s1[66], ciphertext_s0[66]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S13reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4821, new_AGEMA_signal_4817}), .Q ({ciphertext_s1[67], ciphertext_s0[67]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S13reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4829, new_AGEMA_signal_4825}), .Q ({ciphertext_s1[68], ciphertext_s0[68]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S13reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4837, new_AGEMA_signal_4833}), .Q ({ciphertext_s1[69], ciphertext_s0[69]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S13reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4845, new_AGEMA_signal_4841}), .Q ({ciphertext_s1[70], ciphertext_s0[70]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S13reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4853, new_AGEMA_signal_4849}), .Q ({ciphertext_s1[71], ciphertext_s0[71]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S20reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4861, new_AGEMA_signal_4857}), .Q ({ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S20reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4869, new_AGEMA_signal_4865}), .Q ({ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S20reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4877, new_AGEMA_signal_4873}), .Q ({ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S20reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4885, new_AGEMA_signal_4881}), .Q ({ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S20reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4893, new_AGEMA_signal_4889}), .Q ({ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S20reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4901, new_AGEMA_signal_4897}), .Q ({ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S20reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4909, new_AGEMA_signal_4905}), .Q ({ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S20reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4917, new_AGEMA_signal_4913}), .Q ({ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S21reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4925, new_AGEMA_signal_4921}), .Q ({ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S21reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4933, new_AGEMA_signal_4929}), .Q ({ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S21reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4941, new_AGEMA_signal_4937}), .Q ({ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S21reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4949, new_AGEMA_signal_4945}), .Q ({ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S21reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4957, new_AGEMA_signal_4953}), .Q ({ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S21reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4965, new_AGEMA_signal_4961}), .Q ({ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S21reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4973, new_AGEMA_signal_4969}), .Q ({ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S21reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4981, new_AGEMA_signal_4977}), .Q ({ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S22reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4989, new_AGEMA_signal_4985}), .Q ({ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S22reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4997, new_AGEMA_signal_4993}), .Q ({ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S22reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5005, new_AGEMA_signal_5001}), .Q ({ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S22reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5013, new_AGEMA_signal_5009}), .Q ({ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S22reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5021, new_AGEMA_signal_5017}), .Q ({ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S22reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5029, new_AGEMA_signal_5025}), .Q ({ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S22reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5037, new_AGEMA_signal_5033}), .Q ({ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S22reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5045, new_AGEMA_signal_5041}), .Q ({ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S23reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5053, new_AGEMA_signal_5049}), .Q ({ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S23reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5061, new_AGEMA_signal_5057}), .Q ({ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S23reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5069, new_AGEMA_signal_5065}), .Q ({ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S23reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5077, new_AGEMA_signal_5073}), .Q ({ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S23reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5085, new_AGEMA_signal_5081}), .Q ({ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S23reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5093, new_AGEMA_signal_5089}), .Q ({ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S23reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5101, new_AGEMA_signal_5097}), .Q ({ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S23reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5109, new_AGEMA_signal_5105}), .Q ({ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S30reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5117, new_AGEMA_signal_5113}), .Q ({ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S30reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5125, new_AGEMA_signal_5121}), .Q ({ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S30reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5133, new_AGEMA_signal_5129}), .Q ({ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S30reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5141, new_AGEMA_signal_5137}), .Q ({ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S30reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5149, new_AGEMA_signal_5145}), .Q ({ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S30reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5157, new_AGEMA_signal_5153}), .Q ({ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S30reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5165, new_AGEMA_signal_5161}), .Q ({ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S30reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5173, new_AGEMA_signal_5169}), .Q ({ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S31reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5181, new_AGEMA_signal_5177}), .Q ({ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S31reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5189, new_AGEMA_signal_5185}), .Q ({ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S31reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5197, new_AGEMA_signal_5193}), .Q ({ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S31reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5205, new_AGEMA_signal_5201}), .Q ({ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S31reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5213, new_AGEMA_signal_5209}), .Q ({ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S31reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5221, new_AGEMA_signal_5217}), .Q ({ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S31reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5229, new_AGEMA_signal_5225}), .Q ({ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S31reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5237, new_AGEMA_signal_5233}), .Q ({ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S32reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5245, new_AGEMA_signal_5241}), .Q ({ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S32reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5253, new_AGEMA_signal_5249}), .Q ({ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S32reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5261, new_AGEMA_signal_5257}), .Q ({ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S32reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5269, new_AGEMA_signal_5265}), .Q ({ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S32reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5277, new_AGEMA_signal_5273}), .Q ({ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S32reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5285, new_AGEMA_signal_5281}), .Q ({ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S32reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5293, new_AGEMA_signal_5289}), .Q ({ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S32reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5301, new_AGEMA_signal_5297}), .Q ({ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S33reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3497, stateArray_S33reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S33reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3520, stateArray_S33reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S33reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3521, stateArray_S33reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S33reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3522, stateArray_S33reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S33reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3523, stateArray_S33reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S33reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3524, stateArray_S33reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S33reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3525, stateArray_S33reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) stateArray_S33reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3526, stateArray_S33reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S00reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5309, new_AGEMA_signal_5305}), .Q ({new_AGEMA_signal_1983, keyStateIn[0]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S00reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5317, new_AGEMA_signal_5313}), .Q ({new_AGEMA_signal_1986, keyStateIn[1]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S00reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5325, new_AGEMA_signal_5321}), .Q ({new_AGEMA_signal_1989, keyStateIn[2]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S00reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5333, new_AGEMA_signal_5329}), .Q ({new_AGEMA_signal_1992, keyStateIn[3]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S00reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5341, new_AGEMA_signal_5337}), .Q ({new_AGEMA_signal_1995, keyStateIn[4]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S00reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5349, new_AGEMA_signal_5345}), .Q ({new_AGEMA_signal_1998, keyStateIn[5]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S00reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5357, new_AGEMA_signal_5353}), .Q ({new_AGEMA_signal_2001, keyStateIn[6]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S00reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5365, new_AGEMA_signal_5361}), .Q ({new_AGEMA_signal_2004, keyStateIn[7]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S01reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5373, new_AGEMA_signal_5369}), .Q ({new_AGEMA_signal_2020, KeyArray_outS01ser_0_}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S01reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5381, new_AGEMA_signal_5377}), .Q ({new_AGEMA_signal_2018, KeyArray_outS01ser_1_}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S01reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5389, new_AGEMA_signal_5385}), .Q ({new_AGEMA_signal_2016, KeyArray_outS01ser_2_}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S01reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5397, new_AGEMA_signal_5393}), .Q ({new_AGEMA_signal_2014, KeyArray_outS01ser_3_}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S01reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5405, new_AGEMA_signal_5401}), .Q ({new_AGEMA_signal_2012, KeyArray_outS01ser_4_}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S01reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5413, new_AGEMA_signal_5409}), .Q ({new_AGEMA_signal_2010, KeyArray_outS01ser_5_}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S01reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5421, new_AGEMA_signal_5417}), .Q ({new_AGEMA_signal_2008, KeyArray_outS01ser_6_}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S01reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5429, new_AGEMA_signal_5425}), .Q ({new_AGEMA_signal_2006, KeyArray_outS01ser_7_}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S02reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5437, new_AGEMA_signal_5433}), .Q ({new_AGEMA_signal_2443, KeyArray_outS02ser[0]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S02reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5445, new_AGEMA_signal_5441}), .Q ({new_AGEMA_signal_2446, KeyArray_outS02ser[1]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S02reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5453, new_AGEMA_signal_5449}), .Q ({new_AGEMA_signal_2449, KeyArray_outS02ser[2]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S02reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5461, new_AGEMA_signal_5457}), .Q ({new_AGEMA_signal_2452, KeyArray_outS02ser[3]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S02reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5469, new_AGEMA_signal_5465}), .Q ({new_AGEMA_signal_2455, KeyArray_outS02ser[4]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S02reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5477, new_AGEMA_signal_5473}), .Q ({new_AGEMA_signal_2458, KeyArray_outS02ser[5]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S02reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5485, new_AGEMA_signal_5481}), .Q ({new_AGEMA_signal_2461, KeyArray_outS02ser[6]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S02reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5493, new_AGEMA_signal_5489}), .Q ({new_AGEMA_signal_2464, KeyArray_outS02ser[7]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S03reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5501, new_AGEMA_signal_5497}), .Q ({new_AGEMA_signal_2467, KeyArray_outS03ser[0]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S03reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5509, new_AGEMA_signal_5505}), .Q ({new_AGEMA_signal_2470, KeyArray_outS03ser[1]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S03reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5517, new_AGEMA_signal_5513}), .Q ({new_AGEMA_signal_2473, KeyArray_outS03ser[2]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S03reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5525, new_AGEMA_signal_5521}), .Q ({new_AGEMA_signal_2476, KeyArray_outS03ser[3]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S03reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5533, new_AGEMA_signal_5529}), .Q ({new_AGEMA_signal_2479, KeyArray_outS03ser[4]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S03reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5541, new_AGEMA_signal_5537}), .Q ({new_AGEMA_signal_2482, KeyArray_outS03ser[5]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S03reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5549, new_AGEMA_signal_5545}), .Q ({new_AGEMA_signal_2485, KeyArray_outS03ser[6]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S03reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5557, new_AGEMA_signal_5553}), .Q ({new_AGEMA_signal_2488, KeyArray_outS03ser[7]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S10reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5565, new_AGEMA_signal_5561}), .Q ({new_AGEMA_signal_2491, KeyArray_outS10ser[0]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S10reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5573, new_AGEMA_signal_5569}), .Q ({new_AGEMA_signal_2494, KeyArray_outS10ser[1]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S10reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5581, new_AGEMA_signal_5577}), .Q ({new_AGEMA_signal_2497, KeyArray_outS10ser[2]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S10reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5589, new_AGEMA_signal_5585}), .Q ({new_AGEMA_signal_2500, KeyArray_outS10ser[3]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S10reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5597, new_AGEMA_signal_5593}), .Q ({new_AGEMA_signal_2503, KeyArray_outS10ser[4]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S10reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5605, new_AGEMA_signal_5601}), .Q ({new_AGEMA_signal_2506, KeyArray_outS10ser[5]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S10reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5613, new_AGEMA_signal_5609}), .Q ({new_AGEMA_signal_2509, KeyArray_outS10ser[6]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S10reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5621, new_AGEMA_signal_5617}), .Q ({new_AGEMA_signal_2512, KeyArray_outS10ser[7]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S11reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5629, new_AGEMA_signal_5625}), .Q ({new_AGEMA_signal_2515, KeyArray_outS11ser[0]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S11reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5637, new_AGEMA_signal_5633}), .Q ({new_AGEMA_signal_2518, KeyArray_outS11ser[1]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S11reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5645, new_AGEMA_signal_5641}), .Q ({new_AGEMA_signal_2521, KeyArray_outS11ser[2]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S11reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5653, new_AGEMA_signal_5649}), .Q ({new_AGEMA_signal_2524, KeyArray_outS11ser[3]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S11reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5661, new_AGEMA_signal_5657}), .Q ({new_AGEMA_signal_2527, KeyArray_outS11ser[4]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S11reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5669, new_AGEMA_signal_5665}), .Q ({new_AGEMA_signal_2530, KeyArray_outS11ser[5]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S11reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5677, new_AGEMA_signal_5673}), .Q ({new_AGEMA_signal_2533, KeyArray_outS11ser[6]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S11reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5685, new_AGEMA_signal_5681}), .Q ({new_AGEMA_signal_2536, KeyArray_outS11ser[7]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S12reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5693, new_AGEMA_signal_5689}), .Q ({new_AGEMA_signal_2539, KeyArray_outS12ser[0]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S12reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5701, new_AGEMA_signal_5697}), .Q ({new_AGEMA_signal_2542, KeyArray_outS12ser[1]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S12reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5709, new_AGEMA_signal_5705}), .Q ({new_AGEMA_signal_2545, KeyArray_outS12ser[2]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S12reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5717, new_AGEMA_signal_5713}), .Q ({new_AGEMA_signal_2548, KeyArray_outS12ser[3]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S12reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5725, new_AGEMA_signal_5721}), .Q ({new_AGEMA_signal_2551, KeyArray_outS12ser[4]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S12reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5733, new_AGEMA_signal_5729}), .Q ({new_AGEMA_signal_2554, KeyArray_outS12ser[5]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S12reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5741, new_AGEMA_signal_5737}), .Q ({new_AGEMA_signal_2557, KeyArray_outS12ser[6]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S12reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5749, new_AGEMA_signal_5745}), .Q ({new_AGEMA_signal_2560, KeyArray_outS12ser[7]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S13reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5757, new_AGEMA_signal_5753}), .Q ({new_AGEMA_signal_2563, keySBIn[0]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S13reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5765, new_AGEMA_signal_5761}), .Q ({new_AGEMA_signal_2566, keySBIn[1]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S13reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5773, new_AGEMA_signal_5769}), .Q ({new_AGEMA_signal_2569, keySBIn[2]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S13reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5781, new_AGEMA_signal_5777}), .Q ({new_AGEMA_signal_2572, keySBIn[3]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S13reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5789, new_AGEMA_signal_5785}), .Q ({new_AGEMA_signal_2575, keySBIn[4]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S13reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5797, new_AGEMA_signal_5793}), .Q ({new_AGEMA_signal_2578, keySBIn[5]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S13reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5805, new_AGEMA_signal_5801}), .Q ({new_AGEMA_signal_2581, keySBIn[6]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S13reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5813, new_AGEMA_signal_5809}), .Q ({new_AGEMA_signal_2584, keySBIn[7]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S20reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5821, new_AGEMA_signal_5817}), .Q ({new_AGEMA_signal_2587, KeyArray_outS20ser[0]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S20reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5829, new_AGEMA_signal_5825}), .Q ({new_AGEMA_signal_2590, KeyArray_outS20ser[1]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S20reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5837, new_AGEMA_signal_5833}), .Q ({new_AGEMA_signal_2593, KeyArray_outS20ser[2]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S20reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5845, new_AGEMA_signal_5841}), .Q ({new_AGEMA_signal_2596, KeyArray_outS20ser[3]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S20reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5853, new_AGEMA_signal_5849}), .Q ({new_AGEMA_signal_2599, KeyArray_outS20ser[4]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S20reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5861, new_AGEMA_signal_5857}), .Q ({new_AGEMA_signal_2602, KeyArray_outS20ser[5]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S20reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5869, new_AGEMA_signal_5865}), .Q ({new_AGEMA_signal_2605, KeyArray_outS20ser[6]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S20reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5877, new_AGEMA_signal_5873}), .Q ({new_AGEMA_signal_2608, KeyArray_outS20ser[7]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S21reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5885, new_AGEMA_signal_5881}), .Q ({new_AGEMA_signal_2611, KeyArray_outS21ser[0]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S21reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5893, new_AGEMA_signal_5889}), .Q ({new_AGEMA_signal_2614, KeyArray_outS21ser[1]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S21reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5901, new_AGEMA_signal_5897}), .Q ({new_AGEMA_signal_2617, KeyArray_outS21ser[2]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S21reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5909, new_AGEMA_signal_5905}), .Q ({new_AGEMA_signal_2620, KeyArray_outS21ser[3]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S21reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5917, new_AGEMA_signal_5913}), .Q ({new_AGEMA_signal_2623, KeyArray_outS21ser[4]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S21reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5925, new_AGEMA_signal_5921}), .Q ({new_AGEMA_signal_2626, KeyArray_outS21ser[5]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S21reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5933, new_AGEMA_signal_5929}), .Q ({new_AGEMA_signal_2629, KeyArray_outS21ser[6]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S21reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5941, new_AGEMA_signal_5937}), .Q ({new_AGEMA_signal_2632, KeyArray_outS21ser[7]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S22reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5949, new_AGEMA_signal_5945}), .Q ({new_AGEMA_signal_2635, KeyArray_outS22ser[0]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S22reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5957, new_AGEMA_signal_5953}), .Q ({new_AGEMA_signal_2638, KeyArray_outS22ser[1]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S22reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5965, new_AGEMA_signal_5961}), .Q ({new_AGEMA_signal_2641, KeyArray_outS22ser[2]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S22reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5973, new_AGEMA_signal_5969}), .Q ({new_AGEMA_signal_2644, KeyArray_outS22ser[3]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S22reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5981, new_AGEMA_signal_5977}), .Q ({new_AGEMA_signal_2647, KeyArray_outS22ser[4]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S22reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5989, new_AGEMA_signal_5985}), .Q ({new_AGEMA_signal_2650, KeyArray_outS22ser[5]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S22reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_5997, new_AGEMA_signal_5993}), .Q ({new_AGEMA_signal_2653, KeyArray_outS22ser[6]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S22reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6005, new_AGEMA_signal_6001}), .Q ({new_AGEMA_signal_2656, KeyArray_outS22ser[7]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S23reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6013, new_AGEMA_signal_6009}), .Q ({new_AGEMA_signal_2659, KeyArray_outS23ser[0]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S23reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6021, new_AGEMA_signal_6017}), .Q ({new_AGEMA_signal_2662, KeyArray_outS23ser[1]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S23reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6029, new_AGEMA_signal_6025}), .Q ({new_AGEMA_signal_2665, KeyArray_outS23ser[2]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S23reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6037, new_AGEMA_signal_6033}), .Q ({new_AGEMA_signal_2668, KeyArray_outS23ser[3]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S23reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6045, new_AGEMA_signal_6041}), .Q ({new_AGEMA_signal_2671, KeyArray_outS23ser[4]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S23reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6053, new_AGEMA_signal_6049}), .Q ({new_AGEMA_signal_2674, KeyArray_outS23ser[5]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S23reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6061, new_AGEMA_signal_6057}), .Q ({new_AGEMA_signal_2677, KeyArray_outS23ser[6]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S23reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6069, new_AGEMA_signal_6065}), .Q ({new_AGEMA_signal_2680, KeyArray_outS23ser[7]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S30reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3512, KeyArray_S30reg_gff_1_SFF_0_n5}), .Q ({new_AGEMA_signal_2683, KeyArray_outS30ser[0]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S30reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3527, KeyArray_S30reg_gff_1_SFF_1_n5}), .Q ({new_AGEMA_signal_2686, KeyArray_outS30ser[1]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S30reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3528, KeyArray_S30reg_gff_1_SFF_2_n5}), .Q ({new_AGEMA_signal_2689, KeyArray_outS30ser[2]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S30reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3529, KeyArray_S30reg_gff_1_SFF_3_n5}), .Q ({new_AGEMA_signal_2692, KeyArray_outS30ser[3]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S30reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3530, KeyArray_S30reg_gff_1_SFF_4_n5}), .Q ({new_AGEMA_signal_2695, KeyArray_outS30ser[4]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S30reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3531, KeyArray_S30reg_gff_1_SFF_5_n5}), .Q ({new_AGEMA_signal_2698, KeyArray_outS30ser[5]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S30reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3532, KeyArray_S30reg_gff_1_SFF_6_n5}), .Q ({new_AGEMA_signal_2701, KeyArray_outS30ser[6]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S30reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3533, KeyArray_S30reg_gff_1_SFF_7_n5}), .Q ({new_AGEMA_signal_2704, KeyArray_outS30ser[7]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S31reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6077, new_AGEMA_signal_6073}), .Q ({new_AGEMA_signal_2707, KeyArray_outS31ser[0]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S31reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6085, new_AGEMA_signal_6081}), .Q ({new_AGEMA_signal_2710, KeyArray_outS31ser[1]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S31reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6093, new_AGEMA_signal_6089}), .Q ({new_AGEMA_signal_2713, KeyArray_outS31ser[2]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S31reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6101, new_AGEMA_signal_6097}), .Q ({new_AGEMA_signal_2716, KeyArray_outS31ser[3]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S31reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6109, new_AGEMA_signal_6105}), .Q ({new_AGEMA_signal_2719, KeyArray_outS31ser[4]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S31reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6117, new_AGEMA_signal_6113}), .Q ({new_AGEMA_signal_2722, KeyArray_outS31ser[5]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S31reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6125, new_AGEMA_signal_6121}), .Q ({new_AGEMA_signal_2725, KeyArray_outS31ser[6]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S31reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6133, new_AGEMA_signal_6129}), .Q ({new_AGEMA_signal_2728, KeyArray_outS31ser[7]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S32reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6141, new_AGEMA_signal_6137}), .Q ({new_AGEMA_signal_2731, KeyArray_outS32ser[0]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S32reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6149, new_AGEMA_signal_6145}), .Q ({new_AGEMA_signal_2734, KeyArray_outS32ser[1]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S32reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6157, new_AGEMA_signal_6153}), .Q ({new_AGEMA_signal_2737, KeyArray_outS32ser[2]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S32reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6165, new_AGEMA_signal_6161}), .Q ({new_AGEMA_signal_2740, KeyArray_outS32ser[3]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S32reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6173, new_AGEMA_signal_6169}), .Q ({new_AGEMA_signal_2743, KeyArray_outS32ser[4]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S32reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6181, new_AGEMA_signal_6177}), .Q ({new_AGEMA_signal_2746, KeyArray_outS32ser[5]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S32reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6189, new_AGEMA_signal_6185}), .Q ({new_AGEMA_signal_2749, KeyArray_outS32ser[6]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S32reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6197, new_AGEMA_signal_6193}), .Q ({new_AGEMA_signal_2752, KeyArray_outS32ser[7]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S33reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6205, new_AGEMA_signal_6201}), .Q ({new_AGEMA_signal_2755, KeyArray_outS33ser[0]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S33reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6213, new_AGEMA_signal_6209}), .Q ({new_AGEMA_signal_2758, KeyArray_outS33ser[1]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S33reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6221, new_AGEMA_signal_6217}), .Q ({new_AGEMA_signal_2761, KeyArray_outS33ser[2]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S33reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6229, new_AGEMA_signal_6225}), .Q ({new_AGEMA_signal_2764, KeyArray_outS33ser[3]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S33reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6237, new_AGEMA_signal_6233}), .Q ({new_AGEMA_signal_2767, KeyArray_outS33ser[4]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S33reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6245, new_AGEMA_signal_6241}), .Q ({new_AGEMA_signal_2770, KeyArray_outS33ser[5]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S33reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6253, new_AGEMA_signal_6249}), .Q ({new_AGEMA_signal_2773, KeyArray_outS33ser[6]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) KeyArray_S33reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6261, new_AGEMA_signal_6257}), .Q ({new_AGEMA_signal_2776, KeyArray_outS33ser[7]}) ) ;
    DFF_X1 calcRCon_s_current_state_reg_0__FF_FF ( .CK (clk), .D (new_AGEMA_signal_6265), .Q (calcRCon_s_current_state_0_), .QN () ) ;
    DFF_X1 calcRCon_s_current_state_reg_1__FF_FF ( .CK (clk), .D (new_AGEMA_signal_6269), .Q (calcRCon_s_current_state_1_), .QN () ) ;
    DFF_X1 calcRCon_s_current_state_reg_2__FF_FF ( .CK (clk), .D (new_AGEMA_signal_6273), .Q (calcRCon_s_current_state_2_), .QN () ) ;
    DFF_X1 calcRCon_s_current_state_reg_3__FF_FF ( .CK (clk), .D (new_AGEMA_signal_6277), .Q (calcRCon_s_current_state_3_), .QN () ) ;
    DFF_X1 calcRCon_s_current_state_reg_4__FF_FF ( .CK (clk), .D (new_AGEMA_signal_6281), .Q (calcRCon_s_current_state_4_), .QN () ) ;
    DFF_X1 calcRCon_s_current_state_reg_5__FF_FF ( .CK (clk), .D (new_AGEMA_signal_6285), .Q (calcRCon_s_current_state_5_), .QN () ) ;
    DFF_X1 calcRCon_s_current_state_reg_6__FF_FF ( .CK (clk), .D (new_AGEMA_signal_6289), .Q (calcRCon_s_current_state_6_), .QN () ) ;
    DFF_X1 calcRCon_s_current_state_reg_7__FF_FF ( .CK (clk), .D (new_AGEMA_signal_6293), .Q (calcRCon_n3), .QN () ) ;
    DFF_X1 nReset_reg_FF_FF ( .CK (clk), .D (new_AGEMA_signal_6297), .Q (nReset), .QN () ) ;
endmodule
