/* modified netlist. Source: module sbox in file ../sbox_lookup/sbox.v */
/* 12 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 13 register stage(s) in total */

module sbox_HPC2_AIG_Pipeline_d2 (SI_s0, clk, SI_s1, SI_s2, Fresh, SO_s0, SO_s1, SO_s2);
    input [3:0] SI_s0 ;
    input clk ;
    input [3:0] SI_s1 ;
    input [3:0] SI_s2 ;
    input [50:0] Fresh ;
    output [3:0] SO_s0 ;
    output [3:0] SO_s1 ;
    output [3:0] SO_s2 ;
    wire signal_15 ;
    wire signal_16 ;
    wire signal_17 ;
    wire signal_18 ;
    wire signal_34 ;
    wire signal_35 ;
    wire signal_36 ;
    wire signal_37 ;
    wire signal_38 ;
    wire signal_39 ;
    wire signal_40 ;
    wire signal_41 ;
    wire signal_42 ;
    wire signal_43 ;
    wire signal_44 ;
    wire signal_45 ;
    wire signal_46 ;
    wire signal_47 ;
    wire signal_48 ;
    wire signal_49 ;
    wire signal_50 ;
    wire signal_51 ;
    wire signal_52 ;
    wire signal_53 ;
    wire signal_54 ;
    wire signal_55 ;
    wire signal_56 ;
    wire signal_57 ;
    wire signal_58 ;
    wire signal_59 ;
    wire signal_60 ;
    wire signal_61 ;
    wire signal_62 ;
    wire signal_63 ;
    wire signal_64 ;
    wire signal_67 ;
    wire signal_68 ;
    wire signal_71 ;
    wire signal_72 ;
    wire signal_75 ;
    wire signal_76 ;
    wire signal_79 ;
    wire signal_80 ;
    wire signal_81 ;
    wire signal_82 ;
    wire signal_83 ;
    wire signal_84 ;
    wire signal_85 ;
    wire signal_86 ;
    wire signal_87 ;
    wire signal_88 ;
    wire signal_89 ;
    wire signal_90 ;
    wire signal_91 ;
    wire signal_92 ;
    wire signal_93 ;
    wire signal_94 ;
    wire signal_95 ;
    wire signal_96 ;
    wire signal_97 ;
    wire signal_98 ;
    wire signal_99 ;
    wire signal_100 ;
    wire signal_101 ;
    wire signal_102 ;
    wire signal_103 ;
    wire signal_104 ;
    wire signal_105 ;
    wire signal_106 ;
    wire signal_107 ;
    wire signal_108 ;
    wire signal_109 ;
    wire signal_110 ;
    wire signal_111 ;
    wire signal_112 ;
    wire signal_113 ;
    wire signal_114 ;
    wire signal_115 ;
    wire signal_116 ;
    wire signal_117 ;
    wire signal_118 ;
    wire signal_119 ;
    wire signal_120 ;
    wire signal_121 ;
    wire signal_122 ;
    wire signal_123 ;
    wire signal_124 ;
    wire signal_125 ;
    wire signal_126 ;
    wire signal_127 ;
    wire signal_128 ;
    wire signal_129 ;
    wire signal_130 ;
    wire signal_131 ;
    wire signal_132 ;
    wire signal_133 ;
    wire signal_134 ;
    wire signal_135 ;
    wire signal_136 ;
    wire signal_137 ;
    wire signal_138 ;
    wire signal_139 ;
    wire signal_140 ;
    wire signal_141 ;
    wire signal_142 ;
    wire signal_202 ;
    wire signal_203 ;
    wire signal_204 ;
    wire signal_205 ;
    wire signal_206 ;
    wire signal_207 ;
    wire signal_208 ;
    wire signal_209 ;
    wire signal_210 ;
    wire signal_211 ;
    wire signal_212 ;
    wire signal_213 ;
    wire signal_214 ;
    wire signal_215 ;
    wire signal_216 ;
    wire signal_217 ;
    wire signal_218 ;
    wire signal_219 ;
    wire signal_220 ;
    wire signal_221 ;
    wire signal_222 ;
    wire signal_223 ;
    wire signal_224 ;
    wire signal_225 ;
    wire signal_226 ;
    wire signal_227 ;
    wire signal_228 ;
    wire signal_229 ;
    wire signal_230 ;
    wire signal_231 ;
    wire signal_232 ;
    wire signal_233 ;
    wire signal_234 ;
    wire signal_235 ;
    wire signal_236 ;
    wire signal_237 ;
    wire signal_238 ;
    wire signal_239 ;
    wire signal_240 ;
    wire signal_241 ;
    wire signal_242 ;
    wire signal_243 ;
    wire signal_244 ;
    wire signal_245 ;
    wire signal_246 ;
    wire signal_247 ;
    wire signal_248 ;
    wire signal_249 ;
    wire signal_250 ;
    wire signal_251 ;
    wire signal_252 ;
    wire signal_253 ;
    wire signal_254 ;
    wire signal_255 ;
    wire signal_256 ;
    wire signal_257 ;
    wire signal_258 ;
    wire signal_259 ;
    wire signal_260 ;
    wire signal_261 ;
    wire signal_262 ;
    wire signal_263 ;
    wire signal_264 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_285 ;
    wire signal_286 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_295 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_352 ;
    wire signal_353 ;
    wire signal_354 ;
    wire signal_355 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_359 ;
    wire signal_360 ;
    wire signal_361 ;
    wire signal_362 ;
    wire signal_363 ;
    wire signal_364 ;
    wire signal_365 ;
    wire signal_366 ;
    wire signal_367 ;
    wire signal_368 ;
    wire signal_369 ;

    /* cells in depth 0 */
    not_masked #(.security_order(2), .pipeline(1)) cell_23 ( .a ({SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_68, signal_67, signal_34}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_24 ( .a ({SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_72, signal_71, signal_35}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_25 ( .a ({SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({signal_76, signal_75, signal_36}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_26 ( .a ({SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({signal_80, signal_79, signal_37}) ) ;

    /* cells in depth 1 */
    buf_clk cell_58 ( .C ( clk ), .D ( SI_s0[3] ), .Q ( signal_202 ) ) ;
    buf_clk cell_60 ( .C ( clk ), .D ( SI_s1[3] ), .Q ( signal_204 ) ) ;
    buf_clk cell_62 ( .C ( clk ), .D ( SI_s2[3] ), .Q ( signal_206 ) ) ;
    buf_clk cell_64 ( .C ( clk ), .D ( SI_s0[0] ), .Q ( signal_208 ) ) ;
    buf_clk cell_66 ( .C ( clk ), .D ( SI_s1[0] ), .Q ( signal_210 ) ) ;
    buf_clk cell_68 ( .C ( clk ), .D ( SI_s2[0] ), .Q ( signal_212 ) ) ;
    buf_clk cell_70 ( .C ( clk ), .D ( SI_s0[2] ), .Q ( signal_214 ) ) ;
    buf_clk cell_72 ( .C ( clk ), .D ( SI_s1[2] ), .Q ( signal_216 ) ) ;
    buf_clk cell_74 ( .C ( clk ), .D ( SI_s2[2] ), .Q ( signal_218 ) ) ;
    buf_clk cell_76 ( .C ( clk ), .D ( signal_34 ), .Q ( signal_220 ) ) ;
    buf_clk cell_78 ( .C ( clk ), .D ( signal_67 ), .Q ( signal_222 ) ) ;
    buf_clk cell_80 ( .C ( clk ), .D ( signal_68 ), .Q ( signal_224 ) ) ;
    buf_clk cell_82 ( .C ( clk ), .D ( signal_36 ), .Q ( signal_226 ) ) ;
    buf_clk cell_84 ( .C ( clk ), .D ( signal_75 ), .Q ( signal_228 ) ) ;
    buf_clk cell_86 ( .C ( clk ), .D ( signal_76 ), .Q ( signal_230 ) ) ;
    buf_clk cell_106 ( .C ( clk ), .D ( SI_s0[1] ), .Q ( signal_250 ) ) ;
    buf_clk cell_112 ( .C ( clk ), .D ( SI_s1[1] ), .Q ( signal_256 ) ) ;
    buf_clk cell_118 ( .C ( clk ), .D ( SI_s2[1] ), .Q ( signal_262 ) ) ;

    /* cells in depth 2 */
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_27 ( .a ({SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[2], Fresh[1], Fresh[0]}), .c ({signal_82, signal_81, signal_38}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_28 ( .a ({SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ({Fresh[5], Fresh[4], Fresh[3]}), .c ({signal_84, signal_83, signal_39}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_29 ( .a ({signal_82, signal_81, signal_38}), .b ({signal_86, signal_85, signal_40}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_30 ( .a ({signal_84, signal_83, signal_39}), .b ({signal_88, signal_87, signal_41}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_31 ( .a ({signal_72, signal_71, signal_35}), .b ({signal_76, signal_75, signal_36}), .clk ( clk ), .r ({Fresh[8], Fresh[7], Fresh[6]}), .c ({signal_90, signal_89, signal_42}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_32 ( .a ({signal_68, signal_67, signal_34}), .b ({signal_80, signal_79, signal_37}), .clk ( clk ), .r ({Fresh[11], Fresh[10], Fresh[9]}), .c ({signal_92, signal_91, signal_43}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_33 ( .a ({signal_72, signal_71, signal_35}), .b ({signal_80, signal_79, signal_37}), .clk ( clk ), .r ({Fresh[14], Fresh[13], Fresh[12]}), .c ({signal_94, signal_93, signal_44}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_34 ( .a ({SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_72, signal_71, signal_35}), .clk ( clk ), .r ({Fresh[17], Fresh[16], Fresh[15]}), .c ({signal_96, signal_95, signal_45}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_35 ( .a ({signal_68, signal_67, signal_34}), .b ({signal_72, signal_71, signal_35}), .clk ( clk ), .r ({Fresh[20], Fresh[19], Fresh[18]}), .c ({signal_98, signal_97, signal_46}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_36 ( .a ({signal_94, signal_93, signal_44}), .b ({signal_100, signal_99, signal_47}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_39 ( .a ({signal_207, signal_205, signal_203}), .b ({signal_90, signal_89, signal_42}), .c ({signal_106, signal_105, signal_16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_40 ( .a ({signal_213, signal_211, signal_209}), .b ({signal_96, signal_95, signal_45}), .c ({signal_108, signal_107, signal_50}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_41 ( .a ({signal_213, signal_211, signal_209}), .b ({signal_98, signal_97, signal_46}), .c ({signal_110, signal_109, signal_15}) ) ;
    buf_clk cell_59 ( .C ( clk ), .D ( signal_202 ), .Q ( signal_203 ) ) ;
    buf_clk cell_61 ( .C ( clk ), .D ( signal_204 ), .Q ( signal_205 ) ) ;
    buf_clk cell_63 ( .C ( clk ), .D ( signal_206 ), .Q ( signal_207 ) ) ;
    buf_clk cell_65 ( .C ( clk ), .D ( signal_208 ), .Q ( signal_209 ) ) ;
    buf_clk cell_67 ( .C ( clk ), .D ( signal_210 ), .Q ( signal_211 ) ) ;
    buf_clk cell_69 ( .C ( clk ), .D ( signal_212 ), .Q ( signal_213 ) ) ;
    buf_clk cell_71 ( .C ( clk ), .D ( signal_214 ), .Q ( signal_215 ) ) ;
    buf_clk cell_73 ( .C ( clk ), .D ( signal_216 ), .Q ( signal_217 ) ) ;
    buf_clk cell_75 ( .C ( clk ), .D ( signal_218 ), .Q ( signal_219 ) ) ;
    buf_clk cell_77 ( .C ( clk ), .D ( signal_220 ), .Q ( signal_221 ) ) ;
    buf_clk cell_79 ( .C ( clk ), .D ( signal_222 ), .Q ( signal_223 ) ) ;
    buf_clk cell_81 ( .C ( clk ), .D ( signal_224 ), .Q ( signal_225 ) ) ;
    buf_clk cell_83 ( .C ( clk ), .D ( signal_226 ), .Q ( signal_227 ) ) ;
    buf_clk cell_85 ( .C ( clk ), .D ( signal_228 ), .Q ( signal_229 ) ) ;
    buf_clk cell_87 ( .C ( clk ), .D ( signal_230 ), .Q ( signal_231 ) ) ;
    buf_clk cell_107 ( .C ( clk ), .D ( signal_250 ), .Q ( signal_251 ) ) ;
    buf_clk cell_113 ( .C ( clk ), .D ( signal_256 ), .Q ( signal_257 ) ) ;
    buf_clk cell_119 ( .C ( clk ), .D ( signal_262 ), .Q ( signal_263 ) ) ;

    /* cells in depth 3 */
    buf_clk cell_88 ( .C ( clk ), .D ( signal_40 ), .Q ( signal_232 ) ) ;
    buf_clk cell_90 ( .C ( clk ), .D ( signal_85 ), .Q ( signal_234 ) ) ;
    buf_clk cell_92 ( .C ( clk ), .D ( signal_86 ), .Q ( signal_236 ) ) ;
    buf_clk cell_94 ( .C ( clk ), .D ( signal_227 ), .Q ( signal_238 ) ) ;
    buf_clk cell_96 ( .C ( clk ), .D ( signal_229 ), .Q ( signal_240 ) ) ;
    buf_clk cell_98 ( .C ( clk ), .D ( signal_231 ), .Q ( signal_242 ) ) ;
    buf_clk cell_100 ( .C ( clk ), .D ( signal_41 ), .Q ( signal_244 ) ) ;
    buf_clk cell_102 ( .C ( clk ), .D ( signal_87 ), .Q ( signal_246 ) ) ;
    buf_clk cell_104 ( .C ( clk ), .D ( signal_88 ), .Q ( signal_248 ) ) ;
    buf_clk cell_108 ( .C ( clk ), .D ( signal_251 ), .Q ( signal_252 ) ) ;
    buf_clk cell_114 ( .C ( clk ), .D ( signal_257 ), .Q ( signal_258 ) ) ;
    buf_clk cell_120 ( .C ( clk ), .D ( signal_263 ), .Q ( signal_264 ) ) ;
    buf_clk cell_148 ( .C ( clk ), .D ( signal_15 ), .Q ( signal_292 ) ) ;
    buf_clk cell_158 ( .C ( clk ), .D ( signal_109 ), .Q ( signal_302 ) ) ;
    buf_clk cell_168 ( .C ( clk ), .D ( signal_110 ), .Q ( signal_312 ) ) ;
    buf_clk cell_178 ( .C ( clk ), .D ( signal_16 ), .Q ( signal_322 ) ) ;
    buf_clk cell_188 ( .C ( clk ), .D ( signal_105 ), .Q ( signal_332 ) ) ;
    buf_clk cell_198 ( .C ( clk ), .D ( signal_106 ), .Q ( signal_342 ) ) ;

    /* cells in depth 4 */
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_37 ( .a ({signal_219, signal_217, signal_215}), .b ({signal_92, signal_91, signal_43}), .clk ( clk ), .r ({Fresh[23], Fresh[22], Fresh[21]}), .c ({signal_102, signal_101, signal_48}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_38 ( .a ({signal_207, signal_205, signal_203}), .b ({signal_94, signal_93, signal_44}), .clk ( clk ), .r ({Fresh[26], Fresh[25], Fresh[24]}), .c ({signal_104, signal_103, signal_49}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_42 ( .a ({signal_102, signal_101, signal_48}), .b ({signal_112, signal_111, signal_51}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_43 ( .a ({signal_104, signal_103, signal_49}), .b ({signal_114, signal_113, signal_52}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_44 ( .a ({signal_225, signal_223, signal_221}), .b ({signal_100, signal_99, signal_47}), .clk ( clk ), .r ({Fresh[29], Fresh[28], Fresh[27]}), .c ({signal_116, signal_115, signal_53}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_45 ( .a ({signal_231, signal_229, signal_227}), .b ({signal_108, signal_107, signal_50}), .clk ( clk ), .r ({Fresh[32], Fresh[31], Fresh[30]}), .c ({signal_118, signal_117, signal_54}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_46 ( .a ({signal_118, signal_117, signal_54}), .b ({signal_120, signal_119, signal_55}) ) ;
    buf_clk cell_89 ( .C ( clk ), .D ( signal_232 ), .Q ( signal_233 ) ) ;
    buf_clk cell_91 ( .C ( clk ), .D ( signal_234 ), .Q ( signal_235 ) ) ;
    buf_clk cell_93 ( .C ( clk ), .D ( signal_236 ), .Q ( signal_237 ) ) ;
    buf_clk cell_95 ( .C ( clk ), .D ( signal_238 ), .Q ( signal_239 ) ) ;
    buf_clk cell_97 ( .C ( clk ), .D ( signal_240 ), .Q ( signal_241 ) ) ;
    buf_clk cell_99 ( .C ( clk ), .D ( signal_242 ), .Q ( signal_243 ) ) ;
    buf_clk cell_101 ( .C ( clk ), .D ( signal_244 ), .Q ( signal_245 ) ) ;
    buf_clk cell_103 ( .C ( clk ), .D ( signal_246 ), .Q ( signal_247 ) ) ;
    buf_clk cell_105 ( .C ( clk ), .D ( signal_248 ), .Q ( signal_249 ) ) ;
    buf_clk cell_109 ( .C ( clk ), .D ( signal_252 ), .Q ( signal_253 ) ) ;
    buf_clk cell_115 ( .C ( clk ), .D ( signal_258 ), .Q ( signal_259 ) ) ;
    buf_clk cell_121 ( .C ( clk ), .D ( signal_264 ), .Q ( signal_265 ) ) ;
    buf_clk cell_149 ( .C ( clk ), .D ( signal_292 ), .Q ( signal_293 ) ) ;
    buf_clk cell_159 ( .C ( clk ), .D ( signal_302 ), .Q ( signal_303 ) ) ;
    buf_clk cell_169 ( .C ( clk ), .D ( signal_312 ), .Q ( signal_313 ) ) ;
    buf_clk cell_179 ( .C ( clk ), .D ( signal_322 ), .Q ( signal_323 ) ) ;
    buf_clk cell_189 ( .C ( clk ), .D ( signal_332 ), .Q ( signal_333 ) ) ;
    buf_clk cell_199 ( .C ( clk ), .D ( signal_342 ), .Q ( signal_343 ) ) ;

    /* cells in depth 5 */
    buf_clk cell_110 ( .C ( clk ), .D ( signal_253 ), .Q ( signal_254 ) ) ;
    buf_clk cell_116 ( .C ( clk ), .D ( signal_259 ), .Q ( signal_260 ) ) ;
    buf_clk cell_122 ( .C ( clk ), .D ( signal_265 ), .Q ( signal_266 ) ) ;
    buf_clk cell_130 ( .C ( clk ), .D ( signal_52 ), .Q ( signal_274 ) ) ;
    buf_clk cell_136 ( .C ( clk ), .D ( signal_113 ), .Q ( signal_280 ) ) ;
    buf_clk cell_142 ( .C ( clk ), .D ( signal_114 ), .Q ( signal_286 ) ) ;
    buf_clk cell_150 ( .C ( clk ), .D ( signal_293 ), .Q ( signal_294 ) ) ;
    buf_clk cell_160 ( .C ( clk ), .D ( signal_303 ), .Q ( signal_304 ) ) ;
    buf_clk cell_170 ( .C ( clk ), .D ( signal_313 ), .Q ( signal_314 ) ) ;
    buf_clk cell_180 ( .C ( clk ), .D ( signal_323 ), .Q ( signal_324 ) ) ;
    buf_clk cell_190 ( .C ( clk ), .D ( signal_333 ), .Q ( signal_334 ) ) ;
    buf_clk cell_200 ( .C ( clk ), .D ( signal_343 ), .Q ( signal_344 ) ) ;

    /* cells in depth 6 */
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_47 ( .a ({signal_237, signal_235, signal_233}), .b ({signal_116, signal_115, signal_53}), .clk ( clk ), .r ({Fresh[35], Fresh[34], Fresh[33]}), .c ({signal_122, signal_121, signal_56}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_48 ( .a ({signal_243, signal_241, signal_239}), .b ({signal_112, signal_111, signal_51}), .clk ( clk ), .r ({Fresh[38], Fresh[37], Fresh[36]}), .c ({signal_124, signal_123, signal_57}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_49 ( .a ({signal_124, signal_123, signal_57}), .b ({signal_126, signal_125, signal_58}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_50 ( .a ({signal_120, signal_119, signal_55}), .b ({signal_249, signal_247, signal_245}), .clk ( clk ), .r ({Fresh[41], Fresh[40], Fresh[39]}), .c ({signal_128, signal_127, signal_59}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_52 ( .a ({signal_128, signal_127, signal_59}), .b ({signal_132, signal_131, signal_17}) ) ;
    buf_clk cell_111 ( .C ( clk ), .D ( signal_254 ), .Q ( signal_255 ) ) ;
    buf_clk cell_117 ( .C ( clk ), .D ( signal_260 ), .Q ( signal_261 ) ) ;
    buf_clk cell_123 ( .C ( clk ), .D ( signal_266 ), .Q ( signal_267 ) ) ;
    buf_clk cell_131 ( .C ( clk ), .D ( signal_274 ), .Q ( signal_275 ) ) ;
    buf_clk cell_137 ( .C ( clk ), .D ( signal_280 ), .Q ( signal_281 ) ) ;
    buf_clk cell_143 ( .C ( clk ), .D ( signal_286 ), .Q ( signal_287 ) ) ;
    buf_clk cell_151 ( .C ( clk ), .D ( signal_294 ), .Q ( signal_295 ) ) ;
    buf_clk cell_161 ( .C ( clk ), .D ( signal_304 ), .Q ( signal_305 ) ) ;
    buf_clk cell_171 ( .C ( clk ), .D ( signal_314 ), .Q ( signal_315 ) ) ;
    buf_clk cell_181 ( .C ( clk ), .D ( signal_324 ), .Q ( signal_325 ) ) ;
    buf_clk cell_191 ( .C ( clk ), .D ( signal_334 ), .Q ( signal_335 ) ) ;
    buf_clk cell_201 ( .C ( clk ), .D ( signal_344 ), .Q ( signal_345 ) ) ;

    /* cells in depth 7 */
    buf_clk cell_124 ( .C ( clk ), .D ( signal_58 ), .Q ( signal_268 ) ) ;
    buf_clk cell_126 ( .C ( clk ), .D ( signal_125 ), .Q ( signal_270 ) ) ;
    buf_clk cell_128 ( .C ( clk ), .D ( signal_126 ), .Q ( signal_272 ) ) ;
    buf_clk cell_132 ( .C ( clk ), .D ( signal_275 ), .Q ( signal_276 ) ) ;
    buf_clk cell_138 ( .C ( clk ), .D ( signal_281 ), .Q ( signal_282 ) ) ;
    buf_clk cell_144 ( .C ( clk ), .D ( signal_287 ), .Q ( signal_288 ) ) ;
    buf_clk cell_152 ( .C ( clk ), .D ( signal_295 ), .Q ( signal_296 ) ) ;
    buf_clk cell_162 ( .C ( clk ), .D ( signal_305 ), .Q ( signal_306 ) ) ;
    buf_clk cell_172 ( .C ( clk ), .D ( signal_315 ), .Q ( signal_316 ) ) ;
    buf_clk cell_182 ( .C ( clk ), .D ( signal_325 ), .Q ( signal_326 ) ) ;
    buf_clk cell_192 ( .C ( clk ), .D ( signal_335 ), .Q ( signal_336 ) ) ;
    buf_clk cell_202 ( .C ( clk ), .D ( signal_345 ), .Q ( signal_346 ) ) ;
    buf_clk cell_208 ( .C ( clk ), .D ( signal_17 ), .Q ( signal_352 ) ) ;
    buf_clk cell_214 ( .C ( clk ), .D ( signal_131 ), .Q ( signal_358 ) ) ;
    buf_clk cell_220 ( .C ( clk ), .D ( signal_132 ), .Q ( signal_364 ) ) ;

    /* cells in depth 8 */
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_51 ( .a ({signal_267, signal_261, signal_255}), .b ({signal_122, signal_121, signal_56}), .clk ( clk ), .r ({Fresh[44], Fresh[43], Fresh[42]}), .c ({signal_130, signal_129, signal_60}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_53 ( .a ({signal_130, signal_129, signal_60}), .b ({signal_134, signal_133, signal_61}) ) ;
    buf_clk cell_125 ( .C ( clk ), .D ( signal_268 ), .Q ( signal_269 ) ) ;
    buf_clk cell_127 ( .C ( clk ), .D ( signal_270 ), .Q ( signal_271 ) ) ;
    buf_clk cell_129 ( .C ( clk ), .D ( signal_272 ), .Q ( signal_273 ) ) ;
    buf_clk cell_133 ( .C ( clk ), .D ( signal_276 ), .Q ( signal_277 ) ) ;
    buf_clk cell_139 ( .C ( clk ), .D ( signal_282 ), .Q ( signal_283 ) ) ;
    buf_clk cell_145 ( .C ( clk ), .D ( signal_288 ), .Q ( signal_289 ) ) ;
    buf_clk cell_153 ( .C ( clk ), .D ( signal_296 ), .Q ( signal_297 ) ) ;
    buf_clk cell_163 ( .C ( clk ), .D ( signal_306 ), .Q ( signal_307 ) ) ;
    buf_clk cell_173 ( .C ( clk ), .D ( signal_316 ), .Q ( signal_317 ) ) ;
    buf_clk cell_183 ( .C ( clk ), .D ( signal_326 ), .Q ( signal_327 ) ) ;
    buf_clk cell_193 ( .C ( clk ), .D ( signal_336 ), .Q ( signal_337 ) ) ;
    buf_clk cell_203 ( .C ( clk ), .D ( signal_346 ), .Q ( signal_347 ) ) ;
    buf_clk cell_209 ( .C ( clk ), .D ( signal_352 ), .Q ( signal_353 ) ) ;
    buf_clk cell_215 ( .C ( clk ), .D ( signal_358 ), .Q ( signal_359 ) ) ;
    buf_clk cell_221 ( .C ( clk ), .D ( signal_364 ), .Q ( signal_365 ) ) ;

    /* cells in depth 9 */
    buf_clk cell_134 ( .C ( clk ), .D ( signal_277 ), .Q ( signal_278 ) ) ;
    buf_clk cell_140 ( .C ( clk ), .D ( signal_283 ), .Q ( signal_284 ) ) ;
    buf_clk cell_146 ( .C ( clk ), .D ( signal_289 ), .Q ( signal_290 ) ) ;
    buf_clk cell_154 ( .C ( clk ), .D ( signal_297 ), .Q ( signal_298 ) ) ;
    buf_clk cell_164 ( .C ( clk ), .D ( signal_307 ), .Q ( signal_308 ) ) ;
    buf_clk cell_174 ( .C ( clk ), .D ( signal_317 ), .Q ( signal_318 ) ) ;
    buf_clk cell_184 ( .C ( clk ), .D ( signal_327 ), .Q ( signal_328 ) ) ;
    buf_clk cell_194 ( .C ( clk ), .D ( signal_337 ), .Q ( signal_338 ) ) ;
    buf_clk cell_204 ( .C ( clk ), .D ( signal_347 ), .Q ( signal_348 ) ) ;
    buf_clk cell_210 ( .C ( clk ), .D ( signal_353 ), .Q ( signal_354 ) ) ;
    buf_clk cell_216 ( .C ( clk ), .D ( signal_359 ), .Q ( signal_360 ) ) ;
    buf_clk cell_222 ( .C ( clk ), .D ( signal_365 ), .Q ( signal_366 ) ) ;

    /* cells in depth 10 */
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_54 ( .a ({signal_273, signal_271, signal_269}), .b ({signal_134, signal_133, signal_61}), .clk ( clk ), .r ({Fresh[47], Fresh[46], Fresh[45]}), .c ({signal_136, signal_135, signal_62}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_55 ( .a ({signal_136, signal_135, signal_62}), .b ({signal_138, signal_137, signal_63}) ) ;
    buf_clk cell_135 ( .C ( clk ), .D ( signal_278 ), .Q ( signal_279 ) ) ;
    buf_clk cell_141 ( .C ( clk ), .D ( signal_284 ), .Q ( signal_285 ) ) ;
    buf_clk cell_147 ( .C ( clk ), .D ( signal_290 ), .Q ( signal_291 ) ) ;
    buf_clk cell_155 ( .C ( clk ), .D ( signal_298 ), .Q ( signal_299 ) ) ;
    buf_clk cell_165 ( .C ( clk ), .D ( signal_308 ), .Q ( signal_309 ) ) ;
    buf_clk cell_175 ( .C ( clk ), .D ( signal_318 ), .Q ( signal_319 ) ) ;
    buf_clk cell_185 ( .C ( clk ), .D ( signal_328 ), .Q ( signal_329 ) ) ;
    buf_clk cell_195 ( .C ( clk ), .D ( signal_338 ), .Q ( signal_339 ) ) ;
    buf_clk cell_205 ( .C ( clk ), .D ( signal_348 ), .Q ( signal_349 ) ) ;
    buf_clk cell_211 ( .C ( clk ), .D ( signal_354 ), .Q ( signal_355 ) ) ;
    buf_clk cell_217 ( .C ( clk ), .D ( signal_360 ), .Q ( signal_361 ) ) ;
    buf_clk cell_223 ( .C ( clk ), .D ( signal_366 ), .Q ( signal_367 ) ) ;

    /* cells in depth 11 */
    buf_clk cell_156 ( .C ( clk ), .D ( signal_299 ), .Q ( signal_300 ) ) ;
    buf_clk cell_166 ( .C ( clk ), .D ( signal_309 ), .Q ( signal_310 ) ) ;
    buf_clk cell_176 ( .C ( clk ), .D ( signal_319 ), .Q ( signal_320 ) ) ;
    buf_clk cell_186 ( .C ( clk ), .D ( signal_329 ), .Q ( signal_330 ) ) ;
    buf_clk cell_196 ( .C ( clk ), .D ( signal_339 ), .Q ( signal_340 ) ) ;
    buf_clk cell_206 ( .C ( clk ), .D ( signal_349 ), .Q ( signal_350 ) ) ;
    buf_clk cell_212 ( .C ( clk ), .D ( signal_355 ), .Q ( signal_356 ) ) ;
    buf_clk cell_218 ( .C ( clk ), .D ( signal_361 ), .Q ( signal_362 ) ) ;
    buf_clk cell_224 ( .C ( clk ), .D ( signal_367 ), .Q ( signal_368 ) ) ;

    /* cells in depth 12 */
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_56 ( .a ({signal_291, signal_285, signal_279}), .b ({signal_138, signal_137, signal_63}), .clk ( clk ), .r ({Fresh[50], Fresh[49], Fresh[48]}), .c ({signal_140, signal_139, signal_64}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_57 ( .a ({signal_140, signal_139, signal_64}), .b ({signal_142, signal_141, signal_18}) ) ;
    buf_clk cell_157 ( .C ( clk ), .D ( signal_300 ), .Q ( signal_301 ) ) ;
    buf_clk cell_167 ( .C ( clk ), .D ( signal_310 ), .Q ( signal_311 ) ) ;
    buf_clk cell_177 ( .C ( clk ), .D ( signal_320 ), .Q ( signal_321 ) ) ;
    buf_clk cell_187 ( .C ( clk ), .D ( signal_330 ), .Q ( signal_331 ) ) ;
    buf_clk cell_197 ( .C ( clk ), .D ( signal_340 ), .Q ( signal_341 ) ) ;
    buf_clk cell_207 ( .C ( clk ), .D ( signal_350 ), .Q ( signal_351 ) ) ;
    buf_clk cell_213 ( .C ( clk ), .D ( signal_356 ), .Q ( signal_357 ) ) ;
    buf_clk cell_219 ( .C ( clk ), .D ( signal_362 ), .Q ( signal_363 ) ) ;
    buf_clk cell_225 ( .C ( clk ), .D ( signal_368 ), .Q ( signal_369 ) ) ;

    /* register cells */
    reg_masked #(.security_order(2), .pipeline(1)) cell_0 ( .clk ( clk ), .D ({signal_321, signal_311, signal_301}), .Q ({SO_s2[3], SO_s1[3], SO_s0[3]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_1 ( .clk ( clk ), .D ({signal_351, signal_341, signal_331}), .Q ({SO_s2[2], SO_s1[2], SO_s0[2]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_2 ( .clk ( clk ), .D ({signal_369, signal_363, signal_357}), .Q ({SO_s2[1], SO_s1[1], SO_s0[1]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_3 ( .clk ( clk ), .D ({signal_142, signal_141, signal_18}), .Q ({SO_s2[0], SO_s1[0], SO_s0[0]}) ) ;
endmodule
