/* modified netlist. Source: module LED in file /LED_round-based/AGEMA/LED.v */
/* clock gating is added to the circuit, the latency increased 4 time(s)  */

module LED_HPC2_AIG_ClockGating_d1 (IN_plaintext_s0, IN_key_s0, IN_reset, CLK, IN_key_s1, IN_plaintext_s1, Fresh, OUT_ciphertext_s0, OUT_done, OUT_ciphertext_s1, Synch);
    input [63:0] IN_plaintext_s0 ;
    input [127:0] IN_key_s0 ;
    input IN_reset ;
    input CLK ;
    input [127:0] IN_key_s1 ;
    input [63:0] IN_plaintext_s1 ;
    input [63:0] Fresh ;
    output [63:0] OUT_ciphertext_s0 ;
    output OUT_done ;
    output [63:0] OUT_ciphertext_s1 ;
    output Synch ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_285 ;
    wire signal_286 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_295 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_356 ;
    wire signal_375 ;
    wire signal_394 ;
    wire signal_413 ;
    wire signal_432 ;
    wire signal_451 ;
    wire signal_470 ;
    wire signal_489 ;
    wire signal_508 ;
    wire signal_527 ;
    wire signal_546 ;
    wire signal_565 ;
    wire signal_584 ;
    wire signal_603 ;
    wire signal_622 ;
    wire signal_641 ;
    wire signal_656 ;
    wire signal_657 ;
    wire signal_658 ;
    wire signal_659 ;
    wire signal_660 ;
    wire signal_661 ;
    wire signal_662 ;
    wire signal_663 ;
    wire signal_664 ;
    wire signal_665 ;
    wire signal_666 ;
    wire signal_667 ;
    wire signal_668 ;
    wire signal_669 ;
    wire signal_670 ;
    wire signal_671 ;
    wire signal_672 ;
    wire signal_673 ;
    wire signal_674 ;
    wire signal_675 ;
    wire signal_676 ;
    wire signal_677 ;
    wire signal_678 ;
    wire signal_679 ;
    wire signal_680 ;
    wire signal_681 ;
    wire signal_682 ;
    wire signal_683 ;
    wire signal_684 ;
    wire signal_685 ;
    wire signal_686 ;
    wire signal_687 ;
    wire signal_688 ;
    wire signal_689 ;
    wire signal_690 ;
    wire signal_691 ;
    wire signal_692 ;
    wire signal_693 ;
    wire signal_694 ;
    wire signal_695 ;
    wire signal_696 ;
    wire signal_697 ;
    wire signal_698 ;
    wire signal_699 ;
    wire signal_700 ;
    wire signal_701 ;
    wire signal_702 ;
    wire signal_703 ;
    wire signal_704 ;
    wire signal_705 ;
    wire signal_706 ;
    wire signal_707 ;
    wire signal_708 ;
    wire signal_709 ;
    wire signal_710 ;
    wire signal_711 ;
    wire signal_712 ;
    wire signal_713 ;
    wire signal_714 ;
    wire signal_715 ;
    wire signal_716 ;
    wire signal_717 ;
    wire signal_718 ;
    wire signal_719 ;
    wire signal_720 ;
    wire signal_721 ;
    wire signal_722 ;
    wire signal_723 ;
    wire signal_724 ;
    wire signal_725 ;
    wire signal_726 ;
    wire signal_727 ;
    wire signal_728 ;
    wire signal_729 ;
    wire signal_730 ;
    wire signal_731 ;
    wire signal_732 ;
    wire signal_733 ;
    wire signal_734 ;
    wire signal_735 ;
    wire signal_736 ;
    wire signal_737 ;
    wire signal_738 ;
    wire signal_739 ;
    wire signal_740 ;
    wire signal_741 ;
    wire signal_742 ;
    wire signal_743 ;
    wire signal_744 ;
    wire signal_745 ;
    wire signal_746 ;
    wire signal_747 ;
    wire signal_748 ;
    wire signal_749 ;
    wire signal_750 ;
    wire signal_751 ;
    wire signal_752 ;
    wire signal_753 ;
    wire signal_754 ;
    wire signal_755 ;
    wire signal_756 ;
    wire signal_757 ;
    wire signal_758 ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_768 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_771 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_774 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_777 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_780 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_783 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_786 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_789 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_792 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_879 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_885 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_888 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_891 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_894 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_897 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_900 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_903 ;
    wire signal_904 ;
    wire signal_905 ;
    wire signal_906 ;
    wire signal_907 ;
    wire signal_908 ;
    wire signal_909 ;
    wire signal_910 ;
    wire signal_911 ;
    wire signal_912 ;
    wire signal_914 ;
    wire signal_915 ;
    wire signal_916 ;
    wire signal_918 ;
    wire signal_919 ;
    wire signal_920 ;
    wire signal_922 ;
    wire signal_923 ;
    wire signal_924 ;
    wire signal_926 ;
    wire signal_927 ;
    wire signal_928 ;
    wire signal_929 ;
    wire signal_930 ;
    wire signal_932 ;
    wire signal_933 ;
    wire signal_934 ;
    wire signal_936 ;
    wire signal_937 ;
    wire signal_938 ;
    wire signal_940 ;
    wire signal_941 ;
    wire signal_942 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1020 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1023 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1276 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1279 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1282 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1285 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1288 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1294 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1297 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1300 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1303 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1309 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1494 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1499 ;
    wire signal_1500 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1503 ;
    wire signal_1504 ;
    wire signal_1505 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1509 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1512 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1518 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1521 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1527 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1530 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1536 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1539 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1564 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1623 ;
    wire signal_1624 ;
    wire signal_1625 ;
    wire signal_1626 ;
    wire signal_1627 ;
    wire signal_1628 ;
    wire signal_1629 ;
    wire signal_1630 ;
    wire signal_1631 ;
    wire signal_1632 ;
    wire signal_1633 ;
    wire signal_1634 ;
    wire signal_1635 ;
    wire signal_1636 ;
    wire signal_1637 ;
    wire signal_1638 ;
    wire signal_1639 ;
    wire signal_1640 ;
    wire signal_1641 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1658 ;
    wire signal_1661 ;
    wire signal_1664 ;
    wire signal_1667 ;
    wire signal_1670 ;
    wire signal_1673 ;
    wire signal_1676 ;
    wire signal_1679 ;
    wire signal_1682 ;
    wire signal_1685 ;
    wire signal_1688 ;
    wire signal_1691 ;
    wire signal_1694 ;
    wire signal_1696 ;
    wire signal_1698 ;
    wire signal_1700 ;
    wire signal_1702 ;
    wire signal_1704 ;
    wire signal_1706 ;
    wire signal_1708 ;
    wire signal_1710 ;
    wire signal_1712 ;
    wire signal_1714 ;
    wire signal_1716 ;
    wire signal_1718 ;
    wire signal_1720 ;
    wire signal_1723 ;
    wire signal_1726 ;
    wire signal_1729 ;
    wire signal_1732 ;
    wire signal_1735 ;
    wire signal_1738 ;
    wire signal_1741 ;
    wire signal_1744 ;
    wire signal_1747 ;
    wire signal_1750 ;
    wire signal_1753 ;
    wire signal_1756 ;
    wire signal_1759 ;
    wire signal_1762 ;
    wire signal_1765 ;
    wire signal_1768 ;
    wire signal_1771 ;
    wire signal_1774 ;
    wire signal_1777 ;
    wire signal_1780 ;
    wire signal_1783 ;
    wire signal_1786 ;
    wire signal_1789 ;
    wire signal_1792 ;
    wire signal_1795 ;
    wire signal_1798 ;
    wire signal_1801 ;
    wire signal_1804 ;
    wire signal_1807 ;
    wire signal_1810 ;
    wire signal_1813 ;
    wire signal_1816 ;
    wire signal_1819 ;
    wire signal_1822 ;
    wire signal_1825 ;
    wire signal_1828 ;
    wire signal_1831 ;
    wire signal_1834 ;
    wire signal_1837 ;
    wire signal_1840 ;
    wire signal_1843 ;
    wire signal_1846 ;
    wire signal_1849 ;
    wire signal_1852 ;
    wire signal_1855 ;
    wire signal_1858 ;
    wire signal_1861 ;
    wire signal_1864 ;
    wire signal_1867 ;
    wire signal_1870 ;
    wire signal_1873 ;
    wire signal_1874 ;
    wire signal_1875 ;
    wire signal_1876 ;
    wire signal_1877 ;
    wire signal_1878 ;
    wire signal_1879 ;
    wire signal_1880 ;
    wire signal_1882 ;
    wire signal_1884 ;
    wire signal_1886 ;
    wire signal_1888 ;
    wire signal_1890 ;
    wire signal_1892 ;
    wire signal_1894 ;
    wire signal_1896 ;
    wire signal_1898 ;
    wire signal_1900 ;
    wire signal_1902 ;
    wire signal_1904 ;
    wire signal_1906 ;
    wire signal_1908 ;
    wire signal_1910 ;
    wire signal_1912 ;
    wire signal_1914 ;
    wire signal_1916 ;
    wire signal_1918 ;
    wire signal_1920 ;
    wire signal_1922 ;
    wire signal_1924 ;
    wire signal_1926 ;
    wire signal_1928 ;
    wire signal_1930 ;
    wire signal_1932 ;
    wire signal_1934 ;
    wire signal_1936 ;
    wire signal_1938 ;
    wire signal_1940 ;
    wire signal_1942 ;
    wire signal_1944 ;
    wire signal_1946 ;
    wire signal_1948 ;
    wire signal_1950 ;
    wire signal_1952 ;
    wire signal_1954 ;
    wire signal_1956 ;
    wire signal_1958 ;
    wire signal_1960 ;
    wire signal_1962 ;
    wire signal_1964 ;
    wire signal_1966 ;
    wire signal_1968 ;
    wire signal_1970 ;
    wire signal_1972 ;
    wire signal_1974 ;
    wire signal_1976 ;
    wire signal_1978 ;
    wire signal_1980 ;
    wire signal_1982 ;
    wire signal_1983 ;
    wire signal_1984 ;
    wire signal_1985 ;
    wire signal_1986 ;
    wire signal_1987 ;
    wire signal_1988 ;
    wire signal_1989 ;
    wire signal_1990 ;
    wire signal_1991 ;
    wire signal_1992 ;
    wire signal_1993 ;
    wire signal_1994 ;
    wire signal_1995 ;
    wire signal_1996 ;
    wire signal_1997 ;
    wire signal_1998 ;
    wire signal_1999 ;
    wire signal_2000 ;
    wire signal_2001 ;
    wire signal_2002 ;
    wire signal_2003 ;
    wire signal_2004 ;
    wire signal_2005 ;
    wire signal_2006 ;
    wire signal_2007 ;
    wire signal_2008 ;
    wire signal_2009 ;
    wire signal_2010 ;
    wire signal_2011 ;
    wire signal_2012 ;
    wire signal_2013 ;
    wire signal_2014 ;
    wire signal_2015 ;
    wire signal_2016 ;
    wire signal_2017 ;
    wire signal_2018 ;
    wire signal_2019 ;
    wire signal_2020 ;
    wire signal_2021 ;
    wire signal_2022 ;
    wire signal_2023 ;
    wire signal_2024 ;
    wire signal_2025 ;
    wire signal_2026 ;
    wire signal_2027 ;
    wire signal_2028 ;
    wire signal_2029 ;
    wire signal_2030 ;
    wire signal_2031 ;
    wire signal_2032 ;
    wire signal_2033 ;
    wire signal_2034 ;
    wire signal_2035 ;
    wire signal_2036 ;
    wire signal_2037 ;
    wire signal_2038 ;
    wire signal_2039 ;
    wire signal_2040 ;
    wire signal_2041 ;
    wire signal_2042 ;
    wire signal_2043 ;
    wire signal_2044 ;
    wire signal_2045 ;
    wire signal_2046 ;
    wire signal_2047 ;
    wire signal_2048 ;
    wire signal_2049 ;
    wire signal_2050 ;
    wire signal_2051 ;
    wire signal_2052 ;
    wire signal_2053 ;
    wire signal_2054 ;
    wire signal_2055 ;
    wire signal_2056 ;
    wire signal_2057 ;
    wire signal_2058 ;
    wire signal_2059 ;
    wire signal_2060 ;
    wire signal_2061 ;
    wire signal_2062 ;
    wire signal_2063 ;
    wire signal_2064 ;
    wire signal_2065 ;
    wire signal_2066 ;
    wire signal_2067 ;
    wire signal_2068 ;
    wire signal_2069 ;
    wire signal_2070 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2079 ;
    wire signal_2080 ;
    wire signal_2081 ;
    wire signal_2082 ;
    wire signal_2083 ;
    wire signal_2084 ;
    wire signal_2085 ;
    wire signal_2086 ;
    wire signal_2087 ;
    wire signal_2088 ;
    wire signal_2089 ;
    wire signal_2090 ;
    wire signal_2091 ;
    wire signal_2092 ;
    wire signal_2093 ;
    wire signal_2094 ;
    wire signal_2095 ;
    wire signal_2096 ;
    wire signal_2097 ;
    wire signal_2098 ;
    wire signal_2099 ;
    wire signal_2100 ;
    wire signal_2101 ;
    wire signal_2102 ;
    wire signal_2103 ;
    wire signal_2104 ;
    wire signal_2105 ;
    wire signal_2106 ;
    wire signal_2107 ;
    wire signal_2108 ;
    wire signal_2109 ;
    wire signal_2110 ;
    wire signal_2111 ;
    wire signal_2112 ;
    wire signal_2113 ;
    wire signal_2114 ;
    wire signal_2115 ;
    wire signal_2116 ;
    wire signal_2117 ;
    wire signal_2118 ;
    wire signal_2119 ;
    wire signal_2120 ;
    wire signal_2121 ;
    wire signal_2122 ;
    wire signal_2123 ;
    wire signal_2124 ;
    wire signal_2125 ;
    wire signal_2126 ;
    wire signal_2127 ;
    wire signal_2128 ;
    wire signal_2129 ;
    wire signal_2130 ;
    wire signal_2131 ;
    wire signal_2132 ;
    wire signal_2133 ;
    wire signal_2134 ;
    wire signal_2135 ;
    wire signal_2136 ;
    wire signal_2137 ;
    wire signal_2138 ;
    wire signal_2139 ;
    wire signal_2140 ;
    wire signal_2141 ;
    wire signal_2142 ;
    wire signal_2143 ;
    wire signal_2144 ;
    wire signal_2145 ;
    wire signal_2146 ;
    wire signal_2147 ;
    wire signal_2148 ;
    wire signal_2149 ;
    wire signal_2150 ;
    wire signal_2151 ;
    wire signal_2152 ;
    wire signal_2153 ;
    wire signal_2154 ;
    wire signal_2155 ;
    wire signal_2156 ;
    wire signal_2157 ;
    wire signal_2158 ;
    wire signal_2159 ;
    wire signal_2160 ;
    wire signal_2161 ;
    wire signal_2162 ;
    wire signal_2163 ;
    wire signal_2164 ;
    wire signal_2165 ;
    wire signal_2166 ;
    wire signal_2167 ;
    wire signal_2168 ;
    wire signal_2169 ;
    wire signal_2170 ;
    wire signal_2171 ;
    wire signal_2172 ;
    wire signal_2173 ;
    wire signal_2174 ;
    wire signal_2175 ;
    wire signal_2176 ;
    wire signal_2177 ;
    wire signal_2178 ;
    wire signal_2179 ;
    wire signal_2180 ;
    wire signal_2181 ;
    wire signal_2182 ;
    wire signal_2183 ;
    wire signal_2184 ;
    wire signal_2185 ;
    wire signal_2186 ;
    wire signal_2187 ;
    wire signal_2188 ;
    wire signal_2189 ;
    wire signal_2190 ;
    wire signal_2191 ;
    wire signal_2192 ;
    wire signal_2193 ;
    wire signal_2194 ;
    wire signal_2195 ;
    wire signal_2196 ;
    wire signal_2197 ;
    wire signal_2198 ;
    wire signal_2199 ;
    wire signal_2200 ;
    wire signal_2201 ;
    wire signal_2202 ;
    wire signal_2203 ;
    wire signal_2204 ;
    wire signal_2205 ;
    wire signal_2206 ;
    wire signal_2207 ;
    wire signal_2208 ;
    wire signal_2209 ;
    wire signal_2210 ;
    wire signal_2211 ;
    wire signal_2212 ;
    wire signal_2213 ;
    wire signal_2214 ;
    wire signal_2215 ;
    wire signal_2216 ;
    wire signal_2217 ;
    wire signal_2218 ;
    wire signal_2219 ;
    wire signal_2220 ;
    wire signal_2221 ;
    wire signal_2222 ;
    wire signal_2223 ;
    wire signal_2224 ;
    wire signal_2225 ;
    wire signal_2226 ;
    wire signal_2227 ;
    wire signal_2228 ;
    wire signal_2229 ;
    wire signal_2230 ;
    wire signal_2231 ;
    wire signal_2232 ;
    wire signal_2233 ;
    wire signal_2234 ;
    wire signal_2235 ;
    wire signal_2236 ;
    wire signal_2237 ;
    wire signal_2238 ;
    wire signal_2239 ;
    wire signal_2240 ;
    wire signal_2241 ;
    wire signal_2242 ;
    wire signal_2243 ;
    wire signal_2244 ;
    wire signal_2245 ;
    wire signal_2246 ;
    wire signal_2247 ;
    wire signal_2248 ;
    wire signal_2249 ;
    wire signal_2250 ;
    wire signal_2251 ;
    wire signal_2252 ;
    wire signal_2253 ;
    wire signal_2254 ;
    wire signal_2255 ;
    wire signal_2256 ;
    wire signal_2257 ;
    wire signal_2258 ;
    wire signal_2259 ;
    wire signal_2260 ;
    wire signal_2261 ;
    wire signal_2262 ;
    wire signal_2263 ;
    wire signal_2264 ;
    wire signal_2265 ;
    wire signal_2266 ;
    wire signal_2267 ;
    wire signal_2268 ;
    wire signal_2269 ;
    wire signal_2270 ;
    wire signal_2271 ;
    wire signal_2272 ;
    wire signal_2273 ;
    wire signal_2274 ;
    wire signal_2275 ;
    wire signal_2276 ;
    wire signal_2277 ;
    wire signal_2278 ;
    wire signal_2279 ;
    wire signal_2280 ;
    wire signal_2281 ;
    wire signal_2282 ;
    wire signal_2283 ;
    wire signal_2284 ;
    wire signal_2285 ;
    wire signal_2286 ;
    wire signal_2287 ;
    wire signal_2288 ;
    wire signal_2289 ;
    wire signal_2290 ;
    wire signal_2291 ;
    wire signal_2292 ;
    wire signal_2293 ;
    wire signal_2294 ;
    wire signal_2295 ;
    wire signal_2296 ;
    wire signal_2297 ;
    wire signal_2298 ;
    wire signal_2299 ;
    wire signal_2300 ;
    wire signal_2301 ;
    wire signal_2302 ;
    wire signal_2303 ;
    wire signal_2304 ;
    wire signal_2305 ;
    wire signal_2306 ;
    wire signal_2307 ;
    wire signal_2308 ;
    wire signal_2309 ;
    wire signal_2310 ;
    wire signal_2311 ;
    wire signal_2312 ;
    wire signal_2313 ;
    wire signal_2314 ;
    wire signal_2315 ;
    wire signal_2316 ;
    wire signal_2317 ;
    wire signal_2318 ;
    wire signal_2319 ;
    wire signal_2320 ;
    wire signal_2321 ;
    wire signal_2322 ;
    wire signal_2323 ;
    wire signal_2324 ;
    wire signal_2325 ;
    wire signal_2326 ;
    wire signal_2327 ;
    wire signal_2328 ;
    wire signal_2329 ;
    wire signal_2330 ;
    wire signal_2331 ;
    wire signal_2332 ;
    wire signal_2333 ;
    wire signal_2334 ;
    wire signal_2335 ;
    wire signal_2336 ;
    wire signal_2337 ;
    wire signal_2338 ;
    wire signal_2339 ;
    wire signal_2340 ;
    wire signal_2341 ;
    wire signal_2342 ;
    wire signal_2343 ;
    wire signal_2344 ;
    wire signal_2345 ;
    wire signal_2346 ;
    wire signal_2347 ;
    wire signal_2348 ;
    wire signal_2349 ;
    wire signal_2350 ;
    wire signal_2351 ;
    wire signal_2352 ;
    wire signal_2353 ;
    wire signal_2354 ;
    wire signal_2355 ;
    wire signal_2356 ;
    wire signal_2357 ;
    wire signal_2358 ;
    wire signal_2359 ;
    wire signal_2360 ;
    wire signal_2361 ;
    wire signal_2362 ;
    wire signal_2363 ;
    wire signal_2364 ;
    wire signal_2365 ;
    wire signal_2366 ;
    wire signal_2367 ;
    wire signal_2368 ;
    wire signal_2369 ;
    wire signal_2370 ;
    wire signal_2371 ;
    wire signal_2372 ;
    wire signal_2373 ;
    wire signal_2374 ;
    wire signal_2375 ;
    wire signal_2376 ;
    wire signal_2377 ;
    wire signal_2378 ;
    wire signal_2379 ;
    wire signal_2380 ;
    wire signal_2381 ;
    wire signal_2382 ;
    wire signal_2383 ;
    wire signal_2384 ;
    wire signal_2385 ;
    wire signal_2386 ;
    wire signal_2387 ;
    wire signal_2388 ;
    wire signal_2389 ;
    wire signal_2390 ;
    wire signal_2391 ;
    wire signal_2392 ;
    wire signal_2393 ;
    wire signal_2394 ;
    wire signal_2395 ;
    wire signal_2396 ;
    wire signal_2397 ;
    wire signal_2398 ;
    wire signal_2399 ;
    wire signal_2400 ;
    wire signal_2401 ;
    wire signal_2402 ;
    wire signal_2403 ;
    wire signal_2404 ;
    wire signal_2405 ;
    wire signal_2406 ;
    wire signal_2407 ;
    wire signal_2408 ;
    wire signal_2409 ;
    wire signal_2410 ;
    wire signal_2411 ;
    wire signal_2412 ;
    wire signal_2413 ;
    wire signal_2414 ;
    wire signal_2415 ;
    wire signal_2416 ;
    wire signal_2417 ;
    wire signal_2418 ;
    wire signal_2419 ;
    wire signal_2420 ;
    wire signal_2421 ;
    wire signal_2422 ;
    wire signal_2423 ;
    wire signal_2424 ;
    wire signal_2425 ;
    wire signal_2426 ;
    wire signal_2427 ;
    wire signal_2428 ;
    wire signal_2429 ;
    wire signal_2430 ;
    wire signal_2431 ;
    wire signal_2432 ;
    wire signal_2433 ;
    wire signal_2434 ;
    wire signal_2435 ;
    wire signal_2436 ;
    wire signal_2437 ;
    wire signal_2438 ;
    wire signal_2439 ;
    wire signal_2440 ;
    wire signal_2441 ;
    wire signal_2442 ;
    wire signal_2443 ;
    wire signal_2444 ;
    wire signal_2445 ;
    wire signal_2446 ;
    wire signal_2447 ;
    wire signal_2448 ;
    wire signal_2449 ;
    wire signal_2450 ;
    wire signal_2451 ;
    wire signal_2452 ;
    wire signal_2453 ;
    wire signal_2454 ;
    wire signal_2455 ;
    wire signal_2456 ;
    wire signal_2457 ;
    wire signal_2458 ;
    wire signal_2459 ;
    wire signal_2460 ;
    wire signal_2461 ;
    wire signal_2462 ;
    wire signal_2463 ;
    wire signal_2464 ;
    wire signal_2465 ;
    wire signal_2466 ;
    wire signal_2467 ;
    wire signal_2468 ;
    wire signal_2469 ;
    wire signal_2470 ;
    wire signal_2471 ;
    wire signal_2472 ;
    wire signal_2473 ;
    wire signal_2474 ;
    wire signal_2475 ;
    wire signal_2476 ;
    wire signal_2477 ;
    wire signal_2478 ;
    wire signal_2479 ;
    wire signal_2480 ;
    wire signal_2481 ;
    wire signal_2482 ;
    wire signal_2483 ;
    wire signal_2484 ;
    wire signal_2485 ;
    wire signal_2486 ;
    wire signal_2487 ;
    wire signal_2488 ;
    wire signal_2489 ;
    wire signal_2490 ;
    wire signal_2491 ;
    wire signal_2492 ;
    wire signal_2493 ;
    wire signal_2494 ;
    wire signal_2495 ;
    wire signal_2496 ;
    wire signal_2497 ;
    wire signal_2498 ;
    wire signal_2499 ;
    wire signal_2500 ;
    wire signal_2501 ;
    wire signal_2502 ;
    wire signal_2503 ;
    wire signal_2504 ;
    wire signal_2505 ;
    wire signal_2506 ;
    wire signal_2507 ;
    wire signal_2508 ;
    wire signal_2509 ;
    wire signal_2510 ;
    wire signal_2511 ;
    wire signal_2512 ;
    wire signal_2513 ;
    wire signal_2514 ;
    wire signal_2515 ;
    wire signal_2516 ;
    wire signal_2517 ;
    wire signal_2518 ;
    wire signal_2519 ;
    wire signal_2520 ;
    wire signal_2521 ;
    wire signal_2522 ;
    wire signal_2523 ;
    wire signal_2524 ;
    wire signal_2525 ;
    wire signal_2526 ;
    wire signal_2527 ;
    wire signal_2528 ;
    wire signal_2529 ;
    wire signal_2530 ;
    wire signal_2531 ;
    wire signal_2532 ;
    wire signal_2533 ;
    wire signal_2534 ;
    wire signal_2535 ;
    wire signal_2536 ;
    wire signal_2537 ;
    wire signal_2538 ;
    wire signal_2539 ;
    wire signal_2540 ;
    wire signal_2541 ;
    wire signal_2542 ;
    wire signal_2543 ;
    wire signal_2544 ;
    wire signal_2545 ;
    wire signal_2546 ;
    wire signal_2547 ;
    wire signal_2548 ;
    wire signal_2549 ;
    wire signal_2550 ;
    wire signal_2551 ;
    wire signal_2552 ;
    wire signal_2553 ;
    wire signal_2554 ;
    wire signal_2555 ;
    wire signal_2556 ;
    wire signal_2557 ;
    wire signal_2558 ;
    wire signal_2559 ;
    wire signal_2561 ;
    wire signal_2562 ;
    wire signal_2563 ;
    wire signal_2564 ;
    wire signal_2565 ;
    wire signal_2566 ;
    wire signal_2567 ;
    wire signal_2568 ;
    wire signal_2569 ;
    wire signal_2570 ;
    wire signal_2571 ;
    wire signal_2572 ;
    wire signal_2573 ;
    wire signal_2574 ;
    wire signal_2575 ;
    wire signal_2576 ;
    wire signal_2577 ;
    wire signal_2578 ;
    wire signal_2579 ;
    wire signal_2580 ;
    wire signal_2581 ;
    wire signal_2582 ;
    wire signal_2583 ;
    wire signal_2584 ;
    wire signal_2585 ;
    wire signal_2587 ;
    wire signal_2589 ;
    wire signal_2591 ;
    wire signal_2593 ;
    wire signal_2595 ;
    wire signal_2597 ;
    wire signal_2599 ;
    wire signal_2601 ;
    wire signal_2603 ;
    wire signal_2604 ;
    wire signal_2605 ;
    wire signal_2606 ;
    wire signal_2607 ;
    wire signal_2608 ;
    wire signal_2609 ;
    wire signal_2610 ;
    wire signal_2611 ;
    wire signal_2612 ;
    wire signal_2613 ;
    wire signal_2614 ;
    wire signal_2615 ;
    wire signal_2616 ;
    wire signal_2617 ;
    wire signal_2618 ;
    wire signal_2619 ;
    wire signal_2620 ;
    wire signal_2621 ;
    wire signal_2622 ;
    wire signal_2623 ;
    wire signal_2624 ;
    wire signal_2625 ;
    wire signal_2626 ;
    wire signal_2627 ;
    wire signal_2628 ;
    wire signal_2629 ;
    wire signal_2630 ;
    wire signal_2631 ;
    wire signal_2632 ;
    wire signal_2633 ;
    wire signal_2634 ;
    wire signal_2635 ;
    wire signal_2637 ;
    wire signal_2639 ;
    wire signal_2641 ;
    wire signal_2643 ;
    wire signal_2644 ;
    wire signal_2645 ;
    wire signal_2646 ;
    wire signal_2647 ;
    wire signal_2648 ;
    wire signal_2649 ;
    wire signal_2650 ;
    wire signal_2651 ;
    wire signal_2652 ;
    wire signal_2653 ;
    wire signal_2654 ;
    wire signal_2655 ;
    wire signal_2656 ;
    wire signal_2657 ;
    wire signal_2658 ;
    wire signal_2659 ;
    wire signal_2660 ;
    wire signal_2661 ;
    wire signal_2662 ;
    wire signal_2663 ;
    wire signal_2664 ;
    wire signal_2665 ;
    wire signal_2666 ;
    wire signal_2667 ;
    wire signal_2668 ;
    wire signal_2669 ;
    wire signal_2670 ;
    wire signal_2671 ;
    wire signal_2672 ;
    wire signal_2673 ;
    wire signal_2674 ;
    wire signal_2675 ;
    wire signal_2676 ;
    wire signal_2677 ;
    wire signal_2679 ;
    wire signal_2681 ;
    wire signal_2683 ;
    wire signal_2685 ;
    wire signal_2687 ;
    wire signal_2689 ;
    wire signal_2691 ;
    wire signal_2693 ;
    wire signal_2694 ;
    wire signal_2695 ;
    wire signal_2696 ;
    wire signal_2697 ;
    wire signal_2698 ;
    wire signal_2699 ;
    wire signal_2700 ;
    wire signal_2701 ;
    wire signal_2702 ;
    wire signal_2703 ;
    wire signal_2704 ;
    wire signal_2705 ;
    wire signal_2706 ;
    wire signal_2707 ;
    wire signal_2708 ;
    wire signal_2709 ;
    wire signal_2710 ;
    wire signal_2711 ;
    wire signal_2712 ;
    wire signal_2713 ;
    wire signal_2714 ;
    wire signal_2715 ;
    wire signal_2716 ;
    wire signal_2717 ;
    wire signal_2718 ;
    wire signal_2719 ;
    wire signal_2720 ;
    wire signal_2721 ;
    wire signal_2722 ;
    wire signal_2723 ;
    wire signal_2724 ;
    wire signal_2725 ;
    wire signal_2726 ;
    wire signal_2728 ;
    wire signal_2730 ;
    wire signal_2732 ;
    wire signal_2734 ;
    wire signal_2736 ;
    wire signal_2738 ;
    wire signal_2740 ;
    wire signal_2742 ;
    wire signal_2743 ;
    wire signal_2744 ;
    wire signal_2745 ;
    wire signal_2746 ;
    wire signal_2747 ;
    wire signal_2748 ;
    wire signal_2749 ;
    wire signal_2750 ;
    wire signal_2751 ;
    wire signal_2752 ;
    wire signal_2753 ;
    wire signal_2754 ;
    wire signal_2755 ;
    wire signal_2756 ;
    wire signal_2757 ;
    wire signal_2758 ;
    wire signal_2759 ;
    wire signal_2760 ;
    wire signal_2761 ;
    wire signal_2763 ;
    wire signal_2765 ;
    wire signal_2767 ;
    wire signal_2769 ;
    wire signal_2771 ;
    wire signal_2773 ;
    wire signal_2775 ;
    wire signal_2777 ;
    wire signal_2779 ;
    wire signal_2781 ;
    wire signal_2783 ;
    wire signal_2785 ;
    wire signal_2786 ;
    wire signal_2787 ;
    wire signal_2788 ;
    wire signal_2789 ;
    wire signal_2790 ;
    wire signal_2791 ;
    wire signal_2792 ;
    wire signal_2793 ;
    wire signal_2794 ;
    wire signal_2795 ;
    wire signal_2796 ;
    wire signal_2797 ;
    wire signal_2798 ;
    wire signal_2799 ;
    wire signal_2800 ;
    wire signal_2801 ;
    wire signal_2803 ;
    wire signal_2805 ;
    wire signal_2807 ;
    wire signal_2809 ;
    wire signal_2811 ;
    wire signal_2813 ;
    wire signal_2815 ;
    wire signal_2816 ;
    wire signal_2817 ;
    wire signal_2818 ;
    wire signal_2819 ;
    wire signal_2820 ;
    wire signal_2821 ;
    wire signal_2823 ;
    wire signal_2825 ;
    wire signal_2827 ;
    wire signal_2829 ;
    wire signal_2831 ;
    wire signal_2833 ;
    wire signal_2835 ;
    wire signal_2836 ;
    wire signal_2837 ;
    wire signal_2838 ;
    wire signal_2839 ;
    wire signal_2840 ;
    wire signal_2841 ;
    wire signal_2842 ;
    wire signal_2843 ;
    wire signal_2844 ;
    wire signal_2845 ;
    wire signal_2846 ;
    wire signal_2847 ;
    wire signal_2848 ;
    wire signal_2849 ;
    wire signal_2850 ;
    wire signal_2851 ;
    wire signal_2852 ;
    wire signal_2853 ;
    wire signal_2854 ;
    wire signal_2855 ;
    wire signal_2857 ;
    wire signal_2859 ;
    wire signal_2860 ;
    wire signal_2861 ;
    wire signal_2862 ;
    wire signal_2863 ;
    wire signal_2865 ;
    wire signal_2867 ;
    wire signal_2869 ;
    wire signal_2871 ;
    wire signal_2873 ;
    wire signal_2875 ;
    wire signal_2940 ;

    /* cells in depth 0 */
    NOR2_X1 cell_0 ( .A1 (signal_875), .A2 (signal_878), .ZN (signal_266) ) ;
    NAND2_X1 cell_1 ( .A1 (signal_879), .A2 (signal_266), .ZN (signal_267) ) ;
    NOR2_X1 cell_2 ( .A1 (signal_874), .A2 (signal_267), .ZN (signal_268) ) ;
    NAND2_X1 cell_3 ( .A1 (signal_876), .A2 (signal_268), .ZN (signal_269) ) ;
    NOR2_X1 cell_4 ( .A1 (signal_877), .A2 (signal_269), .ZN (signal_270) ) ;
    NOR2_X1 cell_5 ( .A1 (OUT_done), .A2 (signal_270), .ZN (signal_271) ) ;
    NOR2_X1 cell_6 ( .A1 (IN_reset), .A2 (signal_271), .ZN (signal_265) ) ;
    NAND2_X1 cell_7 ( .A1 (signal_273), .A2 (signal_274), .ZN (signal_272) ) ;
    XNOR2_X1 cell_8 ( .A (signal_304), .B (signal_275), .ZN (signal_274) ) ;
    XOR2_X1 cell_9 ( .A (signal_309), .B (signal_307), .Z (signal_275) ) ;
    NAND2_X1 cell_10 ( .A1 (signal_276), .A2 (signal_277), .ZN (signal_273) ) ;
    NAND2_X1 cell_11 ( .A1 (signal_278), .A2 (signal_279), .ZN (signal_277) ) ;
    NOR2_X1 cell_12 ( .A1 (signal_302), .A2 (signal_289), .ZN (signal_279) ) ;
    NOR2_X1 cell_13 ( .A1 (signal_306), .A2 (signal_309), .ZN (signal_278) ) ;
    NAND2_X1 cell_14 ( .A1 (signal_289), .A2 (signal_280), .ZN (signal_276) ) ;
    AND2_X1 cell_15 ( .A1 (signal_306), .A2 (signal_309), .ZN (signal_280) ) ;
    NAND2_X1 cell_16 ( .A1 (signal_298), .A2 (signal_283), .ZN (signal_282) ) ;
    NOR2_X1 cell_17 ( .A1 (signal_300), .A2 (signal_284), .ZN (signal_283) ) ;
    NAND2_X1 cell_18 ( .A1 (signal_296), .A2 (signal_876), .ZN (signal_284) ) ;
    NAND2_X1 cell_19 ( .A1 (signal_292), .A2 (signal_290), .ZN (signal_281) ) ;
    NOR2_X1 cell_20 ( .A1 (signal_292), .A2 (IN_reset), .ZN (signal_291) ) ;
    NOR2_X1 cell_21 ( .A1 (IN_reset), .A2 (signal_294), .ZN (signal_293) ) ;
    NOR2_X1 cell_22 ( .A1 (IN_reset), .A2 (signal_296), .ZN (signal_295) ) ;
    NOR2_X1 cell_23 ( .A1 (IN_reset), .A2 (signal_298), .ZN (signal_297) ) ;
    NOR2_X1 cell_24 ( .A1 (IN_reset), .A2 (signal_300), .ZN (signal_299) ) ;
    NOR2_X1 cell_25 ( .A1 (signal_289), .A2 (IN_reset), .ZN (signal_303) ) ;
    NOR2_X1 cell_26 ( .A1 (signal_306), .A2 (IN_reset), .ZN (signal_305) ) ;
    NOR2_X1 cell_27 ( .A1 (signal_309), .A2 (IN_reset), .ZN (signal_308) ) ;
    NOR2_X1 cell_28 ( .A1 (signal_288), .A2 (IN_reset), .ZN (signal_310) ) ;
    OR2_X1 cell_29 ( .A1 (signal_288), .A2 (signal_276), .ZN (signal_286) ) ;
    NAND2_X1 cell_30 ( .A1 (signal_272), .A2 (signal_286), .ZN (signal_311) ) ;
    NOR2_X1 cell_31 ( .A1 (signal_281), .A2 (signal_282), .ZN (signal_340) ) ;
    INV_X1 cell_32 ( .A (signal_286), .ZN (signal_285) ) ;
    OR2_X1 cell_33 ( .A1 (IN_reset), .A2 (signal_287), .ZN (signal_301) ) ;
    XNOR2_X1 cell_34 ( .A (signal_292), .B (signal_290), .ZN (signal_287) ) ;
    INV_X1 cell_35 ( .A (signal_340), .ZN (signal_341) ) ;
    INV_X1 cell_36 ( .A (signal_341), .ZN (signal_344) ) ;
    INV_X1 cell_37 ( .A (signal_341), .ZN (signal_342) ) ;
    INV_X1 cell_38 ( .A (signal_341), .ZN (signal_343) ) ;
    INV_X1 cell_167 ( .A (signal_345), .ZN (signal_346) ) ;
    INV_X1 cell_168 ( .A (signal_285), .ZN (signal_345) ) ;
    INV_X1 cell_169 ( .A (signal_345), .ZN (signal_348) ) ;
    INV_X1 cell_170 ( .A (signal_345), .ZN (signal_347) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_171 ( .s (signal_285), .b ({IN_key_s1[64], IN_key_s0[64]}), .a ({IN_key_s1[0], IN_key_s0[0]}), .c ({signal_1658, signal_1135}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_172 ( .s (signal_346), .b ({IN_key_s1[65], IN_key_s0[65]}), .a ({IN_key_s1[1], IN_key_s0[1]}), .c ({signal_1723, signal_1134}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_173 ( .s (signal_346), .b ({IN_key_s1[66], IN_key_s0[66]}), .a ({IN_key_s1[2], IN_key_s0[2]}), .c ({signal_1726, signal_1133}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_174 ( .s (signal_285), .b ({IN_key_s1[67], IN_key_s0[67]}), .a ({IN_key_s1[3], IN_key_s0[3]}), .c ({signal_1661, signal_1132}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_175 ( .s (signal_346), .b ({IN_key_s1[68], IN_key_s0[68]}), .a ({IN_key_s1[4], IN_key_s0[4]}), .c ({signal_1729, signal_1131}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_176 ( .s (signal_346), .b ({IN_key_s1[69], IN_key_s0[69]}), .a ({IN_key_s1[5], IN_key_s0[5]}), .c ({signal_1732, signal_1130}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_177 ( .s (signal_346), .b ({IN_key_s1[70], IN_key_s0[70]}), .a ({IN_key_s1[6], IN_key_s0[6]}), .c ({signal_1735, signal_1129}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_178 ( .s (signal_346), .b ({IN_key_s1[71], IN_key_s0[71]}), .a ({IN_key_s1[7], IN_key_s0[7]}), .c ({signal_1738, signal_1128}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_179 ( .s (signal_346), .b ({IN_key_s1[72], IN_key_s0[72]}), .a ({IN_key_s1[8], IN_key_s0[8]}), .c ({signal_1741, signal_1127}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_180 ( .s (signal_346), .b ({IN_key_s1[73], IN_key_s0[73]}), .a ({IN_key_s1[9], IN_key_s0[9]}), .c ({signal_1744, signal_1126}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_181 ( .s (signal_346), .b ({IN_key_s1[74], IN_key_s0[74]}), .a ({IN_key_s1[10], IN_key_s0[10]}), .c ({signal_1747, signal_1125}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_182 ( .s (signal_346), .b ({IN_key_s1[75], IN_key_s0[75]}), .a ({IN_key_s1[11], IN_key_s0[11]}), .c ({signal_1750, signal_1124}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_183 ( .s (signal_346), .b ({IN_key_s1[76], IN_key_s0[76]}), .a ({IN_key_s1[12], IN_key_s0[12]}), .c ({signal_1753, signal_1123}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_184 ( .s (signal_346), .b ({IN_key_s1[77], IN_key_s0[77]}), .a ({IN_key_s1[13], IN_key_s0[13]}), .c ({signal_1756, signal_1122}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_185 ( .s (signal_346), .b ({IN_key_s1[78], IN_key_s0[78]}), .a ({IN_key_s1[14], IN_key_s0[14]}), .c ({signal_1759, signal_1121}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_186 ( .s (signal_346), .b ({IN_key_s1[79], IN_key_s0[79]}), .a ({IN_key_s1[15], IN_key_s0[15]}), .c ({signal_1762, signal_1120}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_187 ( .s (signal_285), .b ({IN_key_s1[80], IN_key_s0[80]}), .a ({IN_key_s1[16], IN_key_s0[16]}), .c ({signal_1664, signal_1119}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_188 ( .s (signal_347), .b ({IN_key_s1[81], IN_key_s0[81]}), .a ({IN_key_s1[17], IN_key_s0[17]}), .c ({signal_1765, signal_1118}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_189 ( .s (signal_348), .b ({IN_key_s1[82], IN_key_s0[82]}), .a ({IN_key_s1[18], IN_key_s0[18]}), .c ({signal_1768, signal_1117}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_190 ( .s (signal_285), .b ({IN_key_s1[83], IN_key_s0[83]}), .a ({IN_key_s1[19], IN_key_s0[19]}), .c ({signal_1667, signal_1116}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_191 ( .s (signal_346), .b ({IN_key_s1[84], IN_key_s0[84]}), .a ({IN_key_s1[20], IN_key_s0[20]}), .c ({signal_1771, signal_1115}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_192 ( .s (signal_348), .b ({IN_key_s1[85], IN_key_s0[85]}), .a ({IN_key_s1[21], IN_key_s0[21]}), .c ({signal_1774, signal_1114}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_193 ( .s (signal_285), .b ({IN_key_s1[86], IN_key_s0[86]}), .a ({IN_key_s1[22], IN_key_s0[22]}), .c ({signal_1670, signal_1113}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_194 ( .s (signal_348), .b ({IN_key_s1[87], IN_key_s0[87]}), .a ({IN_key_s1[23], IN_key_s0[23]}), .c ({signal_1777, signal_1112}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_195 ( .s (signal_285), .b ({IN_key_s1[88], IN_key_s0[88]}), .a ({IN_key_s1[24], IN_key_s0[24]}), .c ({signal_1673, signal_1111}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_196 ( .s (signal_348), .b ({IN_key_s1[89], IN_key_s0[89]}), .a ({IN_key_s1[25], IN_key_s0[25]}), .c ({signal_1780, signal_1110}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_197 ( .s (signal_285), .b ({IN_key_s1[90], IN_key_s0[90]}), .a ({IN_key_s1[26], IN_key_s0[26]}), .c ({signal_1676, signal_1109}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_198 ( .s (signal_348), .b ({IN_key_s1[91], IN_key_s0[91]}), .a ({IN_key_s1[27], IN_key_s0[27]}), .c ({signal_1783, signal_1108}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_199 ( .s (signal_285), .b ({IN_key_s1[92], IN_key_s0[92]}), .a ({IN_key_s1[28], IN_key_s0[28]}), .c ({signal_1679, signal_1107}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_200 ( .s (signal_347), .b ({IN_key_s1[93], IN_key_s0[93]}), .a ({IN_key_s1[29], IN_key_s0[29]}), .c ({signal_1786, signal_1106}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_201 ( .s (signal_347), .b ({IN_key_s1[94], IN_key_s0[94]}), .a ({IN_key_s1[30], IN_key_s0[30]}), .c ({signal_1789, signal_1105}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_202 ( .s (signal_347), .b ({IN_key_s1[95], IN_key_s0[95]}), .a ({IN_key_s1[31], IN_key_s0[31]}), .c ({signal_1792, signal_1104}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_203 ( .s (signal_285), .b ({IN_key_s1[96], IN_key_s0[96]}), .a ({IN_key_s1[32], IN_key_s0[32]}), .c ({signal_1682, signal_1103}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_204 ( .s (signal_348), .b ({IN_key_s1[97], IN_key_s0[97]}), .a ({IN_key_s1[33], IN_key_s0[33]}), .c ({signal_1795, signal_1102}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_205 ( .s (signal_285), .b ({IN_key_s1[98], IN_key_s0[98]}), .a ({IN_key_s1[34], IN_key_s0[34]}), .c ({signal_1685, signal_1101}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_206 ( .s (signal_285), .b ({IN_key_s1[99], IN_key_s0[99]}), .a ({IN_key_s1[35], IN_key_s0[35]}), .c ({signal_1688, signal_1100}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_207 ( .s (signal_285), .b ({IN_key_s1[100], IN_key_s0[100]}), .a ({IN_key_s1[36], IN_key_s0[36]}), .c ({signal_1691, signal_1099}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_208 ( .s (signal_347), .b ({IN_key_s1[101], IN_key_s0[101]}), .a ({IN_key_s1[37], IN_key_s0[37]}), .c ({signal_1798, signal_1098}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_209 ( .s (signal_347), .b ({IN_key_s1[102], IN_key_s0[102]}), .a ({IN_key_s1[38], IN_key_s0[38]}), .c ({signal_1801, signal_1097}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_210 ( .s (signal_285), .b ({IN_key_s1[103], IN_key_s0[103]}), .a ({IN_key_s1[39], IN_key_s0[39]}), .c ({signal_1694, signal_1096}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_211 ( .s (signal_347), .b ({IN_key_s1[104], IN_key_s0[104]}), .a ({IN_key_s1[40], IN_key_s0[40]}), .c ({signal_1804, signal_1095}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_212 ( .s (signal_347), .b ({IN_key_s1[105], IN_key_s0[105]}), .a ({IN_key_s1[41], IN_key_s0[41]}), .c ({signal_1807, signal_1094}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_213 ( .s (signal_347), .b ({IN_key_s1[106], IN_key_s0[106]}), .a ({IN_key_s1[42], IN_key_s0[42]}), .c ({signal_1810, signal_1093}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_214 ( .s (signal_347), .b ({IN_key_s1[107], IN_key_s0[107]}), .a ({IN_key_s1[43], IN_key_s0[43]}), .c ({signal_1813, signal_1092}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_215 ( .s (signal_347), .b ({IN_key_s1[108], IN_key_s0[108]}), .a ({IN_key_s1[44], IN_key_s0[44]}), .c ({signal_1816, signal_1091}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_216 ( .s (signal_347), .b ({IN_key_s1[109], IN_key_s0[109]}), .a ({IN_key_s1[45], IN_key_s0[45]}), .c ({signal_1819, signal_1090}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_217 ( .s (signal_347), .b ({IN_key_s1[110], IN_key_s0[110]}), .a ({IN_key_s1[46], IN_key_s0[46]}), .c ({signal_1822, signal_1089}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_218 ( .s (signal_347), .b ({IN_key_s1[111], IN_key_s0[111]}), .a ({IN_key_s1[47], IN_key_s0[47]}), .c ({signal_1825, signal_1088}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_219 ( .s (signal_347), .b ({IN_key_s1[112], IN_key_s0[112]}), .a ({IN_key_s1[48], IN_key_s0[48]}), .c ({signal_1828, signal_1087}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_220 ( .s (signal_347), .b ({IN_key_s1[113], IN_key_s0[113]}), .a ({IN_key_s1[49], IN_key_s0[49]}), .c ({signal_1831, signal_1086}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_221 ( .s (signal_347), .b ({IN_key_s1[114], IN_key_s0[114]}), .a ({IN_key_s1[50], IN_key_s0[50]}), .c ({signal_1834, signal_1085}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_222 ( .s (signal_347), .b ({IN_key_s1[115], IN_key_s0[115]}), .a ({IN_key_s1[51], IN_key_s0[51]}), .c ({signal_1837, signal_1084}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_223 ( .s (signal_348), .b ({IN_key_s1[116], IN_key_s0[116]}), .a ({IN_key_s1[52], IN_key_s0[52]}), .c ({signal_1840, signal_1083}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_224 ( .s (signal_348), .b ({IN_key_s1[117], IN_key_s0[117]}), .a ({IN_key_s1[53], IN_key_s0[53]}), .c ({signal_1843, signal_1082}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_225 ( .s (signal_348), .b ({IN_key_s1[118], IN_key_s0[118]}), .a ({IN_key_s1[54], IN_key_s0[54]}), .c ({signal_1846, signal_1081}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_226 ( .s (signal_348), .b ({IN_key_s1[119], IN_key_s0[119]}), .a ({IN_key_s1[55], IN_key_s0[55]}), .c ({signal_1849, signal_1080}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_227 ( .s (signal_348), .b ({IN_key_s1[120], IN_key_s0[120]}), .a ({IN_key_s1[56], IN_key_s0[56]}), .c ({signal_1852, signal_1079}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_228 ( .s (signal_348), .b ({IN_key_s1[121], IN_key_s0[121]}), .a ({IN_key_s1[57], IN_key_s0[57]}), .c ({signal_1855, signal_1078}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_229 ( .s (signal_348), .b ({IN_key_s1[122], IN_key_s0[122]}), .a ({IN_key_s1[58], IN_key_s0[58]}), .c ({signal_1858, signal_1077}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_230 ( .s (signal_348), .b ({IN_key_s1[123], IN_key_s0[123]}), .a ({IN_key_s1[59], IN_key_s0[59]}), .c ({signal_1861, signal_1076}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_231 ( .s (signal_348), .b ({IN_key_s1[124], IN_key_s0[124]}), .a ({IN_key_s1[60], IN_key_s0[60]}), .c ({signal_1864, signal_1075}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_232 ( .s (signal_348), .b ({IN_key_s1[125], IN_key_s0[125]}), .a ({IN_key_s1[61], IN_key_s0[61]}), .c ({signal_1867, signal_1074}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_233 ( .s (signal_348), .b ({IN_key_s1[126], IN_key_s0[126]}), .a ({IN_key_s1[62], IN_key_s0[62]}), .c ({signal_1870, signal_1073}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_234 ( .s (signal_348), .b ({IN_key_s1[127], IN_key_s0[127]}), .a ({IN_key_s1[63], IN_key_s0[63]}), .c ({signal_1873, signal_1072}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_235 ( .a ({OUT_ciphertext_s1[9], OUT_ciphertext_s0[9]}), .b ({signal_1744, signal_1126}), .c ({signal_1882, signal_1062}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_236 ( .a ({OUT_ciphertext_s1[8], OUT_ciphertext_s0[8]}), .b ({signal_1741, signal_1127}), .c ({signal_1884, signal_1063}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_237 ( .a ({OUT_ciphertext_s1[7], OUT_ciphertext_s0[7]}), .b ({signal_1738, signal_1128}), .c ({signal_1886, signal_1064}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_238 ( .a ({OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}), .b ({signal_1735, signal_1129}), .c ({signal_1888, signal_1065}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_239 ( .a ({OUT_ciphertext_s1[63], OUT_ciphertext_s0[63]}), .b ({signal_1873, signal_1072}), .c ({signal_1890, signal_1008}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_240 ( .a ({OUT_ciphertext_s1[62], OUT_ciphertext_s0[62]}), .b ({signal_1870, signal_1073}), .c ({signal_1892, signal_1009}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_241 ( .a ({OUT_ciphertext_s1[61], OUT_ciphertext_s0[61]}), .b ({signal_1867, signal_1074}), .c ({signal_1894, signal_1010}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_242 ( .a ({OUT_ciphertext_s1[60], OUT_ciphertext_s0[60]}), .b ({signal_1864, signal_1075}), .c ({signal_1896, signal_1011}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_243 ( .a ({OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}), .b ({signal_1732, signal_1130}), .c ({signal_1898, signal_1066}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_244 ( .a ({OUT_ciphertext_s1[59], OUT_ciphertext_s0[59]}), .b ({signal_1861, signal_1076}), .c ({signal_1900, signal_1012}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_245 ( .a ({OUT_ciphertext_s1[58], OUT_ciphertext_s0[58]}), .b ({signal_1858, signal_1077}), .c ({signal_1902, signal_1013}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_246 ( .a ({OUT_ciphertext_s1[57], OUT_ciphertext_s0[57]}), .b ({signal_1855, signal_1078}), .c ({signal_1904, signal_1014}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_247 ( .a ({OUT_ciphertext_s1[56], OUT_ciphertext_s0[56]}), .b ({signal_1852, signal_1079}), .c ({signal_1906, signal_1015}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_248 ( .a ({OUT_ciphertext_s1[55], OUT_ciphertext_s0[55]}), .b ({signal_1849, signal_1080}), .c ({signal_1908, signal_1016}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_249 ( .a ({OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}), .b ({signal_1846, signal_1081}), .c ({signal_1910, signal_1017}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_250 ( .a ({OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}), .b ({signal_1843, signal_1082}), .c ({signal_1912, signal_1018}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_251 ( .a ({OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}), .b ({signal_1840, signal_1083}), .c ({signal_1914, signal_1019}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_252 ( .a ({OUT_ciphertext_s1[51], OUT_ciphertext_s0[51]}), .b ({signal_1837, signal_1084}), .c ({signal_1916, signal_1020}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_253 ( .a ({OUT_ciphertext_s1[50], OUT_ciphertext_s0[50]}), .b ({signal_1834, signal_1085}), .c ({signal_1918, signal_1021}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_254 ( .a ({OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}), .b ({signal_1729, signal_1131}), .c ({signal_1920, signal_1067}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_255 ( .a ({OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}), .b ({signal_1831, signal_1086}), .c ({signal_1922, signal_1022}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_256 ( .a ({OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}), .b ({signal_1828, signal_1087}), .c ({signal_1924, signal_1023}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_257 ( .a ({OUT_ciphertext_s1[47], OUT_ciphertext_s0[47]}), .b ({signal_1825, signal_1088}), .c ({signal_1926, signal_1024}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_258 ( .a ({OUT_ciphertext_s1[46], OUT_ciphertext_s0[46]}), .b ({signal_1822, signal_1089}), .c ({signal_1928, signal_1025}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_259 ( .a ({OUT_ciphertext_s1[45], OUT_ciphertext_s0[45]}), .b ({signal_1819, signal_1090}), .c ({signal_1930, signal_1026}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_260 ( .a ({OUT_ciphertext_s1[44], OUT_ciphertext_s0[44]}), .b ({signal_1816, signal_1091}), .c ({signal_1932, signal_1027}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_261 ( .a ({OUT_ciphertext_s1[43], OUT_ciphertext_s0[43]}), .b ({signal_1813, signal_1092}), .c ({signal_1934, signal_1028}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_262 ( .a ({OUT_ciphertext_s1[42], OUT_ciphertext_s0[42]}), .b ({signal_1810, signal_1093}), .c ({signal_1936, signal_1029}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_263 ( .a ({OUT_ciphertext_s1[41], OUT_ciphertext_s0[41]}), .b ({signal_1807, signal_1094}), .c ({signal_1938, signal_1030}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_264 ( .a ({OUT_ciphertext_s1[40], OUT_ciphertext_s0[40]}), .b ({signal_1804, signal_1095}), .c ({signal_1940, signal_1031}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_265 ( .a ({OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}), .b ({signal_1661, signal_1132}), .c ({signal_1696, signal_1068}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_266 ( .a ({OUT_ciphertext_s1[39], OUT_ciphertext_s0[39]}), .b ({signal_1694, signal_1096}), .c ({signal_1698, signal_1032}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_267 ( .a ({OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}), .b ({signal_1801, signal_1097}), .c ({signal_1942, signal_1033}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_268 ( .a ({OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}), .b ({signal_1798, signal_1098}), .c ({signal_1944, signal_1034}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_269 ( .a ({OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}), .b ({signal_1691, signal_1099}), .c ({signal_1700, signal_1035}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_270 ( .a ({OUT_ciphertext_s1[35], OUT_ciphertext_s0[35]}), .b ({signal_1688, signal_1100}), .c ({signal_1702, signal_1036}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_271 ( .a ({OUT_ciphertext_s1[34], OUT_ciphertext_s0[34]}), .b ({signal_1685, signal_1101}), .c ({signal_1704, signal_1037}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_272 ( .a ({OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}), .b ({signal_1795, signal_1102}), .c ({signal_1946, signal_1038}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_273 ( .a ({OUT_ciphertext_s1[32], OUT_ciphertext_s0[32]}), .b ({signal_1682, signal_1103}), .c ({signal_1706, signal_1039}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_274 ( .a ({OUT_ciphertext_s1[31], OUT_ciphertext_s0[31]}), .b ({signal_1792, signal_1104}), .c ({signal_1948, signal_1040}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_275 ( .a ({OUT_ciphertext_s1[30], OUT_ciphertext_s0[30]}), .b ({signal_1789, signal_1105}), .c ({signal_1950, signal_1041}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_276 ( .a ({OUT_ciphertext_s1[2], OUT_ciphertext_s0[2]}), .b ({signal_1726, signal_1133}), .c ({signal_1952, signal_1069}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_277 ( .a ({OUT_ciphertext_s1[29], OUT_ciphertext_s0[29]}), .b ({signal_1786, signal_1106}), .c ({signal_1954, signal_1042}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_278 ( .a ({OUT_ciphertext_s1[28], OUT_ciphertext_s0[28]}), .b ({signal_1679, signal_1107}), .c ({signal_1708, signal_1043}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_279 ( .a ({OUT_ciphertext_s1[27], OUT_ciphertext_s0[27]}), .b ({signal_1783, signal_1108}), .c ({signal_1956, signal_1044}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_280 ( .a ({OUT_ciphertext_s1[26], OUT_ciphertext_s0[26]}), .b ({signal_1676, signal_1109}), .c ({signal_1710, signal_1045}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_281 ( .a ({OUT_ciphertext_s1[25], OUT_ciphertext_s0[25]}), .b ({signal_1780, signal_1110}), .c ({signal_1958, signal_1046}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_282 ( .a ({OUT_ciphertext_s1[24], OUT_ciphertext_s0[24]}), .b ({signal_1673, signal_1111}), .c ({signal_1712, signal_1047}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_283 ( .a ({OUT_ciphertext_s1[23], OUT_ciphertext_s0[23]}), .b ({signal_1777, signal_1112}), .c ({signal_1960, signal_1048}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_284 ( .a ({OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}), .b ({signal_1670, signal_1113}), .c ({signal_1714, signal_1049}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_285 ( .a ({OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}), .b ({signal_1774, signal_1114}), .c ({signal_1962, signal_1050}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_286 ( .a ({OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}), .b ({signal_1771, signal_1115}), .c ({signal_1964, signal_1051}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_287 ( .a ({OUT_ciphertext_s1[1], OUT_ciphertext_s0[1]}), .b ({signal_1723, signal_1134}), .c ({signal_1966, signal_1070}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_288 ( .a ({OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}), .b ({signal_1667, signal_1116}), .c ({signal_1716, signal_1052}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_289 ( .a ({OUT_ciphertext_s1[18], OUT_ciphertext_s0[18]}), .b ({signal_1768, signal_1117}), .c ({signal_1968, signal_1053}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_290 ( .a ({OUT_ciphertext_s1[17], OUT_ciphertext_s0[17]}), .b ({signal_1765, signal_1118}), .c ({signal_1970, signal_1054}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_291 ( .a ({OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}), .b ({signal_1664, signal_1119}), .c ({signal_1718, signal_1055}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_292 ( .a ({OUT_ciphertext_s1[15], OUT_ciphertext_s0[15]}), .b ({signal_1762, signal_1120}), .c ({signal_1972, signal_1056}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_293 ( .a ({OUT_ciphertext_s1[14], OUT_ciphertext_s0[14]}), .b ({signal_1759, signal_1121}), .c ({signal_1974, signal_1057}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_294 ( .a ({OUT_ciphertext_s1[13], OUT_ciphertext_s0[13]}), .b ({signal_1756, signal_1122}), .c ({signal_1976, signal_1058}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_295 ( .a ({OUT_ciphertext_s1[12], OUT_ciphertext_s0[12]}), .b ({signal_1753, signal_1123}), .c ({signal_1978, signal_1059}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_296 ( .a ({OUT_ciphertext_s1[11], OUT_ciphertext_s0[11]}), .b ({signal_1750, signal_1124}), .c ({signal_1980, signal_1060}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_297 ( .a ({OUT_ciphertext_s1[10], OUT_ciphertext_s0[10]}), .b ({signal_1747, signal_1125}), .c ({signal_1982, signal_1061}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_298 ( .a ({OUT_ciphertext_s1[0], OUT_ciphertext_s0[0]}), .b ({signal_1658, signal_1135}), .c ({signal_1720, signal_1071}) ) ;
    INV_X1 cell_299 ( .A (signal_349), .ZN (signal_351) ) ;
    INV_X1 cell_300 ( .A (signal_311), .ZN (signal_349) ) ;
    INV_X1 cell_301 ( .A (signal_349), .ZN (signal_350) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_302 ( .s (signal_311), .b ({OUT_ciphertext_s1[0], OUT_ciphertext_s0[0]}), .a ({signal_1720, signal_1071}), .c ({signal_1874, signal_312}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_303 ( .s (signal_311), .b ({OUT_ciphertext_s1[1], OUT_ciphertext_s0[1]}), .a ({signal_1966, signal_1070}), .c ({signal_1994, signal_313}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_304 ( .s (signal_311), .b ({OUT_ciphertext_s1[2], OUT_ciphertext_s0[2]}), .a ({signal_1952, signal_1069}), .c ({signal_1995, signal_314}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_305 ( .s (signal_311), .b ({OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}), .a ({signal_1696, signal_1068}), .c ({signal_1875, signal_315}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_306 ( .s (signal_350), .b ({OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}), .a ({signal_1920, signal_1067}), .c ({signal_1996, signal_316}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_307 ( .s (signal_350), .b ({OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}), .a ({signal_1898, signal_1066}), .c ({signal_1997, signal_317}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_308 ( .s (signal_350), .b ({OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}), .a ({signal_1888, signal_1065}), .c ({signal_1998, signal_318}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_309 ( .s (signal_350), .b ({OUT_ciphertext_s1[7], OUT_ciphertext_s0[7]}), .a ({signal_1886, signal_1064}), .c ({signal_1999, signal_1000}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_310 ( .s (signal_350), .b ({OUT_ciphertext_s1[8], OUT_ciphertext_s0[8]}), .a ({signal_1884, signal_1063}), .c ({signal_2000, signal_999}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_311 ( .s (signal_350), .b ({OUT_ciphertext_s1[9], OUT_ciphertext_s0[9]}), .a ({signal_1882, signal_1062}), .c ({signal_2001, signal_998}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_312 ( .s (signal_350), .b ({OUT_ciphertext_s1[10], OUT_ciphertext_s0[10]}), .a ({signal_1982, signal_1061}), .c ({signal_2002, signal_997}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_313 ( .s (signal_350), .b ({OUT_ciphertext_s1[11], OUT_ciphertext_s0[11]}), .a ({signal_1980, signal_1060}), .c ({signal_2003, signal_996}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_314 ( .s (signal_350), .b ({OUT_ciphertext_s1[12], OUT_ciphertext_s0[12]}), .a ({signal_1978, signal_1059}), .c ({signal_2004, signal_995}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_315 ( .s (signal_350), .b ({OUT_ciphertext_s1[13], OUT_ciphertext_s0[13]}), .a ({signal_1976, signal_1058}), .c ({signal_2005, signal_994}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_316 ( .s (signal_350), .b ({OUT_ciphertext_s1[14], OUT_ciphertext_s0[14]}), .a ({signal_1974, signal_1057}), .c ({signal_2006, signal_993}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_317 ( .s (signal_350), .b ({OUT_ciphertext_s1[15], OUT_ciphertext_s0[15]}), .a ({signal_1972, signal_1056}), .c ({signal_2007, signal_992}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_318 ( .s (signal_311), .b ({OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}), .a ({signal_1718, signal_1055}), .c ({signal_1876, signal_319}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_319 ( .s (signal_311), .b ({OUT_ciphertext_s1[17], OUT_ciphertext_s0[17]}), .a ({signal_1970, signal_1054}), .c ({signal_2008, signal_320}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_320 ( .s (signal_311), .b ({OUT_ciphertext_s1[18], OUT_ciphertext_s0[18]}), .a ({signal_1968, signal_1053}), .c ({signal_2009, signal_321}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_321 ( .s (signal_311), .b ({OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}), .a ({signal_1716, signal_1052}), .c ({signal_1877, signal_322}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_322 ( .s (signal_350), .b ({OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}), .a ({signal_1964, signal_1051}), .c ({signal_2010, signal_323}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_323 ( .s (signal_311), .b ({OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}), .a ({signal_1962, signal_1050}), .c ({signal_2011, signal_324}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_324 ( .s (signal_311), .b ({OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}), .a ({signal_1714, signal_1049}), .c ({signal_1878, signal_325}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_325 ( .s (signal_311), .b ({OUT_ciphertext_s1[23], OUT_ciphertext_s0[23]}), .a ({signal_1960, signal_1048}), .c ({signal_2012, signal_984}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_326 ( .s (signal_311), .b ({OUT_ciphertext_s1[24], OUT_ciphertext_s0[24]}), .a ({signal_1712, signal_1047}), .c ({signal_1879, signal_983}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_327 ( .s (signal_311), .b ({OUT_ciphertext_s1[25], OUT_ciphertext_s0[25]}), .a ({signal_1958, signal_1046}), .c ({signal_2013, signal_982}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_328 ( .s (signal_311), .b ({OUT_ciphertext_s1[26], OUT_ciphertext_s0[26]}), .a ({signal_1710, signal_1045}), .c ({signal_1880, signal_981}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_329 ( .s (signal_311), .b ({OUT_ciphertext_s1[27], OUT_ciphertext_s0[27]}), .a ({signal_1956, signal_1044}), .c ({signal_2014, signal_980}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_330 ( .s (signal_351), .b ({OUT_ciphertext_s1[28], OUT_ciphertext_s0[28]}), .a ({signal_1708, signal_1043}), .c ({signal_1983, signal_979}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_331 ( .s (signal_351), .b ({OUT_ciphertext_s1[29], OUT_ciphertext_s0[29]}), .a ({signal_1954, signal_1042}), .c ({signal_2015, signal_978}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_332 ( .s (signal_351), .b ({OUT_ciphertext_s1[30], OUT_ciphertext_s0[30]}), .a ({signal_1950, signal_1041}), .c ({signal_2016, signal_977}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_333 ( .s (signal_351), .b ({OUT_ciphertext_s1[31], OUT_ciphertext_s0[31]}), .a ({signal_1948, signal_1040}), .c ({signal_2017, signal_976}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_334 ( .s (signal_351), .b ({OUT_ciphertext_s1[32], OUT_ciphertext_s0[32]}), .a ({signal_1706, signal_1039}), .c ({signal_1984, signal_326}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_335 ( .s (signal_351), .b ({OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}), .a ({signal_1946, signal_1038}), .c ({signal_2018, signal_327}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_336 ( .s (signal_351), .b ({OUT_ciphertext_s1[34], OUT_ciphertext_s0[34]}), .a ({signal_1704, signal_1037}), .c ({signal_1985, signal_328}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_337 ( .s (signal_351), .b ({OUT_ciphertext_s1[35], OUT_ciphertext_s0[35]}), .a ({signal_1702, signal_1036}), .c ({signal_1986, signal_329}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_338 ( .s (signal_351), .b ({OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}), .a ({signal_1700, signal_1035}), .c ({signal_1987, signal_330}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_339 ( .s (signal_311), .b ({OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}), .a ({signal_1944, signal_1034}), .c ({signal_2019, signal_331}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_340 ( .s (signal_351), .b ({OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}), .a ({signal_1942, signal_1033}), .c ({signal_2020, signal_332}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_341 ( .s (signal_351), .b ({OUT_ciphertext_s1[39], OUT_ciphertext_s0[39]}), .a ({signal_1698, signal_1032}), .c ({signal_1988, signal_968}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_342 ( .s (signal_351), .b ({OUT_ciphertext_s1[40], OUT_ciphertext_s0[40]}), .a ({signal_1940, signal_1031}), .c ({signal_2021, signal_967}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_343 ( .s (signal_351), .b ({OUT_ciphertext_s1[41], OUT_ciphertext_s0[41]}), .a ({signal_1938, signal_1030}), .c ({signal_2022, signal_966}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_344 ( .s (signal_351), .b ({OUT_ciphertext_s1[42], OUT_ciphertext_s0[42]}), .a ({signal_1936, signal_1029}), .c ({signal_2023, signal_965}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_345 ( .s (signal_351), .b ({OUT_ciphertext_s1[43], OUT_ciphertext_s0[43]}), .a ({signal_1934, signal_1028}), .c ({signal_2024, signal_964}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_346 ( .s (signal_351), .b ({OUT_ciphertext_s1[44], OUT_ciphertext_s0[44]}), .a ({signal_1932, signal_1027}), .c ({signal_2025, signal_963}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_347 ( .s (signal_351), .b ({OUT_ciphertext_s1[45], OUT_ciphertext_s0[45]}), .a ({signal_1930, signal_1026}), .c ({signal_2026, signal_962}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_348 ( .s (signal_351), .b ({OUT_ciphertext_s1[46], OUT_ciphertext_s0[46]}), .a ({signal_1928, signal_1025}), .c ({signal_2027, signal_961}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_349 ( .s (signal_351), .b ({OUT_ciphertext_s1[47], OUT_ciphertext_s0[47]}), .a ({signal_1926, signal_1024}), .c ({signal_2028, signal_960}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_350 ( .s (signal_351), .b ({OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}), .a ({signal_1924, signal_1023}), .c ({signal_2029, signal_333}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_351 ( .s (signal_351), .b ({OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}), .a ({signal_1922, signal_1022}), .c ({signal_2030, signal_334}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_352 ( .s (signal_311), .b ({OUT_ciphertext_s1[50], OUT_ciphertext_s0[50]}), .a ({signal_1918, signal_1021}), .c ({signal_2031, signal_335}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_353 ( .s (signal_351), .b ({OUT_ciphertext_s1[51], OUT_ciphertext_s0[51]}), .a ({signal_1916, signal_1020}), .c ({signal_2032, signal_336}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_354 ( .s (signal_351), .b ({OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}), .a ({signal_1914, signal_1019}), .c ({signal_2033, signal_337}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_355 ( .s (signal_351), .b ({OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}), .a ({signal_1912, signal_1018}), .c ({signal_2034, signal_338}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_356 ( .s (signal_351), .b ({OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}), .a ({signal_1910, signal_1017}), .c ({signal_2035, signal_339}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_357 ( .s (signal_351), .b ({OUT_ciphertext_s1[55], OUT_ciphertext_s0[55]}), .a ({signal_1908, signal_1016}), .c ({signal_2036, signal_952}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_358 ( .s (signal_351), .b ({OUT_ciphertext_s1[56], OUT_ciphertext_s0[56]}), .a ({signal_1906, signal_1015}), .c ({signal_2037, signal_951}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_359 ( .s (signal_351), .b ({OUT_ciphertext_s1[57], OUT_ciphertext_s0[57]}), .a ({signal_1904, signal_1014}), .c ({signal_2038, signal_950}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_360 ( .s (signal_351), .b ({OUT_ciphertext_s1[58], OUT_ciphertext_s0[58]}), .a ({signal_1902, signal_1013}), .c ({signal_2039, signal_949}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_361 ( .s (signal_351), .b ({OUT_ciphertext_s1[59], OUT_ciphertext_s0[59]}), .a ({signal_1900, signal_1012}), .c ({signal_2040, signal_948}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_362 ( .s (signal_351), .b ({OUT_ciphertext_s1[60], OUT_ciphertext_s0[60]}), .a ({signal_1896, signal_1011}), .c ({signal_2041, signal_947}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_363 ( .s (signal_351), .b ({OUT_ciphertext_s1[61], OUT_ciphertext_s0[61]}), .a ({signal_1894, signal_1010}), .c ({signal_2042, signal_946}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_364 ( .s (signal_351), .b ({OUT_ciphertext_s1[62], OUT_ciphertext_s0[62]}), .a ({signal_1892, signal_1009}), .c ({signal_2043, signal_945}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_365 ( .s (signal_351), .b ({OUT_ciphertext_s1[63], OUT_ciphertext_s0[63]}), .a ({signal_1890, signal_1008}), .c ({signal_2044, signal_944}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_366 ( .a ({1'b0, signal_874}), .b ({signal_1998, signal_318}), .c ({signal_2054, signal_1001}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_367 ( .a ({1'b0, signal_875}), .b ({signal_1997, signal_317}), .c ({signal_2055, signal_1002}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_368 ( .a ({1'b0, signal_877}), .b ({signal_2035, signal_339}), .c ({signal_2056, signal_953}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_369 ( .a ({1'b0, signal_878}), .b ({signal_2034, signal_338}), .c ({signal_2057, signal_954}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_370 ( .a ({1'b0, signal_879}), .b ({signal_2033, signal_337}), .c ({signal_2058, signal_955}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_371 ( .a ({1'b0, 1'b0}), .b ({signal_2032, signal_336}), .c ({signal_2059, signal_956}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_372 ( .a ({1'b0, 1'b0}), .b ({signal_2031, signal_335}), .c ({signal_2060, signal_957}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_373 ( .a ({1'b0, signal_876}), .b ({signal_1996, signal_316}), .c ({signal_2061, signal_1003}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_374 ( .a ({1'b0, 1'b0}), .b ({signal_2030, signal_334}), .c ({signal_2062, signal_958}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_375 ( .a ({1'b0, 1'b0}), .b ({signal_2029, signal_333}), .c ({signal_2063, signal_959}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_376 ( .a ({1'b0, 1'b1}), .b ({signal_1875, signal_315}), .c ({signal_1989, signal_1004}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_377 ( .a ({1'b0, signal_874}), .b ({signal_2020, signal_332}), .c ({signal_2064, signal_969}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_378 ( .a ({1'b0, signal_875}), .b ({signal_2019, signal_331}), .c ({signal_2065, signal_970}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_379 ( .a ({1'b0, signal_876}), .b ({signal_1987, signal_330}), .c ({signal_2045, signal_971}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_380 ( .a ({1'b0, 1'b0}), .b ({signal_1986, signal_329}), .c ({signal_2046, signal_972}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_381 ( .a ({1'b0, 1'b0}), .b ({signal_1985, signal_328}), .c ({signal_2047, signal_973}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_382 ( .a ({1'b0, 1'b0}), .b ({signal_2018, signal_327}), .c ({signal_2066, signal_974}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_383 ( .a ({1'b0, 1'b0}), .b ({signal_1984, signal_326}), .c ({signal_2048, signal_975}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_384 ( .a ({1'b0, 1'b0}), .b ({signal_1995, signal_314}), .c ({signal_2067, signal_1005}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_385 ( .a ({1'b0, signal_877}), .b ({signal_1878, signal_325}), .c ({signal_1990, signal_985}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_386 ( .a ({1'b0, signal_878}), .b ({signal_2011, signal_324}), .c ({signal_2068, signal_986}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_387 ( .a ({1'b0, signal_879}), .b ({signal_2010, signal_323}), .c ({signal_2069, signal_987}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_388 ( .a ({1'b0, 1'b0}), .b ({signal_1994, signal_313}), .c ({signal_2070, signal_1006}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_389 ( .a ({1'b0, 1'b1}), .b ({signal_1877, signal_322}), .c ({signal_1991, signal_988}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_390 ( .a ({1'b0, 1'b0}), .b ({signal_2009, signal_321}), .c ({signal_2071, signal_989}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_391 ( .a ({1'b0, 1'b0}), .b ({signal_2008, signal_320}), .c ({signal_2072, signal_990}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_392 ( .a ({1'b0, 1'b0}), .b ({signal_1876, signal_319}), .c ({signal_1992, signal_991}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_393 ( .a ({1'b0, 1'b0}), .b ({signal_1874, signal_312}), .c ({signal_1993, signal_1007}) ) ;
    INV_X1 cell_978 ( .A (signal_808), .ZN (signal_309) ) ;
    INV_X1 cell_980 ( .A (signal_307), .ZN (signal_306) ) ;
    INV_X1 cell_982 ( .A (signal_304), .ZN (signal_289) ) ;
    INV_X1 cell_984 ( .A (signal_288), .ZN (signal_302) ) ;
    INV_X1 cell_986 ( .A (signal_879), .ZN (signal_300) ) ;
    INV_X1 cell_988 ( .A (signal_878), .ZN (signal_298) ) ;
    INV_X1 cell_990 ( .A (signal_877), .ZN (signal_296) ) ;
    INV_X1 cell_992 ( .A (signal_876), .ZN (signal_294) ) ;
    INV_X1 cell_994 ( .A (signal_875), .ZN (signal_292) ) ;
    INV_X1 cell_996 ( .A (signal_874), .ZN (signal_290) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1128 ( .a ({signal_1988, signal_968}), .b ({signal_2049, signal_1328}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1129 ( .a ({signal_1989, signal_1004}), .b ({signal_2050, signal_1329}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1130 ( .a ({signal_1991, signal_988}), .b ({signal_2051, signal_1330}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1131 ( .a ({signal_1999, signal_1000}), .b ({signal_2073, signal_1331}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1132 ( .a ({signal_2001, signal_998}), .b ({signal_2074, signal_1332}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1133 ( .a ({signal_2003, signal_996}), .b ({signal_2075, signal_1333}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1134 ( .a ({signal_2005, signal_994}), .b ({signal_2076, signal_1334}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1135 ( .a ({signal_2007, signal_992}), .b ({signal_2077, signal_1335}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1136 ( .a ({signal_2012, signal_984}), .b ({signal_2078, signal_1336}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1137 ( .a ({signal_2013, signal_982}), .b ({signal_2079, signal_1337}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1138 ( .a ({signal_2014, signal_980}), .b ({signal_2080, signal_1338}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1139 ( .a ({signal_2015, signal_978}), .b ({signal_2081, signal_1339}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1140 ( .a ({signal_2017, signal_976}), .b ({signal_2082, signal_1340}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1141 ( .a ({signal_2022, signal_966}), .b ({signal_2083, signal_1341}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1142 ( .a ({signal_2024, signal_964}), .b ({signal_2084, signal_1342}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1143 ( .a ({signal_2026, signal_962}), .b ({signal_2085, signal_1343}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1144 ( .a ({signal_2028, signal_960}), .b ({signal_2086, signal_1344}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1145 ( .a ({signal_2036, signal_952}), .b ({signal_2087, signal_1345}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1146 ( .a ({signal_2038, signal_950}), .b ({signal_2088, signal_1346}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1147 ( .a ({signal_2040, signal_948}), .b ({signal_2089, signal_1347}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1148 ( .a ({signal_2042, signal_946}), .b ({signal_2090, signal_1348}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1149 ( .a ({signal_2044, signal_944}), .b ({signal_2091, signal_1349}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1150 ( .a ({signal_2046, signal_972}), .b ({signal_2092, signal_1350}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1151 ( .a ({signal_2055, signal_1002}), .b ({signal_2127, signal_1351}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1152 ( .a ({signal_2057, signal_954}), .b ({signal_2128, signal_1352}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1153 ( .a ({signal_2059, signal_956}), .b ({signal_2129, signal_1353}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1154 ( .a ({signal_2062, signal_958}), .b ({signal_2130, signal_1354}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1155 ( .a ({signal_2065, signal_970}), .b ({signal_2131, signal_1355}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1156 ( .a ({signal_2066, signal_974}), .b ({signal_2132, signal_1356}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1157 ( .a ({signal_2068, signal_986}), .b ({signal_2133, signal_1357}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1158 ( .a ({signal_2070, signal_1006}), .b ({signal_2134, signal_1358}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1159 ( .a ({signal_2072, signal_990}), .b ({signal_2135, signal_1359}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1160 ( .a ({signal_2067, signal_1005}), .b ({signal_2070, signal_1006}), .c ({signal_2136, signal_1360}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1161 ( .a ({signal_1993, signal_1007}), .b ({signal_2070, signal_1006}), .c ({signal_2137, signal_1361}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1162 ( .a ({signal_1989, signal_1004}), .b ({signal_1993, signal_1007}), .c ({signal_2052, signal_1362}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1163 ( .a ({signal_1989, signal_1004}), .b ({signal_2070, signal_1006}), .c ({signal_2138, signal_1363}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1164 ( .a ({signal_2054, signal_1001}), .b ({signal_2055, signal_1002}), .c ({signal_2139, signal_1364}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1165 ( .a ({signal_2055, signal_1002}), .b ({signal_2061, signal_1003}), .c ({signal_2140, signal_1365}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1166 ( .a ({signal_1999, signal_1000}), .b ({signal_2061, signal_1003}), .c ({signal_2141, signal_1366}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1167 ( .a ({signal_1999, signal_1000}), .b ({signal_2055, signal_1002}), .c ({signal_2142, signal_1367}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1168 ( .a ({signal_2001, signal_998}), .b ({signal_2002, signal_997}), .c ({signal_2093, signal_1368}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1169 ( .a ({signal_2000, signal_999}), .b ({signal_2001, signal_998}), .c ({signal_2094, signal_1369}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1170 ( .a ({signal_2000, signal_999}), .b ({signal_2003, signal_996}), .c ({signal_2095, signal_1370}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1171 ( .a ({signal_2001, signal_998}), .b ({signal_2003, signal_996}), .c ({signal_2096, signal_1371}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1172 ( .a ({signal_2005, signal_994}), .b ({signal_2006, signal_993}), .c ({signal_2097, signal_1372}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1173 ( .a ({signal_2004, signal_995}), .b ({signal_2005, signal_994}), .c ({signal_2098, signal_1373}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1174 ( .a ({signal_2004, signal_995}), .b ({signal_2007, signal_992}), .c ({signal_2099, signal_1374}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1175 ( .a ({signal_2005, signal_994}), .b ({signal_2007, signal_992}), .c ({signal_2100, signal_1375}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1176 ( .a ({signal_2071, signal_989}), .b ({signal_2072, signal_990}), .c ({signal_2143, signal_1376}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1177 ( .a ({signal_1992, signal_991}), .b ({signal_2072, signal_990}), .c ({signal_2144, signal_1377}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1178 ( .a ({signal_1991, signal_988}), .b ({signal_1992, signal_991}), .c ({signal_2053, signal_1378}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1179 ( .a ({signal_1991, signal_988}), .b ({signal_2072, signal_990}), .c ({signal_2145, signal_1379}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1180 ( .a ({signal_1990, signal_985}), .b ({signal_2068, signal_986}), .c ({signal_2146, signal_1380}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1181 ( .a ({signal_2068, signal_986}), .b ({signal_2069, signal_987}), .c ({signal_2147, signal_1381}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1182 ( .a ({signal_2012, signal_984}), .b ({signal_2069, signal_987}), .c ({signal_2148, signal_1382}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1183 ( .a ({signal_2012, signal_984}), .b ({signal_2068, signal_986}), .c ({signal_2149, signal_1383}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1184 ( .a ({signal_1880, signal_981}), .b ({signal_2013, signal_982}), .c ({signal_2101, signal_1384}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1185 ( .a ({signal_1879, signal_983}), .b ({signal_2013, signal_982}), .c ({signal_2102, signal_1385}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1186 ( .a ({signal_1879, signal_983}), .b ({signal_2014, signal_980}), .c ({signal_2103, signal_1386}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1187 ( .a ({signal_2013, signal_982}), .b ({signal_2014, signal_980}), .c ({signal_2104, signal_1387}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1188 ( .a ({signal_2015, signal_978}), .b ({signal_2016, signal_977}), .c ({signal_2105, signal_1388}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1189 ( .a ({signal_1983, signal_979}), .b ({signal_2015, signal_978}), .c ({signal_2106, signal_1389}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1190 ( .a ({signal_1983, signal_979}), .b ({signal_2017, signal_976}), .c ({signal_2107, signal_1390}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1191 ( .a ({signal_2015, signal_978}), .b ({signal_2017, signal_976}), .c ({signal_2108, signal_1391}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1192 ( .a ({signal_2047, signal_973}), .b ({signal_2066, signal_974}), .c ({signal_2150, signal_1392}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1193 ( .a ({signal_2048, signal_975}), .b ({signal_2066, signal_974}), .c ({signal_2151, signal_1393}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1194 ( .a ({signal_2046, signal_972}), .b ({signal_2048, signal_975}), .c ({signal_2109, signal_1394}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1195 ( .a ({signal_2046, signal_972}), .b ({signal_2066, signal_974}), .c ({signal_2152, signal_1395}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1196 ( .a ({signal_2064, signal_969}), .b ({signal_2065, signal_970}), .c ({signal_2153, signal_1396}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1197 ( .a ({signal_2045, signal_971}), .b ({signal_2065, signal_970}), .c ({signal_2154, signal_1397}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1198 ( .a ({signal_1988, signal_968}), .b ({signal_2045, signal_971}), .c ({signal_2110, signal_1398}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1199 ( .a ({signal_1988, signal_968}), .b ({signal_2065, signal_970}), .c ({signal_2155, signal_1399}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1200 ( .a ({signal_2022, signal_966}), .b ({signal_2023, signal_965}), .c ({signal_2111, signal_1400}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1201 ( .a ({signal_2021, signal_967}), .b ({signal_2022, signal_966}), .c ({signal_2112, signal_1401}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1202 ( .a ({signal_2021, signal_967}), .b ({signal_2024, signal_964}), .c ({signal_2113, signal_1402}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1203 ( .a ({signal_2022, signal_966}), .b ({signal_2024, signal_964}), .c ({signal_2114, signal_1403}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1204 ( .a ({signal_2026, signal_962}), .b ({signal_2027, signal_961}), .c ({signal_2115, signal_1404}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1205 ( .a ({signal_2025, signal_963}), .b ({signal_2026, signal_962}), .c ({signal_2116, signal_1405}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1206 ( .a ({signal_2025, signal_963}), .b ({signal_2028, signal_960}), .c ({signal_2117, signal_1406}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1207 ( .a ({signal_2026, signal_962}), .b ({signal_2028, signal_960}), .c ({signal_2118, signal_1407}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1208 ( .a ({signal_2060, signal_957}), .b ({signal_2062, signal_958}), .c ({signal_2156, signal_1408}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1209 ( .a ({signal_2062, signal_958}), .b ({signal_2063, signal_959}), .c ({signal_2157, signal_1409}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1210 ( .a ({signal_2059, signal_956}), .b ({signal_2063, signal_959}), .c ({signal_2158, signal_1410}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1211 ( .a ({signal_2059, signal_956}), .b ({signal_2062, signal_958}), .c ({signal_2159, signal_1411}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1212 ( .a ({signal_2056, signal_953}), .b ({signal_2057, signal_954}), .c ({signal_2160, signal_1412}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1213 ( .a ({signal_2057, signal_954}), .b ({signal_2058, signal_955}), .c ({signal_2161, signal_1413}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1214 ( .a ({signal_2036, signal_952}), .b ({signal_2058, signal_955}), .c ({signal_2162, signal_1414}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1215 ( .a ({signal_2036, signal_952}), .b ({signal_2057, signal_954}), .c ({signal_2163, signal_1415}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1216 ( .a ({signal_2038, signal_950}), .b ({signal_2039, signal_949}), .c ({signal_2119, signal_1416}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1217 ( .a ({signal_2037, signal_951}), .b ({signal_2038, signal_950}), .c ({signal_2120, signal_1417}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1218 ( .a ({signal_2037, signal_951}), .b ({signal_2040, signal_948}), .c ({signal_2121, signal_1418}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1219 ( .a ({signal_2038, signal_950}), .b ({signal_2040, signal_948}), .c ({signal_2122, signal_1419}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1220 ( .a ({signal_2042, signal_946}), .b ({signal_2043, signal_945}), .c ({signal_2123, signal_1420}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1221 ( .a ({signal_2041, signal_947}), .b ({signal_2042, signal_946}), .c ({signal_2124, signal_1421}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1222 ( .a ({signal_2041, signal_947}), .b ({signal_2044, signal_944}), .c ({signal_2125, signal_1422}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1223 ( .a ({signal_2042, signal_946}), .b ({signal_2044, signal_944}), .c ({signal_2126, signal_1423}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1224 ( .a ({signal_2136, signal_1360}), .b ({signal_2204, signal_1424}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1225 ( .a ({signal_2139, signal_1364}), .b ({signal_2205, signal_1425}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1226 ( .a ({signal_2093, signal_1368}), .b ({signal_2164, signal_1426}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1227 ( .a ({signal_2097, signal_1372}), .b ({signal_2165, signal_1427}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1228 ( .a ({signal_2143, signal_1376}), .b ({signal_2206, signal_1428}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1229 ( .a ({signal_2146, signal_1380}), .b ({signal_2207, signal_1429}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1230 ( .a ({signal_2101, signal_1384}), .b ({signal_2166, signal_1430}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1231 ( .a ({signal_2105, signal_1388}), .b ({signal_2167, signal_1431}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1232 ( .a ({signal_2150, signal_1392}), .b ({signal_2208, signal_1432}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1233 ( .a ({signal_2153, signal_1396}), .b ({signal_2209, signal_1433}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1234 ( .a ({signal_2111, signal_1400}), .b ({signal_2168, signal_1434}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1235 ( .a ({signal_2115, signal_1404}), .b ({signal_2169, signal_1435}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1236 ( .a ({signal_2156, signal_1408}), .b ({signal_2210, signal_1436}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1237 ( .a ({signal_2160, signal_1412}), .b ({signal_2211, signal_1437}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1238 ( .a ({signal_2119, signal_1416}), .b ({signal_2170, signal_1438}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1239 ( .a ({signal_2123, signal_1420}), .b ({signal_2171, signal_1439}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1256 ( .a ({signal_1989, signal_1004}), .b ({signal_2137, signal_1361}), .c ({signal_2220, signal_1456}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1257 ( .a ({signal_2136, signal_1360}), .b ({signal_2052, signal_1362}), .c ({signal_2221, signal_1457}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1258 ( .a ({signal_2067, signal_1005}), .b ({signal_2137, signal_1361}), .c ({signal_2222, signal_1458}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1259 ( .a ({signal_1999, signal_1000}), .b ({signal_2140, signal_1365}), .c ({signal_2223, signal_1459}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1260 ( .a ({signal_2139, signal_1364}), .b ({signal_2141, signal_1366}), .c ({signal_2224, signal_1460}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1261 ( .a ({signal_2054, signal_1001}), .b ({signal_2140, signal_1365}), .c ({signal_2225, signal_1461}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1262 ( .a ({signal_2003, signal_996}), .b ({signal_2094, signal_1369}), .c ({signal_2180, signal_1462}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1263 ( .a ({signal_2093, signal_1368}), .b ({signal_2095, signal_1370}), .c ({signal_2181, signal_1463}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1264 ( .a ({signal_2002, signal_997}), .b ({signal_2094, signal_1369}), .c ({signal_2182, signal_1464}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1265 ( .a ({signal_2007, signal_992}), .b ({signal_2098, signal_1373}), .c ({signal_2183, signal_1465}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1266 ( .a ({signal_2097, signal_1372}), .b ({signal_2099, signal_1374}), .c ({signal_2184, signal_1466}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1267 ( .a ({signal_2006, signal_993}), .b ({signal_2098, signal_1373}), .c ({signal_2185, signal_1467}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1268 ( .a ({signal_1991, signal_988}), .b ({signal_2144, signal_1377}), .c ({signal_2226, signal_1468}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1269 ( .a ({signal_2143, signal_1376}), .b ({signal_2053, signal_1378}), .c ({signal_2227, signal_1469}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1270 ( .a ({signal_2071, signal_989}), .b ({signal_2144, signal_1377}), .c ({signal_2228, signal_1470}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1271 ( .a ({signal_2012, signal_984}), .b ({signal_2147, signal_1381}), .c ({signal_2229, signal_1471}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1272 ( .a ({signal_2146, signal_1380}), .b ({signal_2148, signal_1382}), .c ({signal_2230, signal_1472}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1273 ( .a ({signal_1990, signal_985}), .b ({signal_2147, signal_1381}), .c ({signal_2231, signal_1473}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1274 ( .a ({signal_2014, signal_980}), .b ({signal_2102, signal_1385}), .c ({signal_2186, signal_1474}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1275 ( .a ({signal_2101, signal_1384}), .b ({signal_2103, signal_1386}), .c ({signal_2187, signal_1475}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1276 ( .a ({signal_1880, signal_981}), .b ({signal_2102, signal_1385}), .c ({signal_2188, signal_1476}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1277 ( .a ({signal_2017, signal_976}), .b ({signal_2106, signal_1389}), .c ({signal_2189, signal_1477}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1278 ( .a ({signal_2105, signal_1388}), .b ({signal_2107, signal_1390}), .c ({signal_2190, signal_1478}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1279 ( .a ({signal_2016, signal_977}), .b ({signal_2106, signal_1389}), .c ({signal_2191, signal_1479}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1280 ( .a ({signal_2046, signal_972}), .b ({signal_2151, signal_1393}), .c ({signal_2232, signal_1480}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1281 ( .a ({signal_2150, signal_1392}), .b ({signal_2109, signal_1394}), .c ({signal_2233, signal_1481}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1282 ( .a ({signal_2047, signal_973}), .b ({signal_2151, signal_1393}), .c ({signal_2234, signal_1482}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1283 ( .a ({signal_1988, signal_968}), .b ({signal_2154, signal_1397}), .c ({signal_2235, signal_1483}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1284 ( .a ({signal_2153, signal_1396}), .b ({signal_2110, signal_1398}), .c ({signal_2236, signal_1484}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1285 ( .a ({signal_2064, signal_969}), .b ({signal_2154, signal_1397}), .c ({signal_2237, signal_1485}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1286 ( .a ({signal_2024, signal_964}), .b ({signal_2112, signal_1401}), .c ({signal_2192, signal_1486}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1287 ( .a ({signal_2111, signal_1400}), .b ({signal_2113, signal_1402}), .c ({signal_2193, signal_1487}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1288 ( .a ({signal_2023, signal_965}), .b ({signal_2112, signal_1401}), .c ({signal_2194, signal_1488}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1289 ( .a ({signal_2028, signal_960}), .b ({signal_2116, signal_1405}), .c ({signal_2195, signal_1489}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1290 ( .a ({signal_2115, signal_1404}), .b ({signal_2117, signal_1406}), .c ({signal_2196, signal_1490}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1291 ( .a ({signal_2027, signal_961}), .b ({signal_2116, signal_1405}), .c ({signal_2197, signal_1491}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1292 ( .a ({signal_2059, signal_956}), .b ({signal_2157, signal_1409}), .c ({signal_2238, signal_1492}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1293 ( .a ({signal_2156, signal_1408}), .b ({signal_2158, signal_1410}), .c ({signal_2239, signal_1493}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1294 ( .a ({signal_2060, signal_957}), .b ({signal_2157, signal_1409}), .c ({signal_2240, signal_1494}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1295 ( .a ({signal_2036, signal_952}), .b ({signal_2161, signal_1413}), .c ({signal_2241, signal_1495}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1296 ( .a ({signal_2160, signal_1412}), .b ({signal_2162, signal_1414}), .c ({signal_2242, signal_1496}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1297 ( .a ({signal_2056, signal_953}), .b ({signal_2161, signal_1413}), .c ({signal_2243, signal_1497}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1298 ( .a ({signal_2040, signal_948}), .b ({signal_2120, signal_1417}), .c ({signal_2198, signal_1498}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1299 ( .a ({signal_2119, signal_1416}), .b ({signal_2121, signal_1418}), .c ({signal_2199, signal_1499}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1300 ( .a ({signal_2039, signal_949}), .b ({signal_2120, signal_1417}), .c ({signal_2200, signal_1500}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1301 ( .a ({signal_2044, signal_944}), .b ({signal_2124, signal_1421}), .c ({signal_2201, signal_1501}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1302 ( .a ({signal_2123, signal_1420}), .b ({signal_2125, signal_1422}), .c ({signal_2202, signal_1502}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1303 ( .a ({signal_2043, signal_945}), .b ({signal_2124, signal_1421}), .c ({signal_2203, signal_1503}) ) ;
    ClockGatingController #(5) cell_1528 ( .clk (CLK), .rst (IN_reset), .GatedClk (signal_2940), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1240 ( .a ({signal_2067, signal_1005}), .b ({signal_2134, signal_1358}), .clk (CLK), .r (Fresh[0]), .c ({signal_2212, signal_1440}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1241 ( .a ({signal_2054, signal_1001}), .b ({signal_2127, signal_1351}), .clk (CLK), .r (Fresh[1]), .c ({signal_2213, signal_1441}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1242 ( .a ({signal_2074, signal_1332}), .b ({signal_2002, signal_997}), .clk (CLK), .r (Fresh[2]), .c ({signal_2172, signal_1442}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1243 ( .a ({signal_2076, signal_1334}), .b ({signal_2006, signal_993}), .clk (CLK), .r (Fresh[3]), .c ({signal_2173, signal_1443}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1244 ( .a ({signal_2071, signal_989}), .b ({signal_2135, signal_1359}), .clk (CLK), .r (Fresh[4]), .c ({signal_2214, signal_1444}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1245 ( .a ({signal_1990, signal_985}), .b ({signal_2133, signal_1357}), .clk (CLK), .r (Fresh[5]), .c ({signal_2215, signal_1445}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1246 ( .a ({signal_1880, signal_981}), .b ({signal_2079, signal_1337}), .clk (CLK), .r (Fresh[6]), .c ({signal_2174, signal_1446}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1247 ( .a ({signal_2081, signal_1339}), .b ({signal_2016, signal_977}), .clk (CLK), .r (Fresh[7]), .c ({signal_2175, signal_1447}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1248 ( .a ({signal_2047, signal_973}), .b ({signal_2132, signal_1356}), .clk (CLK), .r (Fresh[8]), .c ({signal_2216, signal_1448}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1249 ( .a ({signal_2064, signal_969}), .b ({signal_2131, signal_1355}), .clk (CLK), .r (Fresh[9]), .c ({signal_2217, signal_1449}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1250 ( .a ({signal_2083, signal_1341}), .b ({signal_2023, signal_965}), .clk (CLK), .r (Fresh[10]), .c ({signal_2176, signal_1450}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1251 ( .a ({signal_2085, signal_1343}), .b ({signal_2027, signal_961}), .clk (CLK), .r (Fresh[11]), .c ({signal_2177, signal_1451}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1252 ( .a ({signal_2060, signal_957}), .b ({signal_2130, signal_1354}), .clk (CLK), .r (Fresh[12]), .c ({signal_2218, signal_1452}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1253 ( .a ({signal_2056, signal_953}), .b ({signal_2128, signal_1352}), .clk (CLK), .r (Fresh[13]), .c ({signal_2219, signal_1453}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1254 ( .a ({signal_2088, signal_1346}), .b ({signal_2039, signal_949}), .clk (CLK), .r (Fresh[14]), .c ({signal_2178, signal_1454}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1255 ( .a ({signal_2090, signal_1348}), .b ({signal_2043, signal_945}), .clk (CLK), .r (Fresh[15]), .c ({signal_2179, signal_1455}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1304 ( .a ({signal_2050, signal_1329}), .b ({signal_2204, signal_1424}), .clk (CLK), .r (Fresh[16]), .c ({signal_2260, signal_1504}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1305 ( .a ({signal_2073, signal_1331}), .b ({signal_2205, signal_1425}), .clk (CLK), .r (Fresh[17]), .c ({signal_2261, signal_1505}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1306 ( .a ({signal_2075, signal_1333}), .b ({signal_2164, signal_1426}), .clk (CLK), .r (Fresh[18]), .c ({signal_2244, signal_1506}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1307 ( .a ({signal_2077, signal_1335}), .b ({signal_2165, signal_1427}), .clk (CLK), .r (Fresh[19]), .c ({signal_2245, signal_1507}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1308 ( .a ({signal_2051, signal_1330}), .b ({signal_2206, signal_1428}), .clk (CLK), .r (Fresh[20]), .c ({signal_2262, signal_1508}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1309 ( .a ({signal_2078, signal_1336}), .b ({signal_2207, signal_1429}), .clk (CLK), .r (Fresh[21]), .c ({signal_2263, signal_1509}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1310 ( .a ({signal_2080, signal_1338}), .b ({signal_2166, signal_1430}), .clk (CLK), .r (Fresh[22]), .c ({signal_2246, signal_1510}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1311 ( .a ({signal_2082, signal_1340}), .b ({signal_2167, signal_1431}), .clk (CLK), .r (Fresh[23]), .c ({signal_2247, signal_1511}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1312 ( .a ({signal_2092, signal_1350}), .b ({signal_2208, signal_1432}), .clk (CLK), .r (Fresh[24]), .c ({signal_2264, signal_1512}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1313 ( .a ({signal_2049, signal_1328}), .b ({signal_2209, signal_1433}), .clk (CLK), .r (Fresh[25]), .c ({signal_2265, signal_1513}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1314 ( .a ({signal_2084, signal_1342}), .b ({signal_2168, signal_1434}), .clk (CLK), .r (Fresh[26]), .c ({signal_2248, signal_1514}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1315 ( .a ({signal_2086, signal_1344}), .b ({signal_2169, signal_1435}), .clk (CLK), .r (Fresh[27]), .c ({signal_2249, signal_1515}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1316 ( .a ({signal_2129, signal_1353}), .b ({signal_2210, signal_1436}), .clk (CLK), .r (Fresh[28]), .c ({signal_2266, signal_1516}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1317 ( .a ({signal_2087, signal_1345}), .b ({signal_2211, signal_1437}), .clk (CLK), .r (Fresh[29]), .c ({signal_2267, signal_1517}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1318 ( .a ({signal_2089, signal_1347}), .b ({signal_2170, signal_1438}), .clk (CLK), .r (Fresh[30]), .c ({signal_2250, signal_1518}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1319 ( .a ({signal_2091, signal_1349}), .b ({signal_2171, signal_1439}), .clk (CLK), .r (Fresh[31]), .c ({signal_2251, signal_1519}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1320 ( .a ({signal_2052, signal_1362}), .b ({signal_2212, signal_1440}), .c ({signal_2268, signal_1520}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1321 ( .a ({signal_2141, signal_1366}), .b ({signal_2213, signal_1441}), .c ({signal_2269, signal_1521}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1322 ( .a ({signal_2095, signal_1370}), .b ({signal_2172, signal_1442}), .c ({signal_2252, signal_1522}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1323 ( .a ({signal_2099, signal_1374}), .b ({signal_2173, signal_1443}), .c ({signal_2253, signal_1523}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1324 ( .a ({signal_2053, signal_1378}), .b ({signal_2214, signal_1444}), .c ({signal_2270, signal_927}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1325 ( .a ({signal_2148, signal_1382}), .b ({signal_2215, signal_1445}), .c ({signal_2271, signal_923}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1326 ( .a ({signal_2103, signal_1386}), .b ({signal_2174, signal_1446}), .c ({signal_2254, signal_919}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1327 ( .a ({signal_2107, signal_1390}), .b ({signal_2175, signal_1447}), .c ({signal_2255, signal_915}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1328 ( .a ({signal_2109, signal_1394}), .b ({signal_2216, signal_1448}), .c ({signal_2272, signal_911}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1329 ( .a ({signal_2110, signal_1398}), .b ({signal_2217, signal_1449}), .c ({signal_2273, signal_907}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1330 ( .a ({signal_2113, signal_1402}), .b ({signal_2176, signal_1450}), .c ({signal_2256, signal_903}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1331 ( .a ({signal_2117, signal_1406}), .b ({signal_2177, signal_1451}), .c ({signal_2257, signal_899}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1332 ( .a ({signal_2158, signal_1410}), .b ({signal_2218, signal_1452}), .c ({signal_2274, signal_895}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1333 ( .a ({signal_2162, signal_1414}), .b ({signal_2219, signal_1453}), .c ({signal_2275, signal_891}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1334 ( .a ({signal_2121, signal_1418}), .b ({signal_2178, signal_1454}), .c ({signal_2258, signal_887}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1335 ( .a ({signal_2125, signal_1422}), .b ({signal_2179, signal_1455}), .c ({signal_2259, signal_883}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1336 ( .a ({signal_2220, signal_1456}), .b ({signal_2260, signal_1504}), .c ({signal_2292, signal_1524}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1337 ( .a ({signal_2212, signal_1440}), .b ({signal_2260, signal_1504}), .c ({signal_2293, signal_1525}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1338 ( .a ({signal_2223, signal_1459}), .b ({signal_2261, signal_1505}), .c ({signal_2294, signal_1526}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1339 ( .a ({signal_2213, signal_1441}), .b ({signal_2261, signal_1505}), .c ({signal_2295, signal_1527}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1340 ( .a ({signal_2180, signal_1462}), .b ({signal_2244, signal_1506}), .c ({signal_2276, signal_1528}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1341 ( .a ({signal_2172, signal_1442}), .b ({signal_2244, signal_1506}), .c ({signal_2277, signal_1529}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1342 ( .a ({signal_2183, signal_1465}), .b ({signal_2245, signal_1507}), .c ({signal_2278, signal_1530}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1343 ( .a ({signal_2173, signal_1443}), .b ({signal_2245, signal_1507}), .c ({signal_2279, signal_1531}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1344 ( .a ({signal_2226, signal_1468}), .b ({signal_2262, signal_1508}), .c ({signal_2296, signal_1532}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1345 ( .a ({signal_2214, signal_1444}), .b ({signal_2262, signal_1508}), .c ({signal_2297, signal_1533}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1346 ( .a ({signal_2229, signal_1471}), .b ({signal_2263, signal_1509}), .c ({signal_2298, signal_1534}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1347 ( .a ({signal_2215, signal_1445}), .b ({signal_2263, signal_1509}), .c ({signal_2299, signal_1535}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1348 ( .a ({signal_2186, signal_1474}), .b ({signal_2246, signal_1510}), .c ({signal_2280, signal_1536}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1349 ( .a ({signal_2174, signal_1446}), .b ({signal_2246, signal_1510}), .c ({signal_2281, signal_1537}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1350 ( .a ({signal_2189, signal_1477}), .b ({signal_2247, signal_1511}), .c ({signal_2282, signal_1538}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1351 ( .a ({signal_2175, signal_1447}), .b ({signal_2247, signal_1511}), .c ({signal_2283, signal_1539}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1352 ( .a ({signal_2232, signal_1480}), .b ({signal_2264, signal_1512}), .c ({signal_2300, signal_1540}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1353 ( .a ({signal_2216, signal_1448}), .b ({signal_2264, signal_1512}), .c ({signal_2301, signal_1541}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1354 ( .a ({signal_2235, signal_1483}), .b ({signal_2265, signal_1513}), .c ({signal_2302, signal_1542}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1355 ( .a ({signal_2217, signal_1449}), .b ({signal_2265, signal_1513}), .c ({signal_2303, signal_1543}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1356 ( .a ({signal_2192, signal_1486}), .b ({signal_2248, signal_1514}), .c ({signal_2284, signal_1544}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1357 ( .a ({signal_2176, signal_1450}), .b ({signal_2248, signal_1514}), .c ({signal_2285, signal_1545}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1358 ( .a ({signal_2195, signal_1489}), .b ({signal_2249, signal_1515}), .c ({signal_2286, signal_1546}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1359 ( .a ({signal_2177, signal_1451}), .b ({signal_2249, signal_1515}), .c ({signal_2287, signal_1547}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1360 ( .a ({signal_2238, signal_1492}), .b ({signal_2266, signal_1516}), .c ({signal_2304, signal_1548}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1361 ( .a ({signal_2218, signal_1452}), .b ({signal_2266, signal_1516}), .c ({signal_2305, signal_1549}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1362 ( .a ({signal_2241, signal_1495}), .b ({signal_2267, signal_1517}), .c ({signal_2306, signal_1550}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1363 ( .a ({signal_2219, signal_1453}), .b ({signal_2267, signal_1517}), .c ({signal_2307, signal_1551}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1364 ( .a ({signal_2198, signal_1498}), .b ({signal_2250, signal_1518}), .c ({signal_2288, signal_1552}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1365 ( .a ({signal_2178, signal_1454}), .b ({signal_2250, signal_1518}), .c ({signal_2289, signal_1553}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1366 ( .a ({signal_2201, signal_1501}), .b ({signal_2251, signal_1519}), .c ({signal_2290, signal_1554}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1367 ( .a ({signal_2179, signal_1455}), .b ({signal_2251, signal_1519}), .c ({signal_2291, signal_1555}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1368 ( .a ({signal_2292, signal_1524}), .b ({signal_2324, signal_1556}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1369 ( .a ({signal_2294, signal_1526}), .b ({signal_2325, signal_1557}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1370 ( .a ({signal_2276, signal_1528}), .b ({signal_2308, signal_1558}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1371 ( .a ({signal_2278, signal_1530}), .b ({signal_2309, signal_1559}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1372 ( .a ({signal_2296, signal_1532}), .b ({signal_2326, signal_1560}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1373 ( .a ({signal_2298, signal_1534}), .b ({signal_2327, signal_1561}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1374 ( .a ({signal_2280, signal_1536}), .b ({signal_2310, signal_1562}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1375 ( .a ({signal_2282, signal_1538}), .b ({signal_2311, signal_1563}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1376 ( .a ({signal_2300, signal_1540}), .b ({signal_2328, signal_1564}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1377 ( .a ({signal_2302, signal_1542}), .b ({signal_2329, signal_1565}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1378 ( .a ({signal_2284, signal_1544}), .b ({signal_2312, signal_1566}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1379 ( .a ({signal_2286, signal_1546}), .b ({signal_2313, signal_1567}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1380 ( .a ({signal_2304, signal_1548}), .b ({signal_2330, signal_1568}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1381 ( .a ({signal_2306, signal_1550}), .b ({signal_2331, signal_1569}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1382 ( .a ({signal_2288, signal_1552}), .b ({signal_2314, signal_1570}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1383 ( .a ({signal_2290, signal_1554}), .b ({signal_2315, signal_1571}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1384 ( .a ({signal_2138, signal_1363}), .b ({signal_2293, signal_1525}), .c ({signal_2332, signal_1572}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1385 ( .a ({signal_2142, signal_1367}), .b ({signal_2295, signal_1527}), .c ({signal_2333, signal_1573}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1386 ( .a ({signal_2096, signal_1371}), .b ({signal_2277, signal_1529}), .c ({signal_2316, signal_1574}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1387 ( .a ({signal_2100, signal_1375}), .b ({signal_2279, signal_1531}), .c ({signal_2317, signal_1575}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1388 ( .a ({signal_2145, signal_1379}), .b ({signal_2297, signal_1533}), .c ({signal_2334, signal_1576}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1389 ( .a ({signal_2149, signal_1383}), .b ({signal_2299, signal_1535}), .c ({signal_2335, signal_1577}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1390 ( .a ({signal_2104, signal_1387}), .b ({signal_2281, signal_1537}), .c ({signal_2318, signal_1578}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1391 ( .a ({signal_2108, signal_1391}), .b ({signal_2283, signal_1539}), .c ({signal_2319, signal_1579}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1392 ( .a ({signal_2152, signal_1395}), .b ({signal_2301, signal_1541}), .c ({signal_2336, signal_1580}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1393 ( .a ({signal_2155, signal_1399}), .b ({signal_2303, signal_1543}), .c ({signal_2337, signal_1581}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1394 ( .a ({signal_2114, signal_1403}), .b ({signal_2285, signal_1545}), .c ({signal_2320, signal_1582}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1395 ( .a ({signal_2118, signal_1407}), .b ({signal_2287, signal_1547}), .c ({signal_2321, signal_1583}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1396 ( .a ({signal_2159, signal_1411}), .b ({signal_2305, signal_1549}), .c ({signal_2338, signal_1584}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1397 ( .a ({signal_2163, signal_1415}), .b ({signal_2307, signal_1551}), .c ({signal_2339, signal_1585}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1398 ( .a ({signal_2122, signal_1419}), .b ({signal_2289, signal_1553}), .c ({signal_2322, signal_1586}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1399 ( .a ({signal_2126, signal_1423}), .b ({signal_2291, signal_1555}), .c ({signal_2323, signal_1587}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1400 ( .a ({signal_2332, signal_1572}), .b ({signal_2356, signal_1588}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1401 ( .a ({signal_2333, signal_1573}), .b ({signal_2357, signal_1589}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1402 ( .a ({signal_2316, signal_1574}), .b ({signal_2340, signal_1590}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1403 ( .a ({signal_2317, signal_1575}), .b ({signal_2341, signal_1591}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1404 ( .a ({signal_2334, signal_1576}), .b ({signal_2358, signal_1592}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1405 ( .a ({signal_2335, signal_1577}), .b ({signal_2359, signal_1593}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1406 ( .a ({signal_2318, signal_1578}), .b ({signal_2342, signal_1594}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1407 ( .a ({signal_2319, signal_1579}), .b ({signal_2343, signal_1595}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1408 ( .a ({signal_2336, signal_1580}), .b ({signal_2360, signal_1596}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1409 ( .a ({signal_2337, signal_1581}), .b ({signal_2361, signal_1597}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1410 ( .a ({signal_2320, signal_1582}), .b ({signal_2344, signal_1598}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1411 ( .a ({signal_2321, signal_1583}), .b ({signal_2345, signal_1599}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1412 ( .a ({signal_2338, signal_1584}), .b ({signal_2362, signal_1600}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1413 ( .a ({signal_2339, signal_1585}), .b ({signal_2363, signal_1601}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1414 ( .a ({signal_2322, signal_1586}), .b ({signal_2346, signal_1602}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1415 ( .a ({signal_2323, signal_1587}), .b ({signal_2347, signal_1603}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    mux2_masked #(.security_order(1), .pipeline(0)) cell_39 ( .s (signal_343), .b ({signal_2503, signal_1327}), .a ({signal_1874, signal_312}), .c ({signal_2531, signal_1263}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_40 ( .s (signal_343), .b ({signal_2606, signal_1326}), .a ({signal_1994, signal_313}), .c ({signal_2628, signal_1262}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_41 ( .s (signal_344), .b ({signal_2534, signal_1325}), .a ({signal_1995, signal_314}), .c ({signal_2551, signal_1261}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_42 ( .s (signal_342), .b ({signal_2565, signal_1324}), .a ({signal_1875, signal_315}), .c ({signal_2582, signal_1260}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_43 ( .s (signal_342), .b ({signal_2538, signal_1323}), .a ({signal_1996, signal_316}), .c ({signal_2552, signal_1259}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_44 ( .s (signal_342), .b ({signal_2610, signal_1322}), .a ({signal_1997, signal_317}), .c ({signal_2629, signal_1258}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_45 ( .s (signal_342), .b ({signal_2537, signal_1321}), .a ({signal_1998, signal_318}), .c ({signal_2553, signal_1257}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_46 ( .s (signal_342), .b ({signal_2539, signal_1320}), .a ({signal_1999, signal_1000}), .c ({signal_2554, signal_1256}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_47 ( .s (signal_342), .b ({signal_2543, signal_1319}), .a ({signal_2000, signal_999}), .c ({signal_2555, signal_1255}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_48 ( .s (signal_342), .b ({signal_2575, signal_1318}), .a ({signal_2001, signal_998}), .c ({signal_2583, signal_1254}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_49 ( .s (signal_342), .b ({signal_2542, signal_1317}), .a ({signal_2002, signal_997}), .c ({signal_2556, signal_1253}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_50 ( .s (signal_342), .b ({signal_2544, signal_1316}), .a ({signal_2003, signal_996}), .c ({signal_2557, signal_1252}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_51 ( .s (signal_342), .b ({signal_2549, signal_1315}), .a ({signal_2004, signal_995}), .c ({signal_2558, signal_1251}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_52 ( .s (signal_342), .b ({signal_2579, signal_1314}), .a ({signal_2005, signal_994}), .c ({signal_2584, signal_1250}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_53 ( .s (signal_342), .b ({signal_2548, signal_1313}), .a ({signal_2006, signal_993}), .c ({signal_2559, signal_1249}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_54 ( .s (signal_342), .b ({signal_2581, signal_1312}), .a ({signal_2007, signal_992}), .c ({signal_2585, signal_1248}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_55 ( .s (signal_343), .b ({signal_2648, signal_1311}), .a ({signal_1876, signal_319}), .c ({signal_2670, signal_1247}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_56 ( .s (signal_343), .b ({signal_2700, signal_1310}), .a ({signal_2008, signal_320}), .c ({signal_2715, signal_1246}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_57 ( .s (signal_343), .b ({signal_2697, signal_1309}), .a ({signal_2009, signal_321}), .c ({signal_2716, signal_1245}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_58 ( .s (signal_343), .b ({signal_2608, signal_1308}), .a ({signal_1877, signal_322}), .c ({signal_2630, signal_1244}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_59 ( .s (signal_343), .b ({signal_2612, signal_1307}), .a ({signal_2010, signal_323}), .c ({signal_2631, signal_1243}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_60 ( .s (signal_343), .b ({signal_2657, signal_1306}), .a ({signal_2011, signal_324}), .c ({signal_2671, signal_1242}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_61 ( .s (signal_343), .b ({signal_2702, signal_1305}), .a ({signal_1878, signal_325}), .c ({signal_2717, signal_1241}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_62 ( .s (signal_343), .b ({signal_2613, signal_1304}), .a ({signal_2012, signal_984}), .c ({signal_2632, signal_1240}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_63 ( .s (signal_343), .b ({signal_2618, signal_1303}), .a ({signal_1879, signal_983}), .c ({signal_2633, signal_1239}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_64 ( .s (signal_343), .b ({signal_2664, signal_1302}), .a ({signal_2013, signal_982}), .c ({signal_2672, signal_1238}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_65 ( .s (signal_343), .b ({signal_2661, signal_1301}), .a ({signal_1880, signal_981}), .c ({signal_2673, signal_1237}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_66 ( .s (signal_343), .b ({signal_2619, signal_1300}), .a ({signal_2014, signal_980}), .c ({signal_2634, signal_1236}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_67 ( .s (signal_344), .b ({signal_2668, signal_1299}), .a ({signal_1983, signal_979}), .c ({signal_2674, signal_1235}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_68 ( .s (signal_344), .b ({signal_2714, signal_1298}), .a ({signal_2015, signal_978}), .c ({signal_2718, signal_1234}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_69 ( .s (signal_344), .b ({signal_2666, signal_1297}), .a ({signal_2016, signal_977}), .c ({signal_2675, signal_1233}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_70 ( .s (signal_344), .b ({signal_2626, signal_1296}), .a ({signal_2017, signal_976}), .c ({signal_2635, signal_1232}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_71 ( .s (signal_344), .b ({signal_2696, signal_1295}), .a ({signal_1984, signal_326}), .c ({signal_2719, signal_1231}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_72 ( .s (signal_344), .b ({signal_2745, signal_1294}), .a ({signal_2018, signal_327}), .c ({signal_2755, signal_1230}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_73 ( .s (signal_344), .b ({signal_2694, signal_1293}), .a ({signal_1985, signal_328}), .c ({signal_2720, signal_1229}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_74 ( .s (signal_344), .b ({signal_2788, signal_1292}), .a ({signal_1986, signal_329}), .c ({signal_2795, signal_1228}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_75 ( .s (signal_344), .b ({signal_2701, signal_1291}), .a ({signal_1987, signal_330}), .c ({signal_2721, signal_1227}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_76 ( .s (signal_344), .b ({signal_2703, signal_1290}), .a ({signal_2019, signal_331}), .c ({signal_2722, signal_1226}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_77 ( .s (signal_344), .b ({signal_2650, signal_1289}), .a ({signal_2020, signal_332}), .c ({signal_2676, signal_1225}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_78 ( .s (signal_344), .b ({signal_2790, signal_1288}), .a ({signal_1988, signal_968}), .c ({signal_2796, signal_1224}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_79 ( .s (signal_344), .b ({signal_2705, signal_1287}), .a ({signal_2021, signal_967}), .c ({signal_2723, signal_1223}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_80 ( .s (signal_343), .b ({signal_2707, signal_1286}), .a ({signal_2022, signal_966}), .c ({signal_2724, signal_1222}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_81 ( .s (signal_342), .b ({signal_2658, signal_1285}), .a ({signal_2023, signal_965}), .c ({signal_2677, signal_1221}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_82 ( .s (signal_340), .b ({signal_2751, signal_1284}), .a ({signal_2024, signal_964}), .c ({signal_2756, signal_1220}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_83 ( .s (signal_343), .b ({signal_2710, signal_1283}), .a ({signal_2025, signal_963}), .c ({signal_2725, signal_1219}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_84 ( .s (signal_342), .b ({signal_2754, signal_1282}), .a ({signal_2026, signal_962}), .c ({signal_2757, signal_1218}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_85 ( .s (signal_344), .b ({signal_2708, signal_1281}), .a ({signal_2027, signal_961}), .c ({signal_2726, signal_1217}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_86 ( .s (signal_340), .b ({signal_2753, signal_1280}), .a ({signal_2028, signal_960}), .c ({signal_2758, signal_1216}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_87 ( .s (signal_340), .b ({signal_2847, signal_1279}), .a ({signal_2029, signal_333}), .c ({signal_2852, signal_1215}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_88 ( .s (signal_340), .b ({signal_2860, signal_1278}), .a ({signal_2030, signal_334}), .c ({signal_2862, signal_1214}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_89 ( .s (signal_340), .b ({signal_2787, signal_1277}), .a ({signal_2031, signal_335}), .c ({signal_2797, signal_1213}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_90 ( .s (signal_340), .b ({signal_2786, signal_1276}), .a ({signal_2032, signal_336}), .c ({signal_2798, signal_1212}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_91 ( .s (signal_340), .b ({signal_2849, signal_1275}), .a ({signal_2033, signal_337}), .c ({signal_2853, signal_1211}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_92 ( .s (signal_340), .b ({signal_2861, signal_1274}), .a ({signal_2034, signal_338}), .c ({signal_2863, signal_1210}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_93 ( .s (signal_344), .b ({signal_2747, signal_1273}), .a ({signal_2035, signal_339}), .c ({signal_2759, signal_1209}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_94 ( .s (signal_343), .b ({signal_2789, signal_1272}), .a ({signal_2036, signal_952}), .c ({signal_2799, signal_1208}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_95 ( .s (signal_342), .b ({signal_2841, signal_1271}), .a ({signal_2037, signal_951}), .c ({signal_2844, signal_1207}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_96 ( .s (signal_344), .b ({signal_2850, signal_1270}), .a ({signal_2038, signal_950}), .c ({signal_2854, signal_1206}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_97 ( .s (signal_343), .b ({signal_2750, signal_1269}), .a ({signal_2039, signal_949}), .c ({signal_2760, signal_1205}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_98 ( .s (signal_342), .b ({signal_2749, signal_1268}), .a ({signal_2040, signal_948}), .c ({signal_2761, signal_1204}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_99 ( .s (signal_343), .b ({signal_2843, signal_1267}), .a ({signal_2041, signal_947}), .c ({signal_2845, signal_1203}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_100 ( .s (signal_342), .b ({signal_2851, signal_1266}), .a ({signal_2042, signal_946}), .c ({signal_2855, signal_1202}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_101 ( .s (signal_344), .b ({signal_2793, signal_1265}), .a ({signal_2043, signal_945}), .c ({signal_2800, signal_1201}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_102 ( .s (signal_344), .b ({signal_2792, signal_1264}), .a ({signal_2044, signal_944}), .c ({signal_2801, signal_1200}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_103 ( .s (IN_reset), .b ({signal_2531, signal_1263}), .a ({IN_plaintext_s1[0], IN_plaintext_s0[0]}), .c ({signal_2561, signal_1199}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_104 ( .s (IN_reset), .b ({signal_2628, signal_1262}), .a ({IN_plaintext_s1[1], IN_plaintext_s0[1]}), .c ({signal_2679, signal_1198}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_105 ( .s (IN_reset), .b ({signal_2551, signal_1261}), .a ({IN_plaintext_s1[2], IN_plaintext_s0[2]}), .c ({signal_2587, signal_1197}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_106 ( .s (IN_reset), .b ({signal_2582, signal_1260}), .a ({IN_plaintext_s1[3], IN_plaintext_s0[3]}), .c ({signal_2637, signal_1196}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_107 ( .s (IN_reset), .b ({signal_2552, signal_1259}), .a ({IN_plaintext_s1[4], IN_plaintext_s0[4]}), .c ({signal_2589, signal_1195}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_108 ( .s (IN_reset), .b ({signal_2629, signal_1258}), .a ({IN_plaintext_s1[5], IN_plaintext_s0[5]}), .c ({signal_2681, signal_1194}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_109 ( .s (IN_reset), .b ({signal_2553, signal_1257}), .a ({IN_plaintext_s1[6], IN_plaintext_s0[6]}), .c ({signal_2591, signal_1193}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_110 ( .s (IN_reset), .b ({signal_2554, signal_1256}), .a ({IN_plaintext_s1[7], IN_plaintext_s0[7]}), .c ({signal_2593, signal_1192}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_111 ( .s (IN_reset), .b ({signal_2555, signal_1255}), .a ({IN_plaintext_s1[8], IN_plaintext_s0[8]}), .c ({signal_2595, signal_1191}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_112 ( .s (IN_reset), .b ({signal_2583, signal_1254}), .a ({IN_plaintext_s1[9], IN_plaintext_s0[9]}), .c ({signal_2639, signal_1190}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_113 ( .s (IN_reset), .b ({signal_2556, signal_1253}), .a ({IN_plaintext_s1[10], IN_plaintext_s0[10]}), .c ({signal_2597, signal_1189}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_114 ( .s (IN_reset), .b ({signal_2557, signal_1252}), .a ({IN_plaintext_s1[11], IN_plaintext_s0[11]}), .c ({signal_2599, signal_1188}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_115 ( .s (IN_reset), .b ({signal_2558, signal_1251}), .a ({IN_plaintext_s1[12], IN_plaintext_s0[12]}), .c ({signal_2601, signal_1187}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_116 ( .s (IN_reset), .b ({signal_2584, signal_1250}), .a ({IN_plaintext_s1[13], IN_plaintext_s0[13]}), .c ({signal_2641, signal_1186}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_117 ( .s (IN_reset), .b ({signal_2559, signal_1249}), .a ({IN_plaintext_s1[14], IN_plaintext_s0[14]}), .c ({signal_2603, signal_1185}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_118 ( .s (IN_reset), .b ({signal_2585, signal_1248}), .a ({IN_plaintext_s1[15], IN_plaintext_s0[15]}), .c ({signal_2643, signal_1184}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_119 ( .s (IN_reset), .b ({signal_2670, signal_1247}), .a ({IN_plaintext_s1[16], IN_plaintext_s0[16]}), .c ({signal_2728, signal_1183}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_120 ( .s (IN_reset), .b ({signal_2715, signal_1246}), .a ({IN_plaintext_s1[17], IN_plaintext_s0[17]}), .c ({signal_2763, signal_1182}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_121 ( .s (IN_reset), .b ({signal_2716, signal_1245}), .a ({IN_plaintext_s1[18], IN_plaintext_s0[18]}), .c ({signal_2765, signal_1181}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_122 ( .s (IN_reset), .b ({signal_2630, signal_1244}), .a ({IN_plaintext_s1[19], IN_plaintext_s0[19]}), .c ({signal_2683, signal_1180}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_123 ( .s (IN_reset), .b ({signal_2631, signal_1243}), .a ({IN_plaintext_s1[20], IN_plaintext_s0[20]}), .c ({signal_2685, signal_1179}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_124 ( .s (IN_reset), .b ({signal_2671, signal_1242}), .a ({IN_plaintext_s1[21], IN_plaintext_s0[21]}), .c ({signal_2730, signal_1178}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_125 ( .s (IN_reset), .b ({signal_2717, signal_1241}), .a ({IN_plaintext_s1[22], IN_plaintext_s0[22]}), .c ({signal_2767, signal_1177}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_126 ( .s (IN_reset), .b ({signal_2632, signal_1240}), .a ({IN_plaintext_s1[23], IN_plaintext_s0[23]}), .c ({signal_2687, signal_1176}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_127 ( .s (IN_reset), .b ({signal_2633, signal_1239}), .a ({IN_plaintext_s1[24], IN_plaintext_s0[24]}), .c ({signal_2689, signal_1175}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_128 ( .s (IN_reset), .b ({signal_2672, signal_1238}), .a ({IN_plaintext_s1[25], IN_plaintext_s0[25]}), .c ({signal_2732, signal_1174}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_129 ( .s (IN_reset), .b ({signal_2673, signal_1237}), .a ({IN_plaintext_s1[26], IN_plaintext_s0[26]}), .c ({signal_2734, signal_1173}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_130 ( .s (IN_reset), .b ({signal_2634, signal_1236}), .a ({IN_plaintext_s1[27], IN_plaintext_s0[27]}), .c ({signal_2691, signal_1172}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_131 ( .s (IN_reset), .b ({signal_2674, signal_1235}), .a ({IN_plaintext_s1[28], IN_plaintext_s0[28]}), .c ({signal_2736, signal_1171}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_132 ( .s (IN_reset), .b ({signal_2718, signal_1234}), .a ({IN_plaintext_s1[29], IN_plaintext_s0[29]}), .c ({signal_2769, signal_1170}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_133 ( .s (IN_reset), .b ({signal_2675, signal_1233}), .a ({IN_plaintext_s1[30], IN_plaintext_s0[30]}), .c ({signal_2738, signal_1169}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_134 ( .s (IN_reset), .b ({signal_2635, signal_1232}), .a ({IN_plaintext_s1[31], IN_plaintext_s0[31]}), .c ({signal_2693, signal_1168}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_135 ( .s (IN_reset), .b ({signal_2719, signal_1231}), .a ({IN_plaintext_s1[32], IN_plaintext_s0[32]}), .c ({signal_2771, signal_1167}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_136 ( .s (IN_reset), .b ({signal_2755, signal_1230}), .a ({IN_plaintext_s1[33], IN_plaintext_s0[33]}), .c ({signal_2803, signal_1166}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_137 ( .s (IN_reset), .b ({signal_2720, signal_1229}), .a ({IN_plaintext_s1[34], IN_plaintext_s0[34]}), .c ({signal_2773, signal_1165}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_138 ( .s (IN_reset), .b ({signal_2795, signal_1228}), .a ({IN_plaintext_s1[35], IN_plaintext_s0[35]}), .c ({signal_2823, signal_1164}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_139 ( .s (IN_reset), .b ({signal_2721, signal_1227}), .a ({IN_plaintext_s1[36], IN_plaintext_s0[36]}), .c ({signal_2775, signal_1163}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_140 ( .s (IN_reset), .b ({signal_2722, signal_1226}), .a ({IN_plaintext_s1[37], IN_plaintext_s0[37]}), .c ({signal_2777, signal_1162}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_141 ( .s (IN_reset), .b ({signal_2676, signal_1225}), .a ({IN_plaintext_s1[38], IN_plaintext_s0[38]}), .c ({signal_2740, signal_1161}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_142 ( .s (IN_reset), .b ({signal_2796, signal_1224}), .a ({IN_plaintext_s1[39], IN_plaintext_s0[39]}), .c ({signal_2825, signal_1160}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_143 ( .s (IN_reset), .b ({signal_2723, signal_1223}), .a ({IN_plaintext_s1[40], IN_plaintext_s0[40]}), .c ({signal_2779, signal_1159}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_144 ( .s (IN_reset), .b ({signal_2724, signal_1222}), .a ({IN_plaintext_s1[41], IN_plaintext_s0[41]}), .c ({signal_2781, signal_1158}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_145 ( .s (IN_reset), .b ({signal_2677, signal_1221}), .a ({IN_plaintext_s1[42], IN_plaintext_s0[42]}), .c ({signal_2742, signal_1157}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_146 ( .s (IN_reset), .b ({signal_2756, signal_1220}), .a ({IN_plaintext_s1[43], IN_plaintext_s0[43]}), .c ({signal_2805, signal_1156}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_147 ( .s (IN_reset), .b ({signal_2725, signal_1219}), .a ({IN_plaintext_s1[44], IN_plaintext_s0[44]}), .c ({signal_2783, signal_1155}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_148 ( .s (IN_reset), .b ({signal_2757, signal_1218}), .a ({IN_plaintext_s1[45], IN_plaintext_s0[45]}), .c ({signal_2807, signal_1154}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_149 ( .s (IN_reset), .b ({signal_2726, signal_1217}), .a ({IN_plaintext_s1[46], IN_plaintext_s0[46]}), .c ({signal_2785, signal_1153}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_150 ( .s (IN_reset), .b ({signal_2758, signal_1216}), .a ({IN_plaintext_s1[47], IN_plaintext_s0[47]}), .c ({signal_2809, signal_1152}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_151 ( .s (IN_reset), .b ({signal_2852, signal_1215}), .a ({IN_plaintext_s1[48], IN_plaintext_s0[48]}), .c ({signal_2865, signal_1151}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_152 ( .s (IN_reset), .b ({signal_2862, signal_1214}), .a ({IN_plaintext_s1[49], IN_plaintext_s0[49]}), .c ({signal_2873, signal_1150}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_153 ( .s (IN_reset), .b ({signal_2797, signal_1213}), .a ({IN_plaintext_s1[50], IN_plaintext_s0[50]}), .c ({signal_2827, signal_1149}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_154 ( .s (IN_reset), .b ({signal_2798, signal_1212}), .a ({IN_plaintext_s1[51], IN_plaintext_s0[51]}), .c ({signal_2829, signal_1148}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_155 ( .s (IN_reset), .b ({signal_2853, signal_1211}), .a ({IN_plaintext_s1[52], IN_plaintext_s0[52]}), .c ({signal_2867, signal_1147}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_156 ( .s (IN_reset), .b ({signal_2863, signal_1210}), .a ({IN_plaintext_s1[53], IN_plaintext_s0[53]}), .c ({signal_2875, signal_1146}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_157 ( .s (IN_reset), .b ({signal_2759, signal_1209}), .a ({IN_plaintext_s1[54], IN_plaintext_s0[54]}), .c ({signal_2811, signal_1145}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_158 ( .s (IN_reset), .b ({signal_2799, signal_1208}), .a ({IN_plaintext_s1[55], IN_plaintext_s0[55]}), .c ({signal_2831, signal_1144}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_159 ( .s (IN_reset), .b ({signal_2844, signal_1207}), .a ({IN_plaintext_s1[56], IN_plaintext_s0[56]}), .c ({signal_2857, signal_1143}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_160 ( .s (IN_reset), .b ({signal_2854, signal_1206}), .a ({IN_plaintext_s1[57], IN_plaintext_s0[57]}), .c ({signal_2869, signal_1142}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_161 ( .s (IN_reset), .b ({signal_2760, signal_1205}), .a ({IN_plaintext_s1[58], IN_plaintext_s0[58]}), .c ({signal_2813, signal_1141}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_162 ( .s (IN_reset), .b ({signal_2761, signal_1204}), .a ({IN_plaintext_s1[59], IN_plaintext_s0[59]}), .c ({signal_2815, signal_1140}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_163 ( .s (IN_reset), .b ({signal_2845, signal_1203}), .a ({IN_plaintext_s1[60], IN_plaintext_s0[60]}), .c ({signal_2859, signal_1139}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_164 ( .s (IN_reset), .b ({signal_2855, signal_1202}), .a ({IN_plaintext_s1[61], IN_plaintext_s0[61]}), .c ({signal_2871, signal_1138}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_165 ( .s (IN_reset), .b ({signal_2800, signal_1201}), .a ({IN_plaintext_s1[62], IN_plaintext_s0[62]}), .c ({signal_2833, signal_1137}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_166 ( .s (IN_reset), .b ({signal_2801, signal_1200}), .a ({IN_plaintext_s1[63], IN_plaintext_s0[63]}), .c ({signal_2835, signal_1136}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_412 ( .a ({signal_1993, signal_1007}), .b ({signal_2436, signal_356}), .c ({signal_2467, signal_940}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_435 ( .a ({signal_2061, signal_1003}), .b ({signal_2439, signal_375}), .c ({signal_2468, signal_936}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_458 ( .a ({signal_2000, signal_999}), .b ({signal_2404, signal_394}), .c ({signal_2428, signal_932}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_481 ( .a ({signal_2004, signal_995}), .b ({signal_2407, signal_413}), .c ({signal_2429, signal_928}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_504 ( .a ({signal_1992, signal_991}), .b ({signal_2442, signal_432}), .c ({signal_2469, signal_924}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_527 ( .a ({signal_2069, signal_987}), .b ({signal_2445, signal_451}), .c ({signal_2470, signal_920}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_550 ( .a ({signal_1879, signal_983}), .b ({signal_2410, signal_470}), .c ({signal_2430, signal_916}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_573 ( .a ({signal_1983, signal_979}), .b ({signal_2413, signal_489}), .c ({signal_2431, signal_912}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_596 ( .a ({signal_2048, signal_975}), .b ({signal_2448, signal_508}), .c ({signal_2471, signal_908}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_619 ( .a ({signal_2045, signal_971}), .b ({signal_2451, signal_527}), .c ({signal_2472, signal_904}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_642 ( .a ({signal_2021, signal_967}), .b ({signal_2416, signal_546}), .c ({signal_2432, signal_900}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_665 ( .a ({signal_2025, signal_963}), .b ({signal_2419, signal_565}), .c ({signal_2433, signal_896}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_688 ( .a ({signal_2063, signal_959}), .b ({signal_2454, signal_584}), .c ({signal_2473, signal_892}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_711 ( .a ({signal_2058, signal_955}), .b ({signal_2457, signal_603}), .c ({signal_2474, signal_888}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_734 ( .a ({signal_2037, signal_951}), .b ({signal_2422, signal_622}), .c ({signal_2434, signal_884}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_757 ( .a ({signal_2041, signal_947}), .b ({signal_2425, signal_641}), .c ({signal_2435, signal_880}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_762 ( .a ({signal_2743, signal_656}), .b ({signal_2604, signal_657}), .c ({signal_2786, signal_1276}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_763 ( .a ({signal_2565, signal_1324}), .b ({signal_2427, signal_882}), .c ({signal_2604, signal_657}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_764 ( .a ({signal_2694, signal_1293}), .b ({signal_2697, signal_1309}), .c ({signal_2743, signal_656}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_765 ( .a ({signal_2562, signal_658}), .b ({signal_2649, signal_659}), .c ({signal_2694, signal_1293}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_766 ( .a ({signal_2426, signal_881}), .b ({signal_2533, signal_660}), .c ({signal_2562, signal_658}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_767 ( .a ({signal_2695, signal_661}), .b ({signal_2745, signal_1294}), .c ({signal_2787, signal_1277}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_768 ( .a ({signal_2534, signal_1325}), .b ({signal_2649, signal_659}), .c ({signal_2695, signal_661}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_769 ( .a ({signal_2846, signal_662}), .b ({signal_2698, signal_663}), .c ({signal_2860, signal_1278}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_770 ( .a ({signal_2836, signal_664}), .b ({signal_2644, signal_665}), .c ({signal_2846, signal_662}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_771 ( .a ({signal_2435, signal_880}), .b ({signal_2606, signal_1326}), .c ({signal_2644, signal_665}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_772 ( .a ({signal_2696, signal_1295}), .b ({signal_2816, signal_666}), .c ({signal_2836, signal_664}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_773 ( .a ({signal_2645, signal_667}), .b ({signal_2605, signal_668}), .c ({signal_2696, signal_1295}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_774 ( .a ({signal_2417, signal_901}), .b ({signal_2565, signal_1324}), .c ({signal_2605, signal_668}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_775 ( .a ({signal_2259, signal_883}), .b ({signal_2608, signal_1308}), .c ({signal_2645, signal_667}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_776 ( .a ({signal_2837, signal_669}), .b ({signal_2503, signal_1327}), .c ({signal_2847, signal_1279}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_777 ( .a ({signal_2608, signal_1308}), .b ({signal_2816, signal_666}), .c ({signal_2837, signal_669}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_778 ( .a ({signal_2426, signal_881}), .b ({signal_2788, signal_1292}), .c ({signal_2816, signal_666}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_779 ( .a ({signal_2744, signal_670}), .b ({signal_2475, signal_671}), .c ({signal_2788, signal_1292}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_780 ( .a ({signal_2435, signal_880}), .b ({signal_2418, signal_902}), .c ({signal_2475, signal_671}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_781 ( .a ({signal_2697, signal_1309}), .b ({signal_2534, signal_1325}), .c ({signal_2744, signal_670}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_782 ( .a ({signal_2646, signal_672}), .b ({signal_2532, signal_673}), .c ({signal_2697, signal_1309}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_783 ( .a ({signal_2504, signal_674}), .b ({signal_2427, signal_882}), .c ({signal_2532, signal_673}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_784 ( .a ({signal_2606, signal_1326}), .b ({signal_2271, signal_923}), .c ({signal_2646, signal_672}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_785 ( .a ({signal_2563, signal_675}), .b ({signal_2476, signal_676}), .c ({signal_2606, signal_1326}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_786 ( .a ({signal_2256, signal_903}), .b ({signal_2432, signal_900}), .c ({signal_2476, signal_676}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_787 ( .a ({signal_2479, signal_677}), .b ({signal_2533, signal_660}), .c ({signal_2563, signal_675}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_788 ( .a ({signal_2500, signal_678}), .b ({signal_2437, signal_941}), .c ({signal_2533, signal_660}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_789 ( .a ({signal_2447, signal_922}), .b ({signal_2467, signal_940}), .c ({signal_2500, signal_678}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_790 ( .a ({signal_2699, signal_679}), .b ({signal_2698, signal_663}), .c ({signal_2745, signal_1294}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_791 ( .a ({signal_2648, signal_1311}), .b ({signal_2608, signal_1308}), .c ({signal_2698, signal_663}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_792 ( .a ({signal_2647, signal_680}), .b ({signal_2477, signal_681}), .c ({signal_2699, signal_679}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_793 ( .a ({signal_2417, signal_901}), .b ({signal_2432, signal_900}), .c ({signal_2477, signal_681}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_794 ( .a ({signal_2609, signal_682}), .b ({signal_2427, signal_882}), .c ({signal_2647, signal_680}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_795 ( .a ({signal_2491, signal_683}), .b ({signal_2607, signal_684}), .c ({signal_2648, signal_1311}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_796 ( .a ({signal_2565, signal_1324}), .b ({signal_2435, signal_880}), .c ({signal_2607, signal_684}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_798 ( .a ({signal_2564, signal_685}), .b ({signal_2478, signal_686}), .c ({signal_2608, signal_1308}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_799 ( .a ({signal_2426, signal_881}), .b ({signal_2432, signal_900}), .c ({signal_2478, signal_686}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_800 ( .a ({signal_2534, signal_1325}), .b ({signal_2447, signal_922}), .c ({signal_2564, signal_685}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_801 ( .a ({signal_2460, signal_687}), .b ({signal_2501, signal_688}), .c ({signal_2534, signal_1325}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_802 ( .a ({signal_2492, signal_689}), .b ({signal_2467, signal_940}), .c ({signal_2501, signal_688}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_804 ( .a ({signal_2479, signal_677}), .b ({signal_2649, signal_659}), .c ({signal_2700, signal_1310}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_805 ( .a ({signal_2502, signal_690}), .b ({signal_2609, signal_682}), .c ({signal_2649, signal_659}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_806 ( .a ({signal_2565, signal_1324}), .b ({signal_2503, signal_1327}), .c ({signal_2609, signal_682}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_807 ( .a ({signal_2470, signal_920}), .b ({signal_2492, signal_689}), .c ({signal_2502, signal_690}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_809 ( .a ({signal_2435, signal_880}), .b ({signal_2259, signal_883}), .c ({signal_2479, signal_677}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_810 ( .a ({signal_2493, signal_691}), .b ({signal_2480, signal_692}), .c ({signal_2503, signal_1327}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_811 ( .a ({signal_2435, signal_880}), .b ({signal_2432, signal_900}), .c ({signal_2480, signal_692}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_813 ( .a ({signal_2535, signal_693}), .b ({signal_2426, signal_881}), .c ({signal_2565, signal_1324}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_814 ( .a ({signal_2504, signal_674}), .b ({signal_2438, signal_942}), .c ({signal_2535, signal_693}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_815 ( .a ({signal_2417, signal_901}), .b ({signal_2470, signal_920}), .c ({signal_2504, signal_674}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_816 ( .a ({signal_2746, signal_694}), .b ({signal_2566, signal_695}), .c ({signal_2789, signal_1272}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_817 ( .a ({signal_2539, signal_1320}), .b ({signal_2456, signal_894}), .c ({signal_2566, signal_695}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_818 ( .a ({signal_2650, signal_1289}), .b ({signal_2702, signal_1305}), .c ({signal_2746, signal_694}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_819 ( .a ({signal_2567, signal_696}), .b ({signal_2614, signal_697}), .c ({signal_2650, signal_1289}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_820 ( .a ({signal_2455, signal_893}), .b ({signal_2536, signal_698}), .c ({signal_2567, signal_696}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_821 ( .a ({signal_2651, signal_699}), .b ({signal_2703, signal_1290}), .c ({signal_2747, signal_1273}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_822 ( .a ({signal_2537, signal_1321}), .b ({signal_2614, signal_697}), .c ({signal_2651, signal_699}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_823 ( .a ({signal_2848, signal_700}), .b ({signal_2655, signal_701}), .c ({signal_2861, signal_1274}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_824 ( .a ({signal_2838, signal_702}), .b ({signal_2652, signal_703}), .c ({signal_2848, signal_700}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_825 ( .a ({signal_2473, signal_892}), .b ({signal_2610, signal_1322}), .c ({signal_2652, signal_703}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_826 ( .a ({signal_2701, signal_1291}), .b ({signal_2817, signal_704}), .c ({signal_2838, signal_702}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_827 ( .a ({signal_2653, signal_705}), .b ({signal_2568, signal_706}), .c ({signal_2701, signal_1291}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_828 ( .a ({signal_2420, signal_897}), .b ({signal_2539, signal_1320}), .c ({signal_2568, signal_706}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_829 ( .a ({signal_2274, signal_895}), .b ({signal_2613, signal_1304}), .c ({signal_2653, signal_705}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_830 ( .a ({signal_2839, signal_707}), .b ({signal_2538, signal_1323}), .c ({signal_2849, signal_1275}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_831 ( .a ({signal_2613, signal_1304}), .b ({signal_2817, signal_704}), .c ({signal_2839, signal_707}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_832 ( .a ({signal_2455, signal_893}), .b ({signal_2790, signal_1288}), .c ({signal_2817, signal_704}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_833 ( .a ({signal_2748, signal_708}), .b ({signal_2505, signal_709}), .c ({signal_2790, signal_1288}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_834 ( .a ({signal_2473, signal_892}), .b ({signal_2421, signal_898}), .c ({signal_2505, signal_709}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_835 ( .a ({signal_2702, signal_1305}), .b ({signal_2537, signal_1321}), .c ({signal_2748, signal_708}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_836 ( .a ({signal_2654, signal_710}), .b ({signal_2506, signal_711}), .c ({signal_2702, signal_1305}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_837 ( .a ({signal_2485, signal_712}), .b ({signal_2456, signal_894}), .c ({signal_2506, signal_711}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_838 ( .a ({signal_2610, signal_1322}), .b ({signal_2254, signal_919}), .c ({signal_2654, signal_710}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_839 ( .a ({signal_2569, signal_713}), .b ({signal_2481, signal_714}), .c ({signal_2610, signal_1322}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_840 ( .a ({signal_2257, signal_899}), .b ({signal_2433, signal_896}), .c ({signal_2481, signal_714}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_841 ( .a ({signal_2509, signal_715}), .b ({signal_2536, signal_698}), .c ({signal_2569, signal_713}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_842 ( .a ({signal_2507, signal_716}), .b ({signal_2440, signal_937}), .c ({signal_2536, signal_698}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_843 ( .a ({signal_2412, signal_918}), .b ({signal_2468, signal_936}), .c ({signal_2507, signal_716}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_844 ( .a ({signal_2656, signal_717}), .b ({signal_2655, signal_701}), .c ({signal_2703, signal_1290}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_845 ( .a ({signal_2612, signal_1307}), .b ({signal_2613, signal_1304}), .c ({signal_2655, signal_701}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_846 ( .a ({signal_2611, signal_718}), .b ({signal_2482, signal_719}), .c ({signal_2656, signal_717}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_847 ( .a ({signal_2420, signal_897}), .b ({signal_2433, signal_896}), .c ({signal_2482, signal_719}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_848 ( .a ({signal_2572, signal_720}), .b ({signal_2456, signal_894}), .c ({signal_2611, signal_718}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_849 ( .a ({signal_2461, signal_721}), .b ({signal_2570, signal_722}), .c ({signal_2612, signal_1307}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_850 ( .a ({signal_2539, signal_1320}), .b ({signal_2473, signal_892}), .c ({signal_2570, signal_722}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_852 ( .a ({signal_2571, signal_723}), .b ({signal_2483, signal_724}), .c ({signal_2613, signal_1304}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_853 ( .a ({signal_2455, signal_893}), .b ({signal_2433, signal_896}), .c ({signal_2483, signal_724}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_854 ( .a ({signal_2537, signal_1321}), .b ({signal_2412, signal_918}), .c ({signal_2571, signal_723}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_855 ( .a ({signal_2494, signal_725}), .b ({signal_2508, signal_726}), .c ({signal_2537, signal_1321}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_856 ( .a ({signal_2462, signal_727}), .b ({signal_2468, signal_936}), .c ({signal_2508, signal_726}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_858 ( .a ({signal_2509, signal_715}), .b ({signal_2614, signal_697}), .c ({signal_2657, signal_1306}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_859 ( .a ({signal_2484, signal_728}), .b ({signal_2572, signal_720}), .c ({signal_2614, signal_697}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_860 ( .a ({signal_2539, signal_1320}), .b ({signal_2538, signal_1323}), .c ({signal_2572, signal_720}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_861 ( .a ({signal_2430, signal_916}), .b ({signal_2462, signal_727}), .c ({signal_2484, signal_728}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_863 ( .a ({signal_2473, signal_892}), .b ({signal_2274, signal_895}), .c ({signal_2509, signal_715}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_864 ( .a ({signal_2495, signal_729}), .b ({signal_2510, signal_730}), .c ({signal_2538, signal_1323}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_865 ( .a ({signal_2473, signal_892}), .b ({signal_2433, signal_896}), .c ({signal_2510, signal_730}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_867 ( .a ({signal_2511, signal_731}), .b ({signal_2455, signal_893}), .c ({signal_2539, signal_1320}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_868 ( .a ({signal_2485, signal_712}), .b ({signal_2441, signal_938}), .c ({signal_2511, signal_731}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_869 ( .a ({signal_2420, signal_897}), .b ({signal_2430, signal_916}), .c ({signal_2485, signal_712}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_870 ( .a ({signal_2704, signal_732}), .b ({signal_2573, signal_733}), .c ({signal_2749, signal_1268}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_871 ( .a ({signal_2544, signal_1316}), .b ({signal_2459, signal_890}), .c ({signal_2573, signal_733}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_872 ( .a ({signal_2658, signal_1285}), .b ({signal_2661, signal_1301}), .c ({signal_2704, signal_732}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_873 ( .a ({signal_2540, signal_734}), .b ({signal_2620, signal_735}), .c ({signal_2658, signal_1285}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_874 ( .a ({signal_2458, signal_889}), .b ({signal_2515, signal_736}), .c ({signal_2540, signal_734}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_875 ( .a ({signal_2659, signal_737}), .b ({signal_2707, signal_1286}), .c ({signal_2750, signal_1269}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_876 ( .a ({signal_2542, signal_1317}), .b ({signal_2620, signal_735}), .c ({signal_2659, signal_737}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_877 ( .a ({signal_2840, signal_738}), .b ({signal_2662, signal_739}), .c ({signal_2850, signal_1270}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_878 ( .a ({signal_2818, signal_740}), .b ({signal_2615, signal_741}), .c ({signal_2840, signal_738}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_879 ( .a ({signal_2474, signal_888}), .b ({signal_2575, signal_1318}), .c ({signal_2615, signal_741}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_880 ( .a ({signal_2705, signal_1287}), .b ({signal_2791, signal_742}), .c ({signal_2818, signal_740}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_881 ( .a ({signal_2660, signal_743}), .b ({signal_2574, signal_744}), .c ({signal_2705, signal_1287}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_882 ( .a ({signal_2449, signal_909}), .b ({signal_2544, signal_1316}), .c ({signal_2574, signal_744}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_883 ( .a ({signal_2275, signal_891}), .b ({signal_2619, signal_1300}), .c ({signal_2660, signal_743}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_884 ( .a ({signal_2819, signal_745}), .b ({signal_2543, signal_1319}), .c ({signal_2841, signal_1271}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_885 ( .a ({signal_2619, signal_1300}), .b ({signal_2791, signal_742}), .c ({signal_2819, signal_745}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_886 ( .a ({signal_2458, signal_889}), .b ({signal_2751, signal_1284}), .c ({signal_2791, signal_742}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_887 ( .a ({signal_2706, signal_746}), .b ({signal_2512, signal_747}), .c ({signal_2751, signal_1284}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_888 ( .a ({signal_2474, signal_888}), .b ({signal_2450, signal_910}), .c ({signal_2512, signal_747}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_889 ( .a ({signal_2661, signal_1301}), .b ({signal_2542, signal_1317}), .c ({signal_2706, signal_746}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_890 ( .a ({signal_2616, signal_748}), .b ({signal_2513, signal_749}), .c ({signal_2661, signal_1301}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_891 ( .a ({signal_2487, signal_750}), .b ({signal_2459, signal_890}), .c ({signal_2513, signal_749}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_892 ( .a ({signal_2575, signal_1318}), .b ({signal_2255, signal_915}), .c ({signal_2616, signal_748}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_893 ( .a ({signal_2541, signal_751}), .b ({signal_2514, signal_752}), .c ({signal_2575, signal_1318}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_894 ( .a ({signal_2272, signal_911}), .b ({signal_2471, signal_908}), .c ({signal_2514, signal_752}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_895 ( .a ({signal_2520, signal_753}), .b ({signal_2515, signal_736}), .c ({signal_2541, signal_751}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_896 ( .a ({signal_2486, signal_754}), .b ({signal_2405, signal_933}), .c ({signal_2515, signal_736}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_897 ( .a ({signal_2415, signal_914}), .b ({signal_2428, signal_932}), .c ({signal_2486, signal_754}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_898 ( .a ({signal_2663, signal_755}), .b ({signal_2662, signal_739}), .c ({signal_2707, signal_1286}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_899 ( .a ({signal_2618, signal_1303}), .b ({signal_2619, signal_1300}), .c ({signal_2662, signal_739}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_900 ( .a ({signal_2617, signal_756}), .b ({signal_2516, signal_757}), .c ({signal_2663, signal_755}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_901 ( .a ({signal_2449, signal_909}), .b ({signal_2471, signal_908}), .c ({signal_2516, signal_757}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_902 ( .a ({signal_2578, signal_758}), .b ({signal_2459, signal_890}), .c ({signal_2617, signal_756}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_903 ( .a ({signal_2463, signal_759}), .b ({signal_2576, signal_760}), .c ({signal_2618, signal_1303}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_904 ( .a ({signal_2544, signal_1316}), .b ({signal_2474, signal_888}), .c ({signal_2576, signal_760}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_906 ( .a ({signal_2577, signal_761}), .b ({signal_2517, signal_762}), .c ({signal_2619, signal_1300}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_907 ( .a ({signal_2458, signal_889}), .b ({signal_2471, signal_908}), .c ({signal_2517, signal_762}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_908 ( .a ({signal_2542, signal_1317}), .b ({signal_2415, signal_914}), .c ({signal_2577, signal_761}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_909 ( .a ({signal_2496, signal_763}), .b ({signal_2518, signal_764}), .c ({signal_2542, signal_1317}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_910 ( .a ({signal_2497, signal_765}), .b ({signal_2428, signal_932}), .c ({signal_2518, signal_764}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_912 ( .a ({signal_2520, signal_753}), .b ({signal_2620, signal_735}), .c ({signal_2664, signal_1302}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_913 ( .a ({signal_2519, signal_766}), .b ({signal_2578, signal_758}), .c ({signal_2620, signal_735}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_914 ( .a ({signal_2544, signal_1316}), .b ({signal_2543, signal_1319}), .c ({signal_2578, signal_758}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_915 ( .a ({signal_2431, signal_912}), .b ({signal_2497, signal_765}), .c ({signal_2519, signal_766}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_917 ( .a ({signal_2474, signal_888}), .b ({signal_2275, signal_891}), .c ({signal_2520, signal_753}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_918 ( .a ({signal_2464, signal_767}), .b ({signal_2521, signal_768}), .c ({signal_2543, signal_1319}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_919 ( .a ({signal_2474, signal_888}), .b ({signal_2471, signal_908}), .c ({signal_2521, signal_768}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_921 ( .a ({signal_2522, signal_769}), .b ({signal_2458, signal_889}), .c ({signal_2544, signal_1316}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_922 ( .a ({signal_2487, signal_750}), .b ({signal_2406, signal_934}), .c ({signal_2522, signal_769}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_923 ( .a ({signal_2449, signal_909}), .b ({signal_2431, signal_912}), .c ({signal_2487, signal_750}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_924 ( .a ({signal_2752, signal_770}), .b ({signal_2621, signal_771}), .c ({signal_2792, signal_1264}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_925 ( .a ({signal_2581, signal_1312}), .b ({signal_2424, signal_886}), .c ({signal_2621, signal_771}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_926 ( .a ({signal_2708, signal_1281}), .b ({signal_2666, signal_1297}), .c ({signal_2752, signal_770}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_927 ( .a ({signal_2545, signal_772}), .b ({signal_2669, signal_773}), .c ({signal_2708, signal_1281}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_928 ( .a ({signal_2423, signal_885}), .b ({signal_2524, signal_774}), .c ({signal_2545, signal_772}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_929 ( .a ({signal_2709, signal_775}), .b ({signal_2754, signal_1282}), .c ({signal_2793, signal_1265}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_930 ( .a ({signal_2548, signal_1313}), .b ({signal_2669, signal_773}), .c ({signal_2709, signal_775}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_931 ( .a ({signal_2842, signal_776}), .b ({signal_2712, signal_777}), .c ({signal_2851, signal_1266}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_932 ( .a ({signal_2820, signal_778}), .b ({signal_2622, signal_779}), .c ({signal_2842, signal_776}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_933 ( .a ({signal_2434, signal_884}), .b ({signal_2579, signal_1314}), .c ({signal_2622, signal_779}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_934 ( .a ({signal_2710, signal_1283}), .b ({signal_2794, signal_780}), .c ({signal_2820, signal_778}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_935 ( .a ({signal_2665, signal_781}), .b ({signal_2623, signal_782}), .c ({signal_2710, signal_1283}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_936 ( .a ({signal_2452, signal_905}), .b ({signal_2581, signal_1312}), .c ({signal_2623, signal_782}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_937 ( .a ({signal_2258, signal_887}), .b ({signal_2626, signal_1296}), .c ({signal_2665, signal_781}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_938 ( .a ({signal_2821, signal_783}), .b ({signal_2549, signal_1315}), .c ({signal_2843, signal_1267}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_939 ( .a ({signal_2626, signal_1296}), .b ({signal_2794, signal_780}), .c ({signal_2821, signal_783}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_940 ( .a ({signal_2423, signal_885}), .b ({signal_2753, signal_1280}), .c ({signal_2794, signal_780}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_941 ( .a ({signal_2711, signal_784}), .b ({signal_2488, signal_785}), .c ({signal_2753, signal_1280}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_942 ( .a ({signal_2434, signal_884}), .b ({signal_2453, signal_906}), .c ({signal_2488, signal_785}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_943 ( .a ({signal_2666, signal_1297}), .b ({signal_2548, signal_1313}), .c ({signal_2711, signal_784}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_944 ( .a ({signal_2624, signal_786}), .b ({signal_2546, signal_787}), .c ({signal_2666, signal_1297}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_945 ( .a ({signal_2530, signal_788}), .b ({signal_2424, signal_886}), .c ({signal_2546, signal_787}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_946 ( .a ({signal_2579, signal_1314}), .b ({signal_2270, signal_927}), .c ({signal_2624, signal_786}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_947 ( .a ({signal_2547, signal_789}), .b ({signal_2523, signal_790}), .c ({signal_2579, signal_1314}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_948 ( .a ({signal_2273, signal_907}), .b ({signal_2472, signal_904}), .c ({signal_2523, signal_790}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_949 ( .a ({signal_2490, signal_791}), .b ({signal_2524, signal_774}), .c ({signal_2547, signal_789}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_950 ( .a ({signal_2489, signal_792}), .b ({signal_2408, signal_929}), .c ({signal_2524, signal_774}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_951 ( .a ({signal_2444, signal_926}), .b ({signal_2429, signal_928}), .c ({signal_2489, signal_792}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_952 ( .a ({signal_2713, signal_793}), .b ({signal_2712, signal_777}), .c ({signal_2754, signal_1282}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_953 ( .a ({signal_2668, signal_1299}), .b ({signal_2626, signal_1296}), .c ({signal_2712, signal_777}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_954 ( .a ({signal_2667, signal_794}), .b ({signal_2525, signal_795}), .c ({signal_2713, signal_793}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_955 ( .a ({signal_2452, signal_905}), .b ({signal_2472, signal_904}), .c ({signal_2525, signal_795}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_956 ( .a ({signal_2627, signal_796}), .b ({signal_2424, signal_886}), .c ({signal_2667, signal_794}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_957 ( .a ({signal_2498, signal_797}), .b ({signal_2625, signal_798}), .c ({signal_2668, signal_1299}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_958 ( .a ({signal_2581, signal_1312}), .b ({signal_2434, signal_884}), .c ({signal_2625, signal_798}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_960 ( .a ({signal_2580, signal_799}), .b ({signal_2526, signal_800}), .c ({signal_2626, signal_1296}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_961 ( .a ({signal_2423, signal_885}), .b ({signal_2472, signal_904}), .c ({signal_2526, signal_800}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_962 ( .a ({signal_2548, signal_1313}), .b ({signal_2444, signal_926}), .c ({signal_2580, signal_799}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_963 ( .a ({signal_2465, signal_801}), .b ({signal_2527, signal_802}), .c ({signal_2548, signal_1313}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_964 ( .a ({signal_2499, signal_803}), .b ({signal_2429, signal_928}), .c ({signal_2527, signal_802}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_966 ( .a ({signal_2490, signal_791}), .b ({signal_2669, signal_773}), .c ({signal_2714, signal_1298}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_967 ( .a ({signal_2528, signal_804}), .b ({signal_2627, signal_796}), .c ({signal_2669, signal_773}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_968 ( .a ({signal_2581, signal_1312}), .b ({signal_2549, signal_1315}), .c ({signal_2627, signal_796}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_969 ( .a ({signal_2469, signal_924}), .b ({signal_2499, signal_803}), .c ({signal_2528, signal_804}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_971 ( .a ({signal_2434, signal_884}), .b ({signal_2258, signal_887}), .c ({signal_2490, signal_791}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_972 ( .a ({signal_2466, signal_805}), .b ({signal_2529, signal_806}), .c ({signal_2549, signal_1315}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_973 ( .a ({signal_2434, signal_884}), .b ({signal_2472, signal_904}), .c ({signal_2529, signal_806}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_975 ( .a ({signal_2550, signal_807}), .b ({signal_2423, signal_885}), .c ({signal_2581, signal_1312}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_976 ( .a ({signal_2530, signal_788}), .b ({signal_2409, signal_930}), .c ({signal_2550, signal_807}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_977 ( .a ({signal_2452, signal_905}), .b ({signal_2469, signal_924}), .c ({signal_2530, signal_788}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1416 ( .a ({signal_2221, signal_1457}), .b ({signal_2324, signal_1556}), .clk (CLK), .r (Fresh[32]), .c ({signal_2364, signal_1604}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1417 ( .a ({signal_2224, signal_1460}), .b ({signal_2325, signal_1557}), .clk (CLK), .r (Fresh[33]), .c ({signal_2365, signal_1605}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1418 ( .a ({signal_2181, signal_1463}), .b ({signal_2308, signal_1558}), .clk (CLK), .r (Fresh[34]), .c ({signal_2348, signal_1606}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1419 ( .a ({signal_2184, signal_1466}), .b ({signal_2309, signal_1559}), .clk (CLK), .r (Fresh[35]), .c ({signal_2349, signal_1607}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1420 ( .a ({signal_2227, signal_1469}), .b ({signal_2326, signal_1560}), .clk (CLK), .r (Fresh[36]), .c ({signal_2366, signal_1608}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1421 ( .a ({signal_2230, signal_1472}), .b ({signal_2327, signal_1561}), .clk (CLK), .r (Fresh[37]), .c ({signal_2367, signal_1609}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1422 ( .a ({signal_2187, signal_1475}), .b ({signal_2310, signal_1562}), .clk (CLK), .r (Fresh[38]), .c ({signal_2350, signal_1610}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1423 ( .a ({signal_2190, signal_1478}), .b ({signal_2311, signal_1563}), .clk (CLK), .r (Fresh[39]), .c ({signal_2351, signal_1611}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1424 ( .a ({signal_2233, signal_1481}), .b ({signal_2328, signal_1564}), .clk (CLK), .r (Fresh[40]), .c ({signal_2368, signal_1612}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1425 ( .a ({signal_2236, signal_1484}), .b ({signal_2329, signal_1565}), .clk (CLK), .r (Fresh[41]), .c ({signal_2369, signal_1613}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1426 ( .a ({signal_2193, signal_1487}), .b ({signal_2312, signal_1566}), .clk (CLK), .r (Fresh[42]), .c ({signal_2352, signal_1614}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1427 ( .a ({signal_2196, signal_1490}), .b ({signal_2313, signal_1567}), .clk (CLK), .r (Fresh[43]), .c ({signal_2353, signal_1615}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1428 ( .a ({signal_2239, signal_1493}), .b ({signal_2330, signal_1568}), .clk (CLK), .r (Fresh[44]), .c ({signal_2370, signal_1616}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1429 ( .a ({signal_2242, signal_1496}), .b ({signal_2331, signal_1569}), .clk (CLK), .r (Fresh[45]), .c ({signal_2371, signal_1617}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1430 ( .a ({signal_2199, signal_1499}), .b ({signal_2314, signal_1570}), .clk (CLK), .r (Fresh[46]), .c ({signal_2354, signal_1618}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1431 ( .a ({signal_2202, signal_1502}), .b ({signal_2315, signal_1571}), .clk (CLK), .r (Fresh[47]), .c ({signal_2355, signal_1619}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1432 ( .a ({signal_2222, signal_1458}), .b ({signal_2356, signal_1588}), .clk (CLK), .r (Fresh[48]), .c ({signal_2388, signal_1620}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1433 ( .a ({signal_2225, signal_1461}), .b ({signal_2357, signal_1589}), .clk (CLK), .r (Fresh[49]), .c ({signal_2389, signal_1621}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1434 ( .a ({signal_2182, signal_1464}), .b ({signal_2340, signal_1590}), .clk (CLK), .r (Fresh[50]), .c ({signal_2372, signal_1622}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1435 ( .a ({signal_2185, signal_1467}), .b ({signal_2341, signal_1591}), .clk (CLK), .r (Fresh[51]), .c ({signal_2373, signal_1623}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1436 ( .a ({signal_2228, signal_1470}), .b ({signal_2358, signal_1592}), .clk (CLK), .r (Fresh[52]), .c ({signal_2390, signal_1624}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1437 ( .a ({signal_2231, signal_1473}), .b ({signal_2359, signal_1593}), .clk (CLK), .r (Fresh[53]), .c ({signal_2391, signal_1625}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1438 ( .a ({signal_2188, signal_1476}), .b ({signal_2342, signal_1594}), .clk (CLK), .r (Fresh[54]), .c ({signal_2374, signal_1626}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1439 ( .a ({signal_2191, signal_1479}), .b ({signal_2343, signal_1595}), .clk (CLK), .r (Fresh[55]), .c ({signal_2375, signal_1627}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1440 ( .a ({signal_2234, signal_1482}), .b ({signal_2360, signal_1596}), .clk (CLK), .r (Fresh[56]), .c ({signal_2392, signal_1628}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1441 ( .a ({signal_2237, signal_1485}), .b ({signal_2361, signal_1597}), .clk (CLK), .r (Fresh[57]), .c ({signal_2393, signal_1629}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1442 ( .a ({signal_2194, signal_1488}), .b ({signal_2344, signal_1598}), .clk (CLK), .r (Fresh[58]), .c ({signal_2376, signal_1630}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1443 ( .a ({signal_2197, signal_1491}), .b ({signal_2345, signal_1599}), .clk (CLK), .r (Fresh[59]), .c ({signal_2377, signal_1631}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1444 ( .a ({signal_2240, signal_1494}), .b ({signal_2362, signal_1600}), .clk (CLK), .r (Fresh[60]), .c ({signal_2394, signal_1632}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1445 ( .a ({signal_2243, signal_1497}), .b ({signal_2363, signal_1601}), .clk (CLK), .r (Fresh[61]), .c ({signal_2395, signal_1633}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1446 ( .a ({signal_2200, signal_1500}), .b ({signal_2346, signal_1602}), .clk (CLK), .r (Fresh[62]), .c ({signal_2378, signal_1634}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1447 ( .a ({signal_2203, signal_1503}), .b ({signal_2347, signal_1603}), .clk (CLK), .r (Fresh[63]), .c ({signal_2379, signal_1635}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1448 ( .a ({signal_2293, signal_1525}), .b ({signal_2364, signal_1604}), .c ({signal_2396, signal_1636}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1449 ( .a ({signal_2295, signal_1527}), .b ({signal_2365, signal_1605}), .c ({signal_2397, signal_1637}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1450 ( .a ({signal_2277, signal_1529}), .b ({signal_2348, signal_1606}), .c ({signal_2380, signal_1638}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1451 ( .a ({signal_2279, signal_1531}), .b ({signal_2349, signal_1607}), .c ({signal_2381, signal_1639}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1452 ( .a ({signal_2297, signal_1533}), .b ({signal_2366, signal_1608}), .c ({signal_2398, signal_1640}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1453 ( .a ({signal_2299, signal_1535}), .b ({signal_2367, signal_1609}), .c ({signal_2399, signal_1641}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1454 ( .a ({signal_2281, signal_1537}), .b ({signal_2350, signal_1610}), .c ({signal_2382, signal_1642}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1455 ( .a ({signal_2283, signal_1539}), .b ({signal_2351, signal_1611}), .c ({signal_2383, signal_1643}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1456 ( .a ({signal_2301, signal_1541}), .b ({signal_2368, signal_1612}), .c ({signal_2400, signal_1644}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1457 ( .a ({signal_2303, signal_1543}), .b ({signal_2369, signal_1613}), .c ({signal_2401, signal_1645}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1458 ( .a ({signal_2285, signal_1545}), .b ({signal_2352, signal_1614}), .c ({signal_2384, signal_1646}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1459 ( .a ({signal_2287, signal_1547}), .b ({signal_2353, signal_1615}), .c ({signal_2385, signal_1647}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1460 ( .a ({signal_2305, signal_1549}), .b ({signal_2370, signal_1616}), .c ({signal_2402, signal_1648}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1461 ( .a ({signal_2307, signal_1551}), .b ({signal_2371, signal_1617}), .c ({signal_2403, signal_1649}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1462 ( .a ({signal_2289, signal_1553}), .b ({signal_2354, signal_1618}), .c ({signal_2386, signal_1650}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1463 ( .a ({signal_2291, signal_1555}), .b ({signal_2355, signal_1619}), .c ({signal_2387, signal_1651}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1464 ( .a ({signal_2293, signal_1525}), .b ({signal_2388, signal_1620}), .c ({signal_2436, signal_356}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1465 ( .a ({signal_2137, signal_1361}), .b ({signal_2396, signal_1636}), .c ({signal_2437, signal_941}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1466 ( .a ({signal_2138, signal_1363}), .b ({signal_2388, signal_1620}), .c ({signal_2438, signal_942}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1467 ( .a ({signal_2295, signal_1527}), .b ({signal_2389, signal_1621}), .c ({signal_2439, signal_375}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1468 ( .a ({signal_2140, signal_1365}), .b ({signal_2397, signal_1637}), .c ({signal_2440, signal_937}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1469 ( .a ({signal_2142, signal_1367}), .b ({signal_2389, signal_1621}), .c ({signal_2441, signal_938}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1470 ( .a ({signal_2277, signal_1529}), .b ({signal_2372, signal_1622}), .c ({signal_2404, signal_394}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1471 ( .a ({signal_2094, signal_1369}), .b ({signal_2380, signal_1638}), .c ({signal_2405, signal_933}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1472 ( .a ({signal_2096, signal_1371}), .b ({signal_2372, signal_1622}), .c ({signal_2406, signal_934}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1473 ( .a ({signal_2279, signal_1531}), .b ({signal_2373, signal_1623}), .c ({signal_2407, signal_413}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1474 ( .a ({signal_2098, signal_1373}), .b ({signal_2381, signal_1639}), .c ({signal_2408, signal_929}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1475 ( .a ({signal_2100, signal_1375}), .b ({signal_2373, signal_1623}), .c ({signal_2409, signal_930}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1476 ( .a ({signal_2297, signal_1533}), .b ({signal_2390, signal_1624}), .c ({signal_2442, signal_432}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1477 ( .a ({signal_2144, signal_1377}), .b ({signal_2398, signal_1640}), .c ({signal_2443, signal_1652}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1478 ( .a ({signal_2145, signal_1379}), .b ({signal_2390, signal_1624}), .c ({signal_2444, signal_926}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1479 ( .a ({signal_2299, signal_1535}), .b ({signal_2391, signal_1625}), .c ({signal_2445, signal_451}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1480 ( .a ({signal_2147, signal_1381}), .b ({signal_2399, signal_1641}), .c ({signal_2446, signal_1653}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1481 ( .a ({signal_2149, signal_1383}), .b ({signal_2391, signal_1625}), .c ({signal_2447, signal_922}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1482 ( .a ({signal_2281, signal_1537}), .b ({signal_2374, signal_1626}), .c ({signal_2410, signal_470}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1483 ( .a ({signal_2102, signal_1385}), .b ({signal_2382, signal_1642}), .c ({signal_2411, signal_1654}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1484 ( .a ({signal_2104, signal_1387}), .b ({signal_2374, signal_1626}), .c ({signal_2412, signal_918}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1485 ( .a ({signal_2283, signal_1539}), .b ({signal_2375, signal_1627}), .c ({signal_2413, signal_489}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1486 ( .a ({signal_2106, signal_1389}), .b ({signal_2383, signal_1643}), .c ({signal_2414, signal_1655}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1487 ( .a ({signal_2108, signal_1391}), .b ({signal_2375, signal_1627}), .c ({signal_2415, signal_914}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1488 ( .a ({signal_2301, signal_1541}), .b ({signal_2392, signal_1628}), .c ({signal_2448, signal_508}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1489 ( .a ({signal_2151, signal_1393}), .b ({signal_2400, signal_1644}), .c ({signal_2449, signal_909}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1490 ( .a ({signal_2152, signal_1395}), .b ({signal_2392, signal_1628}), .c ({signal_2450, signal_910}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1491 ( .a ({signal_2303, signal_1543}), .b ({signal_2393, signal_1629}), .c ({signal_2451, signal_527}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1492 ( .a ({signal_2154, signal_1397}), .b ({signal_2401, signal_1645}), .c ({signal_2452, signal_905}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1493 ( .a ({signal_2155, signal_1399}), .b ({signal_2393, signal_1629}), .c ({signal_2453, signal_906}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1494 ( .a ({signal_2285, signal_1545}), .b ({signal_2376, signal_1630}), .c ({signal_2416, signal_546}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1495 ( .a ({signal_2112, signal_1401}), .b ({signal_2384, signal_1646}), .c ({signal_2417, signal_901}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1496 ( .a ({signal_2114, signal_1403}), .b ({signal_2376, signal_1630}), .c ({signal_2418, signal_902}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1497 ( .a ({signal_2287, signal_1547}), .b ({signal_2377, signal_1631}), .c ({signal_2419, signal_565}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1498 ( .a ({signal_2116, signal_1405}), .b ({signal_2385, signal_1647}), .c ({signal_2420, signal_897}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1499 ( .a ({signal_2118, signal_1407}), .b ({signal_2377, signal_1631}), .c ({signal_2421, signal_898}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1500 ( .a ({signal_2305, signal_1549}), .b ({signal_2394, signal_1632}), .c ({signal_2454, signal_584}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1501 ( .a ({signal_2157, signal_1409}), .b ({signal_2402, signal_1648}), .c ({signal_2455, signal_893}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1502 ( .a ({signal_2159, signal_1411}), .b ({signal_2394, signal_1632}), .c ({signal_2456, signal_894}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1503 ( .a ({signal_2307, signal_1551}), .b ({signal_2395, signal_1633}), .c ({signal_2457, signal_603}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1504 ( .a ({signal_2161, signal_1413}), .b ({signal_2403, signal_1649}), .c ({signal_2458, signal_889}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1505 ( .a ({signal_2163, signal_1415}), .b ({signal_2395, signal_1633}), .c ({signal_2459, signal_890}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1506 ( .a ({signal_2289, signal_1553}), .b ({signal_2378, signal_1634}), .c ({signal_2422, signal_622}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1507 ( .a ({signal_2120, signal_1417}), .b ({signal_2386, signal_1650}), .c ({signal_2423, signal_885}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1508 ( .a ({signal_2122, signal_1419}), .b ({signal_2378, signal_1634}), .c ({signal_2424, signal_886}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1509 ( .a ({signal_2291, signal_1555}), .b ({signal_2379, signal_1635}), .c ({signal_2425, signal_641}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1510 ( .a ({signal_2124, signal_1421}), .b ({signal_2387, signal_1651}), .c ({signal_2426, signal_881}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1511 ( .a ({signal_2126, signal_1423}), .b ({signal_2379, signal_1635}), .c ({signal_2427, signal_882}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1512 ( .a ({signal_2256, signal_903}), .b ({signal_2446, signal_1653}), .c ({signal_2491, signal_683}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1513 ( .a ({signal_2268, signal_1520}), .b ({signal_2427, signal_882}), .c ({signal_2460, signal_687}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1514 ( .a ({signal_2446, signal_1653}), .b ({signal_2418, signal_902}), .c ({signal_2492, signal_689}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1515 ( .a ({signal_2271, signal_923}), .b ({signal_2437, signal_941}), .c ({signal_2493, signal_691}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1516 ( .a ({signal_2257, signal_899}), .b ({signal_2411, signal_1654}), .c ({signal_2461, signal_721}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1517 ( .a ({signal_2269, signal_1521}), .b ({signal_2456, signal_894}), .c ({signal_2494, signal_725}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1518 ( .a ({signal_2411, signal_1654}), .b ({signal_2421, signal_898}), .c ({signal_2462, signal_727}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1519 ( .a ({signal_2254, signal_919}), .b ({signal_2440, signal_937}), .c ({signal_2495, signal_729}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1520 ( .a ({signal_2272, signal_911}), .b ({signal_2414, signal_1655}), .c ({signal_2463, signal_759}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1521 ( .a ({signal_2252, signal_1522}), .b ({signal_2459, signal_890}), .c ({signal_2496, signal_763}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1522 ( .a ({signal_2414, signal_1655}), .b ({signal_2450, signal_910}), .c ({signal_2497, signal_765}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1523 ( .a ({signal_2255, signal_915}), .b ({signal_2405, signal_933}), .c ({signal_2464, signal_767}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1524 ( .a ({signal_2273, signal_907}), .b ({signal_2443, signal_1652}), .c ({signal_2498, signal_797}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1525 ( .a ({signal_2253, signal_1523}), .b ({signal_2424, signal_886}), .c ({signal_2465, signal_801}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1526 ( .a ({signal_2443, signal_1652}), .b ({signal_2453, signal_906}), .c ({signal_2499, signal_803}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1527 ( .a ({signal_2270, signal_927}), .b ({signal_2408, signal_929}), .c ({signal_2466, signal_805}) ) ;

    /* register cells */
    DFF_X1 cell_979 ( .CK (signal_2940), .D (signal_310), .Q (signal_808), .QN () ) ;
    DFF_X1 cell_981 ( .CK (signal_2940), .D (signal_308), .Q (signal_307), .QN () ) ;
    DFF_X1 cell_983 ( .CK (signal_2940), .D (signal_305), .Q (signal_304), .QN () ) ;
    DFF_X1 cell_985 ( .CK (signal_2940), .D (signal_303), .Q (signal_288), .QN () ) ;
    DFF_X1 cell_987 ( .CK (signal_2940), .D (signal_301), .Q (signal_879), .QN () ) ;
    DFF_X1 cell_989 ( .CK (signal_2940), .D (signal_299), .Q (signal_878), .QN () ) ;
    DFF_X1 cell_991 ( .CK (signal_2940), .D (signal_297), .Q (signal_877), .QN () ) ;
    DFF_X1 cell_993 ( .CK (signal_2940), .D (signal_295), .Q (signal_876), .QN () ) ;
    DFF_X1 cell_995 ( .CK (signal_2940), .D (signal_293), .Q (signal_875), .QN () ) ;
    DFF_X1 cell_997 ( .CK (signal_2940), .D (signal_291), .Q (signal_874), .QN () ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_999 ( .clk (signal_2940), .D ({signal_2561, signal_1199}), .Q ({OUT_ciphertext_s1[0], OUT_ciphertext_s0[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1001 ( .clk (signal_2940), .D ({signal_2679, signal_1198}), .Q ({OUT_ciphertext_s1[1], OUT_ciphertext_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1003 ( .clk (signal_2940), .D ({signal_2587, signal_1197}), .Q ({OUT_ciphertext_s1[2], OUT_ciphertext_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1005 ( .clk (signal_2940), .D ({signal_2637, signal_1196}), .Q ({OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1007 ( .clk (signal_2940), .D ({signal_2589, signal_1195}), .Q ({OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1009 ( .clk (signal_2940), .D ({signal_2681, signal_1194}), .Q ({OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1011 ( .clk (signal_2940), .D ({signal_2591, signal_1193}), .Q ({OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1013 ( .clk (signal_2940), .D ({signal_2593, signal_1192}), .Q ({OUT_ciphertext_s1[7], OUT_ciphertext_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1015 ( .clk (signal_2940), .D ({signal_2595, signal_1191}), .Q ({OUT_ciphertext_s1[8], OUT_ciphertext_s0[8]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1017 ( .clk (signal_2940), .D ({signal_2639, signal_1190}), .Q ({OUT_ciphertext_s1[9], OUT_ciphertext_s0[9]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1019 ( .clk (signal_2940), .D ({signal_2597, signal_1189}), .Q ({OUT_ciphertext_s1[10], OUT_ciphertext_s0[10]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1021 ( .clk (signal_2940), .D ({signal_2599, signal_1188}), .Q ({OUT_ciphertext_s1[11], OUT_ciphertext_s0[11]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1023 ( .clk (signal_2940), .D ({signal_2601, signal_1187}), .Q ({OUT_ciphertext_s1[12], OUT_ciphertext_s0[12]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1025 ( .clk (signal_2940), .D ({signal_2641, signal_1186}), .Q ({OUT_ciphertext_s1[13], OUT_ciphertext_s0[13]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1027 ( .clk (signal_2940), .D ({signal_2603, signal_1185}), .Q ({OUT_ciphertext_s1[14], OUT_ciphertext_s0[14]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1029 ( .clk (signal_2940), .D ({signal_2643, signal_1184}), .Q ({OUT_ciphertext_s1[15], OUT_ciphertext_s0[15]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1031 ( .clk (signal_2940), .D ({signal_2728, signal_1183}), .Q ({OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1033 ( .clk (signal_2940), .D ({signal_2763, signal_1182}), .Q ({OUT_ciphertext_s1[17], OUT_ciphertext_s0[17]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1035 ( .clk (signal_2940), .D ({signal_2765, signal_1181}), .Q ({OUT_ciphertext_s1[18], OUT_ciphertext_s0[18]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1037 ( .clk (signal_2940), .D ({signal_2683, signal_1180}), .Q ({OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1039 ( .clk (signal_2940), .D ({signal_2685, signal_1179}), .Q ({OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1041 ( .clk (signal_2940), .D ({signal_2730, signal_1178}), .Q ({OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1043 ( .clk (signal_2940), .D ({signal_2767, signal_1177}), .Q ({OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1045 ( .clk (signal_2940), .D ({signal_2687, signal_1176}), .Q ({OUT_ciphertext_s1[23], OUT_ciphertext_s0[23]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1047 ( .clk (signal_2940), .D ({signal_2689, signal_1175}), .Q ({OUT_ciphertext_s1[24], OUT_ciphertext_s0[24]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1049 ( .clk (signal_2940), .D ({signal_2732, signal_1174}), .Q ({OUT_ciphertext_s1[25], OUT_ciphertext_s0[25]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1051 ( .clk (signal_2940), .D ({signal_2734, signal_1173}), .Q ({OUT_ciphertext_s1[26], OUT_ciphertext_s0[26]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1053 ( .clk (signal_2940), .D ({signal_2691, signal_1172}), .Q ({OUT_ciphertext_s1[27], OUT_ciphertext_s0[27]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1055 ( .clk (signal_2940), .D ({signal_2736, signal_1171}), .Q ({OUT_ciphertext_s1[28], OUT_ciphertext_s0[28]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1057 ( .clk (signal_2940), .D ({signal_2769, signal_1170}), .Q ({OUT_ciphertext_s1[29], OUT_ciphertext_s0[29]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1059 ( .clk (signal_2940), .D ({signal_2738, signal_1169}), .Q ({OUT_ciphertext_s1[30], OUT_ciphertext_s0[30]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1061 ( .clk (signal_2940), .D ({signal_2693, signal_1168}), .Q ({OUT_ciphertext_s1[31], OUT_ciphertext_s0[31]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1063 ( .clk (signal_2940), .D ({signal_2771, signal_1167}), .Q ({OUT_ciphertext_s1[32], OUT_ciphertext_s0[32]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1065 ( .clk (signal_2940), .D ({signal_2803, signal_1166}), .Q ({OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1067 ( .clk (signal_2940), .D ({signal_2773, signal_1165}), .Q ({OUT_ciphertext_s1[34], OUT_ciphertext_s0[34]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1069 ( .clk (signal_2940), .D ({signal_2823, signal_1164}), .Q ({OUT_ciphertext_s1[35], OUT_ciphertext_s0[35]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1071 ( .clk (signal_2940), .D ({signal_2775, signal_1163}), .Q ({OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1073 ( .clk (signal_2940), .D ({signal_2777, signal_1162}), .Q ({OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1075 ( .clk (signal_2940), .D ({signal_2740, signal_1161}), .Q ({OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1077 ( .clk (signal_2940), .D ({signal_2825, signal_1160}), .Q ({OUT_ciphertext_s1[39], OUT_ciphertext_s0[39]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1079 ( .clk (signal_2940), .D ({signal_2779, signal_1159}), .Q ({OUT_ciphertext_s1[40], OUT_ciphertext_s0[40]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1081 ( .clk (signal_2940), .D ({signal_2781, signal_1158}), .Q ({OUT_ciphertext_s1[41], OUT_ciphertext_s0[41]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1083 ( .clk (signal_2940), .D ({signal_2742, signal_1157}), .Q ({OUT_ciphertext_s1[42], OUT_ciphertext_s0[42]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1085 ( .clk (signal_2940), .D ({signal_2805, signal_1156}), .Q ({OUT_ciphertext_s1[43], OUT_ciphertext_s0[43]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1087 ( .clk (signal_2940), .D ({signal_2783, signal_1155}), .Q ({OUT_ciphertext_s1[44], OUT_ciphertext_s0[44]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1089 ( .clk (signal_2940), .D ({signal_2807, signal_1154}), .Q ({OUT_ciphertext_s1[45], OUT_ciphertext_s0[45]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1091 ( .clk (signal_2940), .D ({signal_2785, signal_1153}), .Q ({OUT_ciphertext_s1[46], OUT_ciphertext_s0[46]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1093 ( .clk (signal_2940), .D ({signal_2809, signal_1152}), .Q ({OUT_ciphertext_s1[47], OUT_ciphertext_s0[47]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1095 ( .clk (signal_2940), .D ({signal_2865, signal_1151}), .Q ({OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1097 ( .clk (signal_2940), .D ({signal_2873, signal_1150}), .Q ({OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1099 ( .clk (signal_2940), .D ({signal_2827, signal_1149}), .Q ({OUT_ciphertext_s1[50], OUT_ciphertext_s0[50]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1101 ( .clk (signal_2940), .D ({signal_2829, signal_1148}), .Q ({OUT_ciphertext_s1[51], OUT_ciphertext_s0[51]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1103 ( .clk (signal_2940), .D ({signal_2867, signal_1147}), .Q ({OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1105 ( .clk (signal_2940), .D ({signal_2875, signal_1146}), .Q ({OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1107 ( .clk (signal_2940), .D ({signal_2811, signal_1145}), .Q ({OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1109 ( .clk (signal_2940), .D ({signal_2831, signal_1144}), .Q ({OUT_ciphertext_s1[55], OUT_ciphertext_s0[55]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1111 ( .clk (signal_2940), .D ({signal_2857, signal_1143}), .Q ({OUT_ciphertext_s1[56], OUT_ciphertext_s0[56]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1113 ( .clk (signal_2940), .D ({signal_2869, signal_1142}), .Q ({OUT_ciphertext_s1[57], OUT_ciphertext_s0[57]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1115 ( .clk (signal_2940), .D ({signal_2813, signal_1141}), .Q ({OUT_ciphertext_s1[58], OUT_ciphertext_s0[58]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1117 ( .clk (signal_2940), .D ({signal_2815, signal_1140}), .Q ({OUT_ciphertext_s1[59], OUT_ciphertext_s0[59]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1119 ( .clk (signal_2940), .D ({signal_2859, signal_1139}), .Q ({OUT_ciphertext_s1[60], OUT_ciphertext_s0[60]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1121 ( .clk (signal_2940), .D ({signal_2871, signal_1138}), .Q ({OUT_ciphertext_s1[61], OUT_ciphertext_s0[61]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1123 ( .clk (signal_2940), .D ({signal_2833, signal_1137}), .Q ({OUT_ciphertext_s1[62], OUT_ciphertext_s0[62]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1125 ( .clk (signal_2940), .D ({signal_2835, signal_1136}), .Q ({OUT_ciphertext_s1[63], OUT_ciphertext_s0[63]}) ) ;
    DFF_X1 cell_1127 ( .CK (signal_2940), .D (signal_265), .Q (OUT_done), .QN () ) ;
endmodule
