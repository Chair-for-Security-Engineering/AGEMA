////////////////////////////////////////////////////////////////////////////
// COMPANY : Ruhr University Bochum
// AUTHOR  : David Knichel david.knichel@rub.de and Amir Moradi amir.moradi@rub.de 
// DOCUMENT: [Low-Latency Hardware Private Circuits] https://eprint.iacr.org/2022/507
// /////////////////////////////////////////////////////////////////
//
// Copyright c 2022, David Knichel and  Amir Moradi
//
// All rights reserved.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
// ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
// WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
// DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
// INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
// LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION HOWEVER CAUSED AND
// ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// INCLUDING NEGLIGENCE OR OTHERWISE ARISING IN ANY WAY OUT OF THE USE OF THIS
// SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// Please see LICENSE and README for license and further instructions.
//
/* modified netlist. Source: module AES in file /AGEMA/Designs/AES_round-based/AGEMA/AES.v */
/* 4 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 5 register stage(s) in total */

module AES_HPC3_Pipeline_d1 (plaintext_s0, key_s0, clk, reset, key_s1, plaintext_s1, Fresh, ciphertext_s0, done, ciphertext_s1);
    input [127:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input reset ;
    input [127:0] key_s1 ;
    input [127:0] plaintext_s1 ;
    input [1359:0] Fresh ;
    output [127:0] ciphertext_s0 ;
    output done ;
    output [127:0] ciphertext_s1 ;
    wire n283 ;
    wire n285 ;
    wire n314 ;
    wire n315 ;
    wire n316 ;
    wire n317 ;
    wire n318 ;
    wire n319 ;
    wire n320 ;
    wire n321 ;
    wire n322 ;
    wire n323 ;
    wire n324 ;
    wire n325 ;
    wire n326 ;
    wire n327 ;
    wire n328 ;
    wire n329 ;
    wire n330 ;
    wire n331 ;
    wire n332 ;
    wire n333 ;
    wire n334 ;
    wire n335 ;
    wire n336 ;
    wire n337 ;
    wire n338 ;
    wire n339 ;
    wire RoundReg_Inst_ff_SDE_0_next_state ;
    wire RoundReg_Inst_ff_SDE_1_next_state ;
    wire RoundReg_Inst_ff_SDE_2_next_state ;
    wire RoundReg_Inst_ff_SDE_3_next_state ;
    wire RoundReg_Inst_ff_SDE_4_next_state ;
    wire RoundReg_Inst_ff_SDE_5_next_state ;
    wire RoundReg_Inst_ff_SDE_6_next_state ;
    wire RoundReg_Inst_ff_SDE_7_next_state ;
    wire RoundReg_Inst_ff_SDE_8_next_state ;
    wire RoundReg_Inst_ff_SDE_9_next_state ;
    wire RoundReg_Inst_ff_SDE_10_next_state ;
    wire RoundReg_Inst_ff_SDE_11_next_state ;
    wire RoundReg_Inst_ff_SDE_12_next_state ;
    wire RoundReg_Inst_ff_SDE_13_next_state ;
    wire RoundReg_Inst_ff_SDE_14_next_state ;
    wire RoundReg_Inst_ff_SDE_15_next_state ;
    wire RoundReg_Inst_ff_SDE_16_next_state ;
    wire RoundReg_Inst_ff_SDE_17_next_state ;
    wire RoundReg_Inst_ff_SDE_18_next_state ;
    wire RoundReg_Inst_ff_SDE_19_next_state ;
    wire RoundReg_Inst_ff_SDE_20_next_state ;
    wire RoundReg_Inst_ff_SDE_21_next_state ;
    wire RoundReg_Inst_ff_SDE_22_next_state ;
    wire RoundReg_Inst_ff_SDE_23_next_state ;
    wire RoundReg_Inst_ff_SDE_24_next_state ;
    wire RoundReg_Inst_ff_SDE_25_next_state ;
    wire RoundReg_Inst_ff_SDE_26_next_state ;
    wire RoundReg_Inst_ff_SDE_27_next_state ;
    wire RoundReg_Inst_ff_SDE_28_next_state ;
    wire RoundReg_Inst_ff_SDE_29_next_state ;
    wire RoundReg_Inst_ff_SDE_30_next_state ;
    wire RoundReg_Inst_ff_SDE_31_next_state ;
    wire RoundReg_Inst_ff_SDE_32_next_state ;
    wire RoundReg_Inst_ff_SDE_33_next_state ;
    wire RoundReg_Inst_ff_SDE_34_next_state ;
    wire RoundReg_Inst_ff_SDE_35_next_state ;
    wire RoundReg_Inst_ff_SDE_36_next_state ;
    wire RoundReg_Inst_ff_SDE_37_next_state ;
    wire RoundReg_Inst_ff_SDE_38_next_state ;
    wire RoundReg_Inst_ff_SDE_39_next_state ;
    wire RoundReg_Inst_ff_SDE_40_next_state ;
    wire RoundReg_Inst_ff_SDE_41_next_state ;
    wire RoundReg_Inst_ff_SDE_42_next_state ;
    wire RoundReg_Inst_ff_SDE_43_next_state ;
    wire RoundReg_Inst_ff_SDE_44_next_state ;
    wire RoundReg_Inst_ff_SDE_45_next_state ;
    wire RoundReg_Inst_ff_SDE_46_next_state ;
    wire RoundReg_Inst_ff_SDE_47_next_state ;
    wire RoundReg_Inst_ff_SDE_48_next_state ;
    wire RoundReg_Inst_ff_SDE_49_next_state ;
    wire RoundReg_Inst_ff_SDE_50_next_state ;
    wire RoundReg_Inst_ff_SDE_51_next_state ;
    wire RoundReg_Inst_ff_SDE_52_next_state ;
    wire RoundReg_Inst_ff_SDE_53_next_state ;
    wire RoundReg_Inst_ff_SDE_54_next_state ;
    wire RoundReg_Inst_ff_SDE_55_next_state ;
    wire RoundReg_Inst_ff_SDE_56_next_state ;
    wire RoundReg_Inst_ff_SDE_57_next_state ;
    wire RoundReg_Inst_ff_SDE_58_next_state ;
    wire RoundReg_Inst_ff_SDE_59_next_state ;
    wire RoundReg_Inst_ff_SDE_60_next_state ;
    wire RoundReg_Inst_ff_SDE_61_next_state ;
    wire RoundReg_Inst_ff_SDE_62_next_state ;
    wire RoundReg_Inst_ff_SDE_63_next_state ;
    wire RoundReg_Inst_ff_SDE_64_next_state ;
    wire RoundReg_Inst_ff_SDE_65_next_state ;
    wire RoundReg_Inst_ff_SDE_66_next_state ;
    wire RoundReg_Inst_ff_SDE_67_next_state ;
    wire RoundReg_Inst_ff_SDE_68_next_state ;
    wire RoundReg_Inst_ff_SDE_69_next_state ;
    wire RoundReg_Inst_ff_SDE_70_next_state ;
    wire RoundReg_Inst_ff_SDE_71_next_state ;
    wire RoundReg_Inst_ff_SDE_72_next_state ;
    wire RoundReg_Inst_ff_SDE_73_next_state ;
    wire RoundReg_Inst_ff_SDE_74_next_state ;
    wire RoundReg_Inst_ff_SDE_75_next_state ;
    wire RoundReg_Inst_ff_SDE_76_next_state ;
    wire RoundReg_Inst_ff_SDE_77_next_state ;
    wire RoundReg_Inst_ff_SDE_78_next_state ;
    wire RoundReg_Inst_ff_SDE_79_next_state ;
    wire RoundReg_Inst_ff_SDE_80_next_state ;
    wire RoundReg_Inst_ff_SDE_81_next_state ;
    wire RoundReg_Inst_ff_SDE_82_next_state ;
    wire RoundReg_Inst_ff_SDE_83_next_state ;
    wire RoundReg_Inst_ff_SDE_84_next_state ;
    wire RoundReg_Inst_ff_SDE_85_next_state ;
    wire RoundReg_Inst_ff_SDE_86_next_state ;
    wire RoundReg_Inst_ff_SDE_87_next_state ;
    wire RoundReg_Inst_ff_SDE_88_next_state ;
    wire RoundReg_Inst_ff_SDE_89_next_state ;
    wire RoundReg_Inst_ff_SDE_90_next_state ;
    wire RoundReg_Inst_ff_SDE_91_next_state ;
    wire RoundReg_Inst_ff_SDE_92_next_state ;
    wire RoundReg_Inst_ff_SDE_93_next_state ;
    wire RoundReg_Inst_ff_SDE_94_next_state ;
    wire RoundReg_Inst_ff_SDE_95_next_state ;
    wire RoundReg_Inst_ff_SDE_96_next_state ;
    wire RoundReg_Inst_ff_SDE_97_next_state ;
    wire RoundReg_Inst_ff_SDE_98_next_state ;
    wire RoundReg_Inst_ff_SDE_99_next_state ;
    wire RoundReg_Inst_ff_SDE_100_next_state ;
    wire RoundReg_Inst_ff_SDE_101_next_state ;
    wire RoundReg_Inst_ff_SDE_102_next_state ;
    wire RoundReg_Inst_ff_SDE_103_next_state ;
    wire RoundReg_Inst_ff_SDE_104_next_state ;
    wire RoundReg_Inst_ff_SDE_105_next_state ;
    wire RoundReg_Inst_ff_SDE_106_next_state ;
    wire RoundReg_Inst_ff_SDE_107_next_state ;
    wire RoundReg_Inst_ff_SDE_108_next_state ;
    wire RoundReg_Inst_ff_SDE_109_next_state ;
    wire RoundReg_Inst_ff_SDE_110_next_state ;
    wire RoundReg_Inst_ff_SDE_111_next_state ;
    wire RoundReg_Inst_ff_SDE_112_next_state ;
    wire RoundReg_Inst_ff_SDE_113_next_state ;
    wire RoundReg_Inst_ff_SDE_114_next_state ;
    wire RoundReg_Inst_ff_SDE_115_next_state ;
    wire RoundReg_Inst_ff_SDE_116_next_state ;
    wire RoundReg_Inst_ff_SDE_117_next_state ;
    wire RoundReg_Inst_ff_SDE_118_next_state ;
    wire RoundReg_Inst_ff_SDE_119_next_state ;
    wire RoundReg_Inst_ff_SDE_120_next_state ;
    wire RoundReg_Inst_ff_SDE_121_next_state ;
    wire RoundReg_Inst_ff_SDE_122_next_state ;
    wire RoundReg_Inst_ff_SDE_123_next_state ;
    wire RoundReg_Inst_ff_SDE_124_next_state ;
    wire RoundReg_Inst_ff_SDE_125_next_state ;
    wire RoundReg_Inst_ff_SDE_126_next_state ;
    wire RoundReg_Inst_ff_SDE_127_next_state ;
    wire SubBytesIns_Inst_Sbox_0_L29 ;
    wire SubBytesIns_Inst_Sbox_0_L28 ;
    wire SubBytesIns_Inst_Sbox_0_L27 ;
    wire SubBytesIns_Inst_Sbox_0_L26 ;
    wire SubBytesIns_Inst_Sbox_0_L25 ;
    wire SubBytesIns_Inst_Sbox_0_L24 ;
    wire SubBytesIns_Inst_Sbox_0_L23 ;
    wire SubBytesIns_Inst_Sbox_0_L22 ;
    wire SubBytesIns_Inst_Sbox_0_L21 ;
    wire SubBytesIns_Inst_Sbox_0_L20 ;
    wire SubBytesIns_Inst_Sbox_0_L19 ;
    wire SubBytesIns_Inst_Sbox_0_L18 ;
    wire SubBytesIns_Inst_Sbox_0_L17 ;
    wire SubBytesIns_Inst_Sbox_0_L16 ;
    wire SubBytesIns_Inst_Sbox_0_L15 ;
    wire SubBytesIns_Inst_Sbox_0_L14 ;
    wire SubBytesIns_Inst_Sbox_0_L13 ;
    wire SubBytesIns_Inst_Sbox_0_L12 ;
    wire SubBytesIns_Inst_Sbox_0_L11 ;
    wire SubBytesIns_Inst_Sbox_0_L10 ;
    wire SubBytesIns_Inst_Sbox_0_L9 ;
    wire SubBytesIns_Inst_Sbox_0_L8 ;
    wire SubBytesIns_Inst_Sbox_0_L7 ;
    wire SubBytesIns_Inst_Sbox_0_L6 ;
    wire SubBytesIns_Inst_Sbox_0_L5 ;
    wire SubBytesIns_Inst_Sbox_0_L4 ;
    wire SubBytesIns_Inst_Sbox_0_L3 ;
    wire SubBytesIns_Inst_Sbox_0_L2 ;
    wire SubBytesIns_Inst_Sbox_0_L1 ;
    wire SubBytesIns_Inst_Sbox_0_L0 ;
    wire SubBytesIns_Inst_Sbox_0_M63 ;
    wire SubBytesIns_Inst_Sbox_0_M62 ;
    wire SubBytesIns_Inst_Sbox_0_M61 ;
    wire SubBytesIns_Inst_Sbox_0_M60 ;
    wire SubBytesIns_Inst_Sbox_0_M59 ;
    wire SubBytesIns_Inst_Sbox_0_M58 ;
    wire SubBytesIns_Inst_Sbox_0_M57 ;
    wire SubBytesIns_Inst_Sbox_0_M56 ;
    wire SubBytesIns_Inst_Sbox_0_M55 ;
    wire SubBytesIns_Inst_Sbox_0_M54 ;
    wire SubBytesIns_Inst_Sbox_0_M53 ;
    wire SubBytesIns_Inst_Sbox_0_M52 ;
    wire SubBytesIns_Inst_Sbox_0_M51 ;
    wire SubBytesIns_Inst_Sbox_0_M50 ;
    wire SubBytesIns_Inst_Sbox_0_M49 ;
    wire SubBytesIns_Inst_Sbox_0_M48 ;
    wire SubBytesIns_Inst_Sbox_0_M47 ;
    wire SubBytesIns_Inst_Sbox_0_M46 ;
    wire SubBytesIns_Inst_Sbox_0_M45 ;
    wire SubBytesIns_Inst_Sbox_0_M44 ;
    wire SubBytesIns_Inst_Sbox_0_M43 ;
    wire SubBytesIns_Inst_Sbox_0_M42 ;
    wire SubBytesIns_Inst_Sbox_0_M41 ;
    wire SubBytesIns_Inst_Sbox_0_M40 ;
    wire SubBytesIns_Inst_Sbox_0_M39 ;
    wire SubBytesIns_Inst_Sbox_0_M38 ;
    wire SubBytesIns_Inst_Sbox_0_M37 ;
    wire SubBytesIns_Inst_Sbox_0_M36 ;
    wire SubBytesIns_Inst_Sbox_0_M35 ;
    wire SubBytesIns_Inst_Sbox_0_M34 ;
    wire SubBytesIns_Inst_Sbox_0_M33 ;
    wire SubBytesIns_Inst_Sbox_0_M32 ;
    wire SubBytesIns_Inst_Sbox_0_M31 ;
    wire SubBytesIns_Inst_Sbox_0_M30 ;
    wire SubBytesIns_Inst_Sbox_0_M29 ;
    wire SubBytesIns_Inst_Sbox_0_M28 ;
    wire SubBytesIns_Inst_Sbox_0_M27 ;
    wire SubBytesIns_Inst_Sbox_0_M26 ;
    wire SubBytesIns_Inst_Sbox_0_M25 ;
    wire SubBytesIns_Inst_Sbox_0_M24 ;
    wire SubBytesIns_Inst_Sbox_0_M23 ;
    wire SubBytesIns_Inst_Sbox_0_M22 ;
    wire SubBytesIns_Inst_Sbox_0_M21 ;
    wire SubBytesIns_Inst_Sbox_0_M20 ;
    wire SubBytesIns_Inst_Sbox_0_M19 ;
    wire SubBytesIns_Inst_Sbox_0_M18 ;
    wire SubBytesIns_Inst_Sbox_0_M17 ;
    wire SubBytesIns_Inst_Sbox_0_M16 ;
    wire SubBytesIns_Inst_Sbox_0_M15 ;
    wire SubBytesIns_Inst_Sbox_0_M14 ;
    wire SubBytesIns_Inst_Sbox_0_M13 ;
    wire SubBytesIns_Inst_Sbox_0_M12 ;
    wire SubBytesIns_Inst_Sbox_0_M11 ;
    wire SubBytesIns_Inst_Sbox_0_M10 ;
    wire SubBytesIns_Inst_Sbox_0_M9 ;
    wire SubBytesIns_Inst_Sbox_0_M8 ;
    wire SubBytesIns_Inst_Sbox_0_M7 ;
    wire SubBytesIns_Inst_Sbox_0_M6 ;
    wire SubBytesIns_Inst_Sbox_0_M5 ;
    wire SubBytesIns_Inst_Sbox_0_M4 ;
    wire SubBytesIns_Inst_Sbox_0_M3 ;
    wire SubBytesIns_Inst_Sbox_0_M2 ;
    wire SubBytesIns_Inst_Sbox_0_M1 ;
    wire SubBytesIns_Inst_Sbox_0_T27 ;
    wire SubBytesIns_Inst_Sbox_0_T26 ;
    wire SubBytesIns_Inst_Sbox_0_T25 ;
    wire SubBytesIns_Inst_Sbox_0_T24 ;
    wire SubBytesIns_Inst_Sbox_0_T23 ;
    wire SubBytesIns_Inst_Sbox_0_T22 ;
    wire SubBytesIns_Inst_Sbox_0_T21 ;
    wire SubBytesIns_Inst_Sbox_0_T20 ;
    wire SubBytesIns_Inst_Sbox_0_T19 ;
    wire SubBytesIns_Inst_Sbox_0_T18 ;
    wire SubBytesIns_Inst_Sbox_0_T17 ;
    wire SubBytesIns_Inst_Sbox_0_T16 ;
    wire SubBytesIns_Inst_Sbox_0_T15 ;
    wire SubBytesIns_Inst_Sbox_0_T14 ;
    wire SubBytesIns_Inst_Sbox_0_T13 ;
    wire SubBytesIns_Inst_Sbox_0_T12 ;
    wire SubBytesIns_Inst_Sbox_0_T11 ;
    wire SubBytesIns_Inst_Sbox_0_T10 ;
    wire SubBytesIns_Inst_Sbox_0_T9 ;
    wire SubBytesIns_Inst_Sbox_0_T8 ;
    wire SubBytesIns_Inst_Sbox_0_T7 ;
    wire SubBytesIns_Inst_Sbox_0_T6 ;
    wire SubBytesIns_Inst_Sbox_0_T5 ;
    wire SubBytesIns_Inst_Sbox_0_T4 ;
    wire SubBytesIns_Inst_Sbox_0_T3 ;
    wire SubBytesIns_Inst_Sbox_0_T2 ;
    wire SubBytesIns_Inst_Sbox_0_T1 ;
    wire SubBytesIns_Inst_Sbox_1_L29 ;
    wire SubBytesIns_Inst_Sbox_1_L28 ;
    wire SubBytesIns_Inst_Sbox_1_L27 ;
    wire SubBytesIns_Inst_Sbox_1_L26 ;
    wire SubBytesIns_Inst_Sbox_1_L25 ;
    wire SubBytesIns_Inst_Sbox_1_L24 ;
    wire SubBytesIns_Inst_Sbox_1_L23 ;
    wire SubBytesIns_Inst_Sbox_1_L22 ;
    wire SubBytesIns_Inst_Sbox_1_L21 ;
    wire SubBytesIns_Inst_Sbox_1_L20 ;
    wire SubBytesIns_Inst_Sbox_1_L19 ;
    wire SubBytesIns_Inst_Sbox_1_L18 ;
    wire SubBytesIns_Inst_Sbox_1_L17 ;
    wire SubBytesIns_Inst_Sbox_1_L16 ;
    wire SubBytesIns_Inst_Sbox_1_L15 ;
    wire SubBytesIns_Inst_Sbox_1_L14 ;
    wire SubBytesIns_Inst_Sbox_1_L13 ;
    wire SubBytesIns_Inst_Sbox_1_L12 ;
    wire SubBytesIns_Inst_Sbox_1_L11 ;
    wire SubBytesIns_Inst_Sbox_1_L10 ;
    wire SubBytesIns_Inst_Sbox_1_L9 ;
    wire SubBytesIns_Inst_Sbox_1_L8 ;
    wire SubBytesIns_Inst_Sbox_1_L7 ;
    wire SubBytesIns_Inst_Sbox_1_L6 ;
    wire SubBytesIns_Inst_Sbox_1_L5 ;
    wire SubBytesIns_Inst_Sbox_1_L4 ;
    wire SubBytesIns_Inst_Sbox_1_L3 ;
    wire SubBytesIns_Inst_Sbox_1_L2 ;
    wire SubBytesIns_Inst_Sbox_1_L1 ;
    wire SubBytesIns_Inst_Sbox_1_L0 ;
    wire SubBytesIns_Inst_Sbox_1_M63 ;
    wire SubBytesIns_Inst_Sbox_1_M62 ;
    wire SubBytesIns_Inst_Sbox_1_M61 ;
    wire SubBytesIns_Inst_Sbox_1_M60 ;
    wire SubBytesIns_Inst_Sbox_1_M59 ;
    wire SubBytesIns_Inst_Sbox_1_M58 ;
    wire SubBytesIns_Inst_Sbox_1_M57 ;
    wire SubBytesIns_Inst_Sbox_1_M56 ;
    wire SubBytesIns_Inst_Sbox_1_M55 ;
    wire SubBytesIns_Inst_Sbox_1_M54 ;
    wire SubBytesIns_Inst_Sbox_1_M53 ;
    wire SubBytesIns_Inst_Sbox_1_M52 ;
    wire SubBytesIns_Inst_Sbox_1_M51 ;
    wire SubBytesIns_Inst_Sbox_1_M50 ;
    wire SubBytesIns_Inst_Sbox_1_M49 ;
    wire SubBytesIns_Inst_Sbox_1_M48 ;
    wire SubBytesIns_Inst_Sbox_1_M47 ;
    wire SubBytesIns_Inst_Sbox_1_M46 ;
    wire SubBytesIns_Inst_Sbox_1_M45 ;
    wire SubBytesIns_Inst_Sbox_1_M44 ;
    wire SubBytesIns_Inst_Sbox_1_M43 ;
    wire SubBytesIns_Inst_Sbox_1_M42 ;
    wire SubBytesIns_Inst_Sbox_1_M41 ;
    wire SubBytesIns_Inst_Sbox_1_M40 ;
    wire SubBytesIns_Inst_Sbox_1_M39 ;
    wire SubBytesIns_Inst_Sbox_1_M38 ;
    wire SubBytesIns_Inst_Sbox_1_M37 ;
    wire SubBytesIns_Inst_Sbox_1_M36 ;
    wire SubBytesIns_Inst_Sbox_1_M35 ;
    wire SubBytesIns_Inst_Sbox_1_M34 ;
    wire SubBytesIns_Inst_Sbox_1_M33 ;
    wire SubBytesIns_Inst_Sbox_1_M32 ;
    wire SubBytesIns_Inst_Sbox_1_M31 ;
    wire SubBytesIns_Inst_Sbox_1_M30 ;
    wire SubBytesIns_Inst_Sbox_1_M29 ;
    wire SubBytesIns_Inst_Sbox_1_M28 ;
    wire SubBytesIns_Inst_Sbox_1_M27 ;
    wire SubBytesIns_Inst_Sbox_1_M26 ;
    wire SubBytesIns_Inst_Sbox_1_M25 ;
    wire SubBytesIns_Inst_Sbox_1_M24 ;
    wire SubBytesIns_Inst_Sbox_1_M23 ;
    wire SubBytesIns_Inst_Sbox_1_M22 ;
    wire SubBytesIns_Inst_Sbox_1_M21 ;
    wire SubBytesIns_Inst_Sbox_1_M20 ;
    wire SubBytesIns_Inst_Sbox_1_M19 ;
    wire SubBytesIns_Inst_Sbox_1_M18 ;
    wire SubBytesIns_Inst_Sbox_1_M17 ;
    wire SubBytesIns_Inst_Sbox_1_M16 ;
    wire SubBytesIns_Inst_Sbox_1_M15 ;
    wire SubBytesIns_Inst_Sbox_1_M14 ;
    wire SubBytesIns_Inst_Sbox_1_M13 ;
    wire SubBytesIns_Inst_Sbox_1_M12 ;
    wire SubBytesIns_Inst_Sbox_1_M11 ;
    wire SubBytesIns_Inst_Sbox_1_M10 ;
    wire SubBytesIns_Inst_Sbox_1_M9 ;
    wire SubBytesIns_Inst_Sbox_1_M8 ;
    wire SubBytesIns_Inst_Sbox_1_M7 ;
    wire SubBytesIns_Inst_Sbox_1_M6 ;
    wire SubBytesIns_Inst_Sbox_1_M5 ;
    wire SubBytesIns_Inst_Sbox_1_M4 ;
    wire SubBytesIns_Inst_Sbox_1_M3 ;
    wire SubBytesIns_Inst_Sbox_1_M2 ;
    wire SubBytesIns_Inst_Sbox_1_M1 ;
    wire SubBytesIns_Inst_Sbox_1_T27 ;
    wire SubBytesIns_Inst_Sbox_1_T26 ;
    wire SubBytesIns_Inst_Sbox_1_T25 ;
    wire SubBytesIns_Inst_Sbox_1_T24 ;
    wire SubBytesIns_Inst_Sbox_1_T23 ;
    wire SubBytesIns_Inst_Sbox_1_T22 ;
    wire SubBytesIns_Inst_Sbox_1_T21 ;
    wire SubBytesIns_Inst_Sbox_1_T20 ;
    wire SubBytesIns_Inst_Sbox_1_T19 ;
    wire SubBytesIns_Inst_Sbox_1_T18 ;
    wire SubBytesIns_Inst_Sbox_1_T17 ;
    wire SubBytesIns_Inst_Sbox_1_T16 ;
    wire SubBytesIns_Inst_Sbox_1_T15 ;
    wire SubBytesIns_Inst_Sbox_1_T14 ;
    wire SubBytesIns_Inst_Sbox_1_T13 ;
    wire SubBytesIns_Inst_Sbox_1_T12 ;
    wire SubBytesIns_Inst_Sbox_1_T11 ;
    wire SubBytesIns_Inst_Sbox_1_T10 ;
    wire SubBytesIns_Inst_Sbox_1_T9 ;
    wire SubBytesIns_Inst_Sbox_1_T8 ;
    wire SubBytesIns_Inst_Sbox_1_T7 ;
    wire SubBytesIns_Inst_Sbox_1_T6 ;
    wire SubBytesIns_Inst_Sbox_1_T5 ;
    wire SubBytesIns_Inst_Sbox_1_T4 ;
    wire SubBytesIns_Inst_Sbox_1_T3 ;
    wire SubBytesIns_Inst_Sbox_1_T2 ;
    wire SubBytesIns_Inst_Sbox_1_T1 ;
    wire SubBytesIns_Inst_Sbox_2_L29 ;
    wire SubBytesIns_Inst_Sbox_2_L28 ;
    wire SubBytesIns_Inst_Sbox_2_L27 ;
    wire SubBytesIns_Inst_Sbox_2_L26 ;
    wire SubBytesIns_Inst_Sbox_2_L25 ;
    wire SubBytesIns_Inst_Sbox_2_L24 ;
    wire SubBytesIns_Inst_Sbox_2_L23 ;
    wire SubBytesIns_Inst_Sbox_2_L22 ;
    wire SubBytesIns_Inst_Sbox_2_L21 ;
    wire SubBytesIns_Inst_Sbox_2_L20 ;
    wire SubBytesIns_Inst_Sbox_2_L19 ;
    wire SubBytesIns_Inst_Sbox_2_L18 ;
    wire SubBytesIns_Inst_Sbox_2_L17 ;
    wire SubBytesIns_Inst_Sbox_2_L16 ;
    wire SubBytesIns_Inst_Sbox_2_L15 ;
    wire SubBytesIns_Inst_Sbox_2_L14 ;
    wire SubBytesIns_Inst_Sbox_2_L13 ;
    wire SubBytesIns_Inst_Sbox_2_L12 ;
    wire SubBytesIns_Inst_Sbox_2_L11 ;
    wire SubBytesIns_Inst_Sbox_2_L10 ;
    wire SubBytesIns_Inst_Sbox_2_L9 ;
    wire SubBytesIns_Inst_Sbox_2_L8 ;
    wire SubBytesIns_Inst_Sbox_2_L7 ;
    wire SubBytesIns_Inst_Sbox_2_L6 ;
    wire SubBytesIns_Inst_Sbox_2_L5 ;
    wire SubBytesIns_Inst_Sbox_2_L4 ;
    wire SubBytesIns_Inst_Sbox_2_L3 ;
    wire SubBytesIns_Inst_Sbox_2_L2 ;
    wire SubBytesIns_Inst_Sbox_2_L1 ;
    wire SubBytesIns_Inst_Sbox_2_L0 ;
    wire SubBytesIns_Inst_Sbox_2_M63 ;
    wire SubBytesIns_Inst_Sbox_2_M62 ;
    wire SubBytesIns_Inst_Sbox_2_M61 ;
    wire SubBytesIns_Inst_Sbox_2_M60 ;
    wire SubBytesIns_Inst_Sbox_2_M59 ;
    wire SubBytesIns_Inst_Sbox_2_M58 ;
    wire SubBytesIns_Inst_Sbox_2_M57 ;
    wire SubBytesIns_Inst_Sbox_2_M56 ;
    wire SubBytesIns_Inst_Sbox_2_M55 ;
    wire SubBytesIns_Inst_Sbox_2_M54 ;
    wire SubBytesIns_Inst_Sbox_2_M53 ;
    wire SubBytesIns_Inst_Sbox_2_M52 ;
    wire SubBytesIns_Inst_Sbox_2_M51 ;
    wire SubBytesIns_Inst_Sbox_2_M50 ;
    wire SubBytesIns_Inst_Sbox_2_M49 ;
    wire SubBytesIns_Inst_Sbox_2_M48 ;
    wire SubBytesIns_Inst_Sbox_2_M47 ;
    wire SubBytesIns_Inst_Sbox_2_M46 ;
    wire SubBytesIns_Inst_Sbox_2_M45 ;
    wire SubBytesIns_Inst_Sbox_2_M44 ;
    wire SubBytesIns_Inst_Sbox_2_M43 ;
    wire SubBytesIns_Inst_Sbox_2_M42 ;
    wire SubBytesIns_Inst_Sbox_2_M41 ;
    wire SubBytesIns_Inst_Sbox_2_M40 ;
    wire SubBytesIns_Inst_Sbox_2_M39 ;
    wire SubBytesIns_Inst_Sbox_2_M38 ;
    wire SubBytesIns_Inst_Sbox_2_M37 ;
    wire SubBytesIns_Inst_Sbox_2_M36 ;
    wire SubBytesIns_Inst_Sbox_2_M35 ;
    wire SubBytesIns_Inst_Sbox_2_M34 ;
    wire SubBytesIns_Inst_Sbox_2_M33 ;
    wire SubBytesIns_Inst_Sbox_2_M32 ;
    wire SubBytesIns_Inst_Sbox_2_M31 ;
    wire SubBytesIns_Inst_Sbox_2_M30 ;
    wire SubBytesIns_Inst_Sbox_2_M29 ;
    wire SubBytesIns_Inst_Sbox_2_M28 ;
    wire SubBytesIns_Inst_Sbox_2_M27 ;
    wire SubBytesIns_Inst_Sbox_2_M26 ;
    wire SubBytesIns_Inst_Sbox_2_M25 ;
    wire SubBytesIns_Inst_Sbox_2_M24 ;
    wire SubBytesIns_Inst_Sbox_2_M23 ;
    wire SubBytesIns_Inst_Sbox_2_M22 ;
    wire SubBytesIns_Inst_Sbox_2_M21 ;
    wire SubBytesIns_Inst_Sbox_2_M20 ;
    wire SubBytesIns_Inst_Sbox_2_M19 ;
    wire SubBytesIns_Inst_Sbox_2_M18 ;
    wire SubBytesIns_Inst_Sbox_2_M17 ;
    wire SubBytesIns_Inst_Sbox_2_M16 ;
    wire SubBytesIns_Inst_Sbox_2_M15 ;
    wire SubBytesIns_Inst_Sbox_2_M14 ;
    wire SubBytesIns_Inst_Sbox_2_M13 ;
    wire SubBytesIns_Inst_Sbox_2_M12 ;
    wire SubBytesIns_Inst_Sbox_2_M11 ;
    wire SubBytesIns_Inst_Sbox_2_M10 ;
    wire SubBytesIns_Inst_Sbox_2_M9 ;
    wire SubBytesIns_Inst_Sbox_2_M8 ;
    wire SubBytesIns_Inst_Sbox_2_M7 ;
    wire SubBytesIns_Inst_Sbox_2_M6 ;
    wire SubBytesIns_Inst_Sbox_2_M5 ;
    wire SubBytesIns_Inst_Sbox_2_M4 ;
    wire SubBytesIns_Inst_Sbox_2_M3 ;
    wire SubBytesIns_Inst_Sbox_2_M2 ;
    wire SubBytesIns_Inst_Sbox_2_M1 ;
    wire SubBytesIns_Inst_Sbox_2_T27 ;
    wire SubBytesIns_Inst_Sbox_2_T26 ;
    wire SubBytesIns_Inst_Sbox_2_T25 ;
    wire SubBytesIns_Inst_Sbox_2_T24 ;
    wire SubBytesIns_Inst_Sbox_2_T23 ;
    wire SubBytesIns_Inst_Sbox_2_T22 ;
    wire SubBytesIns_Inst_Sbox_2_T21 ;
    wire SubBytesIns_Inst_Sbox_2_T20 ;
    wire SubBytesIns_Inst_Sbox_2_T19 ;
    wire SubBytesIns_Inst_Sbox_2_T18 ;
    wire SubBytesIns_Inst_Sbox_2_T17 ;
    wire SubBytesIns_Inst_Sbox_2_T16 ;
    wire SubBytesIns_Inst_Sbox_2_T15 ;
    wire SubBytesIns_Inst_Sbox_2_T14 ;
    wire SubBytesIns_Inst_Sbox_2_T13 ;
    wire SubBytesIns_Inst_Sbox_2_T12 ;
    wire SubBytesIns_Inst_Sbox_2_T11 ;
    wire SubBytesIns_Inst_Sbox_2_T10 ;
    wire SubBytesIns_Inst_Sbox_2_T9 ;
    wire SubBytesIns_Inst_Sbox_2_T8 ;
    wire SubBytesIns_Inst_Sbox_2_T7 ;
    wire SubBytesIns_Inst_Sbox_2_T6 ;
    wire SubBytesIns_Inst_Sbox_2_T5 ;
    wire SubBytesIns_Inst_Sbox_2_T4 ;
    wire SubBytesIns_Inst_Sbox_2_T3 ;
    wire SubBytesIns_Inst_Sbox_2_T2 ;
    wire SubBytesIns_Inst_Sbox_2_T1 ;
    wire SubBytesIns_Inst_Sbox_3_L29 ;
    wire SubBytesIns_Inst_Sbox_3_L28 ;
    wire SubBytesIns_Inst_Sbox_3_L27 ;
    wire SubBytesIns_Inst_Sbox_3_L26 ;
    wire SubBytesIns_Inst_Sbox_3_L25 ;
    wire SubBytesIns_Inst_Sbox_3_L24 ;
    wire SubBytesIns_Inst_Sbox_3_L23 ;
    wire SubBytesIns_Inst_Sbox_3_L22 ;
    wire SubBytesIns_Inst_Sbox_3_L21 ;
    wire SubBytesIns_Inst_Sbox_3_L20 ;
    wire SubBytesIns_Inst_Sbox_3_L19 ;
    wire SubBytesIns_Inst_Sbox_3_L18 ;
    wire SubBytesIns_Inst_Sbox_3_L17 ;
    wire SubBytesIns_Inst_Sbox_3_L16 ;
    wire SubBytesIns_Inst_Sbox_3_L15 ;
    wire SubBytesIns_Inst_Sbox_3_L14 ;
    wire SubBytesIns_Inst_Sbox_3_L13 ;
    wire SubBytesIns_Inst_Sbox_3_L12 ;
    wire SubBytesIns_Inst_Sbox_3_L11 ;
    wire SubBytesIns_Inst_Sbox_3_L10 ;
    wire SubBytesIns_Inst_Sbox_3_L9 ;
    wire SubBytesIns_Inst_Sbox_3_L8 ;
    wire SubBytesIns_Inst_Sbox_3_L7 ;
    wire SubBytesIns_Inst_Sbox_3_L6 ;
    wire SubBytesIns_Inst_Sbox_3_L5 ;
    wire SubBytesIns_Inst_Sbox_3_L4 ;
    wire SubBytesIns_Inst_Sbox_3_L3 ;
    wire SubBytesIns_Inst_Sbox_3_L2 ;
    wire SubBytesIns_Inst_Sbox_3_L1 ;
    wire SubBytesIns_Inst_Sbox_3_L0 ;
    wire SubBytesIns_Inst_Sbox_3_M63 ;
    wire SubBytesIns_Inst_Sbox_3_M62 ;
    wire SubBytesIns_Inst_Sbox_3_M61 ;
    wire SubBytesIns_Inst_Sbox_3_M60 ;
    wire SubBytesIns_Inst_Sbox_3_M59 ;
    wire SubBytesIns_Inst_Sbox_3_M58 ;
    wire SubBytesIns_Inst_Sbox_3_M57 ;
    wire SubBytesIns_Inst_Sbox_3_M56 ;
    wire SubBytesIns_Inst_Sbox_3_M55 ;
    wire SubBytesIns_Inst_Sbox_3_M54 ;
    wire SubBytesIns_Inst_Sbox_3_M53 ;
    wire SubBytesIns_Inst_Sbox_3_M52 ;
    wire SubBytesIns_Inst_Sbox_3_M51 ;
    wire SubBytesIns_Inst_Sbox_3_M50 ;
    wire SubBytesIns_Inst_Sbox_3_M49 ;
    wire SubBytesIns_Inst_Sbox_3_M48 ;
    wire SubBytesIns_Inst_Sbox_3_M47 ;
    wire SubBytesIns_Inst_Sbox_3_M46 ;
    wire SubBytesIns_Inst_Sbox_3_M45 ;
    wire SubBytesIns_Inst_Sbox_3_M44 ;
    wire SubBytesIns_Inst_Sbox_3_M43 ;
    wire SubBytesIns_Inst_Sbox_3_M42 ;
    wire SubBytesIns_Inst_Sbox_3_M41 ;
    wire SubBytesIns_Inst_Sbox_3_M40 ;
    wire SubBytesIns_Inst_Sbox_3_M39 ;
    wire SubBytesIns_Inst_Sbox_3_M38 ;
    wire SubBytesIns_Inst_Sbox_3_M37 ;
    wire SubBytesIns_Inst_Sbox_3_M36 ;
    wire SubBytesIns_Inst_Sbox_3_M35 ;
    wire SubBytesIns_Inst_Sbox_3_M34 ;
    wire SubBytesIns_Inst_Sbox_3_M33 ;
    wire SubBytesIns_Inst_Sbox_3_M32 ;
    wire SubBytesIns_Inst_Sbox_3_M31 ;
    wire SubBytesIns_Inst_Sbox_3_M30 ;
    wire SubBytesIns_Inst_Sbox_3_M29 ;
    wire SubBytesIns_Inst_Sbox_3_M28 ;
    wire SubBytesIns_Inst_Sbox_3_M27 ;
    wire SubBytesIns_Inst_Sbox_3_M26 ;
    wire SubBytesIns_Inst_Sbox_3_M25 ;
    wire SubBytesIns_Inst_Sbox_3_M24 ;
    wire SubBytesIns_Inst_Sbox_3_M23 ;
    wire SubBytesIns_Inst_Sbox_3_M22 ;
    wire SubBytesIns_Inst_Sbox_3_M21 ;
    wire SubBytesIns_Inst_Sbox_3_M20 ;
    wire SubBytesIns_Inst_Sbox_3_M19 ;
    wire SubBytesIns_Inst_Sbox_3_M18 ;
    wire SubBytesIns_Inst_Sbox_3_M17 ;
    wire SubBytesIns_Inst_Sbox_3_M16 ;
    wire SubBytesIns_Inst_Sbox_3_M15 ;
    wire SubBytesIns_Inst_Sbox_3_M14 ;
    wire SubBytesIns_Inst_Sbox_3_M13 ;
    wire SubBytesIns_Inst_Sbox_3_M12 ;
    wire SubBytesIns_Inst_Sbox_3_M11 ;
    wire SubBytesIns_Inst_Sbox_3_M10 ;
    wire SubBytesIns_Inst_Sbox_3_M9 ;
    wire SubBytesIns_Inst_Sbox_3_M8 ;
    wire SubBytesIns_Inst_Sbox_3_M7 ;
    wire SubBytesIns_Inst_Sbox_3_M6 ;
    wire SubBytesIns_Inst_Sbox_3_M5 ;
    wire SubBytesIns_Inst_Sbox_3_M4 ;
    wire SubBytesIns_Inst_Sbox_3_M3 ;
    wire SubBytesIns_Inst_Sbox_3_M2 ;
    wire SubBytesIns_Inst_Sbox_3_M1 ;
    wire SubBytesIns_Inst_Sbox_3_T27 ;
    wire SubBytesIns_Inst_Sbox_3_T26 ;
    wire SubBytesIns_Inst_Sbox_3_T25 ;
    wire SubBytesIns_Inst_Sbox_3_T24 ;
    wire SubBytesIns_Inst_Sbox_3_T23 ;
    wire SubBytesIns_Inst_Sbox_3_T22 ;
    wire SubBytesIns_Inst_Sbox_3_T21 ;
    wire SubBytesIns_Inst_Sbox_3_T20 ;
    wire SubBytesIns_Inst_Sbox_3_T19 ;
    wire SubBytesIns_Inst_Sbox_3_T18 ;
    wire SubBytesIns_Inst_Sbox_3_T17 ;
    wire SubBytesIns_Inst_Sbox_3_T16 ;
    wire SubBytesIns_Inst_Sbox_3_T15 ;
    wire SubBytesIns_Inst_Sbox_3_T14 ;
    wire SubBytesIns_Inst_Sbox_3_T13 ;
    wire SubBytesIns_Inst_Sbox_3_T12 ;
    wire SubBytesIns_Inst_Sbox_3_T11 ;
    wire SubBytesIns_Inst_Sbox_3_T10 ;
    wire SubBytesIns_Inst_Sbox_3_T9 ;
    wire SubBytesIns_Inst_Sbox_3_T8 ;
    wire SubBytesIns_Inst_Sbox_3_T7 ;
    wire SubBytesIns_Inst_Sbox_3_T6 ;
    wire SubBytesIns_Inst_Sbox_3_T5 ;
    wire SubBytesIns_Inst_Sbox_3_T4 ;
    wire SubBytesIns_Inst_Sbox_3_T3 ;
    wire SubBytesIns_Inst_Sbox_3_T2 ;
    wire SubBytesIns_Inst_Sbox_3_T1 ;
    wire SubBytesIns_Inst_Sbox_4_L29 ;
    wire SubBytesIns_Inst_Sbox_4_L28 ;
    wire SubBytesIns_Inst_Sbox_4_L27 ;
    wire SubBytesIns_Inst_Sbox_4_L26 ;
    wire SubBytesIns_Inst_Sbox_4_L25 ;
    wire SubBytesIns_Inst_Sbox_4_L24 ;
    wire SubBytesIns_Inst_Sbox_4_L23 ;
    wire SubBytesIns_Inst_Sbox_4_L22 ;
    wire SubBytesIns_Inst_Sbox_4_L21 ;
    wire SubBytesIns_Inst_Sbox_4_L20 ;
    wire SubBytesIns_Inst_Sbox_4_L19 ;
    wire SubBytesIns_Inst_Sbox_4_L18 ;
    wire SubBytesIns_Inst_Sbox_4_L17 ;
    wire SubBytesIns_Inst_Sbox_4_L16 ;
    wire SubBytesIns_Inst_Sbox_4_L15 ;
    wire SubBytesIns_Inst_Sbox_4_L14 ;
    wire SubBytesIns_Inst_Sbox_4_L13 ;
    wire SubBytesIns_Inst_Sbox_4_L12 ;
    wire SubBytesIns_Inst_Sbox_4_L11 ;
    wire SubBytesIns_Inst_Sbox_4_L10 ;
    wire SubBytesIns_Inst_Sbox_4_L9 ;
    wire SubBytesIns_Inst_Sbox_4_L8 ;
    wire SubBytesIns_Inst_Sbox_4_L7 ;
    wire SubBytesIns_Inst_Sbox_4_L6 ;
    wire SubBytesIns_Inst_Sbox_4_L5 ;
    wire SubBytesIns_Inst_Sbox_4_L4 ;
    wire SubBytesIns_Inst_Sbox_4_L3 ;
    wire SubBytesIns_Inst_Sbox_4_L2 ;
    wire SubBytesIns_Inst_Sbox_4_L1 ;
    wire SubBytesIns_Inst_Sbox_4_L0 ;
    wire SubBytesIns_Inst_Sbox_4_M63 ;
    wire SubBytesIns_Inst_Sbox_4_M62 ;
    wire SubBytesIns_Inst_Sbox_4_M61 ;
    wire SubBytesIns_Inst_Sbox_4_M60 ;
    wire SubBytesIns_Inst_Sbox_4_M59 ;
    wire SubBytesIns_Inst_Sbox_4_M58 ;
    wire SubBytesIns_Inst_Sbox_4_M57 ;
    wire SubBytesIns_Inst_Sbox_4_M56 ;
    wire SubBytesIns_Inst_Sbox_4_M55 ;
    wire SubBytesIns_Inst_Sbox_4_M54 ;
    wire SubBytesIns_Inst_Sbox_4_M53 ;
    wire SubBytesIns_Inst_Sbox_4_M52 ;
    wire SubBytesIns_Inst_Sbox_4_M51 ;
    wire SubBytesIns_Inst_Sbox_4_M50 ;
    wire SubBytesIns_Inst_Sbox_4_M49 ;
    wire SubBytesIns_Inst_Sbox_4_M48 ;
    wire SubBytesIns_Inst_Sbox_4_M47 ;
    wire SubBytesIns_Inst_Sbox_4_M46 ;
    wire SubBytesIns_Inst_Sbox_4_M45 ;
    wire SubBytesIns_Inst_Sbox_4_M44 ;
    wire SubBytesIns_Inst_Sbox_4_M43 ;
    wire SubBytesIns_Inst_Sbox_4_M42 ;
    wire SubBytesIns_Inst_Sbox_4_M41 ;
    wire SubBytesIns_Inst_Sbox_4_M40 ;
    wire SubBytesIns_Inst_Sbox_4_M39 ;
    wire SubBytesIns_Inst_Sbox_4_M38 ;
    wire SubBytesIns_Inst_Sbox_4_M37 ;
    wire SubBytesIns_Inst_Sbox_4_M36 ;
    wire SubBytesIns_Inst_Sbox_4_M35 ;
    wire SubBytesIns_Inst_Sbox_4_M34 ;
    wire SubBytesIns_Inst_Sbox_4_M33 ;
    wire SubBytesIns_Inst_Sbox_4_M32 ;
    wire SubBytesIns_Inst_Sbox_4_M31 ;
    wire SubBytesIns_Inst_Sbox_4_M30 ;
    wire SubBytesIns_Inst_Sbox_4_M29 ;
    wire SubBytesIns_Inst_Sbox_4_M28 ;
    wire SubBytesIns_Inst_Sbox_4_M27 ;
    wire SubBytesIns_Inst_Sbox_4_M26 ;
    wire SubBytesIns_Inst_Sbox_4_M25 ;
    wire SubBytesIns_Inst_Sbox_4_M24 ;
    wire SubBytesIns_Inst_Sbox_4_M23 ;
    wire SubBytesIns_Inst_Sbox_4_M22 ;
    wire SubBytesIns_Inst_Sbox_4_M21 ;
    wire SubBytesIns_Inst_Sbox_4_M20 ;
    wire SubBytesIns_Inst_Sbox_4_M19 ;
    wire SubBytesIns_Inst_Sbox_4_M18 ;
    wire SubBytesIns_Inst_Sbox_4_M17 ;
    wire SubBytesIns_Inst_Sbox_4_M16 ;
    wire SubBytesIns_Inst_Sbox_4_M15 ;
    wire SubBytesIns_Inst_Sbox_4_M14 ;
    wire SubBytesIns_Inst_Sbox_4_M13 ;
    wire SubBytesIns_Inst_Sbox_4_M12 ;
    wire SubBytesIns_Inst_Sbox_4_M11 ;
    wire SubBytesIns_Inst_Sbox_4_M10 ;
    wire SubBytesIns_Inst_Sbox_4_M9 ;
    wire SubBytesIns_Inst_Sbox_4_M8 ;
    wire SubBytesIns_Inst_Sbox_4_M7 ;
    wire SubBytesIns_Inst_Sbox_4_M6 ;
    wire SubBytesIns_Inst_Sbox_4_M5 ;
    wire SubBytesIns_Inst_Sbox_4_M4 ;
    wire SubBytesIns_Inst_Sbox_4_M3 ;
    wire SubBytesIns_Inst_Sbox_4_M2 ;
    wire SubBytesIns_Inst_Sbox_4_M1 ;
    wire SubBytesIns_Inst_Sbox_4_T27 ;
    wire SubBytesIns_Inst_Sbox_4_T26 ;
    wire SubBytesIns_Inst_Sbox_4_T25 ;
    wire SubBytesIns_Inst_Sbox_4_T24 ;
    wire SubBytesIns_Inst_Sbox_4_T23 ;
    wire SubBytesIns_Inst_Sbox_4_T22 ;
    wire SubBytesIns_Inst_Sbox_4_T21 ;
    wire SubBytesIns_Inst_Sbox_4_T20 ;
    wire SubBytesIns_Inst_Sbox_4_T19 ;
    wire SubBytesIns_Inst_Sbox_4_T18 ;
    wire SubBytesIns_Inst_Sbox_4_T17 ;
    wire SubBytesIns_Inst_Sbox_4_T16 ;
    wire SubBytesIns_Inst_Sbox_4_T15 ;
    wire SubBytesIns_Inst_Sbox_4_T14 ;
    wire SubBytesIns_Inst_Sbox_4_T13 ;
    wire SubBytesIns_Inst_Sbox_4_T12 ;
    wire SubBytesIns_Inst_Sbox_4_T11 ;
    wire SubBytesIns_Inst_Sbox_4_T10 ;
    wire SubBytesIns_Inst_Sbox_4_T9 ;
    wire SubBytesIns_Inst_Sbox_4_T8 ;
    wire SubBytesIns_Inst_Sbox_4_T7 ;
    wire SubBytesIns_Inst_Sbox_4_T6 ;
    wire SubBytesIns_Inst_Sbox_4_T5 ;
    wire SubBytesIns_Inst_Sbox_4_T4 ;
    wire SubBytesIns_Inst_Sbox_4_T3 ;
    wire SubBytesIns_Inst_Sbox_4_T2 ;
    wire SubBytesIns_Inst_Sbox_4_T1 ;
    wire SubBytesIns_Inst_Sbox_5_L29 ;
    wire SubBytesIns_Inst_Sbox_5_L28 ;
    wire SubBytesIns_Inst_Sbox_5_L27 ;
    wire SubBytesIns_Inst_Sbox_5_L26 ;
    wire SubBytesIns_Inst_Sbox_5_L25 ;
    wire SubBytesIns_Inst_Sbox_5_L24 ;
    wire SubBytesIns_Inst_Sbox_5_L23 ;
    wire SubBytesIns_Inst_Sbox_5_L22 ;
    wire SubBytesIns_Inst_Sbox_5_L21 ;
    wire SubBytesIns_Inst_Sbox_5_L20 ;
    wire SubBytesIns_Inst_Sbox_5_L19 ;
    wire SubBytesIns_Inst_Sbox_5_L18 ;
    wire SubBytesIns_Inst_Sbox_5_L17 ;
    wire SubBytesIns_Inst_Sbox_5_L16 ;
    wire SubBytesIns_Inst_Sbox_5_L15 ;
    wire SubBytesIns_Inst_Sbox_5_L14 ;
    wire SubBytesIns_Inst_Sbox_5_L13 ;
    wire SubBytesIns_Inst_Sbox_5_L12 ;
    wire SubBytesIns_Inst_Sbox_5_L11 ;
    wire SubBytesIns_Inst_Sbox_5_L10 ;
    wire SubBytesIns_Inst_Sbox_5_L9 ;
    wire SubBytesIns_Inst_Sbox_5_L8 ;
    wire SubBytesIns_Inst_Sbox_5_L7 ;
    wire SubBytesIns_Inst_Sbox_5_L6 ;
    wire SubBytesIns_Inst_Sbox_5_L5 ;
    wire SubBytesIns_Inst_Sbox_5_L4 ;
    wire SubBytesIns_Inst_Sbox_5_L3 ;
    wire SubBytesIns_Inst_Sbox_5_L2 ;
    wire SubBytesIns_Inst_Sbox_5_L1 ;
    wire SubBytesIns_Inst_Sbox_5_L0 ;
    wire SubBytesIns_Inst_Sbox_5_M63 ;
    wire SubBytesIns_Inst_Sbox_5_M62 ;
    wire SubBytesIns_Inst_Sbox_5_M61 ;
    wire SubBytesIns_Inst_Sbox_5_M60 ;
    wire SubBytesIns_Inst_Sbox_5_M59 ;
    wire SubBytesIns_Inst_Sbox_5_M58 ;
    wire SubBytesIns_Inst_Sbox_5_M57 ;
    wire SubBytesIns_Inst_Sbox_5_M56 ;
    wire SubBytesIns_Inst_Sbox_5_M55 ;
    wire SubBytesIns_Inst_Sbox_5_M54 ;
    wire SubBytesIns_Inst_Sbox_5_M53 ;
    wire SubBytesIns_Inst_Sbox_5_M52 ;
    wire SubBytesIns_Inst_Sbox_5_M51 ;
    wire SubBytesIns_Inst_Sbox_5_M50 ;
    wire SubBytesIns_Inst_Sbox_5_M49 ;
    wire SubBytesIns_Inst_Sbox_5_M48 ;
    wire SubBytesIns_Inst_Sbox_5_M47 ;
    wire SubBytesIns_Inst_Sbox_5_M46 ;
    wire SubBytesIns_Inst_Sbox_5_M45 ;
    wire SubBytesIns_Inst_Sbox_5_M44 ;
    wire SubBytesIns_Inst_Sbox_5_M43 ;
    wire SubBytesIns_Inst_Sbox_5_M42 ;
    wire SubBytesIns_Inst_Sbox_5_M41 ;
    wire SubBytesIns_Inst_Sbox_5_M40 ;
    wire SubBytesIns_Inst_Sbox_5_M39 ;
    wire SubBytesIns_Inst_Sbox_5_M38 ;
    wire SubBytesIns_Inst_Sbox_5_M37 ;
    wire SubBytesIns_Inst_Sbox_5_M36 ;
    wire SubBytesIns_Inst_Sbox_5_M35 ;
    wire SubBytesIns_Inst_Sbox_5_M34 ;
    wire SubBytesIns_Inst_Sbox_5_M33 ;
    wire SubBytesIns_Inst_Sbox_5_M32 ;
    wire SubBytesIns_Inst_Sbox_5_M31 ;
    wire SubBytesIns_Inst_Sbox_5_M30 ;
    wire SubBytesIns_Inst_Sbox_5_M29 ;
    wire SubBytesIns_Inst_Sbox_5_M28 ;
    wire SubBytesIns_Inst_Sbox_5_M27 ;
    wire SubBytesIns_Inst_Sbox_5_M26 ;
    wire SubBytesIns_Inst_Sbox_5_M25 ;
    wire SubBytesIns_Inst_Sbox_5_M24 ;
    wire SubBytesIns_Inst_Sbox_5_M23 ;
    wire SubBytesIns_Inst_Sbox_5_M22 ;
    wire SubBytesIns_Inst_Sbox_5_M21 ;
    wire SubBytesIns_Inst_Sbox_5_M20 ;
    wire SubBytesIns_Inst_Sbox_5_M19 ;
    wire SubBytesIns_Inst_Sbox_5_M18 ;
    wire SubBytesIns_Inst_Sbox_5_M17 ;
    wire SubBytesIns_Inst_Sbox_5_M16 ;
    wire SubBytesIns_Inst_Sbox_5_M15 ;
    wire SubBytesIns_Inst_Sbox_5_M14 ;
    wire SubBytesIns_Inst_Sbox_5_M13 ;
    wire SubBytesIns_Inst_Sbox_5_M12 ;
    wire SubBytesIns_Inst_Sbox_5_M11 ;
    wire SubBytesIns_Inst_Sbox_5_M10 ;
    wire SubBytesIns_Inst_Sbox_5_M9 ;
    wire SubBytesIns_Inst_Sbox_5_M8 ;
    wire SubBytesIns_Inst_Sbox_5_M7 ;
    wire SubBytesIns_Inst_Sbox_5_M6 ;
    wire SubBytesIns_Inst_Sbox_5_M5 ;
    wire SubBytesIns_Inst_Sbox_5_M4 ;
    wire SubBytesIns_Inst_Sbox_5_M3 ;
    wire SubBytesIns_Inst_Sbox_5_M2 ;
    wire SubBytesIns_Inst_Sbox_5_M1 ;
    wire SubBytesIns_Inst_Sbox_5_T27 ;
    wire SubBytesIns_Inst_Sbox_5_T26 ;
    wire SubBytesIns_Inst_Sbox_5_T25 ;
    wire SubBytesIns_Inst_Sbox_5_T24 ;
    wire SubBytesIns_Inst_Sbox_5_T23 ;
    wire SubBytesIns_Inst_Sbox_5_T22 ;
    wire SubBytesIns_Inst_Sbox_5_T21 ;
    wire SubBytesIns_Inst_Sbox_5_T20 ;
    wire SubBytesIns_Inst_Sbox_5_T19 ;
    wire SubBytesIns_Inst_Sbox_5_T18 ;
    wire SubBytesIns_Inst_Sbox_5_T17 ;
    wire SubBytesIns_Inst_Sbox_5_T16 ;
    wire SubBytesIns_Inst_Sbox_5_T15 ;
    wire SubBytesIns_Inst_Sbox_5_T14 ;
    wire SubBytesIns_Inst_Sbox_5_T13 ;
    wire SubBytesIns_Inst_Sbox_5_T12 ;
    wire SubBytesIns_Inst_Sbox_5_T11 ;
    wire SubBytesIns_Inst_Sbox_5_T10 ;
    wire SubBytesIns_Inst_Sbox_5_T9 ;
    wire SubBytesIns_Inst_Sbox_5_T8 ;
    wire SubBytesIns_Inst_Sbox_5_T7 ;
    wire SubBytesIns_Inst_Sbox_5_T6 ;
    wire SubBytesIns_Inst_Sbox_5_T5 ;
    wire SubBytesIns_Inst_Sbox_5_T4 ;
    wire SubBytesIns_Inst_Sbox_5_T3 ;
    wire SubBytesIns_Inst_Sbox_5_T2 ;
    wire SubBytesIns_Inst_Sbox_5_T1 ;
    wire SubBytesIns_Inst_Sbox_6_L29 ;
    wire SubBytesIns_Inst_Sbox_6_L28 ;
    wire SubBytesIns_Inst_Sbox_6_L27 ;
    wire SubBytesIns_Inst_Sbox_6_L26 ;
    wire SubBytesIns_Inst_Sbox_6_L25 ;
    wire SubBytesIns_Inst_Sbox_6_L24 ;
    wire SubBytesIns_Inst_Sbox_6_L23 ;
    wire SubBytesIns_Inst_Sbox_6_L22 ;
    wire SubBytesIns_Inst_Sbox_6_L21 ;
    wire SubBytesIns_Inst_Sbox_6_L20 ;
    wire SubBytesIns_Inst_Sbox_6_L19 ;
    wire SubBytesIns_Inst_Sbox_6_L18 ;
    wire SubBytesIns_Inst_Sbox_6_L17 ;
    wire SubBytesIns_Inst_Sbox_6_L16 ;
    wire SubBytesIns_Inst_Sbox_6_L15 ;
    wire SubBytesIns_Inst_Sbox_6_L14 ;
    wire SubBytesIns_Inst_Sbox_6_L13 ;
    wire SubBytesIns_Inst_Sbox_6_L12 ;
    wire SubBytesIns_Inst_Sbox_6_L11 ;
    wire SubBytesIns_Inst_Sbox_6_L10 ;
    wire SubBytesIns_Inst_Sbox_6_L9 ;
    wire SubBytesIns_Inst_Sbox_6_L8 ;
    wire SubBytesIns_Inst_Sbox_6_L7 ;
    wire SubBytesIns_Inst_Sbox_6_L6 ;
    wire SubBytesIns_Inst_Sbox_6_L5 ;
    wire SubBytesIns_Inst_Sbox_6_L4 ;
    wire SubBytesIns_Inst_Sbox_6_L3 ;
    wire SubBytesIns_Inst_Sbox_6_L2 ;
    wire SubBytesIns_Inst_Sbox_6_L1 ;
    wire SubBytesIns_Inst_Sbox_6_L0 ;
    wire SubBytesIns_Inst_Sbox_6_M63 ;
    wire SubBytesIns_Inst_Sbox_6_M62 ;
    wire SubBytesIns_Inst_Sbox_6_M61 ;
    wire SubBytesIns_Inst_Sbox_6_M60 ;
    wire SubBytesIns_Inst_Sbox_6_M59 ;
    wire SubBytesIns_Inst_Sbox_6_M58 ;
    wire SubBytesIns_Inst_Sbox_6_M57 ;
    wire SubBytesIns_Inst_Sbox_6_M56 ;
    wire SubBytesIns_Inst_Sbox_6_M55 ;
    wire SubBytesIns_Inst_Sbox_6_M54 ;
    wire SubBytesIns_Inst_Sbox_6_M53 ;
    wire SubBytesIns_Inst_Sbox_6_M52 ;
    wire SubBytesIns_Inst_Sbox_6_M51 ;
    wire SubBytesIns_Inst_Sbox_6_M50 ;
    wire SubBytesIns_Inst_Sbox_6_M49 ;
    wire SubBytesIns_Inst_Sbox_6_M48 ;
    wire SubBytesIns_Inst_Sbox_6_M47 ;
    wire SubBytesIns_Inst_Sbox_6_M46 ;
    wire SubBytesIns_Inst_Sbox_6_M45 ;
    wire SubBytesIns_Inst_Sbox_6_M44 ;
    wire SubBytesIns_Inst_Sbox_6_M43 ;
    wire SubBytesIns_Inst_Sbox_6_M42 ;
    wire SubBytesIns_Inst_Sbox_6_M41 ;
    wire SubBytesIns_Inst_Sbox_6_M40 ;
    wire SubBytesIns_Inst_Sbox_6_M39 ;
    wire SubBytesIns_Inst_Sbox_6_M38 ;
    wire SubBytesIns_Inst_Sbox_6_M37 ;
    wire SubBytesIns_Inst_Sbox_6_M36 ;
    wire SubBytesIns_Inst_Sbox_6_M35 ;
    wire SubBytesIns_Inst_Sbox_6_M34 ;
    wire SubBytesIns_Inst_Sbox_6_M33 ;
    wire SubBytesIns_Inst_Sbox_6_M32 ;
    wire SubBytesIns_Inst_Sbox_6_M31 ;
    wire SubBytesIns_Inst_Sbox_6_M30 ;
    wire SubBytesIns_Inst_Sbox_6_M29 ;
    wire SubBytesIns_Inst_Sbox_6_M28 ;
    wire SubBytesIns_Inst_Sbox_6_M27 ;
    wire SubBytesIns_Inst_Sbox_6_M26 ;
    wire SubBytesIns_Inst_Sbox_6_M25 ;
    wire SubBytesIns_Inst_Sbox_6_M24 ;
    wire SubBytesIns_Inst_Sbox_6_M23 ;
    wire SubBytesIns_Inst_Sbox_6_M22 ;
    wire SubBytesIns_Inst_Sbox_6_M21 ;
    wire SubBytesIns_Inst_Sbox_6_M20 ;
    wire SubBytesIns_Inst_Sbox_6_M19 ;
    wire SubBytesIns_Inst_Sbox_6_M18 ;
    wire SubBytesIns_Inst_Sbox_6_M17 ;
    wire SubBytesIns_Inst_Sbox_6_M16 ;
    wire SubBytesIns_Inst_Sbox_6_M15 ;
    wire SubBytesIns_Inst_Sbox_6_M14 ;
    wire SubBytesIns_Inst_Sbox_6_M13 ;
    wire SubBytesIns_Inst_Sbox_6_M12 ;
    wire SubBytesIns_Inst_Sbox_6_M11 ;
    wire SubBytesIns_Inst_Sbox_6_M10 ;
    wire SubBytesIns_Inst_Sbox_6_M9 ;
    wire SubBytesIns_Inst_Sbox_6_M8 ;
    wire SubBytesIns_Inst_Sbox_6_M7 ;
    wire SubBytesIns_Inst_Sbox_6_M6 ;
    wire SubBytesIns_Inst_Sbox_6_M5 ;
    wire SubBytesIns_Inst_Sbox_6_M4 ;
    wire SubBytesIns_Inst_Sbox_6_M3 ;
    wire SubBytesIns_Inst_Sbox_6_M2 ;
    wire SubBytesIns_Inst_Sbox_6_M1 ;
    wire SubBytesIns_Inst_Sbox_6_T27 ;
    wire SubBytesIns_Inst_Sbox_6_T26 ;
    wire SubBytesIns_Inst_Sbox_6_T25 ;
    wire SubBytesIns_Inst_Sbox_6_T24 ;
    wire SubBytesIns_Inst_Sbox_6_T23 ;
    wire SubBytesIns_Inst_Sbox_6_T22 ;
    wire SubBytesIns_Inst_Sbox_6_T21 ;
    wire SubBytesIns_Inst_Sbox_6_T20 ;
    wire SubBytesIns_Inst_Sbox_6_T19 ;
    wire SubBytesIns_Inst_Sbox_6_T18 ;
    wire SubBytesIns_Inst_Sbox_6_T17 ;
    wire SubBytesIns_Inst_Sbox_6_T16 ;
    wire SubBytesIns_Inst_Sbox_6_T15 ;
    wire SubBytesIns_Inst_Sbox_6_T14 ;
    wire SubBytesIns_Inst_Sbox_6_T13 ;
    wire SubBytesIns_Inst_Sbox_6_T12 ;
    wire SubBytesIns_Inst_Sbox_6_T11 ;
    wire SubBytesIns_Inst_Sbox_6_T10 ;
    wire SubBytesIns_Inst_Sbox_6_T9 ;
    wire SubBytesIns_Inst_Sbox_6_T8 ;
    wire SubBytesIns_Inst_Sbox_6_T7 ;
    wire SubBytesIns_Inst_Sbox_6_T6 ;
    wire SubBytesIns_Inst_Sbox_6_T5 ;
    wire SubBytesIns_Inst_Sbox_6_T4 ;
    wire SubBytesIns_Inst_Sbox_6_T3 ;
    wire SubBytesIns_Inst_Sbox_6_T2 ;
    wire SubBytesIns_Inst_Sbox_6_T1 ;
    wire SubBytesIns_Inst_Sbox_7_L29 ;
    wire SubBytesIns_Inst_Sbox_7_L28 ;
    wire SubBytesIns_Inst_Sbox_7_L27 ;
    wire SubBytesIns_Inst_Sbox_7_L26 ;
    wire SubBytesIns_Inst_Sbox_7_L25 ;
    wire SubBytesIns_Inst_Sbox_7_L24 ;
    wire SubBytesIns_Inst_Sbox_7_L23 ;
    wire SubBytesIns_Inst_Sbox_7_L22 ;
    wire SubBytesIns_Inst_Sbox_7_L21 ;
    wire SubBytesIns_Inst_Sbox_7_L20 ;
    wire SubBytesIns_Inst_Sbox_7_L19 ;
    wire SubBytesIns_Inst_Sbox_7_L18 ;
    wire SubBytesIns_Inst_Sbox_7_L17 ;
    wire SubBytesIns_Inst_Sbox_7_L16 ;
    wire SubBytesIns_Inst_Sbox_7_L15 ;
    wire SubBytesIns_Inst_Sbox_7_L14 ;
    wire SubBytesIns_Inst_Sbox_7_L13 ;
    wire SubBytesIns_Inst_Sbox_7_L12 ;
    wire SubBytesIns_Inst_Sbox_7_L11 ;
    wire SubBytesIns_Inst_Sbox_7_L10 ;
    wire SubBytesIns_Inst_Sbox_7_L9 ;
    wire SubBytesIns_Inst_Sbox_7_L8 ;
    wire SubBytesIns_Inst_Sbox_7_L7 ;
    wire SubBytesIns_Inst_Sbox_7_L6 ;
    wire SubBytesIns_Inst_Sbox_7_L5 ;
    wire SubBytesIns_Inst_Sbox_7_L4 ;
    wire SubBytesIns_Inst_Sbox_7_L3 ;
    wire SubBytesIns_Inst_Sbox_7_L2 ;
    wire SubBytesIns_Inst_Sbox_7_L1 ;
    wire SubBytesIns_Inst_Sbox_7_L0 ;
    wire SubBytesIns_Inst_Sbox_7_M63 ;
    wire SubBytesIns_Inst_Sbox_7_M62 ;
    wire SubBytesIns_Inst_Sbox_7_M61 ;
    wire SubBytesIns_Inst_Sbox_7_M60 ;
    wire SubBytesIns_Inst_Sbox_7_M59 ;
    wire SubBytesIns_Inst_Sbox_7_M58 ;
    wire SubBytesIns_Inst_Sbox_7_M57 ;
    wire SubBytesIns_Inst_Sbox_7_M56 ;
    wire SubBytesIns_Inst_Sbox_7_M55 ;
    wire SubBytesIns_Inst_Sbox_7_M54 ;
    wire SubBytesIns_Inst_Sbox_7_M53 ;
    wire SubBytesIns_Inst_Sbox_7_M52 ;
    wire SubBytesIns_Inst_Sbox_7_M51 ;
    wire SubBytesIns_Inst_Sbox_7_M50 ;
    wire SubBytesIns_Inst_Sbox_7_M49 ;
    wire SubBytesIns_Inst_Sbox_7_M48 ;
    wire SubBytesIns_Inst_Sbox_7_M47 ;
    wire SubBytesIns_Inst_Sbox_7_M46 ;
    wire SubBytesIns_Inst_Sbox_7_M45 ;
    wire SubBytesIns_Inst_Sbox_7_M44 ;
    wire SubBytesIns_Inst_Sbox_7_M43 ;
    wire SubBytesIns_Inst_Sbox_7_M42 ;
    wire SubBytesIns_Inst_Sbox_7_M41 ;
    wire SubBytesIns_Inst_Sbox_7_M40 ;
    wire SubBytesIns_Inst_Sbox_7_M39 ;
    wire SubBytesIns_Inst_Sbox_7_M38 ;
    wire SubBytesIns_Inst_Sbox_7_M37 ;
    wire SubBytesIns_Inst_Sbox_7_M36 ;
    wire SubBytesIns_Inst_Sbox_7_M35 ;
    wire SubBytesIns_Inst_Sbox_7_M34 ;
    wire SubBytesIns_Inst_Sbox_7_M33 ;
    wire SubBytesIns_Inst_Sbox_7_M32 ;
    wire SubBytesIns_Inst_Sbox_7_M31 ;
    wire SubBytesIns_Inst_Sbox_7_M30 ;
    wire SubBytesIns_Inst_Sbox_7_M29 ;
    wire SubBytesIns_Inst_Sbox_7_M28 ;
    wire SubBytesIns_Inst_Sbox_7_M27 ;
    wire SubBytesIns_Inst_Sbox_7_M26 ;
    wire SubBytesIns_Inst_Sbox_7_M25 ;
    wire SubBytesIns_Inst_Sbox_7_M24 ;
    wire SubBytesIns_Inst_Sbox_7_M23 ;
    wire SubBytesIns_Inst_Sbox_7_M22 ;
    wire SubBytesIns_Inst_Sbox_7_M21 ;
    wire SubBytesIns_Inst_Sbox_7_M20 ;
    wire SubBytesIns_Inst_Sbox_7_M19 ;
    wire SubBytesIns_Inst_Sbox_7_M18 ;
    wire SubBytesIns_Inst_Sbox_7_M17 ;
    wire SubBytesIns_Inst_Sbox_7_M16 ;
    wire SubBytesIns_Inst_Sbox_7_M15 ;
    wire SubBytesIns_Inst_Sbox_7_M14 ;
    wire SubBytesIns_Inst_Sbox_7_M13 ;
    wire SubBytesIns_Inst_Sbox_7_M12 ;
    wire SubBytesIns_Inst_Sbox_7_M11 ;
    wire SubBytesIns_Inst_Sbox_7_M10 ;
    wire SubBytesIns_Inst_Sbox_7_M9 ;
    wire SubBytesIns_Inst_Sbox_7_M8 ;
    wire SubBytesIns_Inst_Sbox_7_M7 ;
    wire SubBytesIns_Inst_Sbox_7_M6 ;
    wire SubBytesIns_Inst_Sbox_7_M5 ;
    wire SubBytesIns_Inst_Sbox_7_M4 ;
    wire SubBytesIns_Inst_Sbox_7_M3 ;
    wire SubBytesIns_Inst_Sbox_7_M2 ;
    wire SubBytesIns_Inst_Sbox_7_M1 ;
    wire SubBytesIns_Inst_Sbox_7_T27 ;
    wire SubBytesIns_Inst_Sbox_7_T26 ;
    wire SubBytesIns_Inst_Sbox_7_T25 ;
    wire SubBytesIns_Inst_Sbox_7_T24 ;
    wire SubBytesIns_Inst_Sbox_7_T23 ;
    wire SubBytesIns_Inst_Sbox_7_T22 ;
    wire SubBytesIns_Inst_Sbox_7_T21 ;
    wire SubBytesIns_Inst_Sbox_7_T20 ;
    wire SubBytesIns_Inst_Sbox_7_T19 ;
    wire SubBytesIns_Inst_Sbox_7_T18 ;
    wire SubBytesIns_Inst_Sbox_7_T17 ;
    wire SubBytesIns_Inst_Sbox_7_T16 ;
    wire SubBytesIns_Inst_Sbox_7_T15 ;
    wire SubBytesIns_Inst_Sbox_7_T14 ;
    wire SubBytesIns_Inst_Sbox_7_T13 ;
    wire SubBytesIns_Inst_Sbox_7_T12 ;
    wire SubBytesIns_Inst_Sbox_7_T11 ;
    wire SubBytesIns_Inst_Sbox_7_T10 ;
    wire SubBytesIns_Inst_Sbox_7_T9 ;
    wire SubBytesIns_Inst_Sbox_7_T8 ;
    wire SubBytesIns_Inst_Sbox_7_T7 ;
    wire SubBytesIns_Inst_Sbox_7_T6 ;
    wire SubBytesIns_Inst_Sbox_7_T5 ;
    wire SubBytesIns_Inst_Sbox_7_T4 ;
    wire SubBytesIns_Inst_Sbox_7_T3 ;
    wire SubBytesIns_Inst_Sbox_7_T2 ;
    wire SubBytesIns_Inst_Sbox_7_T1 ;
    wire SubBytesIns_Inst_Sbox_8_L29 ;
    wire SubBytesIns_Inst_Sbox_8_L28 ;
    wire SubBytesIns_Inst_Sbox_8_L27 ;
    wire SubBytesIns_Inst_Sbox_8_L26 ;
    wire SubBytesIns_Inst_Sbox_8_L25 ;
    wire SubBytesIns_Inst_Sbox_8_L24 ;
    wire SubBytesIns_Inst_Sbox_8_L23 ;
    wire SubBytesIns_Inst_Sbox_8_L22 ;
    wire SubBytesIns_Inst_Sbox_8_L21 ;
    wire SubBytesIns_Inst_Sbox_8_L20 ;
    wire SubBytesIns_Inst_Sbox_8_L19 ;
    wire SubBytesIns_Inst_Sbox_8_L18 ;
    wire SubBytesIns_Inst_Sbox_8_L17 ;
    wire SubBytesIns_Inst_Sbox_8_L16 ;
    wire SubBytesIns_Inst_Sbox_8_L15 ;
    wire SubBytesIns_Inst_Sbox_8_L14 ;
    wire SubBytesIns_Inst_Sbox_8_L13 ;
    wire SubBytesIns_Inst_Sbox_8_L12 ;
    wire SubBytesIns_Inst_Sbox_8_L11 ;
    wire SubBytesIns_Inst_Sbox_8_L10 ;
    wire SubBytesIns_Inst_Sbox_8_L9 ;
    wire SubBytesIns_Inst_Sbox_8_L8 ;
    wire SubBytesIns_Inst_Sbox_8_L7 ;
    wire SubBytesIns_Inst_Sbox_8_L6 ;
    wire SubBytesIns_Inst_Sbox_8_L5 ;
    wire SubBytesIns_Inst_Sbox_8_L4 ;
    wire SubBytesIns_Inst_Sbox_8_L3 ;
    wire SubBytesIns_Inst_Sbox_8_L2 ;
    wire SubBytesIns_Inst_Sbox_8_L1 ;
    wire SubBytesIns_Inst_Sbox_8_L0 ;
    wire SubBytesIns_Inst_Sbox_8_M63 ;
    wire SubBytesIns_Inst_Sbox_8_M62 ;
    wire SubBytesIns_Inst_Sbox_8_M61 ;
    wire SubBytesIns_Inst_Sbox_8_M60 ;
    wire SubBytesIns_Inst_Sbox_8_M59 ;
    wire SubBytesIns_Inst_Sbox_8_M58 ;
    wire SubBytesIns_Inst_Sbox_8_M57 ;
    wire SubBytesIns_Inst_Sbox_8_M56 ;
    wire SubBytesIns_Inst_Sbox_8_M55 ;
    wire SubBytesIns_Inst_Sbox_8_M54 ;
    wire SubBytesIns_Inst_Sbox_8_M53 ;
    wire SubBytesIns_Inst_Sbox_8_M52 ;
    wire SubBytesIns_Inst_Sbox_8_M51 ;
    wire SubBytesIns_Inst_Sbox_8_M50 ;
    wire SubBytesIns_Inst_Sbox_8_M49 ;
    wire SubBytesIns_Inst_Sbox_8_M48 ;
    wire SubBytesIns_Inst_Sbox_8_M47 ;
    wire SubBytesIns_Inst_Sbox_8_M46 ;
    wire SubBytesIns_Inst_Sbox_8_M45 ;
    wire SubBytesIns_Inst_Sbox_8_M44 ;
    wire SubBytesIns_Inst_Sbox_8_M43 ;
    wire SubBytesIns_Inst_Sbox_8_M42 ;
    wire SubBytesIns_Inst_Sbox_8_M41 ;
    wire SubBytesIns_Inst_Sbox_8_M40 ;
    wire SubBytesIns_Inst_Sbox_8_M39 ;
    wire SubBytesIns_Inst_Sbox_8_M38 ;
    wire SubBytesIns_Inst_Sbox_8_M37 ;
    wire SubBytesIns_Inst_Sbox_8_M36 ;
    wire SubBytesIns_Inst_Sbox_8_M35 ;
    wire SubBytesIns_Inst_Sbox_8_M34 ;
    wire SubBytesIns_Inst_Sbox_8_M33 ;
    wire SubBytesIns_Inst_Sbox_8_M32 ;
    wire SubBytesIns_Inst_Sbox_8_M31 ;
    wire SubBytesIns_Inst_Sbox_8_M30 ;
    wire SubBytesIns_Inst_Sbox_8_M29 ;
    wire SubBytesIns_Inst_Sbox_8_M28 ;
    wire SubBytesIns_Inst_Sbox_8_M27 ;
    wire SubBytesIns_Inst_Sbox_8_M26 ;
    wire SubBytesIns_Inst_Sbox_8_M25 ;
    wire SubBytesIns_Inst_Sbox_8_M24 ;
    wire SubBytesIns_Inst_Sbox_8_M23 ;
    wire SubBytesIns_Inst_Sbox_8_M22 ;
    wire SubBytesIns_Inst_Sbox_8_M21 ;
    wire SubBytesIns_Inst_Sbox_8_M20 ;
    wire SubBytesIns_Inst_Sbox_8_M19 ;
    wire SubBytesIns_Inst_Sbox_8_M18 ;
    wire SubBytesIns_Inst_Sbox_8_M17 ;
    wire SubBytesIns_Inst_Sbox_8_M16 ;
    wire SubBytesIns_Inst_Sbox_8_M15 ;
    wire SubBytesIns_Inst_Sbox_8_M14 ;
    wire SubBytesIns_Inst_Sbox_8_M13 ;
    wire SubBytesIns_Inst_Sbox_8_M12 ;
    wire SubBytesIns_Inst_Sbox_8_M11 ;
    wire SubBytesIns_Inst_Sbox_8_M10 ;
    wire SubBytesIns_Inst_Sbox_8_M9 ;
    wire SubBytesIns_Inst_Sbox_8_M8 ;
    wire SubBytesIns_Inst_Sbox_8_M7 ;
    wire SubBytesIns_Inst_Sbox_8_M6 ;
    wire SubBytesIns_Inst_Sbox_8_M5 ;
    wire SubBytesIns_Inst_Sbox_8_M4 ;
    wire SubBytesIns_Inst_Sbox_8_M3 ;
    wire SubBytesIns_Inst_Sbox_8_M2 ;
    wire SubBytesIns_Inst_Sbox_8_M1 ;
    wire SubBytesIns_Inst_Sbox_8_T27 ;
    wire SubBytesIns_Inst_Sbox_8_T26 ;
    wire SubBytesIns_Inst_Sbox_8_T25 ;
    wire SubBytesIns_Inst_Sbox_8_T24 ;
    wire SubBytesIns_Inst_Sbox_8_T23 ;
    wire SubBytesIns_Inst_Sbox_8_T22 ;
    wire SubBytesIns_Inst_Sbox_8_T21 ;
    wire SubBytesIns_Inst_Sbox_8_T20 ;
    wire SubBytesIns_Inst_Sbox_8_T19 ;
    wire SubBytesIns_Inst_Sbox_8_T18 ;
    wire SubBytesIns_Inst_Sbox_8_T17 ;
    wire SubBytesIns_Inst_Sbox_8_T16 ;
    wire SubBytesIns_Inst_Sbox_8_T15 ;
    wire SubBytesIns_Inst_Sbox_8_T14 ;
    wire SubBytesIns_Inst_Sbox_8_T13 ;
    wire SubBytesIns_Inst_Sbox_8_T12 ;
    wire SubBytesIns_Inst_Sbox_8_T11 ;
    wire SubBytesIns_Inst_Sbox_8_T10 ;
    wire SubBytesIns_Inst_Sbox_8_T9 ;
    wire SubBytesIns_Inst_Sbox_8_T8 ;
    wire SubBytesIns_Inst_Sbox_8_T7 ;
    wire SubBytesIns_Inst_Sbox_8_T6 ;
    wire SubBytesIns_Inst_Sbox_8_T5 ;
    wire SubBytesIns_Inst_Sbox_8_T4 ;
    wire SubBytesIns_Inst_Sbox_8_T3 ;
    wire SubBytesIns_Inst_Sbox_8_T2 ;
    wire SubBytesIns_Inst_Sbox_8_T1 ;
    wire SubBytesIns_Inst_Sbox_9_L29 ;
    wire SubBytesIns_Inst_Sbox_9_L28 ;
    wire SubBytesIns_Inst_Sbox_9_L27 ;
    wire SubBytesIns_Inst_Sbox_9_L26 ;
    wire SubBytesIns_Inst_Sbox_9_L25 ;
    wire SubBytesIns_Inst_Sbox_9_L24 ;
    wire SubBytesIns_Inst_Sbox_9_L23 ;
    wire SubBytesIns_Inst_Sbox_9_L22 ;
    wire SubBytesIns_Inst_Sbox_9_L21 ;
    wire SubBytesIns_Inst_Sbox_9_L20 ;
    wire SubBytesIns_Inst_Sbox_9_L19 ;
    wire SubBytesIns_Inst_Sbox_9_L18 ;
    wire SubBytesIns_Inst_Sbox_9_L17 ;
    wire SubBytesIns_Inst_Sbox_9_L16 ;
    wire SubBytesIns_Inst_Sbox_9_L15 ;
    wire SubBytesIns_Inst_Sbox_9_L14 ;
    wire SubBytesIns_Inst_Sbox_9_L13 ;
    wire SubBytesIns_Inst_Sbox_9_L12 ;
    wire SubBytesIns_Inst_Sbox_9_L11 ;
    wire SubBytesIns_Inst_Sbox_9_L10 ;
    wire SubBytesIns_Inst_Sbox_9_L9 ;
    wire SubBytesIns_Inst_Sbox_9_L8 ;
    wire SubBytesIns_Inst_Sbox_9_L7 ;
    wire SubBytesIns_Inst_Sbox_9_L6 ;
    wire SubBytesIns_Inst_Sbox_9_L5 ;
    wire SubBytesIns_Inst_Sbox_9_L4 ;
    wire SubBytesIns_Inst_Sbox_9_L3 ;
    wire SubBytesIns_Inst_Sbox_9_L2 ;
    wire SubBytesIns_Inst_Sbox_9_L1 ;
    wire SubBytesIns_Inst_Sbox_9_L0 ;
    wire SubBytesIns_Inst_Sbox_9_M63 ;
    wire SubBytesIns_Inst_Sbox_9_M62 ;
    wire SubBytesIns_Inst_Sbox_9_M61 ;
    wire SubBytesIns_Inst_Sbox_9_M60 ;
    wire SubBytesIns_Inst_Sbox_9_M59 ;
    wire SubBytesIns_Inst_Sbox_9_M58 ;
    wire SubBytesIns_Inst_Sbox_9_M57 ;
    wire SubBytesIns_Inst_Sbox_9_M56 ;
    wire SubBytesIns_Inst_Sbox_9_M55 ;
    wire SubBytesIns_Inst_Sbox_9_M54 ;
    wire SubBytesIns_Inst_Sbox_9_M53 ;
    wire SubBytesIns_Inst_Sbox_9_M52 ;
    wire SubBytesIns_Inst_Sbox_9_M51 ;
    wire SubBytesIns_Inst_Sbox_9_M50 ;
    wire SubBytesIns_Inst_Sbox_9_M49 ;
    wire SubBytesIns_Inst_Sbox_9_M48 ;
    wire SubBytesIns_Inst_Sbox_9_M47 ;
    wire SubBytesIns_Inst_Sbox_9_M46 ;
    wire SubBytesIns_Inst_Sbox_9_M45 ;
    wire SubBytesIns_Inst_Sbox_9_M44 ;
    wire SubBytesIns_Inst_Sbox_9_M43 ;
    wire SubBytesIns_Inst_Sbox_9_M42 ;
    wire SubBytesIns_Inst_Sbox_9_M41 ;
    wire SubBytesIns_Inst_Sbox_9_M40 ;
    wire SubBytesIns_Inst_Sbox_9_M39 ;
    wire SubBytesIns_Inst_Sbox_9_M38 ;
    wire SubBytesIns_Inst_Sbox_9_M37 ;
    wire SubBytesIns_Inst_Sbox_9_M36 ;
    wire SubBytesIns_Inst_Sbox_9_M35 ;
    wire SubBytesIns_Inst_Sbox_9_M34 ;
    wire SubBytesIns_Inst_Sbox_9_M33 ;
    wire SubBytesIns_Inst_Sbox_9_M32 ;
    wire SubBytesIns_Inst_Sbox_9_M31 ;
    wire SubBytesIns_Inst_Sbox_9_M30 ;
    wire SubBytesIns_Inst_Sbox_9_M29 ;
    wire SubBytesIns_Inst_Sbox_9_M28 ;
    wire SubBytesIns_Inst_Sbox_9_M27 ;
    wire SubBytesIns_Inst_Sbox_9_M26 ;
    wire SubBytesIns_Inst_Sbox_9_M25 ;
    wire SubBytesIns_Inst_Sbox_9_M24 ;
    wire SubBytesIns_Inst_Sbox_9_M23 ;
    wire SubBytesIns_Inst_Sbox_9_M22 ;
    wire SubBytesIns_Inst_Sbox_9_M21 ;
    wire SubBytesIns_Inst_Sbox_9_M20 ;
    wire SubBytesIns_Inst_Sbox_9_M19 ;
    wire SubBytesIns_Inst_Sbox_9_M18 ;
    wire SubBytesIns_Inst_Sbox_9_M17 ;
    wire SubBytesIns_Inst_Sbox_9_M16 ;
    wire SubBytesIns_Inst_Sbox_9_M15 ;
    wire SubBytesIns_Inst_Sbox_9_M14 ;
    wire SubBytesIns_Inst_Sbox_9_M13 ;
    wire SubBytesIns_Inst_Sbox_9_M12 ;
    wire SubBytesIns_Inst_Sbox_9_M11 ;
    wire SubBytesIns_Inst_Sbox_9_M10 ;
    wire SubBytesIns_Inst_Sbox_9_M9 ;
    wire SubBytesIns_Inst_Sbox_9_M8 ;
    wire SubBytesIns_Inst_Sbox_9_M7 ;
    wire SubBytesIns_Inst_Sbox_9_M6 ;
    wire SubBytesIns_Inst_Sbox_9_M5 ;
    wire SubBytesIns_Inst_Sbox_9_M4 ;
    wire SubBytesIns_Inst_Sbox_9_M3 ;
    wire SubBytesIns_Inst_Sbox_9_M2 ;
    wire SubBytesIns_Inst_Sbox_9_M1 ;
    wire SubBytesIns_Inst_Sbox_9_T27 ;
    wire SubBytesIns_Inst_Sbox_9_T26 ;
    wire SubBytesIns_Inst_Sbox_9_T25 ;
    wire SubBytesIns_Inst_Sbox_9_T24 ;
    wire SubBytesIns_Inst_Sbox_9_T23 ;
    wire SubBytesIns_Inst_Sbox_9_T22 ;
    wire SubBytesIns_Inst_Sbox_9_T21 ;
    wire SubBytesIns_Inst_Sbox_9_T20 ;
    wire SubBytesIns_Inst_Sbox_9_T19 ;
    wire SubBytesIns_Inst_Sbox_9_T18 ;
    wire SubBytesIns_Inst_Sbox_9_T17 ;
    wire SubBytesIns_Inst_Sbox_9_T16 ;
    wire SubBytesIns_Inst_Sbox_9_T15 ;
    wire SubBytesIns_Inst_Sbox_9_T14 ;
    wire SubBytesIns_Inst_Sbox_9_T13 ;
    wire SubBytesIns_Inst_Sbox_9_T12 ;
    wire SubBytesIns_Inst_Sbox_9_T11 ;
    wire SubBytesIns_Inst_Sbox_9_T10 ;
    wire SubBytesIns_Inst_Sbox_9_T9 ;
    wire SubBytesIns_Inst_Sbox_9_T8 ;
    wire SubBytesIns_Inst_Sbox_9_T7 ;
    wire SubBytesIns_Inst_Sbox_9_T6 ;
    wire SubBytesIns_Inst_Sbox_9_T5 ;
    wire SubBytesIns_Inst_Sbox_9_T4 ;
    wire SubBytesIns_Inst_Sbox_9_T3 ;
    wire SubBytesIns_Inst_Sbox_9_T2 ;
    wire SubBytesIns_Inst_Sbox_9_T1 ;
    wire SubBytesIns_Inst_Sbox_10_L29 ;
    wire SubBytesIns_Inst_Sbox_10_L28 ;
    wire SubBytesIns_Inst_Sbox_10_L27 ;
    wire SubBytesIns_Inst_Sbox_10_L26 ;
    wire SubBytesIns_Inst_Sbox_10_L25 ;
    wire SubBytesIns_Inst_Sbox_10_L24 ;
    wire SubBytesIns_Inst_Sbox_10_L23 ;
    wire SubBytesIns_Inst_Sbox_10_L22 ;
    wire SubBytesIns_Inst_Sbox_10_L21 ;
    wire SubBytesIns_Inst_Sbox_10_L20 ;
    wire SubBytesIns_Inst_Sbox_10_L19 ;
    wire SubBytesIns_Inst_Sbox_10_L18 ;
    wire SubBytesIns_Inst_Sbox_10_L17 ;
    wire SubBytesIns_Inst_Sbox_10_L16 ;
    wire SubBytesIns_Inst_Sbox_10_L15 ;
    wire SubBytesIns_Inst_Sbox_10_L14 ;
    wire SubBytesIns_Inst_Sbox_10_L13 ;
    wire SubBytesIns_Inst_Sbox_10_L12 ;
    wire SubBytesIns_Inst_Sbox_10_L11 ;
    wire SubBytesIns_Inst_Sbox_10_L10 ;
    wire SubBytesIns_Inst_Sbox_10_L9 ;
    wire SubBytesIns_Inst_Sbox_10_L8 ;
    wire SubBytesIns_Inst_Sbox_10_L7 ;
    wire SubBytesIns_Inst_Sbox_10_L6 ;
    wire SubBytesIns_Inst_Sbox_10_L5 ;
    wire SubBytesIns_Inst_Sbox_10_L4 ;
    wire SubBytesIns_Inst_Sbox_10_L3 ;
    wire SubBytesIns_Inst_Sbox_10_L2 ;
    wire SubBytesIns_Inst_Sbox_10_L1 ;
    wire SubBytesIns_Inst_Sbox_10_L0 ;
    wire SubBytesIns_Inst_Sbox_10_M63 ;
    wire SubBytesIns_Inst_Sbox_10_M62 ;
    wire SubBytesIns_Inst_Sbox_10_M61 ;
    wire SubBytesIns_Inst_Sbox_10_M60 ;
    wire SubBytesIns_Inst_Sbox_10_M59 ;
    wire SubBytesIns_Inst_Sbox_10_M58 ;
    wire SubBytesIns_Inst_Sbox_10_M57 ;
    wire SubBytesIns_Inst_Sbox_10_M56 ;
    wire SubBytesIns_Inst_Sbox_10_M55 ;
    wire SubBytesIns_Inst_Sbox_10_M54 ;
    wire SubBytesIns_Inst_Sbox_10_M53 ;
    wire SubBytesIns_Inst_Sbox_10_M52 ;
    wire SubBytesIns_Inst_Sbox_10_M51 ;
    wire SubBytesIns_Inst_Sbox_10_M50 ;
    wire SubBytesIns_Inst_Sbox_10_M49 ;
    wire SubBytesIns_Inst_Sbox_10_M48 ;
    wire SubBytesIns_Inst_Sbox_10_M47 ;
    wire SubBytesIns_Inst_Sbox_10_M46 ;
    wire SubBytesIns_Inst_Sbox_10_M45 ;
    wire SubBytesIns_Inst_Sbox_10_M44 ;
    wire SubBytesIns_Inst_Sbox_10_M43 ;
    wire SubBytesIns_Inst_Sbox_10_M42 ;
    wire SubBytesIns_Inst_Sbox_10_M41 ;
    wire SubBytesIns_Inst_Sbox_10_M40 ;
    wire SubBytesIns_Inst_Sbox_10_M39 ;
    wire SubBytesIns_Inst_Sbox_10_M38 ;
    wire SubBytesIns_Inst_Sbox_10_M37 ;
    wire SubBytesIns_Inst_Sbox_10_M36 ;
    wire SubBytesIns_Inst_Sbox_10_M35 ;
    wire SubBytesIns_Inst_Sbox_10_M34 ;
    wire SubBytesIns_Inst_Sbox_10_M33 ;
    wire SubBytesIns_Inst_Sbox_10_M32 ;
    wire SubBytesIns_Inst_Sbox_10_M31 ;
    wire SubBytesIns_Inst_Sbox_10_M30 ;
    wire SubBytesIns_Inst_Sbox_10_M29 ;
    wire SubBytesIns_Inst_Sbox_10_M28 ;
    wire SubBytesIns_Inst_Sbox_10_M27 ;
    wire SubBytesIns_Inst_Sbox_10_M26 ;
    wire SubBytesIns_Inst_Sbox_10_M25 ;
    wire SubBytesIns_Inst_Sbox_10_M24 ;
    wire SubBytesIns_Inst_Sbox_10_M23 ;
    wire SubBytesIns_Inst_Sbox_10_M22 ;
    wire SubBytesIns_Inst_Sbox_10_M21 ;
    wire SubBytesIns_Inst_Sbox_10_M20 ;
    wire SubBytesIns_Inst_Sbox_10_M19 ;
    wire SubBytesIns_Inst_Sbox_10_M18 ;
    wire SubBytesIns_Inst_Sbox_10_M17 ;
    wire SubBytesIns_Inst_Sbox_10_M16 ;
    wire SubBytesIns_Inst_Sbox_10_M15 ;
    wire SubBytesIns_Inst_Sbox_10_M14 ;
    wire SubBytesIns_Inst_Sbox_10_M13 ;
    wire SubBytesIns_Inst_Sbox_10_M12 ;
    wire SubBytesIns_Inst_Sbox_10_M11 ;
    wire SubBytesIns_Inst_Sbox_10_M10 ;
    wire SubBytesIns_Inst_Sbox_10_M9 ;
    wire SubBytesIns_Inst_Sbox_10_M8 ;
    wire SubBytesIns_Inst_Sbox_10_M7 ;
    wire SubBytesIns_Inst_Sbox_10_M6 ;
    wire SubBytesIns_Inst_Sbox_10_M5 ;
    wire SubBytesIns_Inst_Sbox_10_M4 ;
    wire SubBytesIns_Inst_Sbox_10_M3 ;
    wire SubBytesIns_Inst_Sbox_10_M2 ;
    wire SubBytesIns_Inst_Sbox_10_M1 ;
    wire SubBytesIns_Inst_Sbox_10_T27 ;
    wire SubBytesIns_Inst_Sbox_10_T26 ;
    wire SubBytesIns_Inst_Sbox_10_T25 ;
    wire SubBytesIns_Inst_Sbox_10_T24 ;
    wire SubBytesIns_Inst_Sbox_10_T23 ;
    wire SubBytesIns_Inst_Sbox_10_T22 ;
    wire SubBytesIns_Inst_Sbox_10_T21 ;
    wire SubBytesIns_Inst_Sbox_10_T20 ;
    wire SubBytesIns_Inst_Sbox_10_T19 ;
    wire SubBytesIns_Inst_Sbox_10_T18 ;
    wire SubBytesIns_Inst_Sbox_10_T17 ;
    wire SubBytesIns_Inst_Sbox_10_T16 ;
    wire SubBytesIns_Inst_Sbox_10_T15 ;
    wire SubBytesIns_Inst_Sbox_10_T14 ;
    wire SubBytesIns_Inst_Sbox_10_T13 ;
    wire SubBytesIns_Inst_Sbox_10_T12 ;
    wire SubBytesIns_Inst_Sbox_10_T11 ;
    wire SubBytesIns_Inst_Sbox_10_T10 ;
    wire SubBytesIns_Inst_Sbox_10_T9 ;
    wire SubBytesIns_Inst_Sbox_10_T8 ;
    wire SubBytesIns_Inst_Sbox_10_T7 ;
    wire SubBytesIns_Inst_Sbox_10_T6 ;
    wire SubBytesIns_Inst_Sbox_10_T5 ;
    wire SubBytesIns_Inst_Sbox_10_T4 ;
    wire SubBytesIns_Inst_Sbox_10_T3 ;
    wire SubBytesIns_Inst_Sbox_10_T2 ;
    wire SubBytesIns_Inst_Sbox_10_T1 ;
    wire SubBytesIns_Inst_Sbox_11_L29 ;
    wire SubBytesIns_Inst_Sbox_11_L28 ;
    wire SubBytesIns_Inst_Sbox_11_L27 ;
    wire SubBytesIns_Inst_Sbox_11_L26 ;
    wire SubBytesIns_Inst_Sbox_11_L25 ;
    wire SubBytesIns_Inst_Sbox_11_L24 ;
    wire SubBytesIns_Inst_Sbox_11_L23 ;
    wire SubBytesIns_Inst_Sbox_11_L22 ;
    wire SubBytesIns_Inst_Sbox_11_L21 ;
    wire SubBytesIns_Inst_Sbox_11_L20 ;
    wire SubBytesIns_Inst_Sbox_11_L19 ;
    wire SubBytesIns_Inst_Sbox_11_L18 ;
    wire SubBytesIns_Inst_Sbox_11_L17 ;
    wire SubBytesIns_Inst_Sbox_11_L16 ;
    wire SubBytesIns_Inst_Sbox_11_L15 ;
    wire SubBytesIns_Inst_Sbox_11_L14 ;
    wire SubBytesIns_Inst_Sbox_11_L13 ;
    wire SubBytesIns_Inst_Sbox_11_L12 ;
    wire SubBytesIns_Inst_Sbox_11_L11 ;
    wire SubBytesIns_Inst_Sbox_11_L10 ;
    wire SubBytesIns_Inst_Sbox_11_L9 ;
    wire SubBytesIns_Inst_Sbox_11_L8 ;
    wire SubBytesIns_Inst_Sbox_11_L7 ;
    wire SubBytesIns_Inst_Sbox_11_L6 ;
    wire SubBytesIns_Inst_Sbox_11_L5 ;
    wire SubBytesIns_Inst_Sbox_11_L4 ;
    wire SubBytesIns_Inst_Sbox_11_L3 ;
    wire SubBytesIns_Inst_Sbox_11_L2 ;
    wire SubBytesIns_Inst_Sbox_11_L1 ;
    wire SubBytesIns_Inst_Sbox_11_L0 ;
    wire SubBytesIns_Inst_Sbox_11_M63 ;
    wire SubBytesIns_Inst_Sbox_11_M62 ;
    wire SubBytesIns_Inst_Sbox_11_M61 ;
    wire SubBytesIns_Inst_Sbox_11_M60 ;
    wire SubBytesIns_Inst_Sbox_11_M59 ;
    wire SubBytesIns_Inst_Sbox_11_M58 ;
    wire SubBytesIns_Inst_Sbox_11_M57 ;
    wire SubBytesIns_Inst_Sbox_11_M56 ;
    wire SubBytesIns_Inst_Sbox_11_M55 ;
    wire SubBytesIns_Inst_Sbox_11_M54 ;
    wire SubBytesIns_Inst_Sbox_11_M53 ;
    wire SubBytesIns_Inst_Sbox_11_M52 ;
    wire SubBytesIns_Inst_Sbox_11_M51 ;
    wire SubBytesIns_Inst_Sbox_11_M50 ;
    wire SubBytesIns_Inst_Sbox_11_M49 ;
    wire SubBytesIns_Inst_Sbox_11_M48 ;
    wire SubBytesIns_Inst_Sbox_11_M47 ;
    wire SubBytesIns_Inst_Sbox_11_M46 ;
    wire SubBytesIns_Inst_Sbox_11_M45 ;
    wire SubBytesIns_Inst_Sbox_11_M44 ;
    wire SubBytesIns_Inst_Sbox_11_M43 ;
    wire SubBytesIns_Inst_Sbox_11_M42 ;
    wire SubBytesIns_Inst_Sbox_11_M41 ;
    wire SubBytesIns_Inst_Sbox_11_M40 ;
    wire SubBytesIns_Inst_Sbox_11_M39 ;
    wire SubBytesIns_Inst_Sbox_11_M38 ;
    wire SubBytesIns_Inst_Sbox_11_M37 ;
    wire SubBytesIns_Inst_Sbox_11_M36 ;
    wire SubBytesIns_Inst_Sbox_11_M35 ;
    wire SubBytesIns_Inst_Sbox_11_M34 ;
    wire SubBytesIns_Inst_Sbox_11_M33 ;
    wire SubBytesIns_Inst_Sbox_11_M32 ;
    wire SubBytesIns_Inst_Sbox_11_M31 ;
    wire SubBytesIns_Inst_Sbox_11_M30 ;
    wire SubBytesIns_Inst_Sbox_11_M29 ;
    wire SubBytesIns_Inst_Sbox_11_M28 ;
    wire SubBytesIns_Inst_Sbox_11_M27 ;
    wire SubBytesIns_Inst_Sbox_11_M26 ;
    wire SubBytesIns_Inst_Sbox_11_M25 ;
    wire SubBytesIns_Inst_Sbox_11_M24 ;
    wire SubBytesIns_Inst_Sbox_11_M23 ;
    wire SubBytesIns_Inst_Sbox_11_M22 ;
    wire SubBytesIns_Inst_Sbox_11_M21 ;
    wire SubBytesIns_Inst_Sbox_11_M20 ;
    wire SubBytesIns_Inst_Sbox_11_M19 ;
    wire SubBytesIns_Inst_Sbox_11_M18 ;
    wire SubBytesIns_Inst_Sbox_11_M17 ;
    wire SubBytesIns_Inst_Sbox_11_M16 ;
    wire SubBytesIns_Inst_Sbox_11_M15 ;
    wire SubBytesIns_Inst_Sbox_11_M14 ;
    wire SubBytesIns_Inst_Sbox_11_M13 ;
    wire SubBytesIns_Inst_Sbox_11_M12 ;
    wire SubBytesIns_Inst_Sbox_11_M11 ;
    wire SubBytesIns_Inst_Sbox_11_M10 ;
    wire SubBytesIns_Inst_Sbox_11_M9 ;
    wire SubBytesIns_Inst_Sbox_11_M8 ;
    wire SubBytesIns_Inst_Sbox_11_M7 ;
    wire SubBytesIns_Inst_Sbox_11_M6 ;
    wire SubBytesIns_Inst_Sbox_11_M5 ;
    wire SubBytesIns_Inst_Sbox_11_M4 ;
    wire SubBytesIns_Inst_Sbox_11_M3 ;
    wire SubBytesIns_Inst_Sbox_11_M2 ;
    wire SubBytesIns_Inst_Sbox_11_M1 ;
    wire SubBytesIns_Inst_Sbox_11_T27 ;
    wire SubBytesIns_Inst_Sbox_11_T26 ;
    wire SubBytesIns_Inst_Sbox_11_T25 ;
    wire SubBytesIns_Inst_Sbox_11_T24 ;
    wire SubBytesIns_Inst_Sbox_11_T23 ;
    wire SubBytesIns_Inst_Sbox_11_T22 ;
    wire SubBytesIns_Inst_Sbox_11_T21 ;
    wire SubBytesIns_Inst_Sbox_11_T20 ;
    wire SubBytesIns_Inst_Sbox_11_T19 ;
    wire SubBytesIns_Inst_Sbox_11_T18 ;
    wire SubBytesIns_Inst_Sbox_11_T17 ;
    wire SubBytesIns_Inst_Sbox_11_T16 ;
    wire SubBytesIns_Inst_Sbox_11_T15 ;
    wire SubBytesIns_Inst_Sbox_11_T14 ;
    wire SubBytesIns_Inst_Sbox_11_T13 ;
    wire SubBytesIns_Inst_Sbox_11_T12 ;
    wire SubBytesIns_Inst_Sbox_11_T11 ;
    wire SubBytesIns_Inst_Sbox_11_T10 ;
    wire SubBytesIns_Inst_Sbox_11_T9 ;
    wire SubBytesIns_Inst_Sbox_11_T8 ;
    wire SubBytesIns_Inst_Sbox_11_T7 ;
    wire SubBytesIns_Inst_Sbox_11_T6 ;
    wire SubBytesIns_Inst_Sbox_11_T5 ;
    wire SubBytesIns_Inst_Sbox_11_T4 ;
    wire SubBytesIns_Inst_Sbox_11_T3 ;
    wire SubBytesIns_Inst_Sbox_11_T2 ;
    wire SubBytesIns_Inst_Sbox_11_T1 ;
    wire SubBytesIns_Inst_Sbox_12_L29 ;
    wire SubBytesIns_Inst_Sbox_12_L28 ;
    wire SubBytesIns_Inst_Sbox_12_L27 ;
    wire SubBytesIns_Inst_Sbox_12_L26 ;
    wire SubBytesIns_Inst_Sbox_12_L25 ;
    wire SubBytesIns_Inst_Sbox_12_L24 ;
    wire SubBytesIns_Inst_Sbox_12_L23 ;
    wire SubBytesIns_Inst_Sbox_12_L22 ;
    wire SubBytesIns_Inst_Sbox_12_L21 ;
    wire SubBytesIns_Inst_Sbox_12_L20 ;
    wire SubBytesIns_Inst_Sbox_12_L19 ;
    wire SubBytesIns_Inst_Sbox_12_L18 ;
    wire SubBytesIns_Inst_Sbox_12_L17 ;
    wire SubBytesIns_Inst_Sbox_12_L16 ;
    wire SubBytesIns_Inst_Sbox_12_L15 ;
    wire SubBytesIns_Inst_Sbox_12_L14 ;
    wire SubBytesIns_Inst_Sbox_12_L13 ;
    wire SubBytesIns_Inst_Sbox_12_L12 ;
    wire SubBytesIns_Inst_Sbox_12_L11 ;
    wire SubBytesIns_Inst_Sbox_12_L10 ;
    wire SubBytesIns_Inst_Sbox_12_L9 ;
    wire SubBytesIns_Inst_Sbox_12_L8 ;
    wire SubBytesIns_Inst_Sbox_12_L7 ;
    wire SubBytesIns_Inst_Sbox_12_L6 ;
    wire SubBytesIns_Inst_Sbox_12_L5 ;
    wire SubBytesIns_Inst_Sbox_12_L4 ;
    wire SubBytesIns_Inst_Sbox_12_L3 ;
    wire SubBytesIns_Inst_Sbox_12_L2 ;
    wire SubBytesIns_Inst_Sbox_12_L1 ;
    wire SubBytesIns_Inst_Sbox_12_L0 ;
    wire SubBytesIns_Inst_Sbox_12_M63 ;
    wire SubBytesIns_Inst_Sbox_12_M62 ;
    wire SubBytesIns_Inst_Sbox_12_M61 ;
    wire SubBytesIns_Inst_Sbox_12_M60 ;
    wire SubBytesIns_Inst_Sbox_12_M59 ;
    wire SubBytesIns_Inst_Sbox_12_M58 ;
    wire SubBytesIns_Inst_Sbox_12_M57 ;
    wire SubBytesIns_Inst_Sbox_12_M56 ;
    wire SubBytesIns_Inst_Sbox_12_M55 ;
    wire SubBytesIns_Inst_Sbox_12_M54 ;
    wire SubBytesIns_Inst_Sbox_12_M53 ;
    wire SubBytesIns_Inst_Sbox_12_M52 ;
    wire SubBytesIns_Inst_Sbox_12_M51 ;
    wire SubBytesIns_Inst_Sbox_12_M50 ;
    wire SubBytesIns_Inst_Sbox_12_M49 ;
    wire SubBytesIns_Inst_Sbox_12_M48 ;
    wire SubBytesIns_Inst_Sbox_12_M47 ;
    wire SubBytesIns_Inst_Sbox_12_M46 ;
    wire SubBytesIns_Inst_Sbox_12_M45 ;
    wire SubBytesIns_Inst_Sbox_12_M44 ;
    wire SubBytesIns_Inst_Sbox_12_M43 ;
    wire SubBytesIns_Inst_Sbox_12_M42 ;
    wire SubBytesIns_Inst_Sbox_12_M41 ;
    wire SubBytesIns_Inst_Sbox_12_M40 ;
    wire SubBytesIns_Inst_Sbox_12_M39 ;
    wire SubBytesIns_Inst_Sbox_12_M38 ;
    wire SubBytesIns_Inst_Sbox_12_M37 ;
    wire SubBytesIns_Inst_Sbox_12_M36 ;
    wire SubBytesIns_Inst_Sbox_12_M35 ;
    wire SubBytesIns_Inst_Sbox_12_M34 ;
    wire SubBytesIns_Inst_Sbox_12_M33 ;
    wire SubBytesIns_Inst_Sbox_12_M32 ;
    wire SubBytesIns_Inst_Sbox_12_M31 ;
    wire SubBytesIns_Inst_Sbox_12_M30 ;
    wire SubBytesIns_Inst_Sbox_12_M29 ;
    wire SubBytesIns_Inst_Sbox_12_M28 ;
    wire SubBytesIns_Inst_Sbox_12_M27 ;
    wire SubBytesIns_Inst_Sbox_12_M26 ;
    wire SubBytesIns_Inst_Sbox_12_M25 ;
    wire SubBytesIns_Inst_Sbox_12_M24 ;
    wire SubBytesIns_Inst_Sbox_12_M23 ;
    wire SubBytesIns_Inst_Sbox_12_M22 ;
    wire SubBytesIns_Inst_Sbox_12_M21 ;
    wire SubBytesIns_Inst_Sbox_12_M20 ;
    wire SubBytesIns_Inst_Sbox_12_M19 ;
    wire SubBytesIns_Inst_Sbox_12_M18 ;
    wire SubBytesIns_Inst_Sbox_12_M17 ;
    wire SubBytesIns_Inst_Sbox_12_M16 ;
    wire SubBytesIns_Inst_Sbox_12_M15 ;
    wire SubBytesIns_Inst_Sbox_12_M14 ;
    wire SubBytesIns_Inst_Sbox_12_M13 ;
    wire SubBytesIns_Inst_Sbox_12_M12 ;
    wire SubBytesIns_Inst_Sbox_12_M11 ;
    wire SubBytesIns_Inst_Sbox_12_M10 ;
    wire SubBytesIns_Inst_Sbox_12_M9 ;
    wire SubBytesIns_Inst_Sbox_12_M8 ;
    wire SubBytesIns_Inst_Sbox_12_M7 ;
    wire SubBytesIns_Inst_Sbox_12_M6 ;
    wire SubBytesIns_Inst_Sbox_12_M5 ;
    wire SubBytesIns_Inst_Sbox_12_M4 ;
    wire SubBytesIns_Inst_Sbox_12_M3 ;
    wire SubBytesIns_Inst_Sbox_12_M2 ;
    wire SubBytesIns_Inst_Sbox_12_M1 ;
    wire SubBytesIns_Inst_Sbox_12_T27 ;
    wire SubBytesIns_Inst_Sbox_12_T26 ;
    wire SubBytesIns_Inst_Sbox_12_T25 ;
    wire SubBytesIns_Inst_Sbox_12_T24 ;
    wire SubBytesIns_Inst_Sbox_12_T23 ;
    wire SubBytesIns_Inst_Sbox_12_T22 ;
    wire SubBytesIns_Inst_Sbox_12_T21 ;
    wire SubBytesIns_Inst_Sbox_12_T20 ;
    wire SubBytesIns_Inst_Sbox_12_T19 ;
    wire SubBytesIns_Inst_Sbox_12_T18 ;
    wire SubBytesIns_Inst_Sbox_12_T17 ;
    wire SubBytesIns_Inst_Sbox_12_T16 ;
    wire SubBytesIns_Inst_Sbox_12_T15 ;
    wire SubBytesIns_Inst_Sbox_12_T14 ;
    wire SubBytesIns_Inst_Sbox_12_T13 ;
    wire SubBytesIns_Inst_Sbox_12_T12 ;
    wire SubBytesIns_Inst_Sbox_12_T11 ;
    wire SubBytesIns_Inst_Sbox_12_T10 ;
    wire SubBytesIns_Inst_Sbox_12_T9 ;
    wire SubBytesIns_Inst_Sbox_12_T8 ;
    wire SubBytesIns_Inst_Sbox_12_T7 ;
    wire SubBytesIns_Inst_Sbox_12_T6 ;
    wire SubBytesIns_Inst_Sbox_12_T5 ;
    wire SubBytesIns_Inst_Sbox_12_T4 ;
    wire SubBytesIns_Inst_Sbox_12_T3 ;
    wire SubBytesIns_Inst_Sbox_12_T2 ;
    wire SubBytesIns_Inst_Sbox_12_T1 ;
    wire SubBytesIns_Inst_Sbox_13_L29 ;
    wire SubBytesIns_Inst_Sbox_13_L28 ;
    wire SubBytesIns_Inst_Sbox_13_L27 ;
    wire SubBytesIns_Inst_Sbox_13_L26 ;
    wire SubBytesIns_Inst_Sbox_13_L25 ;
    wire SubBytesIns_Inst_Sbox_13_L24 ;
    wire SubBytesIns_Inst_Sbox_13_L23 ;
    wire SubBytesIns_Inst_Sbox_13_L22 ;
    wire SubBytesIns_Inst_Sbox_13_L21 ;
    wire SubBytesIns_Inst_Sbox_13_L20 ;
    wire SubBytesIns_Inst_Sbox_13_L19 ;
    wire SubBytesIns_Inst_Sbox_13_L18 ;
    wire SubBytesIns_Inst_Sbox_13_L17 ;
    wire SubBytesIns_Inst_Sbox_13_L16 ;
    wire SubBytesIns_Inst_Sbox_13_L15 ;
    wire SubBytesIns_Inst_Sbox_13_L14 ;
    wire SubBytesIns_Inst_Sbox_13_L13 ;
    wire SubBytesIns_Inst_Sbox_13_L12 ;
    wire SubBytesIns_Inst_Sbox_13_L11 ;
    wire SubBytesIns_Inst_Sbox_13_L10 ;
    wire SubBytesIns_Inst_Sbox_13_L9 ;
    wire SubBytesIns_Inst_Sbox_13_L8 ;
    wire SubBytesIns_Inst_Sbox_13_L7 ;
    wire SubBytesIns_Inst_Sbox_13_L6 ;
    wire SubBytesIns_Inst_Sbox_13_L5 ;
    wire SubBytesIns_Inst_Sbox_13_L4 ;
    wire SubBytesIns_Inst_Sbox_13_L3 ;
    wire SubBytesIns_Inst_Sbox_13_L2 ;
    wire SubBytesIns_Inst_Sbox_13_L1 ;
    wire SubBytesIns_Inst_Sbox_13_L0 ;
    wire SubBytesIns_Inst_Sbox_13_M63 ;
    wire SubBytesIns_Inst_Sbox_13_M62 ;
    wire SubBytesIns_Inst_Sbox_13_M61 ;
    wire SubBytesIns_Inst_Sbox_13_M60 ;
    wire SubBytesIns_Inst_Sbox_13_M59 ;
    wire SubBytesIns_Inst_Sbox_13_M58 ;
    wire SubBytesIns_Inst_Sbox_13_M57 ;
    wire SubBytesIns_Inst_Sbox_13_M56 ;
    wire SubBytesIns_Inst_Sbox_13_M55 ;
    wire SubBytesIns_Inst_Sbox_13_M54 ;
    wire SubBytesIns_Inst_Sbox_13_M53 ;
    wire SubBytesIns_Inst_Sbox_13_M52 ;
    wire SubBytesIns_Inst_Sbox_13_M51 ;
    wire SubBytesIns_Inst_Sbox_13_M50 ;
    wire SubBytesIns_Inst_Sbox_13_M49 ;
    wire SubBytesIns_Inst_Sbox_13_M48 ;
    wire SubBytesIns_Inst_Sbox_13_M47 ;
    wire SubBytesIns_Inst_Sbox_13_M46 ;
    wire SubBytesIns_Inst_Sbox_13_M45 ;
    wire SubBytesIns_Inst_Sbox_13_M44 ;
    wire SubBytesIns_Inst_Sbox_13_M43 ;
    wire SubBytesIns_Inst_Sbox_13_M42 ;
    wire SubBytesIns_Inst_Sbox_13_M41 ;
    wire SubBytesIns_Inst_Sbox_13_M40 ;
    wire SubBytesIns_Inst_Sbox_13_M39 ;
    wire SubBytesIns_Inst_Sbox_13_M38 ;
    wire SubBytesIns_Inst_Sbox_13_M37 ;
    wire SubBytesIns_Inst_Sbox_13_M36 ;
    wire SubBytesIns_Inst_Sbox_13_M35 ;
    wire SubBytesIns_Inst_Sbox_13_M34 ;
    wire SubBytesIns_Inst_Sbox_13_M33 ;
    wire SubBytesIns_Inst_Sbox_13_M32 ;
    wire SubBytesIns_Inst_Sbox_13_M31 ;
    wire SubBytesIns_Inst_Sbox_13_M30 ;
    wire SubBytesIns_Inst_Sbox_13_M29 ;
    wire SubBytesIns_Inst_Sbox_13_M28 ;
    wire SubBytesIns_Inst_Sbox_13_M27 ;
    wire SubBytesIns_Inst_Sbox_13_M26 ;
    wire SubBytesIns_Inst_Sbox_13_M25 ;
    wire SubBytesIns_Inst_Sbox_13_M24 ;
    wire SubBytesIns_Inst_Sbox_13_M23 ;
    wire SubBytesIns_Inst_Sbox_13_M22 ;
    wire SubBytesIns_Inst_Sbox_13_M21 ;
    wire SubBytesIns_Inst_Sbox_13_M20 ;
    wire SubBytesIns_Inst_Sbox_13_M19 ;
    wire SubBytesIns_Inst_Sbox_13_M18 ;
    wire SubBytesIns_Inst_Sbox_13_M17 ;
    wire SubBytesIns_Inst_Sbox_13_M16 ;
    wire SubBytesIns_Inst_Sbox_13_M15 ;
    wire SubBytesIns_Inst_Sbox_13_M14 ;
    wire SubBytesIns_Inst_Sbox_13_M13 ;
    wire SubBytesIns_Inst_Sbox_13_M12 ;
    wire SubBytesIns_Inst_Sbox_13_M11 ;
    wire SubBytesIns_Inst_Sbox_13_M10 ;
    wire SubBytesIns_Inst_Sbox_13_M9 ;
    wire SubBytesIns_Inst_Sbox_13_M8 ;
    wire SubBytesIns_Inst_Sbox_13_M7 ;
    wire SubBytesIns_Inst_Sbox_13_M6 ;
    wire SubBytesIns_Inst_Sbox_13_M5 ;
    wire SubBytesIns_Inst_Sbox_13_M4 ;
    wire SubBytesIns_Inst_Sbox_13_M3 ;
    wire SubBytesIns_Inst_Sbox_13_M2 ;
    wire SubBytesIns_Inst_Sbox_13_M1 ;
    wire SubBytesIns_Inst_Sbox_13_T27 ;
    wire SubBytesIns_Inst_Sbox_13_T26 ;
    wire SubBytesIns_Inst_Sbox_13_T25 ;
    wire SubBytesIns_Inst_Sbox_13_T24 ;
    wire SubBytesIns_Inst_Sbox_13_T23 ;
    wire SubBytesIns_Inst_Sbox_13_T22 ;
    wire SubBytesIns_Inst_Sbox_13_T21 ;
    wire SubBytesIns_Inst_Sbox_13_T20 ;
    wire SubBytesIns_Inst_Sbox_13_T19 ;
    wire SubBytesIns_Inst_Sbox_13_T18 ;
    wire SubBytesIns_Inst_Sbox_13_T17 ;
    wire SubBytesIns_Inst_Sbox_13_T16 ;
    wire SubBytesIns_Inst_Sbox_13_T15 ;
    wire SubBytesIns_Inst_Sbox_13_T14 ;
    wire SubBytesIns_Inst_Sbox_13_T13 ;
    wire SubBytesIns_Inst_Sbox_13_T12 ;
    wire SubBytesIns_Inst_Sbox_13_T11 ;
    wire SubBytesIns_Inst_Sbox_13_T10 ;
    wire SubBytesIns_Inst_Sbox_13_T9 ;
    wire SubBytesIns_Inst_Sbox_13_T8 ;
    wire SubBytesIns_Inst_Sbox_13_T7 ;
    wire SubBytesIns_Inst_Sbox_13_T6 ;
    wire SubBytesIns_Inst_Sbox_13_T5 ;
    wire SubBytesIns_Inst_Sbox_13_T4 ;
    wire SubBytesIns_Inst_Sbox_13_T3 ;
    wire SubBytesIns_Inst_Sbox_13_T2 ;
    wire SubBytesIns_Inst_Sbox_13_T1 ;
    wire SubBytesIns_Inst_Sbox_14_L29 ;
    wire SubBytesIns_Inst_Sbox_14_L28 ;
    wire SubBytesIns_Inst_Sbox_14_L27 ;
    wire SubBytesIns_Inst_Sbox_14_L26 ;
    wire SubBytesIns_Inst_Sbox_14_L25 ;
    wire SubBytesIns_Inst_Sbox_14_L24 ;
    wire SubBytesIns_Inst_Sbox_14_L23 ;
    wire SubBytesIns_Inst_Sbox_14_L22 ;
    wire SubBytesIns_Inst_Sbox_14_L21 ;
    wire SubBytesIns_Inst_Sbox_14_L20 ;
    wire SubBytesIns_Inst_Sbox_14_L19 ;
    wire SubBytesIns_Inst_Sbox_14_L18 ;
    wire SubBytesIns_Inst_Sbox_14_L17 ;
    wire SubBytesIns_Inst_Sbox_14_L16 ;
    wire SubBytesIns_Inst_Sbox_14_L15 ;
    wire SubBytesIns_Inst_Sbox_14_L14 ;
    wire SubBytesIns_Inst_Sbox_14_L13 ;
    wire SubBytesIns_Inst_Sbox_14_L12 ;
    wire SubBytesIns_Inst_Sbox_14_L11 ;
    wire SubBytesIns_Inst_Sbox_14_L10 ;
    wire SubBytesIns_Inst_Sbox_14_L9 ;
    wire SubBytesIns_Inst_Sbox_14_L8 ;
    wire SubBytesIns_Inst_Sbox_14_L7 ;
    wire SubBytesIns_Inst_Sbox_14_L6 ;
    wire SubBytesIns_Inst_Sbox_14_L5 ;
    wire SubBytesIns_Inst_Sbox_14_L4 ;
    wire SubBytesIns_Inst_Sbox_14_L3 ;
    wire SubBytesIns_Inst_Sbox_14_L2 ;
    wire SubBytesIns_Inst_Sbox_14_L1 ;
    wire SubBytesIns_Inst_Sbox_14_L0 ;
    wire SubBytesIns_Inst_Sbox_14_M63 ;
    wire SubBytesIns_Inst_Sbox_14_M62 ;
    wire SubBytesIns_Inst_Sbox_14_M61 ;
    wire SubBytesIns_Inst_Sbox_14_M60 ;
    wire SubBytesIns_Inst_Sbox_14_M59 ;
    wire SubBytesIns_Inst_Sbox_14_M58 ;
    wire SubBytesIns_Inst_Sbox_14_M57 ;
    wire SubBytesIns_Inst_Sbox_14_M56 ;
    wire SubBytesIns_Inst_Sbox_14_M55 ;
    wire SubBytesIns_Inst_Sbox_14_M54 ;
    wire SubBytesIns_Inst_Sbox_14_M53 ;
    wire SubBytesIns_Inst_Sbox_14_M52 ;
    wire SubBytesIns_Inst_Sbox_14_M51 ;
    wire SubBytesIns_Inst_Sbox_14_M50 ;
    wire SubBytesIns_Inst_Sbox_14_M49 ;
    wire SubBytesIns_Inst_Sbox_14_M48 ;
    wire SubBytesIns_Inst_Sbox_14_M47 ;
    wire SubBytesIns_Inst_Sbox_14_M46 ;
    wire SubBytesIns_Inst_Sbox_14_M45 ;
    wire SubBytesIns_Inst_Sbox_14_M44 ;
    wire SubBytesIns_Inst_Sbox_14_M43 ;
    wire SubBytesIns_Inst_Sbox_14_M42 ;
    wire SubBytesIns_Inst_Sbox_14_M41 ;
    wire SubBytesIns_Inst_Sbox_14_M40 ;
    wire SubBytesIns_Inst_Sbox_14_M39 ;
    wire SubBytesIns_Inst_Sbox_14_M38 ;
    wire SubBytesIns_Inst_Sbox_14_M37 ;
    wire SubBytesIns_Inst_Sbox_14_M36 ;
    wire SubBytesIns_Inst_Sbox_14_M35 ;
    wire SubBytesIns_Inst_Sbox_14_M34 ;
    wire SubBytesIns_Inst_Sbox_14_M33 ;
    wire SubBytesIns_Inst_Sbox_14_M32 ;
    wire SubBytesIns_Inst_Sbox_14_M31 ;
    wire SubBytesIns_Inst_Sbox_14_M30 ;
    wire SubBytesIns_Inst_Sbox_14_M29 ;
    wire SubBytesIns_Inst_Sbox_14_M28 ;
    wire SubBytesIns_Inst_Sbox_14_M27 ;
    wire SubBytesIns_Inst_Sbox_14_M26 ;
    wire SubBytesIns_Inst_Sbox_14_M25 ;
    wire SubBytesIns_Inst_Sbox_14_M24 ;
    wire SubBytesIns_Inst_Sbox_14_M23 ;
    wire SubBytesIns_Inst_Sbox_14_M22 ;
    wire SubBytesIns_Inst_Sbox_14_M21 ;
    wire SubBytesIns_Inst_Sbox_14_M20 ;
    wire SubBytesIns_Inst_Sbox_14_M19 ;
    wire SubBytesIns_Inst_Sbox_14_M18 ;
    wire SubBytesIns_Inst_Sbox_14_M17 ;
    wire SubBytesIns_Inst_Sbox_14_M16 ;
    wire SubBytesIns_Inst_Sbox_14_M15 ;
    wire SubBytesIns_Inst_Sbox_14_M14 ;
    wire SubBytesIns_Inst_Sbox_14_M13 ;
    wire SubBytesIns_Inst_Sbox_14_M12 ;
    wire SubBytesIns_Inst_Sbox_14_M11 ;
    wire SubBytesIns_Inst_Sbox_14_M10 ;
    wire SubBytesIns_Inst_Sbox_14_M9 ;
    wire SubBytesIns_Inst_Sbox_14_M8 ;
    wire SubBytesIns_Inst_Sbox_14_M7 ;
    wire SubBytesIns_Inst_Sbox_14_M6 ;
    wire SubBytesIns_Inst_Sbox_14_M5 ;
    wire SubBytesIns_Inst_Sbox_14_M4 ;
    wire SubBytesIns_Inst_Sbox_14_M3 ;
    wire SubBytesIns_Inst_Sbox_14_M2 ;
    wire SubBytesIns_Inst_Sbox_14_M1 ;
    wire SubBytesIns_Inst_Sbox_14_T27 ;
    wire SubBytesIns_Inst_Sbox_14_T26 ;
    wire SubBytesIns_Inst_Sbox_14_T25 ;
    wire SubBytesIns_Inst_Sbox_14_T24 ;
    wire SubBytesIns_Inst_Sbox_14_T23 ;
    wire SubBytesIns_Inst_Sbox_14_T22 ;
    wire SubBytesIns_Inst_Sbox_14_T21 ;
    wire SubBytesIns_Inst_Sbox_14_T20 ;
    wire SubBytesIns_Inst_Sbox_14_T19 ;
    wire SubBytesIns_Inst_Sbox_14_T18 ;
    wire SubBytesIns_Inst_Sbox_14_T17 ;
    wire SubBytesIns_Inst_Sbox_14_T16 ;
    wire SubBytesIns_Inst_Sbox_14_T15 ;
    wire SubBytesIns_Inst_Sbox_14_T14 ;
    wire SubBytesIns_Inst_Sbox_14_T13 ;
    wire SubBytesIns_Inst_Sbox_14_T12 ;
    wire SubBytesIns_Inst_Sbox_14_T11 ;
    wire SubBytesIns_Inst_Sbox_14_T10 ;
    wire SubBytesIns_Inst_Sbox_14_T9 ;
    wire SubBytesIns_Inst_Sbox_14_T8 ;
    wire SubBytesIns_Inst_Sbox_14_T7 ;
    wire SubBytesIns_Inst_Sbox_14_T6 ;
    wire SubBytesIns_Inst_Sbox_14_T5 ;
    wire SubBytesIns_Inst_Sbox_14_T4 ;
    wire SubBytesIns_Inst_Sbox_14_T3 ;
    wire SubBytesIns_Inst_Sbox_14_T2 ;
    wire SubBytesIns_Inst_Sbox_14_T1 ;
    wire SubBytesIns_Inst_Sbox_15_L29 ;
    wire SubBytesIns_Inst_Sbox_15_L28 ;
    wire SubBytesIns_Inst_Sbox_15_L27 ;
    wire SubBytesIns_Inst_Sbox_15_L26 ;
    wire SubBytesIns_Inst_Sbox_15_L25 ;
    wire SubBytesIns_Inst_Sbox_15_L24 ;
    wire SubBytesIns_Inst_Sbox_15_L23 ;
    wire SubBytesIns_Inst_Sbox_15_L22 ;
    wire SubBytesIns_Inst_Sbox_15_L21 ;
    wire SubBytesIns_Inst_Sbox_15_L20 ;
    wire SubBytesIns_Inst_Sbox_15_L19 ;
    wire SubBytesIns_Inst_Sbox_15_L18 ;
    wire SubBytesIns_Inst_Sbox_15_L17 ;
    wire SubBytesIns_Inst_Sbox_15_L16 ;
    wire SubBytesIns_Inst_Sbox_15_L15 ;
    wire SubBytesIns_Inst_Sbox_15_L14 ;
    wire SubBytesIns_Inst_Sbox_15_L13 ;
    wire SubBytesIns_Inst_Sbox_15_L12 ;
    wire SubBytesIns_Inst_Sbox_15_L11 ;
    wire SubBytesIns_Inst_Sbox_15_L10 ;
    wire SubBytesIns_Inst_Sbox_15_L9 ;
    wire SubBytesIns_Inst_Sbox_15_L8 ;
    wire SubBytesIns_Inst_Sbox_15_L7 ;
    wire SubBytesIns_Inst_Sbox_15_L6 ;
    wire SubBytesIns_Inst_Sbox_15_L5 ;
    wire SubBytesIns_Inst_Sbox_15_L4 ;
    wire SubBytesIns_Inst_Sbox_15_L3 ;
    wire SubBytesIns_Inst_Sbox_15_L2 ;
    wire SubBytesIns_Inst_Sbox_15_L1 ;
    wire SubBytesIns_Inst_Sbox_15_L0 ;
    wire SubBytesIns_Inst_Sbox_15_M63 ;
    wire SubBytesIns_Inst_Sbox_15_M62 ;
    wire SubBytesIns_Inst_Sbox_15_M61 ;
    wire SubBytesIns_Inst_Sbox_15_M60 ;
    wire SubBytesIns_Inst_Sbox_15_M59 ;
    wire SubBytesIns_Inst_Sbox_15_M58 ;
    wire SubBytesIns_Inst_Sbox_15_M57 ;
    wire SubBytesIns_Inst_Sbox_15_M56 ;
    wire SubBytesIns_Inst_Sbox_15_M55 ;
    wire SubBytesIns_Inst_Sbox_15_M54 ;
    wire SubBytesIns_Inst_Sbox_15_M53 ;
    wire SubBytesIns_Inst_Sbox_15_M52 ;
    wire SubBytesIns_Inst_Sbox_15_M51 ;
    wire SubBytesIns_Inst_Sbox_15_M50 ;
    wire SubBytesIns_Inst_Sbox_15_M49 ;
    wire SubBytesIns_Inst_Sbox_15_M48 ;
    wire SubBytesIns_Inst_Sbox_15_M47 ;
    wire SubBytesIns_Inst_Sbox_15_M46 ;
    wire SubBytesIns_Inst_Sbox_15_M45 ;
    wire SubBytesIns_Inst_Sbox_15_M44 ;
    wire SubBytesIns_Inst_Sbox_15_M43 ;
    wire SubBytesIns_Inst_Sbox_15_M42 ;
    wire SubBytesIns_Inst_Sbox_15_M41 ;
    wire SubBytesIns_Inst_Sbox_15_M40 ;
    wire SubBytesIns_Inst_Sbox_15_M39 ;
    wire SubBytesIns_Inst_Sbox_15_M38 ;
    wire SubBytesIns_Inst_Sbox_15_M37 ;
    wire SubBytesIns_Inst_Sbox_15_M36 ;
    wire SubBytesIns_Inst_Sbox_15_M35 ;
    wire SubBytesIns_Inst_Sbox_15_M34 ;
    wire SubBytesIns_Inst_Sbox_15_M33 ;
    wire SubBytesIns_Inst_Sbox_15_M32 ;
    wire SubBytesIns_Inst_Sbox_15_M31 ;
    wire SubBytesIns_Inst_Sbox_15_M30 ;
    wire SubBytesIns_Inst_Sbox_15_M29 ;
    wire SubBytesIns_Inst_Sbox_15_M28 ;
    wire SubBytesIns_Inst_Sbox_15_M27 ;
    wire SubBytesIns_Inst_Sbox_15_M26 ;
    wire SubBytesIns_Inst_Sbox_15_M25 ;
    wire SubBytesIns_Inst_Sbox_15_M24 ;
    wire SubBytesIns_Inst_Sbox_15_M23 ;
    wire SubBytesIns_Inst_Sbox_15_M22 ;
    wire SubBytesIns_Inst_Sbox_15_M21 ;
    wire SubBytesIns_Inst_Sbox_15_M20 ;
    wire SubBytesIns_Inst_Sbox_15_M19 ;
    wire SubBytesIns_Inst_Sbox_15_M18 ;
    wire SubBytesIns_Inst_Sbox_15_M17 ;
    wire SubBytesIns_Inst_Sbox_15_M16 ;
    wire SubBytesIns_Inst_Sbox_15_M15 ;
    wire SubBytesIns_Inst_Sbox_15_M14 ;
    wire SubBytesIns_Inst_Sbox_15_M13 ;
    wire SubBytesIns_Inst_Sbox_15_M12 ;
    wire SubBytesIns_Inst_Sbox_15_M11 ;
    wire SubBytesIns_Inst_Sbox_15_M10 ;
    wire SubBytesIns_Inst_Sbox_15_M9 ;
    wire SubBytesIns_Inst_Sbox_15_M8 ;
    wire SubBytesIns_Inst_Sbox_15_M7 ;
    wire SubBytesIns_Inst_Sbox_15_M6 ;
    wire SubBytesIns_Inst_Sbox_15_M5 ;
    wire SubBytesIns_Inst_Sbox_15_M4 ;
    wire SubBytesIns_Inst_Sbox_15_M3 ;
    wire SubBytesIns_Inst_Sbox_15_M2 ;
    wire SubBytesIns_Inst_Sbox_15_M1 ;
    wire SubBytesIns_Inst_Sbox_15_T27 ;
    wire SubBytesIns_Inst_Sbox_15_T26 ;
    wire SubBytesIns_Inst_Sbox_15_T25 ;
    wire SubBytesIns_Inst_Sbox_15_T24 ;
    wire SubBytesIns_Inst_Sbox_15_T23 ;
    wire SubBytesIns_Inst_Sbox_15_T22 ;
    wire SubBytesIns_Inst_Sbox_15_T21 ;
    wire SubBytesIns_Inst_Sbox_15_T20 ;
    wire SubBytesIns_Inst_Sbox_15_T19 ;
    wire SubBytesIns_Inst_Sbox_15_T18 ;
    wire SubBytesIns_Inst_Sbox_15_T17 ;
    wire SubBytesIns_Inst_Sbox_15_T16 ;
    wire SubBytesIns_Inst_Sbox_15_T15 ;
    wire SubBytesIns_Inst_Sbox_15_T14 ;
    wire SubBytesIns_Inst_Sbox_15_T13 ;
    wire SubBytesIns_Inst_Sbox_15_T12 ;
    wire SubBytesIns_Inst_Sbox_15_T11 ;
    wire SubBytesIns_Inst_Sbox_15_T10 ;
    wire SubBytesIns_Inst_Sbox_15_T9 ;
    wire SubBytesIns_Inst_Sbox_15_T8 ;
    wire SubBytesIns_Inst_Sbox_15_T7 ;
    wire SubBytesIns_Inst_Sbox_15_T6 ;
    wire SubBytesIns_Inst_Sbox_15_T5 ;
    wire SubBytesIns_Inst_Sbox_15_T4 ;
    wire SubBytesIns_Inst_Sbox_15_T3 ;
    wire SubBytesIns_Inst_Sbox_15_T2 ;
    wire SubBytesIns_Inst_Sbox_15_T1 ;
    wire MixColumnsIns_MixOneColumnInst_0_n64 ;
    wire MixColumnsIns_MixOneColumnInst_0_n63 ;
    wire MixColumnsIns_MixOneColumnInst_0_n62 ;
    wire MixColumnsIns_MixOneColumnInst_0_n61 ;
    wire MixColumnsIns_MixOneColumnInst_0_n60 ;
    wire MixColumnsIns_MixOneColumnInst_0_n59 ;
    wire MixColumnsIns_MixOneColumnInst_0_n58 ;
    wire MixColumnsIns_MixOneColumnInst_0_n57 ;
    wire MixColumnsIns_MixOneColumnInst_0_n56 ;
    wire MixColumnsIns_MixOneColumnInst_0_n55 ;
    wire MixColumnsIns_MixOneColumnInst_0_n54 ;
    wire MixColumnsIns_MixOneColumnInst_0_n53 ;
    wire MixColumnsIns_MixOneColumnInst_0_n52 ;
    wire MixColumnsIns_MixOneColumnInst_0_n51 ;
    wire MixColumnsIns_MixOneColumnInst_0_n50 ;
    wire MixColumnsIns_MixOneColumnInst_0_n49 ;
    wire MixColumnsIns_MixOneColumnInst_0_n48 ;
    wire MixColumnsIns_MixOneColumnInst_0_n47 ;
    wire MixColumnsIns_MixOneColumnInst_0_n46 ;
    wire MixColumnsIns_MixOneColumnInst_0_n45 ;
    wire MixColumnsIns_MixOneColumnInst_0_n44 ;
    wire MixColumnsIns_MixOneColumnInst_0_n43 ;
    wire MixColumnsIns_MixOneColumnInst_0_n42 ;
    wire MixColumnsIns_MixOneColumnInst_0_n41 ;
    wire MixColumnsIns_MixOneColumnInst_0_n40 ;
    wire MixColumnsIns_MixOneColumnInst_0_n39 ;
    wire MixColumnsIns_MixOneColumnInst_0_n38 ;
    wire MixColumnsIns_MixOneColumnInst_0_n37 ;
    wire MixColumnsIns_MixOneColumnInst_0_n36 ;
    wire MixColumnsIns_MixOneColumnInst_0_n35 ;
    wire MixColumnsIns_MixOneColumnInst_0_n34 ;
    wire MixColumnsIns_MixOneColumnInst_0_n33 ;
    wire MixColumnsIns_MixOneColumnInst_0_n32 ;
    wire MixColumnsIns_MixOneColumnInst_0_n31 ;
    wire MixColumnsIns_MixOneColumnInst_0_n30 ;
    wire MixColumnsIns_MixOneColumnInst_0_n29 ;
    wire MixColumnsIns_MixOneColumnInst_0_n28 ;
    wire MixColumnsIns_MixOneColumnInst_0_n27 ;
    wire MixColumnsIns_MixOneColumnInst_0_n26 ;
    wire MixColumnsIns_MixOneColumnInst_0_n25 ;
    wire MixColumnsIns_MixOneColumnInst_0_n24 ;
    wire MixColumnsIns_MixOneColumnInst_0_n23 ;
    wire MixColumnsIns_MixOneColumnInst_0_n22 ;
    wire MixColumnsIns_MixOneColumnInst_0_n21 ;
    wire MixColumnsIns_MixOneColumnInst_0_n20 ;
    wire MixColumnsIns_MixOneColumnInst_0_n19 ;
    wire MixColumnsIns_MixOneColumnInst_0_n18 ;
    wire MixColumnsIns_MixOneColumnInst_0_n17 ;
    wire MixColumnsIns_MixOneColumnInst_0_n16 ;
    wire MixColumnsIns_MixOneColumnInst_0_n15 ;
    wire MixColumnsIns_MixOneColumnInst_0_n14 ;
    wire MixColumnsIns_MixOneColumnInst_0_n13 ;
    wire MixColumnsIns_MixOneColumnInst_0_n12 ;
    wire MixColumnsIns_MixOneColumnInst_0_n11 ;
    wire MixColumnsIns_MixOneColumnInst_0_n10 ;
    wire MixColumnsIns_MixOneColumnInst_0_n9 ;
    wire MixColumnsIns_MixOneColumnInst_0_n8 ;
    wire MixColumnsIns_MixOneColumnInst_0_n7 ;
    wire MixColumnsIns_MixOneColumnInst_0_n6 ;
    wire MixColumnsIns_MixOneColumnInst_0_n5 ;
    wire MixColumnsIns_MixOneColumnInst_0_n4 ;
    wire MixColumnsIns_MixOneColumnInst_0_n3 ;
    wire MixColumnsIns_MixOneColumnInst_0_n2 ;
    wire MixColumnsIns_MixOneColumnInst_0_n1 ;
    wire MixColumnsIns_MixOneColumnInst_1_n64 ;
    wire MixColumnsIns_MixOneColumnInst_1_n63 ;
    wire MixColumnsIns_MixOneColumnInst_1_n62 ;
    wire MixColumnsIns_MixOneColumnInst_1_n61 ;
    wire MixColumnsIns_MixOneColumnInst_1_n60 ;
    wire MixColumnsIns_MixOneColumnInst_1_n59 ;
    wire MixColumnsIns_MixOneColumnInst_1_n58 ;
    wire MixColumnsIns_MixOneColumnInst_1_n57 ;
    wire MixColumnsIns_MixOneColumnInst_1_n56 ;
    wire MixColumnsIns_MixOneColumnInst_1_n55 ;
    wire MixColumnsIns_MixOneColumnInst_1_n54 ;
    wire MixColumnsIns_MixOneColumnInst_1_n53 ;
    wire MixColumnsIns_MixOneColumnInst_1_n52 ;
    wire MixColumnsIns_MixOneColumnInst_1_n51 ;
    wire MixColumnsIns_MixOneColumnInst_1_n50 ;
    wire MixColumnsIns_MixOneColumnInst_1_n49 ;
    wire MixColumnsIns_MixOneColumnInst_1_n48 ;
    wire MixColumnsIns_MixOneColumnInst_1_n47 ;
    wire MixColumnsIns_MixOneColumnInst_1_n46 ;
    wire MixColumnsIns_MixOneColumnInst_1_n45 ;
    wire MixColumnsIns_MixOneColumnInst_1_n44 ;
    wire MixColumnsIns_MixOneColumnInst_1_n43 ;
    wire MixColumnsIns_MixOneColumnInst_1_n42 ;
    wire MixColumnsIns_MixOneColumnInst_1_n41 ;
    wire MixColumnsIns_MixOneColumnInst_1_n40 ;
    wire MixColumnsIns_MixOneColumnInst_1_n39 ;
    wire MixColumnsIns_MixOneColumnInst_1_n38 ;
    wire MixColumnsIns_MixOneColumnInst_1_n37 ;
    wire MixColumnsIns_MixOneColumnInst_1_n36 ;
    wire MixColumnsIns_MixOneColumnInst_1_n35 ;
    wire MixColumnsIns_MixOneColumnInst_1_n34 ;
    wire MixColumnsIns_MixOneColumnInst_1_n33 ;
    wire MixColumnsIns_MixOneColumnInst_1_n32 ;
    wire MixColumnsIns_MixOneColumnInst_1_n31 ;
    wire MixColumnsIns_MixOneColumnInst_1_n30 ;
    wire MixColumnsIns_MixOneColumnInst_1_n29 ;
    wire MixColumnsIns_MixOneColumnInst_1_n28 ;
    wire MixColumnsIns_MixOneColumnInst_1_n27 ;
    wire MixColumnsIns_MixOneColumnInst_1_n26 ;
    wire MixColumnsIns_MixOneColumnInst_1_n25 ;
    wire MixColumnsIns_MixOneColumnInst_1_n24 ;
    wire MixColumnsIns_MixOneColumnInst_1_n23 ;
    wire MixColumnsIns_MixOneColumnInst_1_n22 ;
    wire MixColumnsIns_MixOneColumnInst_1_n21 ;
    wire MixColumnsIns_MixOneColumnInst_1_n20 ;
    wire MixColumnsIns_MixOneColumnInst_1_n19 ;
    wire MixColumnsIns_MixOneColumnInst_1_n18 ;
    wire MixColumnsIns_MixOneColumnInst_1_n17 ;
    wire MixColumnsIns_MixOneColumnInst_1_n16 ;
    wire MixColumnsIns_MixOneColumnInst_1_n15 ;
    wire MixColumnsIns_MixOneColumnInst_1_n14 ;
    wire MixColumnsIns_MixOneColumnInst_1_n13 ;
    wire MixColumnsIns_MixOneColumnInst_1_n12 ;
    wire MixColumnsIns_MixOneColumnInst_1_n11 ;
    wire MixColumnsIns_MixOneColumnInst_1_n10 ;
    wire MixColumnsIns_MixOneColumnInst_1_n9 ;
    wire MixColumnsIns_MixOneColumnInst_1_n8 ;
    wire MixColumnsIns_MixOneColumnInst_1_n7 ;
    wire MixColumnsIns_MixOneColumnInst_1_n6 ;
    wire MixColumnsIns_MixOneColumnInst_1_n5 ;
    wire MixColumnsIns_MixOneColumnInst_1_n4 ;
    wire MixColumnsIns_MixOneColumnInst_1_n3 ;
    wire MixColumnsIns_MixOneColumnInst_1_n2 ;
    wire MixColumnsIns_MixOneColumnInst_1_n1 ;
    wire MixColumnsIns_MixOneColumnInst_2_n64 ;
    wire MixColumnsIns_MixOneColumnInst_2_n63 ;
    wire MixColumnsIns_MixOneColumnInst_2_n62 ;
    wire MixColumnsIns_MixOneColumnInst_2_n61 ;
    wire MixColumnsIns_MixOneColumnInst_2_n60 ;
    wire MixColumnsIns_MixOneColumnInst_2_n59 ;
    wire MixColumnsIns_MixOneColumnInst_2_n58 ;
    wire MixColumnsIns_MixOneColumnInst_2_n57 ;
    wire MixColumnsIns_MixOneColumnInst_2_n56 ;
    wire MixColumnsIns_MixOneColumnInst_2_n55 ;
    wire MixColumnsIns_MixOneColumnInst_2_n54 ;
    wire MixColumnsIns_MixOneColumnInst_2_n53 ;
    wire MixColumnsIns_MixOneColumnInst_2_n52 ;
    wire MixColumnsIns_MixOneColumnInst_2_n51 ;
    wire MixColumnsIns_MixOneColumnInst_2_n50 ;
    wire MixColumnsIns_MixOneColumnInst_2_n49 ;
    wire MixColumnsIns_MixOneColumnInst_2_n48 ;
    wire MixColumnsIns_MixOneColumnInst_2_n47 ;
    wire MixColumnsIns_MixOneColumnInst_2_n46 ;
    wire MixColumnsIns_MixOneColumnInst_2_n45 ;
    wire MixColumnsIns_MixOneColumnInst_2_n44 ;
    wire MixColumnsIns_MixOneColumnInst_2_n43 ;
    wire MixColumnsIns_MixOneColumnInst_2_n42 ;
    wire MixColumnsIns_MixOneColumnInst_2_n41 ;
    wire MixColumnsIns_MixOneColumnInst_2_n40 ;
    wire MixColumnsIns_MixOneColumnInst_2_n39 ;
    wire MixColumnsIns_MixOneColumnInst_2_n38 ;
    wire MixColumnsIns_MixOneColumnInst_2_n37 ;
    wire MixColumnsIns_MixOneColumnInst_2_n36 ;
    wire MixColumnsIns_MixOneColumnInst_2_n35 ;
    wire MixColumnsIns_MixOneColumnInst_2_n34 ;
    wire MixColumnsIns_MixOneColumnInst_2_n33 ;
    wire MixColumnsIns_MixOneColumnInst_2_n32 ;
    wire MixColumnsIns_MixOneColumnInst_2_n31 ;
    wire MixColumnsIns_MixOneColumnInst_2_n30 ;
    wire MixColumnsIns_MixOneColumnInst_2_n29 ;
    wire MixColumnsIns_MixOneColumnInst_2_n28 ;
    wire MixColumnsIns_MixOneColumnInst_2_n27 ;
    wire MixColumnsIns_MixOneColumnInst_2_n26 ;
    wire MixColumnsIns_MixOneColumnInst_2_n25 ;
    wire MixColumnsIns_MixOneColumnInst_2_n24 ;
    wire MixColumnsIns_MixOneColumnInst_2_n23 ;
    wire MixColumnsIns_MixOneColumnInst_2_n22 ;
    wire MixColumnsIns_MixOneColumnInst_2_n21 ;
    wire MixColumnsIns_MixOneColumnInst_2_n20 ;
    wire MixColumnsIns_MixOneColumnInst_2_n19 ;
    wire MixColumnsIns_MixOneColumnInst_2_n18 ;
    wire MixColumnsIns_MixOneColumnInst_2_n17 ;
    wire MixColumnsIns_MixOneColumnInst_2_n16 ;
    wire MixColumnsIns_MixOneColumnInst_2_n15 ;
    wire MixColumnsIns_MixOneColumnInst_2_n14 ;
    wire MixColumnsIns_MixOneColumnInst_2_n13 ;
    wire MixColumnsIns_MixOneColumnInst_2_n12 ;
    wire MixColumnsIns_MixOneColumnInst_2_n11 ;
    wire MixColumnsIns_MixOneColumnInst_2_n10 ;
    wire MixColumnsIns_MixOneColumnInst_2_n9 ;
    wire MixColumnsIns_MixOneColumnInst_2_n8 ;
    wire MixColumnsIns_MixOneColumnInst_2_n7 ;
    wire MixColumnsIns_MixOneColumnInst_2_n6 ;
    wire MixColumnsIns_MixOneColumnInst_2_n5 ;
    wire MixColumnsIns_MixOneColumnInst_2_n4 ;
    wire MixColumnsIns_MixOneColumnInst_2_n3 ;
    wire MixColumnsIns_MixOneColumnInst_2_n2 ;
    wire MixColumnsIns_MixOneColumnInst_2_n1 ;
    wire MixColumnsIns_MixOneColumnInst_3_n64 ;
    wire MixColumnsIns_MixOneColumnInst_3_n63 ;
    wire MixColumnsIns_MixOneColumnInst_3_n62 ;
    wire MixColumnsIns_MixOneColumnInst_3_n61 ;
    wire MixColumnsIns_MixOneColumnInst_3_n60 ;
    wire MixColumnsIns_MixOneColumnInst_3_n59 ;
    wire MixColumnsIns_MixOneColumnInst_3_n58 ;
    wire MixColumnsIns_MixOneColumnInst_3_n57 ;
    wire MixColumnsIns_MixOneColumnInst_3_n56 ;
    wire MixColumnsIns_MixOneColumnInst_3_n55 ;
    wire MixColumnsIns_MixOneColumnInst_3_n54 ;
    wire MixColumnsIns_MixOneColumnInst_3_n53 ;
    wire MixColumnsIns_MixOneColumnInst_3_n52 ;
    wire MixColumnsIns_MixOneColumnInst_3_n51 ;
    wire MixColumnsIns_MixOneColumnInst_3_n50 ;
    wire MixColumnsIns_MixOneColumnInst_3_n49 ;
    wire MixColumnsIns_MixOneColumnInst_3_n48 ;
    wire MixColumnsIns_MixOneColumnInst_3_n47 ;
    wire MixColumnsIns_MixOneColumnInst_3_n46 ;
    wire MixColumnsIns_MixOneColumnInst_3_n45 ;
    wire MixColumnsIns_MixOneColumnInst_3_n44 ;
    wire MixColumnsIns_MixOneColumnInst_3_n43 ;
    wire MixColumnsIns_MixOneColumnInst_3_n42 ;
    wire MixColumnsIns_MixOneColumnInst_3_n41 ;
    wire MixColumnsIns_MixOneColumnInst_3_n40 ;
    wire MixColumnsIns_MixOneColumnInst_3_n39 ;
    wire MixColumnsIns_MixOneColumnInst_3_n38 ;
    wire MixColumnsIns_MixOneColumnInst_3_n37 ;
    wire MixColumnsIns_MixOneColumnInst_3_n36 ;
    wire MixColumnsIns_MixOneColumnInst_3_n35 ;
    wire MixColumnsIns_MixOneColumnInst_3_n34 ;
    wire MixColumnsIns_MixOneColumnInst_3_n33 ;
    wire MixColumnsIns_MixOneColumnInst_3_n32 ;
    wire MixColumnsIns_MixOneColumnInst_3_n31 ;
    wire MixColumnsIns_MixOneColumnInst_3_n30 ;
    wire MixColumnsIns_MixOneColumnInst_3_n29 ;
    wire MixColumnsIns_MixOneColumnInst_3_n28 ;
    wire MixColumnsIns_MixOneColumnInst_3_n27 ;
    wire MixColumnsIns_MixOneColumnInst_3_n26 ;
    wire MixColumnsIns_MixOneColumnInst_3_n25 ;
    wire MixColumnsIns_MixOneColumnInst_3_n24 ;
    wire MixColumnsIns_MixOneColumnInst_3_n23 ;
    wire MixColumnsIns_MixOneColumnInst_3_n22 ;
    wire MixColumnsIns_MixOneColumnInst_3_n21 ;
    wire MixColumnsIns_MixOneColumnInst_3_n20 ;
    wire MixColumnsIns_MixOneColumnInst_3_n19 ;
    wire MixColumnsIns_MixOneColumnInst_3_n18 ;
    wire MixColumnsIns_MixOneColumnInst_3_n17 ;
    wire MixColumnsIns_MixOneColumnInst_3_n16 ;
    wire MixColumnsIns_MixOneColumnInst_3_n15 ;
    wire MixColumnsIns_MixOneColumnInst_3_n14 ;
    wire MixColumnsIns_MixOneColumnInst_3_n13 ;
    wire MixColumnsIns_MixOneColumnInst_3_n12 ;
    wire MixColumnsIns_MixOneColumnInst_3_n11 ;
    wire MixColumnsIns_MixOneColumnInst_3_n10 ;
    wire MixColumnsIns_MixOneColumnInst_3_n9 ;
    wire MixColumnsIns_MixOneColumnInst_3_n8 ;
    wire MixColumnsIns_MixOneColumnInst_3_n7 ;
    wire MixColumnsIns_MixOneColumnInst_3_n6 ;
    wire MixColumnsIns_MixOneColumnInst_3_n5 ;
    wire MixColumnsIns_MixOneColumnInst_3_n4 ;
    wire MixColumnsIns_MixOneColumnInst_3_n3 ;
    wire MixColumnsIns_MixOneColumnInst_3_n2 ;
    wire MixColumnsIns_MixOneColumnInst_3_n1 ;
    wire KeyReg_Inst_ff_SDE_0_next_state ;
    wire KeyReg_Inst_ff_SDE_1_next_state ;
    wire KeyReg_Inst_ff_SDE_2_next_state ;
    wire KeyReg_Inst_ff_SDE_3_next_state ;
    wire KeyReg_Inst_ff_SDE_4_next_state ;
    wire KeyReg_Inst_ff_SDE_5_next_state ;
    wire KeyReg_Inst_ff_SDE_6_next_state ;
    wire KeyReg_Inst_ff_SDE_7_next_state ;
    wire KeyReg_Inst_ff_SDE_8_next_state ;
    wire KeyReg_Inst_ff_SDE_9_next_state ;
    wire KeyReg_Inst_ff_SDE_10_next_state ;
    wire KeyReg_Inst_ff_SDE_11_next_state ;
    wire KeyReg_Inst_ff_SDE_12_next_state ;
    wire KeyReg_Inst_ff_SDE_13_next_state ;
    wire KeyReg_Inst_ff_SDE_14_next_state ;
    wire KeyReg_Inst_ff_SDE_15_next_state ;
    wire KeyReg_Inst_ff_SDE_16_next_state ;
    wire KeyReg_Inst_ff_SDE_17_next_state ;
    wire KeyReg_Inst_ff_SDE_18_next_state ;
    wire KeyReg_Inst_ff_SDE_19_next_state ;
    wire KeyReg_Inst_ff_SDE_20_next_state ;
    wire KeyReg_Inst_ff_SDE_21_next_state ;
    wire KeyReg_Inst_ff_SDE_22_next_state ;
    wire KeyReg_Inst_ff_SDE_23_next_state ;
    wire KeyReg_Inst_ff_SDE_24_next_state ;
    wire KeyReg_Inst_ff_SDE_25_next_state ;
    wire KeyReg_Inst_ff_SDE_26_next_state ;
    wire KeyReg_Inst_ff_SDE_27_next_state ;
    wire KeyReg_Inst_ff_SDE_28_next_state ;
    wire KeyReg_Inst_ff_SDE_29_next_state ;
    wire KeyReg_Inst_ff_SDE_30_next_state ;
    wire KeyReg_Inst_ff_SDE_31_next_state ;
    wire KeyReg_Inst_ff_SDE_32_next_state ;
    wire KeyReg_Inst_ff_SDE_33_next_state ;
    wire KeyReg_Inst_ff_SDE_34_next_state ;
    wire KeyReg_Inst_ff_SDE_35_next_state ;
    wire KeyReg_Inst_ff_SDE_36_next_state ;
    wire KeyReg_Inst_ff_SDE_37_next_state ;
    wire KeyReg_Inst_ff_SDE_38_next_state ;
    wire KeyReg_Inst_ff_SDE_39_next_state ;
    wire KeyReg_Inst_ff_SDE_40_next_state ;
    wire KeyReg_Inst_ff_SDE_41_next_state ;
    wire KeyReg_Inst_ff_SDE_42_next_state ;
    wire KeyReg_Inst_ff_SDE_43_next_state ;
    wire KeyReg_Inst_ff_SDE_44_next_state ;
    wire KeyReg_Inst_ff_SDE_45_next_state ;
    wire KeyReg_Inst_ff_SDE_46_next_state ;
    wire KeyReg_Inst_ff_SDE_47_next_state ;
    wire KeyReg_Inst_ff_SDE_48_next_state ;
    wire KeyReg_Inst_ff_SDE_49_next_state ;
    wire KeyReg_Inst_ff_SDE_50_next_state ;
    wire KeyReg_Inst_ff_SDE_51_next_state ;
    wire KeyReg_Inst_ff_SDE_52_next_state ;
    wire KeyReg_Inst_ff_SDE_53_next_state ;
    wire KeyReg_Inst_ff_SDE_54_next_state ;
    wire KeyReg_Inst_ff_SDE_55_next_state ;
    wire KeyReg_Inst_ff_SDE_56_next_state ;
    wire KeyReg_Inst_ff_SDE_57_next_state ;
    wire KeyReg_Inst_ff_SDE_58_next_state ;
    wire KeyReg_Inst_ff_SDE_59_next_state ;
    wire KeyReg_Inst_ff_SDE_60_next_state ;
    wire KeyReg_Inst_ff_SDE_61_next_state ;
    wire KeyReg_Inst_ff_SDE_62_next_state ;
    wire KeyReg_Inst_ff_SDE_63_next_state ;
    wire KeyReg_Inst_ff_SDE_64_next_state ;
    wire KeyReg_Inst_ff_SDE_65_next_state ;
    wire KeyReg_Inst_ff_SDE_66_next_state ;
    wire KeyReg_Inst_ff_SDE_67_next_state ;
    wire KeyReg_Inst_ff_SDE_68_next_state ;
    wire KeyReg_Inst_ff_SDE_69_next_state ;
    wire KeyReg_Inst_ff_SDE_70_next_state ;
    wire KeyReg_Inst_ff_SDE_71_next_state ;
    wire KeyReg_Inst_ff_SDE_72_next_state ;
    wire KeyReg_Inst_ff_SDE_73_next_state ;
    wire KeyReg_Inst_ff_SDE_74_next_state ;
    wire KeyReg_Inst_ff_SDE_75_next_state ;
    wire KeyReg_Inst_ff_SDE_76_next_state ;
    wire KeyReg_Inst_ff_SDE_77_next_state ;
    wire KeyReg_Inst_ff_SDE_78_next_state ;
    wire KeyReg_Inst_ff_SDE_79_next_state ;
    wire KeyReg_Inst_ff_SDE_80_next_state ;
    wire KeyReg_Inst_ff_SDE_81_next_state ;
    wire KeyReg_Inst_ff_SDE_82_next_state ;
    wire KeyReg_Inst_ff_SDE_83_next_state ;
    wire KeyReg_Inst_ff_SDE_84_next_state ;
    wire KeyReg_Inst_ff_SDE_85_next_state ;
    wire KeyReg_Inst_ff_SDE_86_next_state ;
    wire KeyReg_Inst_ff_SDE_87_next_state ;
    wire KeyReg_Inst_ff_SDE_88_next_state ;
    wire KeyReg_Inst_ff_SDE_89_next_state ;
    wire KeyReg_Inst_ff_SDE_90_next_state ;
    wire KeyReg_Inst_ff_SDE_91_next_state ;
    wire KeyReg_Inst_ff_SDE_92_next_state ;
    wire KeyReg_Inst_ff_SDE_93_next_state ;
    wire KeyReg_Inst_ff_SDE_94_next_state ;
    wire KeyReg_Inst_ff_SDE_95_next_state ;
    wire KeyReg_Inst_ff_SDE_96_next_state ;
    wire KeyReg_Inst_ff_SDE_97_next_state ;
    wire KeyReg_Inst_ff_SDE_98_next_state ;
    wire KeyReg_Inst_ff_SDE_99_next_state ;
    wire KeyReg_Inst_ff_SDE_100_next_state ;
    wire KeyReg_Inst_ff_SDE_101_next_state ;
    wire KeyReg_Inst_ff_SDE_102_next_state ;
    wire KeyReg_Inst_ff_SDE_103_next_state ;
    wire KeyReg_Inst_ff_SDE_104_next_state ;
    wire KeyReg_Inst_ff_SDE_105_next_state ;
    wire KeyReg_Inst_ff_SDE_106_next_state ;
    wire KeyReg_Inst_ff_SDE_107_next_state ;
    wire KeyReg_Inst_ff_SDE_108_next_state ;
    wire KeyReg_Inst_ff_SDE_109_next_state ;
    wire KeyReg_Inst_ff_SDE_110_next_state ;
    wire KeyReg_Inst_ff_SDE_111_next_state ;
    wire KeyReg_Inst_ff_SDE_112_next_state ;
    wire KeyReg_Inst_ff_SDE_113_next_state ;
    wire KeyReg_Inst_ff_SDE_114_next_state ;
    wire KeyReg_Inst_ff_SDE_115_next_state ;
    wire KeyReg_Inst_ff_SDE_116_next_state ;
    wire KeyReg_Inst_ff_SDE_117_next_state ;
    wire KeyReg_Inst_ff_SDE_118_next_state ;
    wire KeyReg_Inst_ff_SDE_119_next_state ;
    wire KeyReg_Inst_ff_SDE_120_next_state ;
    wire KeyReg_Inst_ff_SDE_121_next_state ;
    wire KeyReg_Inst_ff_SDE_122_next_state ;
    wire KeyReg_Inst_ff_SDE_123_next_state ;
    wire KeyReg_Inst_ff_SDE_124_next_state ;
    wire KeyReg_Inst_ff_SDE_125_next_state ;
    wire KeyReg_Inst_ff_SDE_126_next_state ;
    wire KeyReg_Inst_ff_SDE_127_next_state ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__0_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__1_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__2_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__3_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__4_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__5_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__6_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__7_ ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M63 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M60 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M59 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M57 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M54 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M49 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M47 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M36 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M35 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M34 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M33 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M32 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M31 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M30 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M63 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M60 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M59 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M57 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M54 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M49 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M47 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M36 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M35 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M34 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M33 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M32 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M31 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M30 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M63 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M60 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M59 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M57 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M54 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M49 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M47 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M36 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M35 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M34 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M33 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M32 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M31 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M30 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M63 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M60 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M59 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M57 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M54 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M49 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M47 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M36 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M35 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M34 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M33 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M32 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M31 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M30 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1 ;
    wire RoundCounterIns_n13 ;
    wire RoundCounterIns_n12 ;
    wire RoundCounterIns_n11 ;
    wire RoundCounterIns_n10 ;
    wire RoundCounterIns_n9 ;
    wire RoundCounterIns_n8 ;
    wire RoundCounterIns_n7 ;
    wire RoundCounterIns_n4 ;
    wire RoundCounterIns_n3 ;
    wire RoundCounterIns_n2 ;
    wire RoundCounterIns_n1 ;
    wire RoundCounterIns_N10 ;
    wire RoundCounterIns_n5 ;
    wire RoundCounterIns_N8 ;
    wire RoundCounterIns_n6 ;
    wire RoundCounterIns_N7 ;
    wire [127:0] RoundOutput ;
    wire [127:0] RoundInput ;
    wire [123:0] MixColumnsInput ;
    wire [127:0] MixColumnsOutput ;
    wire [127:0] KeyExpansionOutput ;
    wire [127:0] RoundKey ;
    wire [5:0] Rcon ;
    wire [3:0] RoundCounter ;
    wire [31:0] MixColumnsIns_MixOneColumnInst_0_DoubleBytes ;
    wire [31:0] MixColumnsIns_MixOneColumnInst_1_DoubleBytes ;
    wire [31:0] MixColumnsIns_MixOneColumnInst_2_DoubleBytes ;
    wire [31:0] MixColumnsIns_MixOneColumnInst_3_DoubleBytes ;
    wire [31:0] KeyExpansionIns_tmp ;
    wire new_AGEMA_signal_4549 ;
    wire new_AGEMA_signal_4550 ;
    wire new_AGEMA_signal_4552 ;
    wire new_AGEMA_signal_4553 ;
    wire new_AGEMA_signal_4555 ;
    wire new_AGEMA_signal_4556 ;
    wire new_AGEMA_signal_4558 ;
    wire new_AGEMA_signal_4559 ;
    wire new_AGEMA_signal_4561 ;
    wire new_AGEMA_signal_4562 ;
    wire new_AGEMA_signal_4564 ;
    wire new_AGEMA_signal_4565 ;
    wire new_AGEMA_signal_4567 ;
    wire new_AGEMA_signal_4568 ;
    wire new_AGEMA_signal_4570 ;
    wire new_AGEMA_signal_4571 ;
    wire new_AGEMA_signal_4573 ;
    wire new_AGEMA_signal_4574 ;
    wire new_AGEMA_signal_4576 ;
    wire new_AGEMA_signal_4577 ;
    wire new_AGEMA_signal_4579 ;
    wire new_AGEMA_signal_4580 ;
    wire new_AGEMA_signal_4582 ;
    wire new_AGEMA_signal_4583 ;
    wire new_AGEMA_signal_4585 ;
    wire new_AGEMA_signal_4586 ;
    wire new_AGEMA_signal_4588 ;
    wire new_AGEMA_signal_4589 ;
    wire new_AGEMA_signal_4591 ;
    wire new_AGEMA_signal_4592 ;
    wire new_AGEMA_signal_4594 ;
    wire new_AGEMA_signal_4595 ;
    wire new_AGEMA_signal_4597 ;
    wire new_AGEMA_signal_4598 ;
    wire new_AGEMA_signal_4600 ;
    wire new_AGEMA_signal_4601 ;
    wire new_AGEMA_signal_4603 ;
    wire new_AGEMA_signal_4604 ;
    wire new_AGEMA_signal_4606 ;
    wire new_AGEMA_signal_4607 ;
    wire new_AGEMA_signal_4609 ;
    wire new_AGEMA_signal_4610 ;
    wire new_AGEMA_signal_4612 ;
    wire new_AGEMA_signal_4613 ;
    wire new_AGEMA_signal_4615 ;
    wire new_AGEMA_signal_4616 ;
    wire new_AGEMA_signal_4618 ;
    wire new_AGEMA_signal_4619 ;
    wire new_AGEMA_signal_4621 ;
    wire new_AGEMA_signal_4622 ;
    wire new_AGEMA_signal_4624 ;
    wire new_AGEMA_signal_4625 ;
    wire new_AGEMA_signal_4627 ;
    wire new_AGEMA_signal_4628 ;
    wire new_AGEMA_signal_4630 ;
    wire new_AGEMA_signal_4631 ;
    wire new_AGEMA_signal_4633 ;
    wire new_AGEMA_signal_4634 ;
    wire new_AGEMA_signal_4636 ;
    wire new_AGEMA_signal_4637 ;
    wire new_AGEMA_signal_4639 ;
    wire new_AGEMA_signal_4640 ;
    wire new_AGEMA_signal_4642 ;
    wire new_AGEMA_signal_4643 ;
    wire new_AGEMA_signal_4645 ;
    wire new_AGEMA_signal_4646 ;
    wire new_AGEMA_signal_4648 ;
    wire new_AGEMA_signal_4649 ;
    wire new_AGEMA_signal_4651 ;
    wire new_AGEMA_signal_4652 ;
    wire new_AGEMA_signal_4654 ;
    wire new_AGEMA_signal_4655 ;
    wire new_AGEMA_signal_4657 ;
    wire new_AGEMA_signal_4658 ;
    wire new_AGEMA_signal_4660 ;
    wire new_AGEMA_signal_4661 ;
    wire new_AGEMA_signal_4663 ;
    wire new_AGEMA_signal_4664 ;
    wire new_AGEMA_signal_4666 ;
    wire new_AGEMA_signal_4667 ;
    wire new_AGEMA_signal_4669 ;
    wire new_AGEMA_signal_4670 ;
    wire new_AGEMA_signal_4672 ;
    wire new_AGEMA_signal_4673 ;
    wire new_AGEMA_signal_4675 ;
    wire new_AGEMA_signal_4676 ;
    wire new_AGEMA_signal_4678 ;
    wire new_AGEMA_signal_4679 ;
    wire new_AGEMA_signal_4681 ;
    wire new_AGEMA_signal_4682 ;
    wire new_AGEMA_signal_4684 ;
    wire new_AGEMA_signal_4685 ;
    wire new_AGEMA_signal_4687 ;
    wire new_AGEMA_signal_4688 ;
    wire new_AGEMA_signal_4690 ;
    wire new_AGEMA_signal_4691 ;
    wire new_AGEMA_signal_4693 ;
    wire new_AGEMA_signal_4694 ;
    wire new_AGEMA_signal_4696 ;
    wire new_AGEMA_signal_4697 ;
    wire new_AGEMA_signal_4699 ;
    wire new_AGEMA_signal_4700 ;
    wire new_AGEMA_signal_4702 ;
    wire new_AGEMA_signal_4703 ;
    wire new_AGEMA_signal_4705 ;
    wire new_AGEMA_signal_4706 ;
    wire new_AGEMA_signal_4708 ;
    wire new_AGEMA_signal_4709 ;
    wire new_AGEMA_signal_4711 ;
    wire new_AGEMA_signal_4712 ;
    wire new_AGEMA_signal_4714 ;
    wire new_AGEMA_signal_4715 ;
    wire new_AGEMA_signal_4717 ;
    wire new_AGEMA_signal_4718 ;
    wire new_AGEMA_signal_4720 ;
    wire new_AGEMA_signal_4721 ;
    wire new_AGEMA_signal_4723 ;
    wire new_AGEMA_signal_4724 ;
    wire new_AGEMA_signal_4726 ;
    wire new_AGEMA_signal_4727 ;
    wire new_AGEMA_signal_4729 ;
    wire new_AGEMA_signal_4730 ;
    wire new_AGEMA_signal_4732 ;
    wire new_AGEMA_signal_4733 ;
    wire new_AGEMA_signal_4735 ;
    wire new_AGEMA_signal_4736 ;
    wire new_AGEMA_signal_4738 ;
    wire new_AGEMA_signal_4739 ;
    wire new_AGEMA_signal_4741 ;
    wire new_AGEMA_signal_4742 ;
    wire new_AGEMA_signal_4744 ;
    wire new_AGEMA_signal_4745 ;
    wire new_AGEMA_signal_4747 ;
    wire new_AGEMA_signal_4748 ;
    wire new_AGEMA_signal_4750 ;
    wire new_AGEMA_signal_4751 ;
    wire new_AGEMA_signal_4753 ;
    wire new_AGEMA_signal_4754 ;
    wire new_AGEMA_signal_4756 ;
    wire new_AGEMA_signal_4757 ;
    wire new_AGEMA_signal_4759 ;
    wire new_AGEMA_signal_4760 ;
    wire new_AGEMA_signal_4762 ;
    wire new_AGEMA_signal_4763 ;
    wire new_AGEMA_signal_4765 ;
    wire new_AGEMA_signal_4766 ;
    wire new_AGEMA_signal_4768 ;
    wire new_AGEMA_signal_4769 ;
    wire new_AGEMA_signal_4771 ;
    wire new_AGEMA_signal_4772 ;
    wire new_AGEMA_signal_4774 ;
    wire new_AGEMA_signal_4775 ;
    wire new_AGEMA_signal_4777 ;
    wire new_AGEMA_signal_4778 ;
    wire new_AGEMA_signal_4780 ;
    wire new_AGEMA_signal_4781 ;
    wire new_AGEMA_signal_4783 ;
    wire new_AGEMA_signal_4784 ;
    wire new_AGEMA_signal_4786 ;
    wire new_AGEMA_signal_4787 ;
    wire new_AGEMA_signal_4789 ;
    wire new_AGEMA_signal_4790 ;
    wire new_AGEMA_signal_4792 ;
    wire new_AGEMA_signal_4793 ;
    wire new_AGEMA_signal_4795 ;
    wire new_AGEMA_signal_4796 ;
    wire new_AGEMA_signal_4798 ;
    wire new_AGEMA_signal_4799 ;
    wire new_AGEMA_signal_4801 ;
    wire new_AGEMA_signal_4802 ;
    wire new_AGEMA_signal_4804 ;
    wire new_AGEMA_signal_4805 ;
    wire new_AGEMA_signal_4807 ;
    wire new_AGEMA_signal_4808 ;
    wire new_AGEMA_signal_4810 ;
    wire new_AGEMA_signal_4811 ;
    wire new_AGEMA_signal_4813 ;
    wire new_AGEMA_signal_4814 ;
    wire new_AGEMA_signal_4816 ;
    wire new_AGEMA_signal_4817 ;
    wire new_AGEMA_signal_4819 ;
    wire new_AGEMA_signal_4820 ;
    wire new_AGEMA_signal_4822 ;
    wire new_AGEMA_signal_4823 ;
    wire new_AGEMA_signal_4825 ;
    wire new_AGEMA_signal_4826 ;
    wire new_AGEMA_signal_4828 ;
    wire new_AGEMA_signal_4829 ;
    wire new_AGEMA_signal_4831 ;
    wire new_AGEMA_signal_4832 ;
    wire new_AGEMA_signal_4834 ;
    wire new_AGEMA_signal_4835 ;
    wire new_AGEMA_signal_4837 ;
    wire new_AGEMA_signal_4838 ;
    wire new_AGEMA_signal_4840 ;
    wire new_AGEMA_signal_4841 ;
    wire new_AGEMA_signal_4843 ;
    wire new_AGEMA_signal_4844 ;
    wire new_AGEMA_signal_4846 ;
    wire new_AGEMA_signal_4847 ;
    wire new_AGEMA_signal_4849 ;
    wire new_AGEMA_signal_4850 ;
    wire new_AGEMA_signal_4852 ;
    wire new_AGEMA_signal_4853 ;
    wire new_AGEMA_signal_4855 ;
    wire new_AGEMA_signal_4856 ;
    wire new_AGEMA_signal_4858 ;
    wire new_AGEMA_signal_4859 ;
    wire new_AGEMA_signal_4861 ;
    wire new_AGEMA_signal_4862 ;
    wire new_AGEMA_signal_4864 ;
    wire new_AGEMA_signal_4865 ;
    wire new_AGEMA_signal_4867 ;
    wire new_AGEMA_signal_4868 ;
    wire new_AGEMA_signal_4870 ;
    wire new_AGEMA_signal_4871 ;
    wire new_AGEMA_signal_4873 ;
    wire new_AGEMA_signal_4874 ;
    wire new_AGEMA_signal_4876 ;
    wire new_AGEMA_signal_4877 ;
    wire new_AGEMA_signal_4879 ;
    wire new_AGEMA_signal_4880 ;
    wire new_AGEMA_signal_4882 ;
    wire new_AGEMA_signal_4883 ;
    wire new_AGEMA_signal_4885 ;
    wire new_AGEMA_signal_4886 ;
    wire new_AGEMA_signal_4888 ;
    wire new_AGEMA_signal_4889 ;
    wire new_AGEMA_signal_4891 ;
    wire new_AGEMA_signal_4892 ;
    wire new_AGEMA_signal_4894 ;
    wire new_AGEMA_signal_4895 ;
    wire new_AGEMA_signal_4897 ;
    wire new_AGEMA_signal_4898 ;
    wire new_AGEMA_signal_4900 ;
    wire new_AGEMA_signal_4901 ;
    wire new_AGEMA_signal_4903 ;
    wire new_AGEMA_signal_4904 ;
    wire new_AGEMA_signal_4906 ;
    wire new_AGEMA_signal_4907 ;
    wire new_AGEMA_signal_4909 ;
    wire new_AGEMA_signal_4910 ;
    wire new_AGEMA_signal_4912 ;
    wire new_AGEMA_signal_4913 ;
    wire new_AGEMA_signal_4915 ;
    wire new_AGEMA_signal_4916 ;
    wire new_AGEMA_signal_4918 ;
    wire new_AGEMA_signal_4919 ;
    wire new_AGEMA_signal_4921 ;
    wire new_AGEMA_signal_4922 ;
    wire new_AGEMA_signal_4924 ;
    wire new_AGEMA_signal_4925 ;
    wire new_AGEMA_signal_4927 ;
    wire new_AGEMA_signal_4928 ;
    wire new_AGEMA_signal_4930 ;
    wire new_AGEMA_signal_4931 ;
    wire new_AGEMA_signal_4933 ;
    wire new_AGEMA_signal_4934 ;
    wire new_AGEMA_signal_4935 ;
    wire new_AGEMA_signal_4936 ;
    wire new_AGEMA_signal_4937 ;
    wire new_AGEMA_signal_4938 ;
    wire new_AGEMA_signal_4939 ;
    wire new_AGEMA_signal_4940 ;
    wire new_AGEMA_signal_4941 ;
    wire new_AGEMA_signal_4942 ;
    wire new_AGEMA_signal_4943 ;
    wire new_AGEMA_signal_4944 ;
    wire new_AGEMA_signal_4945 ;
    wire new_AGEMA_signal_4946 ;
    wire new_AGEMA_signal_4947 ;
    wire new_AGEMA_signal_4948 ;
    wire new_AGEMA_signal_4949 ;
    wire new_AGEMA_signal_4950 ;
    wire new_AGEMA_signal_4951 ;
    wire new_AGEMA_signal_4952 ;
    wire new_AGEMA_signal_4953 ;
    wire new_AGEMA_signal_4954 ;
    wire new_AGEMA_signal_4955 ;
    wire new_AGEMA_signal_4956 ;
    wire new_AGEMA_signal_4957 ;
    wire new_AGEMA_signal_4958 ;
    wire new_AGEMA_signal_4959 ;
    wire new_AGEMA_signal_4960 ;
    wire new_AGEMA_signal_4961 ;
    wire new_AGEMA_signal_4962 ;
    wire new_AGEMA_signal_4963 ;
    wire new_AGEMA_signal_4964 ;
    wire new_AGEMA_signal_4965 ;
    wire new_AGEMA_signal_4966 ;
    wire new_AGEMA_signal_4967 ;
    wire new_AGEMA_signal_4968 ;
    wire new_AGEMA_signal_4969 ;
    wire new_AGEMA_signal_4970 ;
    wire new_AGEMA_signal_4971 ;
    wire new_AGEMA_signal_4972 ;
    wire new_AGEMA_signal_4973 ;
    wire new_AGEMA_signal_4974 ;
    wire new_AGEMA_signal_4975 ;
    wire new_AGEMA_signal_4976 ;
    wire new_AGEMA_signal_4977 ;
    wire new_AGEMA_signal_4978 ;
    wire new_AGEMA_signal_4979 ;
    wire new_AGEMA_signal_4980 ;
    wire new_AGEMA_signal_4981 ;
    wire new_AGEMA_signal_4982 ;
    wire new_AGEMA_signal_4983 ;
    wire new_AGEMA_signal_4984 ;
    wire new_AGEMA_signal_4985 ;
    wire new_AGEMA_signal_4986 ;
    wire new_AGEMA_signal_4987 ;
    wire new_AGEMA_signal_4988 ;
    wire new_AGEMA_signal_4989 ;
    wire new_AGEMA_signal_4990 ;
    wire new_AGEMA_signal_4991 ;
    wire new_AGEMA_signal_4992 ;
    wire new_AGEMA_signal_4993 ;
    wire new_AGEMA_signal_4994 ;
    wire new_AGEMA_signal_4995 ;
    wire new_AGEMA_signal_4996 ;
    wire new_AGEMA_signal_4997 ;
    wire new_AGEMA_signal_4998 ;
    wire new_AGEMA_signal_4999 ;
    wire new_AGEMA_signal_5000 ;
    wire new_AGEMA_signal_5001 ;
    wire new_AGEMA_signal_5002 ;
    wire new_AGEMA_signal_5003 ;
    wire new_AGEMA_signal_5004 ;
    wire new_AGEMA_signal_5005 ;
    wire new_AGEMA_signal_5006 ;
    wire new_AGEMA_signal_5007 ;
    wire new_AGEMA_signal_5008 ;
    wire new_AGEMA_signal_5009 ;
    wire new_AGEMA_signal_5010 ;
    wire new_AGEMA_signal_5011 ;
    wire new_AGEMA_signal_5012 ;
    wire new_AGEMA_signal_5013 ;
    wire new_AGEMA_signal_5014 ;
    wire new_AGEMA_signal_5015 ;
    wire new_AGEMA_signal_5016 ;
    wire new_AGEMA_signal_5017 ;
    wire new_AGEMA_signal_5018 ;
    wire new_AGEMA_signal_5019 ;
    wire new_AGEMA_signal_5020 ;
    wire new_AGEMA_signal_5021 ;
    wire new_AGEMA_signal_5022 ;
    wire new_AGEMA_signal_5023 ;
    wire new_AGEMA_signal_5024 ;
    wire new_AGEMA_signal_5025 ;
    wire new_AGEMA_signal_5026 ;
    wire new_AGEMA_signal_5027 ;
    wire new_AGEMA_signal_5028 ;
    wire new_AGEMA_signal_5029 ;
    wire new_AGEMA_signal_5030 ;
    wire new_AGEMA_signal_5031 ;
    wire new_AGEMA_signal_5032 ;
    wire new_AGEMA_signal_5033 ;
    wire new_AGEMA_signal_5034 ;
    wire new_AGEMA_signal_5035 ;
    wire new_AGEMA_signal_5036 ;
    wire new_AGEMA_signal_5037 ;
    wire new_AGEMA_signal_5038 ;
    wire new_AGEMA_signal_5039 ;
    wire new_AGEMA_signal_5040 ;
    wire new_AGEMA_signal_5041 ;
    wire new_AGEMA_signal_5042 ;
    wire new_AGEMA_signal_5043 ;
    wire new_AGEMA_signal_5044 ;
    wire new_AGEMA_signal_5045 ;
    wire new_AGEMA_signal_5046 ;
    wire new_AGEMA_signal_5047 ;
    wire new_AGEMA_signal_5048 ;
    wire new_AGEMA_signal_5049 ;
    wire new_AGEMA_signal_5050 ;
    wire new_AGEMA_signal_5051 ;
    wire new_AGEMA_signal_5052 ;
    wire new_AGEMA_signal_5053 ;
    wire new_AGEMA_signal_5054 ;
    wire new_AGEMA_signal_5055 ;
    wire new_AGEMA_signal_5056 ;
    wire new_AGEMA_signal_5057 ;
    wire new_AGEMA_signal_5058 ;
    wire new_AGEMA_signal_5059 ;
    wire new_AGEMA_signal_5060 ;
    wire new_AGEMA_signal_5061 ;
    wire new_AGEMA_signal_5062 ;
    wire new_AGEMA_signal_5063 ;
    wire new_AGEMA_signal_5064 ;
    wire new_AGEMA_signal_5065 ;
    wire new_AGEMA_signal_5066 ;
    wire new_AGEMA_signal_5067 ;
    wire new_AGEMA_signal_5068 ;
    wire new_AGEMA_signal_5069 ;
    wire new_AGEMA_signal_5070 ;
    wire new_AGEMA_signal_5071 ;
    wire new_AGEMA_signal_5072 ;
    wire new_AGEMA_signal_5073 ;
    wire new_AGEMA_signal_5074 ;
    wire new_AGEMA_signal_5075 ;
    wire new_AGEMA_signal_5076 ;
    wire new_AGEMA_signal_5077 ;
    wire new_AGEMA_signal_5078 ;
    wire new_AGEMA_signal_5079 ;
    wire new_AGEMA_signal_5080 ;
    wire new_AGEMA_signal_5081 ;
    wire new_AGEMA_signal_5082 ;
    wire new_AGEMA_signal_5083 ;
    wire new_AGEMA_signal_5084 ;
    wire new_AGEMA_signal_5085 ;
    wire new_AGEMA_signal_5086 ;
    wire new_AGEMA_signal_5087 ;
    wire new_AGEMA_signal_5088 ;
    wire new_AGEMA_signal_5089 ;
    wire new_AGEMA_signal_5090 ;
    wire new_AGEMA_signal_5091 ;
    wire new_AGEMA_signal_5092 ;
    wire new_AGEMA_signal_5093 ;
    wire new_AGEMA_signal_5094 ;
    wire new_AGEMA_signal_5095 ;
    wire new_AGEMA_signal_5096 ;
    wire new_AGEMA_signal_5097 ;
    wire new_AGEMA_signal_5098 ;
    wire new_AGEMA_signal_5099 ;
    wire new_AGEMA_signal_5100 ;
    wire new_AGEMA_signal_5101 ;
    wire new_AGEMA_signal_5102 ;
    wire new_AGEMA_signal_5103 ;
    wire new_AGEMA_signal_5104 ;
    wire new_AGEMA_signal_5105 ;
    wire new_AGEMA_signal_5106 ;
    wire new_AGEMA_signal_5107 ;
    wire new_AGEMA_signal_5108 ;
    wire new_AGEMA_signal_5109 ;
    wire new_AGEMA_signal_5110 ;
    wire new_AGEMA_signal_5111 ;
    wire new_AGEMA_signal_5112 ;
    wire new_AGEMA_signal_5113 ;
    wire new_AGEMA_signal_5114 ;
    wire new_AGEMA_signal_5115 ;
    wire new_AGEMA_signal_5116 ;
    wire new_AGEMA_signal_5117 ;
    wire new_AGEMA_signal_5118 ;
    wire new_AGEMA_signal_5119 ;
    wire new_AGEMA_signal_5120 ;
    wire new_AGEMA_signal_5121 ;
    wire new_AGEMA_signal_5122 ;
    wire new_AGEMA_signal_5123 ;
    wire new_AGEMA_signal_5124 ;
    wire new_AGEMA_signal_5125 ;
    wire new_AGEMA_signal_5126 ;
    wire new_AGEMA_signal_5127 ;
    wire new_AGEMA_signal_5128 ;
    wire new_AGEMA_signal_5129 ;
    wire new_AGEMA_signal_5130 ;
    wire new_AGEMA_signal_5131 ;
    wire new_AGEMA_signal_5132 ;
    wire new_AGEMA_signal_5133 ;
    wire new_AGEMA_signal_5134 ;
    wire new_AGEMA_signal_5135 ;
    wire new_AGEMA_signal_5136 ;
    wire new_AGEMA_signal_5137 ;
    wire new_AGEMA_signal_5138 ;
    wire new_AGEMA_signal_5139 ;
    wire new_AGEMA_signal_5140 ;
    wire new_AGEMA_signal_5141 ;
    wire new_AGEMA_signal_5142 ;
    wire new_AGEMA_signal_5143 ;
    wire new_AGEMA_signal_5144 ;
    wire new_AGEMA_signal_5145 ;
    wire new_AGEMA_signal_5146 ;
    wire new_AGEMA_signal_5147 ;
    wire new_AGEMA_signal_5148 ;
    wire new_AGEMA_signal_5149 ;
    wire new_AGEMA_signal_5150 ;
    wire new_AGEMA_signal_5151 ;
    wire new_AGEMA_signal_5152 ;
    wire new_AGEMA_signal_5153 ;
    wire new_AGEMA_signal_5154 ;
    wire new_AGEMA_signal_5155 ;
    wire new_AGEMA_signal_5156 ;
    wire new_AGEMA_signal_5157 ;
    wire new_AGEMA_signal_5158 ;
    wire new_AGEMA_signal_5159 ;
    wire new_AGEMA_signal_5160 ;
    wire new_AGEMA_signal_5161 ;
    wire new_AGEMA_signal_5162 ;
    wire new_AGEMA_signal_5163 ;
    wire new_AGEMA_signal_5164 ;
    wire new_AGEMA_signal_5165 ;
    wire new_AGEMA_signal_5166 ;
    wire new_AGEMA_signal_5167 ;
    wire new_AGEMA_signal_5168 ;
    wire new_AGEMA_signal_5169 ;
    wire new_AGEMA_signal_5170 ;
    wire new_AGEMA_signal_5171 ;
    wire new_AGEMA_signal_5172 ;
    wire new_AGEMA_signal_5173 ;
    wire new_AGEMA_signal_5174 ;
    wire new_AGEMA_signal_5175 ;
    wire new_AGEMA_signal_5176 ;
    wire new_AGEMA_signal_5177 ;
    wire new_AGEMA_signal_5178 ;
    wire new_AGEMA_signal_5179 ;
    wire new_AGEMA_signal_5180 ;
    wire new_AGEMA_signal_5181 ;
    wire new_AGEMA_signal_5182 ;
    wire new_AGEMA_signal_5183 ;
    wire new_AGEMA_signal_5184 ;
    wire new_AGEMA_signal_5185 ;
    wire new_AGEMA_signal_5186 ;
    wire new_AGEMA_signal_5187 ;
    wire new_AGEMA_signal_5188 ;
    wire new_AGEMA_signal_5189 ;
    wire new_AGEMA_signal_5190 ;
    wire new_AGEMA_signal_5191 ;
    wire new_AGEMA_signal_5192 ;
    wire new_AGEMA_signal_5193 ;
    wire new_AGEMA_signal_5194 ;
    wire new_AGEMA_signal_5195 ;
    wire new_AGEMA_signal_5196 ;
    wire new_AGEMA_signal_5197 ;
    wire new_AGEMA_signal_5198 ;
    wire new_AGEMA_signal_5199 ;
    wire new_AGEMA_signal_5200 ;
    wire new_AGEMA_signal_5201 ;
    wire new_AGEMA_signal_5202 ;
    wire new_AGEMA_signal_5203 ;
    wire new_AGEMA_signal_5204 ;
    wire new_AGEMA_signal_5205 ;
    wire new_AGEMA_signal_5206 ;
    wire new_AGEMA_signal_5207 ;
    wire new_AGEMA_signal_5208 ;
    wire new_AGEMA_signal_5209 ;
    wire new_AGEMA_signal_5210 ;
    wire new_AGEMA_signal_5211 ;
    wire new_AGEMA_signal_5212 ;
    wire new_AGEMA_signal_5213 ;
    wire new_AGEMA_signal_5214 ;
    wire new_AGEMA_signal_5215 ;
    wire new_AGEMA_signal_5216 ;
    wire new_AGEMA_signal_5217 ;
    wire new_AGEMA_signal_5218 ;
    wire new_AGEMA_signal_5219 ;
    wire new_AGEMA_signal_5220 ;
    wire new_AGEMA_signal_5221 ;
    wire new_AGEMA_signal_5222 ;
    wire new_AGEMA_signal_5223 ;
    wire new_AGEMA_signal_5224 ;
    wire new_AGEMA_signal_5225 ;
    wire new_AGEMA_signal_5226 ;
    wire new_AGEMA_signal_5227 ;
    wire new_AGEMA_signal_5228 ;
    wire new_AGEMA_signal_5229 ;
    wire new_AGEMA_signal_5230 ;
    wire new_AGEMA_signal_5231 ;
    wire new_AGEMA_signal_5232 ;
    wire new_AGEMA_signal_5233 ;
    wire new_AGEMA_signal_5234 ;
    wire new_AGEMA_signal_5235 ;
    wire new_AGEMA_signal_5236 ;
    wire new_AGEMA_signal_5237 ;
    wire new_AGEMA_signal_5238 ;
    wire new_AGEMA_signal_5239 ;
    wire new_AGEMA_signal_5240 ;
    wire new_AGEMA_signal_5241 ;
    wire new_AGEMA_signal_5242 ;
    wire new_AGEMA_signal_5243 ;
    wire new_AGEMA_signal_5244 ;
    wire new_AGEMA_signal_5245 ;
    wire new_AGEMA_signal_5246 ;
    wire new_AGEMA_signal_5247 ;
    wire new_AGEMA_signal_5248 ;
    wire new_AGEMA_signal_5249 ;
    wire new_AGEMA_signal_5250 ;
    wire new_AGEMA_signal_5251 ;
    wire new_AGEMA_signal_5252 ;
    wire new_AGEMA_signal_5253 ;
    wire new_AGEMA_signal_5254 ;
    wire new_AGEMA_signal_5255 ;
    wire new_AGEMA_signal_5256 ;
    wire new_AGEMA_signal_5257 ;
    wire new_AGEMA_signal_5258 ;
    wire new_AGEMA_signal_5259 ;
    wire new_AGEMA_signal_5260 ;
    wire new_AGEMA_signal_5261 ;
    wire new_AGEMA_signal_5262 ;
    wire new_AGEMA_signal_5263 ;
    wire new_AGEMA_signal_5264 ;
    wire new_AGEMA_signal_5265 ;
    wire new_AGEMA_signal_5266 ;
    wire new_AGEMA_signal_5267 ;
    wire new_AGEMA_signal_5268 ;
    wire new_AGEMA_signal_5269 ;
    wire new_AGEMA_signal_5270 ;
    wire new_AGEMA_signal_5271 ;
    wire new_AGEMA_signal_5272 ;
    wire new_AGEMA_signal_5273 ;
    wire new_AGEMA_signal_5274 ;
    wire new_AGEMA_signal_5275 ;
    wire new_AGEMA_signal_5276 ;
    wire new_AGEMA_signal_5277 ;
    wire new_AGEMA_signal_5278 ;
    wire new_AGEMA_signal_5279 ;
    wire new_AGEMA_signal_5280 ;
    wire new_AGEMA_signal_5281 ;
    wire new_AGEMA_signal_5282 ;
    wire new_AGEMA_signal_5283 ;
    wire new_AGEMA_signal_5284 ;
    wire new_AGEMA_signal_5285 ;
    wire new_AGEMA_signal_5286 ;
    wire new_AGEMA_signal_5287 ;
    wire new_AGEMA_signal_5288 ;
    wire new_AGEMA_signal_5289 ;
    wire new_AGEMA_signal_5290 ;
    wire new_AGEMA_signal_5291 ;
    wire new_AGEMA_signal_5292 ;
    wire new_AGEMA_signal_5293 ;
    wire new_AGEMA_signal_5294 ;
    wire new_AGEMA_signal_5295 ;
    wire new_AGEMA_signal_5296 ;
    wire new_AGEMA_signal_5297 ;
    wire new_AGEMA_signal_5298 ;
    wire new_AGEMA_signal_5299 ;
    wire new_AGEMA_signal_5300 ;
    wire new_AGEMA_signal_5301 ;
    wire new_AGEMA_signal_5302 ;
    wire new_AGEMA_signal_5303 ;
    wire new_AGEMA_signal_5304 ;
    wire new_AGEMA_signal_5305 ;
    wire new_AGEMA_signal_5306 ;
    wire new_AGEMA_signal_5307 ;
    wire new_AGEMA_signal_5308 ;
    wire new_AGEMA_signal_5309 ;
    wire new_AGEMA_signal_5310 ;
    wire new_AGEMA_signal_5311 ;
    wire new_AGEMA_signal_5312 ;
    wire new_AGEMA_signal_5313 ;
    wire new_AGEMA_signal_5314 ;
    wire new_AGEMA_signal_5315 ;
    wire new_AGEMA_signal_5316 ;
    wire new_AGEMA_signal_5317 ;
    wire new_AGEMA_signal_5318 ;
    wire new_AGEMA_signal_5319 ;
    wire new_AGEMA_signal_5320 ;
    wire new_AGEMA_signal_5321 ;
    wire new_AGEMA_signal_5322 ;
    wire new_AGEMA_signal_5323 ;
    wire new_AGEMA_signal_5324 ;
    wire new_AGEMA_signal_5325 ;
    wire new_AGEMA_signal_5326 ;
    wire new_AGEMA_signal_5327 ;
    wire new_AGEMA_signal_5328 ;
    wire new_AGEMA_signal_5329 ;
    wire new_AGEMA_signal_5330 ;
    wire new_AGEMA_signal_5331 ;
    wire new_AGEMA_signal_5332 ;
    wire new_AGEMA_signal_5333 ;
    wire new_AGEMA_signal_5334 ;
    wire new_AGEMA_signal_5335 ;
    wire new_AGEMA_signal_5336 ;
    wire new_AGEMA_signal_5337 ;
    wire new_AGEMA_signal_5338 ;
    wire new_AGEMA_signal_5339 ;
    wire new_AGEMA_signal_5340 ;
    wire new_AGEMA_signal_5341 ;
    wire new_AGEMA_signal_5342 ;
    wire new_AGEMA_signal_5343 ;
    wire new_AGEMA_signal_5344 ;
    wire new_AGEMA_signal_5345 ;
    wire new_AGEMA_signal_5346 ;
    wire new_AGEMA_signal_5347 ;
    wire new_AGEMA_signal_5348 ;
    wire new_AGEMA_signal_5349 ;
    wire new_AGEMA_signal_5350 ;
    wire new_AGEMA_signal_5351 ;
    wire new_AGEMA_signal_5352 ;
    wire new_AGEMA_signal_5353 ;
    wire new_AGEMA_signal_5354 ;
    wire new_AGEMA_signal_5355 ;
    wire new_AGEMA_signal_5356 ;
    wire new_AGEMA_signal_5357 ;
    wire new_AGEMA_signal_5358 ;
    wire new_AGEMA_signal_5359 ;
    wire new_AGEMA_signal_5360 ;
    wire new_AGEMA_signal_5361 ;
    wire new_AGEMA_signal_5362 ;
    wire new_AGEMA_signal_5363 ;
    wire new_AGEMA_signal_5364 ;
    wire new_AGEMA_signal_5365 ;
    wire new_AGEMA_signal_5366 ;
    wire new_AGEMA_signal_5367 ;
    wire new_AGEMA_signal_5368 ;
    wire new_AGEMA_signal_5369 ;
    wire new_AGEMA_signal_5370 ;
    wire new_AGEMA_signal_5371 ;
    wire new_AGEMA_signal_5372 ;
    wire new_AGEMA_signal_5373 ;
    wire new_AGEMA_signal_5374 ;
    wire new_AGEMA_signal_5375 ;
    wire new_AGEMA_signal_5376 ;
    wire new_AGEMA_signal_5377 ;
    wire new_AGEMA_signal_5378 ;
    wire new_AGEMA_signal_5379 ;
    wire new_AGEMA_signal_5380 ;
    wire new_AGEMA_signal_5381 ;
    wire new_AGEMA_signal_5382 ;
    wire new_AGEMA_signal_5383 ;
    wire new_AGEMA_signal_5384 ;
    wire new_AGEMA_signal_5385 ;
    wire new_AGEMA_signal_5386 ;
    wire new_AGEMA_signal_5387 ;
    wire new_AGEMA_signal_5388 ;
    wire new_AGEMA_signal_5389 ;
    wire new_AGEMA_signal_5390 ;
    wire new_AGEMA_signal_5391 ;
    wire new_AGEMA_signal_5392 ;
    wire new_AGEMA_signal_5393 ;
    wire new_AGEMA_signal_5394 ;
    wire new_AGEMA_signal_5395 ;
    wire new_AGEMA_signal_5396 ;
    wire new_AGEMA_signal_5397 ;
    wire new_AGEMA_signal_5398 ;
    wire new_AGEMA_signal_5399 ;
    wire new_AGEMA_signal_5400 ;
    wire new_AGEMA_signal_5401 ;
    wire new_AGEMA_signal_5402 ;
    wire new_AGEMA_signal_5403 ;
    wire new_AGEMA_signal_5404 ;
    wire new_AGEMA_signal_5405 ;
    wire new_AGEMA_signal_5406 ;
    wire new_AGEMA_signal_5407 ;
    wire new_AGEMA_signal_5408 ;
    wire new_AGEMA_signal_5409 ;
    wire new_AGEMA_signal_5410 ;
    wire new_AGEMA_signal_5411 ;
    wire new_AGEMA_signal_5412 ;
    wire new_AGEMA_signal_5413 ;
    wire new_AGEMA_signal_5414 ;
    wire new_AGEMA_signal_5415 ;
    wire new_AGEMA_signal_5416 ;
    wire new_AGEMA_signal_5417 ;
    wire new_AGEMA_signal_5418 ;
    wire new_AGEMA_signal_5419 ;
    wire new_AGEMA_signal_5420 ;
    wire new_AGEMA_signal_5421 ;
    wire new_AGEMA_signal_5422 ;
    wire new_AGEMA_signal_5423 ;
    wire new_AGEMA_signal_5424 ;
    wire new_AGEMA_signal_5425 ;
    wire new_AGEMA_signal_5426 ;
    wire new_AGEMA_signal_5427 ;
    wire new_AGEMA_signal_5428 ;
    wire new_AGEMA_signal_5429 ;
    wire new_AGEMA_signal_5430 ;
    wire new_AGEMA_signal_5431 ;
    wire new_AGEMA_signal_5432 ;
    wire new_AGEMA_signal_5433 ;
    wire new_AGEMA_signal_5434 ;
    wire new_AGEMA_signal_5435 ;
    wire new_AGEMA_signal_5436 ;
    wire new_AGEMA_signal_5437 ;
    wire new_AGEMA_signal_5438 ;
    wire new_AGEMA_signal_5439 ;
    wire new_AGEMA_signal_5440 ;
    wire new_AGEMA_signal_5441 ;
    wire new_AGEMA_signal_5442 ;
    wire new_AGEMA_signal_5443 ;
    wire new_AGEMA_signal_5444 ;
    wire new_AGEMA_signal_5445 ;
    wire new_AGEMA_signal_5446 ;
    wire new_AGEMA_signal_5447 ;
    wire new_AGEMA_signal_5448 ;
    wire new_AGEMA_signal_5449 ;
    wire new_AGEMA_signal_5450 ;
    wire new_AGEMA_signal_5451 ;
    wire new_AGEMA_signal_5452 ;
    wire new_AGEMA_signal_5453 ;
    wire new_AGEMA_signal_5454 ;
    wire new_AGEMA_signal_5455 ;
    wire new_AGEMA_signal_5456 ;
    wire new_AGEMA_signal_5457 ;
    wire new_AGEMA_signal_5458 ;
    wire new_AGEMA_signal_5459 ;
    wire new_AGEMA_signal_5460 ;
    wire new_AGEMA_signal_5461 ;
    wire new_AGEMA_signal_5462 ;
    wire new_AGEMA_signal_5463 ;
    wire new_AGEMA_signal_5464 ;
    wire new_AGEMA_signal_5465 ;
    wire new_AGEMA_signal_5466 ;
    wire new_AGEMA_signal_5467 ;
    wire new_AGEMA_signal_5468 ;
    wire new_AGEMA_signal_5469 ;
    wire new_AGEMA_signal_5470 ;
    wire new_AGEMA_signal_5471 ;
    wire new_AGEMA_signal_5472 ;
    wire new_AGEMA_signal_5473 ;
    wire new_AGEMA_signal_5474 ;
    wire new_AGEMA_signal_5475 ;
    wire new_AGEMA_signal_5476 ;
    wire new_AGEMA_signal_5477 ;
    wire new_AGEMA_signal_5478 ;
    wire new_AGEMA_signal_5479 ;
    wire new_AGEMA_signal_5480 ;
    wire new_AGEMA_signal_5481 ;
    wire new_AGEMA_signal_5482 ;
    wire new_AGEMA_signal_5483 ;
    wire new_AGEMA_signal_5484 ;
    wire new_AGEMA_signal_5485 ;
    wire new_AGEMA_signal_5486 ;
    wire new_AGEMA_signal_5487 ;
    wire new_AGEMA_signal_5488 ;
    wire new_AGEMA_signal_5489 ;
    wire new_AGEMA_signal_5490 ;
    wire new_AGEMA_signal_5491 ;
    wire new_AGEMA_signal_5492 ;
    wire new_AGEMA_signal_5493 ;
    wire new_AGEMA_signal_5494 ;
    wire new_AGEMA_signal_5495 ;
    wire new_AGEMA_signal_5496 ;
    wire new_AGEMA_signal_5497 ;
    wire new_AGEMA_signal_5498 ;
    wire new_AGEMA_signal_5499 ;
    wire new_AGEMA_signal_5500 ;
    wire new_AGEMA_signal_5501 ;
    wire new_AGEMA_signal_5502 ;
    wire new_AGEMA_signal_5503 ;
    wire new_AGEMA_signal_5504 ;
    wire new_AGEMA_signal_5505 ;
    wire new_AGEMA_signal_5506 ;
    wire new_AGEMA_signal_5507 ;
    wire new_AGEMA_signal_5508 ;
    wire new_AGEMA_signal_5509 ;
    wire new_AGEMA_signal_5510 ;
    wire new_AGEMA_signal_5511 ;
    wire new_AGEMA_signal_5512 ;
    wire new_AGEMA_signal_5513 ;
    wire new_AGEMA_signal_5514 ;
    wire new_AGEMA_signal_5515 ;
    wire new_AGEMA_signal_5516 ;
    wire new_AGEMA_signal_5517 ;
    wire new_AGEMA_signal_5518 ;
    wire new_AGEMA_signal_5519 ;
    wire new_AGEMA_signal_5520 ;
    wire new_AGEMA_signal_5521 ;
    wire new_AGEMA_signal_5522 ;
    wire new_AGEMA_signal_5523 ;
    wire new_AGEMA_signal_5524 ;
    wire new_AGEMA_signal_5525 ;
    wire new_AGEMA_signal_5526 ;
    wire new_AGEMA_signal_5527 ;
    wire new_AGEMA_signal_5528 ;
    wire new_AGEMA_signal_5529 ;
    wire new_AGEMA_signal_5530 ;
    wire new_AGEMA_signal_5531 ;
    wire new_AGEMA_signal_5532 ;
    wire new_AGEMA_signal_5533 ;
    wire new_AGEMA_signal_5534 ;
    wire new_AGEMA_signal_5535 ;
    wire new_AGEMA_signal_5536 ;
    wire new_AGEMA_signal_5537 ;
    wire new_AGEMA_signal_5538 ;
    wire new_AGEMA_signal_5539 ;
    wire new_AGEMA_signal_5540 ;
    wire new_AGEMA_signal_5541 ;
    wire new_AGEMA_signal_5542 ;
    wire new_AGEMA_signal_5543 ;
    wire new_AGEMA_signal_5544 ;
    wire new_AGEMA_signal_5545 ;
    wire new_AGEMA_signal_5546 ;
    wire new_AGEMA_signal_5547 ;
    wire new_AGEMA_signal_5548 ;
    wire new_AGEMA_signal_5549 ;
    wire new_AGEMA_signal_5550 ;
    wire new_AGEMA_signal_5551 ;
    wire new_AGEMA_signal_5552 ;
    wire new_AGEMA_signal_5553 ;
    wire new_AGEMA_signal_5554 ;
    wire new_AGEMA_signal_5555 ;
    wire new_AGEMA_signal_5556 ;
    wire new_AGEMA_signal_5557 ;
    wire new_AGEMA_signal_5558 ;
    wire new_AGEMA_signal_5559 ;
    wire new_AGEMA_signal_5560 ;
    wire new_AGEMA_signal_5561 ;
    wire new_AGEMA_signal_5562 ;
    wire new_AGEMA_signal_5563 ;
    wire new_AGEMA_signal_5564 ;
    wire new_AGEMA_signal_5565 ;
    wire new_AGEMA_signal_5566 ;
    wire new_AGEMA_signal_5567 ;
    wire new_AGEMA_signal_5568 ;
    wire new_AGEMA_signal_5569 ;
    wire new_AGEMA_signal_5570 ;
    wire new_AGEMA_signal_5571 ;
    wire new_AGEMA_signal_5572 ;
    wire new_AGEMA_signal_5573 ;
    wire new_AGEMA_signal_5574 ;
    wire new_AGEMA_signal_5575 ;
    wire new_AGEMA_signal_5576 ;
    wire new_AGEMA_signal_5577 ;
    wire new_AGEMA_signal_5578 ;
    wire new_AGEMA_signal_5579 ;
    wire new_AGEMA_signal_5580 ;
    wire new_AGEMA_signal_5581 ;
    wire new_AGEMA_signal_5582 ;
    wire new_AGEMA_signal_5583 ;
    wire new_AGEMA_signal_5584 ;
    wire new_AGEMA_signal_5585 ;
    wire new_AGEMA_signal_5586 ;
    wire new_AGEMA_signal_5587 ;
    wire new_AGEMA_signal_5588 ;
    wire new_AGEMA_signal_5589 ;
    wire new_AGEMA_signal_5590 ;
    wire new_AGEMA_signal_5591 ;
    wire new_AGEMA_signal_5592 ;
    wire new_AGEMA_signal_5593 ;
    wire new_AGEMA_signal_5594 ;
    wire new_AGEMA_signal_5595 ;
    wire new_AGEMA_signal_5596 ;
    wire new_AGEMA_signal_5597 ;
    wire new_AGEMA_signal_5598 ;
    wire new_AGEMA_signal_5599 ;
    wire new_AGEMA_signal_5600 ;
    wire new_AGEMA_signal_5601 ;
    wire new_AGEMA_signal_5602 ;
    wire new_AGEMA_signal_5603 ;
    wire new_AGEMA_signal_5604 ;
    wire new_AGEMA_signal_5605 ;
    wire new_AGEMA_signal_5606 ;
    wire new_AGEMA_signal_5607 ;
    wire new_AGEMA_signal_5608 ;
    wire new_AGEMA_signal_5609 ;
    wire new_AGEMA_signal_5610 ;
    wire new_AGEMA_signal_5611 ;
    wire new_AGEMA_signal_5612 ;
    wire new_AGEMA_signal_5613 ;
    wire new_AGEMA_signal_5614 ;
    wire new_AGEMA_signal_5615 ;
    wire new_AGEMA_signal_5616 ;
    wire new_AGEMA_signal_5617 ;
    wire new_AGEMA_signal_5618 ;
    wire new_AGEMA_signal_5619 ;
    wire new_AGEMA_signal_5620 ;
    wire new_AGEMA_signal_5621 ;
    wire new_AGEMA_signal_5622 ;
    wire new_AGEMA_signal_5623 ;
    wire new_AGEMA_signal_5624 ;
    wire new_AGEMA_signal_5625 ;
    wire new_AGEMA_signal_5626 ;
    wire new_AGEMA_signal_5627 ;
    wire new_AGEMA_signal_5628 ;
    wire new_AGEMA_signal_5629 ;
    wire new_AGEMA_signal_5630 ;
    wire new_AGEMA_signal_5631 ;
    wire new_AGEMA_signal_5632 ;
    wire new_AGEMA_signal_5633 ;
    wire new_AGEMA_signal_5634 ;
    wire new_AGEMA_signal_5635 ;
    wire new_AGEMA_signal_5636 ;
    wire new_AGEMA_signal_5637 ;
    wire new_AGEMA_signal_5638 ;
    wire new_AGEMA_signal_5639 ;
    wire new_AGEMA_signal_5640 ;
    wire new_AGEMA_signal_5641 ;
    wire new_AGEMA_signal_5642 ;
    wire new_AGEMA_signal_5643 ;
    wire new_AGEMA_signal_5644 ;
    wire new_AGEMA_signal_5645 ;
    wire new_AGEMA_signal_5646 ;
    wire new_AGEMA_signal_5647 ;
    wire new_AGEMA_signal_5648 ;
    wire new_AGEMA_signal_5649 ;
    wire new_AGEMA_signal_5650 ;
    wire new_AGEMA_signal_5651 ;
    wire new_AGEMA_signal_5652 ;
    wire new_AGEMA_signal_5653 ;
    wire new_AGEMA_signal_5654 ;
    wire new_AGEMA_signal_5655 ;
    wire new_AGEMA_signal_5656 ;
    wire new_AGEMA_signal_5657 ;
    wire new_AGEMA_signal_5658 ;
    wire new_AGEMA_signal_5659 ;
    wire new_AGEMA_signal_5660 ;
    wire new_AGEMA_signal_5661 ;
    wire new_AGEMA_signal_5662 ;
    wire new_AGEMA_signal_5663 ;
    wire new_AGEMA_signal_5664 ;
    wire new_AGEMA_signal_5665 ;
    wire new_AGEMA_signal_5666 ;
    wire new_AGEMA_signal_5667 ;
    wire new_AGEMA_signal_5668 ;
    wire new_AGEMA_signal_5669 ;
    wire new_AGEMA_signal_5670 ;
    wire new_AGEMA_signal_5671 ;
    wire new_AGEMA_signal_5672 ;
    wire new_AGEMA_signal_5673 ;
    wire new_AGEMA_signal_5674 ;
    wire new_AGEMA_signal_5675 ;
    wire new_AGEMA_signal_5676 ;
    wire new_AGEMA_signal_5677 ;
    wire new_AGEMA_signal_5678 ;
    wire new_AGEMA_signal_5679 ;
    wire new_AGEMA_signal_5680 ;
    wire new_AGEMA_signal_5681 ;
    wire new_AGEMA_signal_5682 ;
    wire new_AGEMA_signal_5683 ;
    wire new_AGEMA_signal_5684 ;
    wire new_AGEMA_signal_5685 ;
    wire new_AGEMA_signal_5686 ;
    wire new_AGEMA_signal_5687 ;
    wire new_AGEMA_signal_5688 ;
    wire new_AGEMA_signal_5689 ;
    wire new_AGEMA_signal_5690 ;
    wire new_AGEMA_signal_5691 ;
    wire new_AGEMA_signal_5692 ;
    wire new_AGEMA_signal_5693 ;
    wire new_AGEMA_signal_5694 ;
    wire new_AGEMA_signal_5695 ;
    wire new_AGEMA_signal_5696 ;
    wire new_AGEMA_signal_5697 ;
    wire new_AGEMA_signal_5698 ;
    wire new_AGEMA_signal_5699 ;
    wire new_AGEMA_signal_5700 ;
    wire new_AGEMA_signal_5701 ;
    wire new_AGEMA_signal_5702 ;
    wire new_AGEMA_signal_5703 ;
    wire new_AGEMA_signal_5704 ;
    wire new_AGEMA_signal_5705 ;
    wire new_AGEMA_signal_5706 ;
    wire new_AGEMA_signal_5707 ;
    wire new_AGEMA_signal_5708 ;
    wire new_AGEMA_signal_5709 ;
    wire new_AGEMA_signal_5710 ;
    wire new_AGEMA_signal_5711 ;
    wire new_AGEMA_signal_5712 ;
    wire new_AGEMA_signal_5713 ;
    wire new_AGEMA_signal_5714 ;
    wire new_AGEMA_signal_5715 ;
    wire new_AGEMA_signal_5716 ;
    wire new_AGEMA_signal_5717 ;
    wire new_AGEMA_signal_5718 ;
    wire new_AGEMA_signal_5719 ;
    wire new_AGEMA_signal_5720 ;
    wire new_AGEMA_signal_5721 ;
    wire new_AGEMA_signal_5722 ;
    wire new_AGEMA_signal_5723 ;
    wire new_AGEMA_signal_5724 ;
    wire new_AGEMA_signal_5725 ;
    wire new_AGEMA_signal_5726 ;
    wire new_AGEMA_signal_5727 ;
    wire new_AGEMA_signal_5728 ;
    wire new_AGEMA_signal_5729 ;
    wire new_AGEMA_signal_5730 ;
    wire new_AGEMA_signal_5731 ;
    wire new_AGEMA_signal_5732 ;
    wire new_AGEMA_signal_5733 ;
    wire new_AGEMA_signal_5734 ;
    wire new_AGEMA_signal_5735 ;
    wire new_AGEMA_signal_5736 ;
    wire new_AGEMA_signal_5737 ;
    wire new_AGEMA_signal_5738 ;
    wire new_AGEMA_signal_5739 ;
    wire new_AGEMA_signal_5740 ;
    wire new_AGEMA_signal_5741 ;
    wire new_AGEMA_signal_5742 ;
    wire new_AGEMA_signal_5743 ;
    wire new_AGEMA_signal_5744 ;
    wire new_AGEMA_signal_5745 ;
    wire new_AGEMA_signal_5746 ;
    wire new_AGEMA_signal_5747 ;
    wire new_AGEMA_signal_5748 ;
    wire new_AGEMA_signal_5749 ;
    wire new_AGEMA_signal_5750 ;
    wire new_AGEMA_signal_5751 ;
    wire new_AGEMA_signal_5752 ;
    wire new_AGEMA_signal_5753 ;
    wire new_AGEMA_signal_5754 ;
    wire new_AGEMA_signal_5755 ;
    wire new_AGEMA_signal_5756 ;
    wire new_AGEMA_signal_5757 ;
    wire new_AGEMA_signal_5758 ;
    wire new_AGEMA_signal_5759 ;
    wire new_AGEMA_signal_5760 ;
    wire new_AGEMA_signal_5761 ;
    wire new_AGEMA_signal_5762 ;
    wire new_AGEMA_signal_5763 ;
    wire new_AGEMA_signal_5764 ;
    wire new_AGEMA_signal_5765 ;
    wire new_AGEMA_signal_5766 ;
    wire new_AGEMA_signal_5767 ;
    wire new_AGEMA_signal_5768 ;
    wire new_AGEMA_signal_5769 ;
    wire new_AGEMA_signal_5770 ;
    wire new_AGEMA_signal_5771 ;
    wire new_AGEMA_signal_5772 ;
    wire new_AGEMA_signal_5773 ;
    wire new_AGEMA_signal_5774 ;
    wire new_AGEMA_signal_5775 ;
    wire new_AGEMA_signal_5776 ;
    wire new_AGEMA_signal_5777 ;
    wire new_AGEMA_signal_5778 ;
    wire new_AGEMA_signal_5779 ;
    wire new_AGEMA_signal_5780 ;
    wire new_AGEMA_signal_5781 ;
    wire new_AGEMA_signal_5782 ;
    wire new_AGEMA_signal_5783 ;
    wire new_AGEMA_signal_5784 ;
    wire new_AGEMA_signal_5785 ;
    wire new_AGEMA_signal_5786 ;
    wire new_AGEMA_signal_5787 ;
    wire new_AGEMA_signal_5788 ;
    wire new_AGEMA_signal_5789 ;
    wire new_AGEMA_signal_5790 ;
    wire new_AGEMA_signal_5791 ;
    wire new_AGEMA_signal_5792 ;
    wire new_AGEMA_signal_5793 ;
    wire new_AGEMA_signal_5794 ;
    wire new_AGEMA_signal_5795 ;
    wire new_AGEMA_signal_5796 ;
    wire new_AGEMA_signal_5797 ;
    wire new_AGEMA_signal_5798 ;
    wire new_AGEMA_signal_5799 ;
    wire new_AGEMA_signal_5800 ;
    wire new_AGEMA_signal_5801 ;
    wire new_AGEMA_signal_5802 ;
    wire new_AGEMA_signal_5803 ;
    wire new_AGEMA_signal_5804 ;
    wire new_AGEMA_signal_5805 ;
    wire new_AGEMA_signal_5806 ;
    wire new_AGEMA_signal_5807 ;
    wire new_AGEMA_signal_5808 ;
    wire new_AGEMA_signal_5809 ;
    wire new_AGEMA_signal_5810 ;
    wire new_AGEMA_signal_5811 ;
    wire new_AGEMA_signal_5812 ;
    wire new_AGEMA_signal_5813 ;
    wire new_AGEMA_signal_5814 ;
    wire new_AGEMA_signal_5815 ;
    wire new_AGEMA_signal_5816 ;
    wire new_AGEMA_signal_5817 ;
    wire new_AGEMA_signal_5818 ;
    wire new_AGEMA_signal_5819 ;
    wire new_AGEMA_signal_5820 ;
    wire new_AGEMA_signal_5821 ;
    wire new_AGEMA_signal_5822 ;
    wire new_AGEMA_signal_5823 ;
    wire new_AGEMA_signal_5824 ;
    wire new_AGEMA_signal_5825 ;
    wire new_AGEMA_signal_5826 ;
    wire new_AGEMA_signal_5827 ;
    wire new_AGEMA_signal_5828 ;
    wire new_AGEMA_signal_5829 ;
    wire new_AGEMA_signal_5830 ;
    wire new_AGEMA_signal_5831 ;
    wire new_AGEMA_signal_5832 ;
    wire new_AGEMA_signal_5833 ;
    wire new_AGEMA_signal_5834 ;
    wire new_AGEMA_signal_5835 ;
    wire new_AGEMA_signal_5836 ;
    wire new_AGEMA_signal_5837 ;
    wire new_AGEMA_signal_5838 ;
    wire new_AGEMA_signal_5839 ;
    wire new_AGEMA_signal_5840 ;
    wire new_AGEMA_signal_5841 ;
    wire new_AGEMA_signal_5842 ;
    wire new_AGEMA_signal_5843 ;
    wire new_AGEMA_signal_5844 ;
    wire new_AGEMA_signal_5845 ;
    wire new_AGEMA_signal_5846 ;
    wire new_AGEMA_signal_5847 ;
    wire new_AGEMA_signal_5848 ;
    wire new_AGEMA_signal_5849 ;
    wire new_AGEMA_signal_5850 ;
    wire new_AGEMA_signal_5851 ;
    wire new_AGEMA_signal_5852 ;
    wire new_AGEMA_signal_5853 ;
    wire new_AGEMA_signal_5854 ;
    wire new_AGEMA_signal_5855 ;
    wire new_AGEMA_signal_5856 ;
    wire new_AGEMA_signal_5857 ;
    wire new_AGEMA_signal_5858 ;
    wire new_AGEMA_signal_5859 ;
    wire new_AGEMA_signal_5860 ;
    wire new_AGEMA_signal_5861 ;
    wire new_AGEMA_signal_5862 ;
    wire new_AGEMA_signal_5863 ;
    wire new_AGEMA_signal_5864 ;
    wire new_AGEMA_signal_5865 ;
    wire new_AGEMA_signal_5866 ;
    wire new_AGEMA_signal_5867 ;
    wire new_AGEMA_signal_5868 ;
    wire new_AGEMA_signal_5869 ;
    wire new_AGEMA_signal_5870 ;
    wire new_AGEMA_signal_5871 ;
    wire new_AGEMA_signal_5872 ;
    wire new_AGEMA_signal_5873 ;
    wire new_AGEMA_signal_5874 ;
    wire new_AGEMA_signal_5875 ;
    wire new_AGEMA_signal_5876 ;
    wire new_AGEMA_signal_5877 ;
    wire new_AGEMA_signal_5878 ;
    wire new_AGEMA_signal_5879 ;
    wire new_AGEMA_signal_5880 ;
    wire new_AGEMA_signal_5881 ;
    wire new_AGEMA_signal_5882 ;
    wire new_AGEMA_signal_5883 ;
    wire new_AGEMA_signal_5884 ;
    wire new_AGEMA_signal_5885 ;
    wire new_AGEMA_signal_5886 ;
    wire new_AGEMA_signal_5887 ;
    wire new_AGEMA_signal_5888 ;
    wire new_AGEMA_signal_5889 ;
    wire new_AGEMA_signal_5890 ;
    wire new_AGEMA_signal_5891 ;
    wire new_AGEMA_signal_5892 ;
    wire new_AGEMA_signal_5893 ;
    wire new_AGEMA_signal_5894 ;
    wire new_AGEMA_signal_5895 ;
    wire new_AGEMA_signal_5896 ;
    wire new_AGEMA_signal_5897 ;
    wire new_AGEMA_signal_5898 ;
    wire new_AGEMA_signal_5899 ;
    wire new_AGEMA_signal_5900 ;
    wire new_AGEMA_signal_5901 ;
    wire new_AGEMA_signal_5902 ;
    wire new_AGEMA_signal_5903 ;
    wire new_AGEMA_signal_5904 ;
    wire new_AGEMA_signal_5905 ;
    wire new_AGEMA_signal_5906 ;
    wire new_AGEMA_signal_5907 ;
    wire new_AGEMA_signal_5908 ;
    wire new_AGEMA_signal_5909 ;
    wire new_AGEMA_signal_5910 ;
    wire new_AGEMA_signal_5911 ;
    wire new_AGEMA_signal_5912 ;
    wire new_AGEMA_signal_5913 ;
    wire new_AGEMA_signal_5914 ;
    wire new_AGEMA_signal_5915 ;
    wire new_AGEMA_signal_5916 ;
    wire new_AGEMA_signal_5917 ;
    wire new_AGEMA_signal_5918 ;
    wire new_AGEMA_signal_5919 ;
    wire new_AGEMA_signal_5920 ;
    wire new_AGEMA_signal_5921 ;
    wire new_AGEMA_signal_5922 ;
    wire new_AGEMA_signal_5923 ;
    wire new_AGEMA_signal_5924 ;
    wire new_AGEMA_signal_5925 ;
    wire new_AGEMA_signal_5926 ;
    wire new_AGEMA_signal_5927 ;
    wire new_AGEMA_signal_5928 ;
    wire new_AGEMA_signal_5929 ;
    wire new_AGEMA_signal_5930 ;
    wire new_AGEMA_signal_5931 ;
    wire new_AGEMA_signal_5932 ;
    wire new_AGEMA_signal_5933 ;
    wire new_AGEMA_signal_5934 ;
    wire new_AGEMA_signal_5935 ;
    wire new_AGEMA_signal_5936 ;
    wire new_AGEMA_signal_5937 ;
    wire new_AGEMA_signal_5938 ;
    wire new_AGEMA_signal_5939 ;
    wire new_AGEMA_signal_5940 ;
    wire new_AGEMA_signal_5941 ;
    wire new_AGEMA_signal_5942 ;
    wire new_AGEMA_signal_5943 ;
    wire new_AGEMA_signal_5944 ;
    wire new_AGEMA_signal_5945 ;
    wire new_AGEMA_signal_5946 ;
    wire new_AGEMA_signal_5947 ;
    wire new_AGEMA_signal_5948 ;
    wire new_AGEMA_signal_5949 ;
    wire new_AGEMA_signal_5950 ;
    wire new_AGEMA_signal_5951 ;
    wire new_AGEMA_signal_5952 ;
    wire new_AGEMA_signal_5953 ;
    wire new_AGEMA_signal_5954 ;
    wire new_AGEMA_signal_5955 ;
    wire new_AGEMA_signal_5956 ;
    wire new_AGEMA_signal_5957 ;
    wire new_AGEMA_signal_5958 ;
    wire new_AGEMA_signal_5959 ;
    wire new_AGEMA_signal_5960 ;
    wire new_AGEMA_signal_5961 ;
    wire new_AGEMA_signal_5962 ;
    wire new_AGEMA_signal_5963 ;
    wire new_AGEMA_signal_5964 ;
    wire new_AGEMA_signal_5965 ;
    wire new_AGEMA_signal_5966 ;
    wire new_AGEMA_signal_5967 ;
    wire new_AGEMA_signal_5968 ;
    wire new_AGEMA_signal_5969 ;
    wire new_AGEMA_signal_5970 ;
    wire new_AGEMA_signal_5971 ;
    wire new_AGEMA_signal_5972 ;
    wire new_AGEMA_signal_5973 ;
    wire new_AGEMA_signal_5974 ;
    wire new_AGEMA_signal_5975 ;
    wire new_AGEMA_signal_5976 ;
    wire new_AGEMA_signal_5977 ;
    wire new_AGEMA_signal_5978 ;
    wire new_AGEMA_signal_5979 ;
    wire new_AGEMA_signal_5980 ;
    wire new_AGEMA_signal_5981 ;
    wire new_AGEMA_signal_5982 ;
    wire new_AGEMA_signal_5983 ;
    wire new_AGEMA_signal_5984 ;
    wire new_AGEMA_signal_5985 ;
    wire new_AGEMA_signal_5986 ;
    wire new_AGEMA_signal_5987 ;
    wire new_AGEMA_signal_5988 ;
    wire new_AGEMA_signal_5989 ;
    wire new_AGEMA_signal_5990 ;
    wire new_AGEMA_signal_5991 ;
    wire new_AGEMA_signal_5992 ;
    wire new_AGEMA_signal_5993 ;
    wire new_AGEMA_signal_5994 ;
    wire new_AGEMA_signal_5995 ;
    wire new_AGEMA_signal_5996 ;
    wire new_AGEMA_signal_5997 ;
    wire new_AGEMA_signal_5998 ;
    wire new_AGEMA_signal_5999 ;
    wire new_AGEMA_signal_6000 ;
    wire new_AGEMA_signal_6001 ;
    wire new_AGEMA_signal_6002 ;
    wire new_AGEMA_signal_6003 ;
    wire new_AGEMA_signal_6004 ;
    wire new_AGEMA_signal_6005 ;
    wire new_AGEMA_signal_6006 ;
    wire new_AGEMA_signal_6007 ;
    wire new_AGEMA_signal_6008 ;
    wire new_AGEMA_signal_6009 ;
    wire new_AGEMA_signal_6010 ;
    wire new_AGEMA_signal_6011 ;
    wire new_AGEMA_signal_6012 ;
    wire new_AGEMA_signal_6013 ;
    wire new_AGEMA_signal_6014 ;
    wire new_AGEMA_signal_6015 ;
    wire new_AGEMA_signal_6016 ;
    wire new_AGEMA_signal_6017 ;
    wire new_AGEMA_signal_6018 ;
    wire new_AGEMA_signal_6019 ;
    wire new_AGEMA_signal_6020 ;
    wire new_AGEMA_signal_6021 ;
    wire new_AGEMA_signal_6022 ;
    wire new_AGEMA_signal_6023 ;
    wire new_AGEMA_signal_6024 ;
    wire new_AGEMA_signal_6025 ;
    wire new_AGEMA_signal_6026 ;
    wire new_AGEMA_signal_6027 ;
    wire new_AGEMA_signal_6028 ;
    wire new_AGEMA_signal_6029 ;
    wire new_AGEMA_signal_6030 ;
    wire new_AGEMA_signal_6031 ;
    wire new_AGEMA_signal_6032 ;
    wire new_AGEMA_signal_6033 ;
    wire new_AGEMA_signal_6034 ;
    wire new_AGEMA_signal_6035 ;
    wire new_AGEMA_signal_6036 ;
    wire new_AGEMA_signal_6037 ;
    wire new_AGEMA_signal_6038 ;
    wire new_AGEMA_signal_6039 ;
    wire new_AGEMA_signal_6040 ;
    wire new_AGEMA_signal_6041 ;
    wire new_AGEMA_signal_6042 ;
    wire new_AGEMA_signal_6043 ;
    wire new_AGEMA_signal_6044 ;
    wire new_AGEMA_signal_6045 ;
    wire new_AGEMA_signal_6046 ;
    wire new_AGEMA_signal_6047 ;
    wire new_AGEMA_signal_6048 ;
    wire new_AGEMA_signal_6049 ;
    wire new_AGEMA_signal_6050 ;
    wire new_AGEMA_signal_6051 ;
    wire new_AGEMA_signal_6052 ;
    wire new_AGEMA_signal_6053 ;
    wire new_AGEMA_signal_6054 ;
    wire new_AGEMA_signal_6055 ;
    wire new_AGEMA_signal_6056 ;
    wire new_AGEMA_signal_6057 ;
    wire new_AGEMA_signal_6058 ;
    wire new_AGEMA_signal_6059 ;
    wire new_AGEMA_signal_6060 ;
    wire new_AGEMA_signal_6061 ;
    wire new_AGEMA_signal_6062 ;
    wire new_AGEMA_signal_6063 ;
    wire new_AGEMA_signal_6064 ;
    wire new_AGEMA_signal_6065 ;
    wire new_AGEMA_signal_6066 ;
    wire new_AGEMA_signal_6067 ;
    wire new_AGEMA_signal_6068 ;
    wire new_AGEMA_signal_6069 ;
    wire new_AGEMA_signal_6070 ;
    wire new_AGEMA_signal_6071 ;
    wire new_AGEMA_signal_6072 ;
    wire new_AGEMA_signal_6073 ;
    wire new_AGEMA_signal_6074 ;
    wire new_AGEMA_signal_6075 ;
    wire new_AGEMA_signal_6076 ;
    wire new_AGEMA_signal_6077 ;
    wire new_AGEMA_signal_6078 ;
    wire new_AGEMA_signal_6079 ;
    wire new_AGEMA_signal_6080 ;
    wire new_AGEMA_signal_6081 ;
    wire new_AGEMA_signal_6082 ;
    wire new_AGEMA_signal_6083 ;
    wire new_AGEMA_signal_6084 ;
    wire new_AGEMA_signal_6085 ;
    wire new_AGEMA_signal_6086 ;
    wire new_AGEMA_signal_6087 ;
    wire new_AGEMA_signal_6088 ;
    wire new_AGEMA_signal_6089 ;
    wire new_AGEMA_signal_6090 ;
    wire new_AGEMA_signal_6091 ;
    wire new_AGEMA_signal_6092 ;
    wire new_AGEMA_signal_6093 ;
    wire new_AGEMA_signal_6094 ;
    wire new_AGEMA_signal_6095 ;
    wire new_AGEMA_signal_6096 ;
    wire new_AGEMA_signal_6097 ;
    wire new_AGEMA_signal_6098 ;
    wire new_AGEMA_signal_6099 ;
    wire new_AGEMA_signal_6100 ;
    wire new_AGEMA_signal_6101 ;
    wire new_AGEMA_signal_6102 ;
    wire new_AGEMA_signal_6103 ;
    wire new_AGEMA_signal_6104 ;
    wire new_AGEMA_signal_6105 ;
    wire new_AGEMA_signal_6106 ;
    wire new_AGEMA_signal_6107 ;
    wire new_AGEMA_signal_6108 ;
    wire new_AGEMA_signal_6109 ;
    wire new_AGEMA_signal_6110 ;
    wire new_AGEMA_signal_6111 ;
    wire new_AGEMA_signal_6112 ;
    wire new_AGEMA_signal_6113 ;
    wire new_AGEMA_signal_6114 ;
    wire new_AGEMA_signal_6115 ;
    wire new_AGEMA_signal_6116 ;
    wire new_AGEMA_signal_6117 ;
    wire new_AGEMA_signal_6118 ;
    wire new_AGEMA_signal_6119 ;
    wire new_AGEMA_signal_6120 ;
    wire new_AGEMA_signal_6121 ;
    wire new_AGEMA_signal_6122 ;
    wire new_AGEMA_signal_6123 ;
    wire new_AGEMA_signal_6124 ;
    wire new_AGEMA_signal_6125 ;
    wire new_AGEMA_signal_6126 ;
    wire new_AGEMA_signal_6127 ;
    wire new_AGEMA_signal_6128 ;
    wire new_AGEMA_signal_6129 ;
    wire new_AGEMA_signal_6130 ;
    wire new_AGEMA_signal_6131 ;
    wire new_AGEMA_signal_6132 ;
    wire new_AGEMA_signal_6133 ;
    wire new_AGEMA_signal_6134 ;
    wire new_AGEMA_signal_6135 ;
    wire new_AGEMA_signal_6136 ;
    wire new_AGEMA_signal_6137 ;
    wire new_AGEMA_signal_6138 ;
    wire new_AGEMA_signal_6139 ;
    wire new_AGEMA_signal_6140 ;
    wire new_AGEMA_signal_6141 ;
    wire new_AGEMA_signal_6142 ;
    wire new_AGEMA_signal_6143 ;
    wire new_AGEMA_signal_6144 ;
    wire new_AGEMA_signal_6145 ;
    wire new_AGEMA_signal_6146 ;
    wire new_AGEMA_signal_6147 ;
    wire new_AGEMA_signal_6148 ;
    wire new_AGEMA_signal_6149 ;
    wire new_AGEMA_signal_6150 ;
    wire new_AGEMA_signal_6151 ;
    wire new_AGEMA_signal_6152 ;
    wire new_AGEMA_signal_6153 ;
    wire new_AGEMA_signal_6154 ;
    wire new_AGEMA_signal_6155 ;
    wire new_AGEMA_signal_6156 ;
    wire new_AGEMA_signal_6157 ;
    wire new_AGEMA_signal_6158 ;
    wire new_AGEMA_signal_6159 ;
    wire new_AGEMA_signal_6160 ;
    wire new_AGEMA_signal_6161 ;
    wire new_AGEMA_signal_6162 ;
    wire new_AGEMA_signal_6163 ;
    wire new_AGEMA_signal_6164 ;
    wire new_AGEMA_signal_6165 ;
    wire new_AGEMA_signal_6166 ;
    wire new_AGEMA_signal_6167 ;
    wire new_AGEMA_signal_6168 ;
    wire new_AGEMA_signal_6169 ;
    wire new_AGEMA_signal_6170 ;
    wire new_AGEMA_signal_6171 ;
    wire new_AGEMA_signal_6172 ;
    wire new_AGEMA_signal_6173 ;
    wire new_AGEMA_signal_6174 ;
    wire new_AGEMA_signal_6175 ;
    wire new_AGEMA_signal_6176 ;
    wire new_AGEMA_signal_6177 ;
    wire new_AGEMA_signal_6178 ;
    wire new_AGEMA_signal_6179 ;
    wire new_AGEMA_signal_6180 ;
    wire new_AGEMA_signal_6181 ;
    wire new_AGEMA_signal_6182 ;
    wire new_AGEMA_signal_6183 ;
    wire new_AGEMA_signal_6184 ;
    wire new_AGEMA_signal_6185 ;
    wire new_AGEMA_signal_6186 ;
    wire new_AGEMA_signal_6187 ;
    wire new_AGEMA_signal_6188 ;
    wire new_AGEMA_signal_6189 ;
    wire new_AGEMA_signal_6190 ;
    wire new_AGEMA_signal_6191 ;
    wire new_AGEMA_signal_6192 ;
    wire new_AGEMA_signal_6193 ;
    wire new_AGEMA_signal_6194 ;
    wire new_AGEMA_signal_6195 ;
    wire new_AGEMA_signal_6196 ;
    wire new_AGEMA_signal_6197 ;
    wire new_AGEMA_signal_6198 ;
    wire new_AGEMA_signal_6199 ;
    wire new_AGEMA_signal_6200 ;
    wire new_AGEMA_signal_6201 ;
    wire new_AGEMA_signal_6202 ;
    wire new_AGEMA_signal_6203 ;
    wire new_AGEMA_signal_6204 ;
    wire new_AGEMA_signal_6205 ;
    wire new_AGEMA_signal_6206 ;
    wire new_AGEMA_signal_6207 ;
    wire new_AGEMA_signal_6208 ;
    wire new_AGEMA_signal_6209 ;
    wire new_AGEMA_signal_6210 ;
    wire new_AGEMA_signal_6211 ;
    wire new_AGEMA_signal_6212 ;
    wire new_AGEMA_signal_6213 ;
    wire new_AGEMA_signal_6214 ;
    wire new_AGEMA_signal_6215 ;
    wire new_AGEMA_signal_6216 ;
    wire new_AGEMA_signal_6217 ;
    wire new_AGEMA_signal_6218 ;
    wire new_AGEMA_signal_6219 ;
    wire new_AGEMA_signal_6220 ;
    wire new_AGEMA_signal_6221 ;
    wire new_AGEMA_signal_6222 ;
    wire new_AGEMA_signal_6223 ;
    wire new_AGEMA_signal_6224 ;
    wire new_AGEMA_signal_6225 ;
    wire new_AGEMA_signal_6226 ;
    wire new_AGEMA_signal_6227 ;
    wire new_AGEMA_signal_6228 ;
    wire new_AGEMA_signal_6229 ;
    wire new_AGEMA_signal_6230 ;
    wire new_AGEMA_signal_6231 ;
    wire new_AGEMA_signal_6232 ;
    wire new_AGEMA_signal_6233 ;
    wire new_AGEMA_signal_6234 ;
    wire new_AGEMA_signal_6235 ;
    wire new_AGEMA_signal_6236 ;
    wire new_AGEMA_signal_6237 ;
    wire new_AGEMA_signal_6238 ;
    wire new_AGEMA_signal_6239 ;
    wire new_AGEMA_signal_6240 ;
    wire new_AGEMA_signal_6241 ;
    wire new_AGEMA_signal_6242 ;
    wire new_AGEMA_signal_6243 ;
    wire new_AGEMA_signal_6244 ;
    wire new_AGEMA_signal_6245 ;
    wire new_AGEMA_signal_6246 ;
    wire new_AGEMA_signal_6247 ;
    wire new_AGEMA_signal_6248 ;
    wire new_AGEMA_signal_6249 ;
    wire new_AGEMA_signal_6250 ;
    wire new_AGEMA_signal_6251 ;
    wire new_AGEMA_signal_6252 ;
    wire new_AGEMA_signal_6253 ;
    wire new_AGEMA_signal_6254 ;
    wire new_AGEMA_signal_6255 ;
    wire new_AGEMA_signal_6256 ;
    wire new_AGEMA_signal_6257 ;
    wire new_AGEMA_signal_6258 ;
    wire new_AGEMA_signal_6259 ;
    wire new_AGEMA_signal_6260 ;
    wire new_AGEMA_signal_6261 ;
    wire new_AGEMA_signal_6262 ;
    wire new_AGEMA_signal_6263 ;
    wire new_AGEMA_signal_6264 ;
    wire new_AGEMA_signal_6265 ;
    wire new_AGEMA_signal_6266 ;
    wire new_AGEMA_signal_6267 ;
    wire new_AGEMA_signal_6268 ;
    wire new_AGEMA_signal_6269 ;
    wire new_AGEMA_signal_6270 ;
    wire new_AGEMA_signal_6271 ;
    wire new_AGEMA_signal_6272 ;
    wire new_AGEMA_signal_6273 ;
    wire new_AGEMA_signal_6274 ;
    wire new_AGEMA_signal_6275 ;
    wire new_AGEMA_signal_6276 ;
    wire new_AGEMA_signal_6277 ;
    wire new_AGEMA_signal_6278 ;
    wire new_AGEMA_signal_6279 ;
    wire new_AGEMA_signal_6280 ;
    wire new_AGEMA_signal_6281 ;
    wire new_AGEMA_signal_6282 ;
    wire new_AGEMA_signal_6283 ;
    wire new_AGEMA_signal_6284 ;
    wire new_AGEMA_signal_6285 ;
    wire new_AGEMA_signal_6286 ;
    wire new_AGEMA_signal_6287 ;
    wire new_AGEMA_signal_6288 ;
    wire new_AGEMA_signal_6289 ;
    wire new_AGEMA_signal_6290 ;
    wire new_AGEMA_signal_6291 ;
    wire new_AGEMA_signal_6292 ;
    wire new_AGEMA_signal_6293 ;
    wire new_AGEMA_signal_6294 ;
    wire new_AGEMA_signal_6295 ;
    wire new_AGEMA_signal_6296 ;
    wire new_AGEMA_signal_6297 ;
    wire new_AGEMA_signal_6298 ;
    wire new_AGEMA_signal_6299 ;
    wire new_AGEMA_signal_6300 ;
    wire new_AGEMA_signal_6301 ;
    wire new_AGEMA_signal_6302 ;
    wire new_AGEMA_signal_6303 ;
    wire new_AGEMA_signal_6304 ;
    wire new_AGEMA_signal_6305 ;
    wire new_AGEMA_signal_6306 ;
    wire new_AGEMA_signal_6307 ;
    wire new_AGEMA_signal_6308 ;
    wire new_AGEMA_signal_6309 ;
    wire new_AGEMA_signal_6310 ;
    wire new_AGEMA_signal_6311 ;
    wire new_AGEMA_signal_6312 ;
    wire new_AGEMA_signal_6313 ;
    wire new_AGEMA_signal_6314 ;
    wire new_AGEMA_signal_6315 ;
    wire new_AGEMA_signal_6316 ;
    wire new_AGEMA_signal_6317 ;
    wire new_AGEMA_signal_6318 ;
    wire new_AGEMA_signal_6319 ;
    wire new_AGEMA_signal_6320 ;
    wire new_AGEMA_signal_6321 ;
    wire new_AGEMA_signal_6322 ;
    wire new_AGEMA_signal_6323 ;
    wire new_AGEMA_signal_6324 ;
    wire new_AGEMA_signal_6325 ;
    wire new_AGEMA_signal_6326 ;
    wire new_AGEMA_signal_6327 ;
    wire new_AGEMA_signal_6328 ;
    wire new_AGEMA_signal_6329 ;
    wire new_AGEMA_signal_6330 ;
    wire new_AGEMA_signal_6331 ;
    wire new_AGEMA_signal_6332 ;
    wire new_AGEMA_signal_6333 ;
    wire new_AGEMA_signal_6334 ;
    wire new_AGEMA_signal_6335 ;
    wire new_AGEMA_signal_6336 ;
    wire new_AGEMA_signal_6337 ;
    wire new_AGEMA_signal_6338 ;
    wire new_AGEMA_signal_6339 ;
    wire new_AGEMA_signal_6340 ;
    wire new_AGEMA_signal_6341 ;
    wire new_AGEMA_signal_6342 ;
    wire new_AGEMA_signal_6343 ;
    wire new_AGEMA_signal_6344 ;
    wire new_AGEMA_signal_6345 ;
    wire new_AGEMA_signal_6346 ;
    wire new_AGEMA_signal_6347 ;
    wire new_AGEMA_signal_6348 ;
    wire new_AGEMA_signal_6349 ;
    wire new_AGEMA_signal_6350 ;
    wire new_AGEMA_signal_6351 ;
    wire new_AGEMA_signal_6352 ;
    wire new_AGEMA_signal_6353 ;
    wire new_AGEMA_signal_6354 ;
    wire new_AGEMA_signal_6355 ;
    wire new_AGEMA_signal_6356 ;
    wire new_AGEMA_signal_6357 ;
    wire new_AGEMA_signal_6358 ;
    wire new_AGEMA_signal_6359 ;
    wire new_AGEMA_signal_6360 ;
    wire new_AGEMA_signal_6361 ;
    wire new_AGEMA_signal_6362 ;
    wire new_AGEMA_signal_6363 ;
    wire new_AGEMA_signal_6364 ;
    wire new_AGEMA_signal_6365 ;
    wire new_AGEMA_signal_6366 ;
    wire new_AGEMA_signal_6367 ;
    wire new_AGEMA_signal_6368 ;
    wire new_AGEMA_signal_6369 ;
    wire new_AGEMA_signal_6370 ;
    wire new_AGEMA_signal_6371 ;
    wire new_AGEMA_signal_6372 ;
    wire new_AGEMA_signal_6373 ;
    wire new_AGEMA_signal_6374 ;
    wire new_AGEMA_signal_6375 ;
    wire new_AGEMA_signal_6376 ;
    wire new_AGEMA_signal_6377 ;
    wire new_AGEMA_signal_6378 ;
    wire new_AGEMA_signal_6379 ;
    wire new_AGEMA_signal_6380 ;
    wire new_AGEMA_signal_6381 ;
    wire new_AGEMA_signal_6382 ;
    wire new_AGEMA_signal_6383 ;
    wire new_AGEMA_signal_6384 ;
    wire new_AGEMA_signal_6385 ;
    wire new_AGEMA_signal_6386 ;
    wire new_AGEMA_signal_6387 ;
    wire new_AGEMA_signal_6388 ;
    wire new_AGEMA_signal_6389 ;
    wire new_AGEMA_signal_6390 ;
    wire new_AGEMA_signal_6391 ;
    wire new_AGEMA_signal_6392 ;
    wire new_AGEMA_signal_6393 ;
    wire new_AGEMA_signal_6394 ;
    wire new_AGEMA_signal_6395 ;
    wire new_AGEMA_signal_6396 ;
    wire new_AGEMA_signal_6397 ;
    wire new_AGEMA_signal_6398 ;
    wire new_AGEMA_signal_6399 ;
    wire new_AGEMA_signal_6400 ;
    wire new_AGEMA_signal_6401 ;
    wire new_AGEMA_signal_6402 ;
    wire new_AGEMA_signal_6403 ;
    wire new_AGEMA_signal_6404 ;
    wire new_AGEMA_signal_6405 ;
    wire new_AGEMA_signal_6406 ;
    wire new_AGEMA_signal_6407 ;
    wire new_AGEMA_signal_6408 ;
    wire new_AGEMA_signal_6409 ;
    wire new_AGEMA_signal_6410 ;
    wire new_AGEMA_signal_6411 ;
    wire new_AGEMA_signal_6412 ;
    wire new_AGEMA_signal_6413 ;
    wire new_AGEMA_signal_6414 ;
    wire new_AGEMA_signal_6415 ;
    wire new_AGEMA_signal_6416 ;
    wire new_AGEMA_signal_6417 ;
    wire new_AGEMA_signal_6418 ;
    wire new_AGEMA_signal_6419 ;
    wire new_AGEMA_signal_6420 ;
    wire new_AGEMA_signal_6421 ;
    wire new_AGEMA_signal_6422 ;
    wire new_AGEMA_signal_6423 ;
    wire new_AGEMA_signal_6424 ;
    wire new_AGEMA_signal_6425 ;
    wire new_AGEMA_signal_6426 ;
    wire new_AGEMA_signal_6427 ;
    wire new_AGEMA_signal_6428 ;
    wire new_AGEMA_signal_6429 ;
    wire new_AGEMA_signal_6430 ;
    wire new_AGEMA_signal_6431 ;
    wire new_AGEMA_signal_6432 ;
    wire new_AGEMA_signal_6433 ;
    wire new_AGEMA_signal_6434 ;
    wire new_AGEMA_signal_6435 ;
    wire new_AGEMA_signal_6436 ;
    wire new_AGEMA_signal_6437 ;
    wire new_AGEMA_signal_6438 ;
    wire new_AGEMA_signal_6439 ;
    wire new_AGEMA_signal_6440 ;
    wire new_AGEMA_signal_6441 ;
    wire new_AGEMA_signal_6442 ;
    wire new_AGEMA_signal_6443 ;
    wire new_AGEMA_signal_6444 ;
    wire new_AGEMA_signal_6445 ;
    wire new_AGEMA_signal_6446 ;
    wire new_AGEMA_signal_6447 ;
    wire new_AGEMA_signal_6448 ;
    wire new_AGEMA_signal_6449 ;
    wire new_AGEMA_signal_6450 ;
    wire new_AGEMA_signal_6451 ;
    wire new_AGEMA_signal_6452 ;
    wire new_AGEMA_signal_6453 ;
    wire new_AGEMA_signal_6454 ;
    wire new_AGEMA_signal_6455 ;
    wire new_AGEMA_signal_6456 ;
    wire new_AGEMA_signal_6457 ;
    wire new_AGEMA_signal_6458 ;
    wire new_AGEMA_signal_6459 ;
    wire new_AGEMA_signal_6460 ;
    wire new_AGEMA_signal_6461 ;
    wire new_AGEMA_signal_6462 ;
    wire new_AGEMA_signal_6463 ;
    wire new_AGEMA_signal_6464 ;
    wire new_AGEMA_signal_6465 ;
    wire new_AGEMA_signal_6466 ;
    wire new_AGEMA_signal_6467 ;
    wire new_AGEMA_signal_6468 ;
    wire new_AGEMA_signal_6469 ;
    wire new_AGEMA_signal_6470 ;
    wire new_AGEMA_signal_6471 ;
    wire new_AGEMA_signal_6472 ;
    wire new_AGEMA_signal_6473 ;
    wire new_AGEMA_signal_6474 ;
    wire new_AGEMA_signal_6475 ;
    wire new_AGEMA_signal_6476 ;
    wire new_AGEMA_signal_6477 ;
    wire new_AGEMA_signal_6478 ;
    wire new_AGEMA_signal_6479 ;
    wire new_AGEMA_signal_6480 ;
    wire new_AGEMA_signal_6481 ;
    wire new_AGEMA_signal_6482 ;
    wire new_AGEMA_signal_6483 ;
    wire new_AGEMA_signal_6484 ;
    wire new_AGEMA_signal_6485 ;
    wire new_AGEMA_signal_6486 ;
    wire new_AGEMA_signal_6487 ;
    wire new_AGEMA_signal_6488 ;
    wire new_AGEMA_signal_6489 ;
    wire new_AGEMA_signal_6490 ;
    wire new_AGEMA_signal_6491 ;
    wire new_AGEMA_signal_6492 ;
    wire new_AGEMA_signal_6493 ;
    wire new_AGEMA_signal_6494 ;
    wire new_AGEMA_signal_6495 ;
    wire new_AGEMA_signal_6496 ;
    wire new_AGEMA_signal_6497 ;
    wire new_AGEMA_signal_6498 ;
    wire new_AGEMA_signal_6499 ;
    wire new_AGEMA_signal_6500 ;
    wire new_AGEMA_signal_6501 ;
    wire new_AGEMA_signal_6502 ;
    wire new_AGEMA_signal_6503 ;
    wire new_AGEMA_signal_6504 ;
    wire new_AGEMA_signal_6505 ;
    wire new_AGEMA_signal_6506 ;
    wire new_AGEMA_signal_6507 ;
    wire new_AGEMA_signal_6508 ;
    wire new_AGEMA_signal_6509 ;
    wire new_AGEMA_signal_6510 ;
    wire new_AGEMA_signal_6511 ;
    wire new_AGEMA_signal_6512 ;
    wire new_AGEMA_signal_6513 ;
    wire new_AGEMA_signal_6514 ;
    wire new_AGEMA_signal_6515 ;
    wire new_AGEMA_signal_6516 ;
    wire new_AGEMA_signal_6517 ;
    wire new_AGEMA_signal_6518 ;
    wire new_AGEMA_signal_6519 ;
    wire new_AGEMA_signal_6520 ;
    wire new_AGEMA_signal_6521 ;
    wire new_AGEMA_signal_6522 ;
    wire new_AGEMA_signal_6523 ;
    wire new_AGEMA_signal_6524 ;
    wire new_AGEMA_signal_6525 ;
    wire new_AGEMA_signal_6526 ;
    wire new_AGEMA_signal_6527 ;
    wire new_AGEMA_signal_6528 ;
    wire new_AGEMA_signal_6529 ;
    wire new_AGEMA_signal_6530 ;
    wire new_AGEMA_signal_6531 ;
    wire new_AGEMA_signal_6532 ;
    wire new_AGEMA_signal_6533 ;
    wire new_AGEMA_signal_6534 ;
    wire new_AGEMA_signal_6535 ;
    wire new_AGEMA_signal_6536 ;
    wire new_AGEMA_signal_6537 ;
    wire new_AGEMA_signal_6538 ;
    wire new_AGEMA_signal_6539 ;
    wire new_AGEMA_signal_6540 ;
    wire new_AGEMA_signal_6541 ;
    wire new_AGEMA_signal_6542 ;
    wire new_AGEMA_signal_6543 ;
    wire new_AGEMA_signal_6544 ;
    wire new_AGEMA_signal_6545 ;
    wire new_AGEMA_signal_6546 ;
    wire new_AGEMA_signal_6547 ;
    wire new_AGEMA_signal_6548 ;
    wire new_AGEMA_signal_6549 ;
    wire new_AGEMA_signal_6550 ;
    wire new_AGEMA_signal_6551 ;
    wire new_AGEMA_signal_6552 ;
    wire new_AGEMA_signal_6553 ;
    wire new_AGEMA_signal_6554 ;
    wire new_AGEMA_signal_6555 ;
    wire new_AGEMA_signal_6556 ;
    wire new_AGEMA_signal_6557 ;
    wire new_AGEMA_signal_6558 ;
    wire new_AGEMA_signal_6559 ;
    wire new_AGEMA_signal_6560 ;
    wire new_AGEMA_signal_6561 ;
    wire new_AGEMA_signal_6562 ;
    wire new_AGEMA_signal_6563 ;
    wire new_AGEMA_signal_6564 ;
    wire new_AGEMA_signal_6565 ;
    wire new_AGEMA_signal_6566 ;
    wire new_AGEMA_signal_6567 ;
    wire new_AGEMA_signal_6568 ;
    wire new_AGEMA_signal_6569 ;
    wire new_AGEMA_signal_6570 ;
    wire new_AGEMA_signal_6571 ;
    wire new_AGEMA_signal_6572 ;
    wire new_AGEMA_signal_6573 ;
    wire new_AGEMA_signal_6574 ;
    wire new_AGEMA_signal_6575 ;
    wire new_AGEMA_signal_6576 ;
    wire new_AGEMA_signal_6577 ;
    wire new_AGEMA_signal_6578 ;
    wire new_AGEMA_signal_6579 ;
    wire new_AGEMA_signal_6580 ;
    wire new_AGEMA_signal_6581 ;
    wire new_AGEMA_signal_6582 ;
    wire new_AGEMA_signal_6583 ;
    wire new_AGEMA_signal_6584 ;
    wire new_AGEMA_signal_6585 ;
    wire new_AGEMA_signal_6586 ;
    wire new_AGEMA_signal_6587 ;
    wire new_AGEMA_signal_6588 ;
    wire new_AGEMA_signal_6589 ;
    wire new_AGEMA_signal_6590 ;
    wire new_AGEMA_signal_6591 ;
    wire new_AGEMA_signal_6592 ;
    wire new_AGEMA_signal_6593 ;
    wire new_AGEMA_signal_6594 ;
    wire new_AGEMA_signal_6595 ;
    wire new_AGEMA_signal_6596 ;
    wire new_AGEMA_signal_6597 ;
    wire new_AGEMA_signal_6598 ;
    wire new_AGEMA_signal_6599 ;
    wire new_AGEMA_signal_6600 ;
    wire new_AGEMA_signal_6601 ;
    wire new_AGEMA_signal_6602 ;
    wire new_AGEMA_signal_6603 ;
    wire new_AGEMA_signal_6604 ;
    wire new_AGEMA_signal_6605 ;
    wire new_AGEMA_signal_6606 ;
    wire new_AGEMA_signal_6607 ;
    wire new_AGEMA_signal_6608 ;
    wire new_AGEMA_signal_6609 ;
    wire new_AGEMA_signal_6610 ;
    wire new_AGEMA_signal_6611 ;
    wire new_AGEMA_signal_6612 ;
    wire new_AGEMA_signal_6613 ;
    wire new_AGEMA_signal_6614 ;
    wire new_AGEMA_signal_6615 ;
    wire new_AGEMA_signal_6616 ;
    wire new_AGEMA_signal_6617 ;
    wire new_AGEMA_signal_6618 ;
    wire new_AGEMA_signal_6619 ;
    wire new_AGEMA_signal_6620 ;
    wire new_AGEMA_signal_6621 ;
    wire new_AGEMA_signal_6622 ;
    wire new_AGEMA_signal_6623 ;
    wire new_AGEMA_signal_6624 ;
    wire new_AGEMA_signal_6625 ;
    wire new_AGEMA_signal_6626 ;
    wire new_AGEMA_signal_6627 ;
    wire new_AGEMA_signal_6628 ;
    wire new_AGEMA_signal_6629 ;
    wire new_AGEMA_signal_6630 ;
    wire new_AGEMA_signal_6631 ;
    wire new_AGEMA_signal_6632 ;
    wire new_AGEMA_signal_6633 ;
    wire new_AGEMA_signal_6634 ;
    wire new_AGEMA_signal_6635 ;
    wire new_AGEMA_signal_6636 ;
    wire new_AGEMA_signal_6637 ;
    wire new_AGEMA_signal_6638 ;
    wire new_AGEMA_signal_6639 ;
    wire new_AGEMA_signal_6640 ;
    wire new_AGEMA_signal_6641 ;
    wire new_AGEMA_signal_6642 ;
    wire new_AGEMA_signal_6643 ;
    wire new_AGEMA_signal_6644 ;
    wire new_AGEMA_signal_6645 ;
    wire new_AGEMA_signal_6646 ;
    wire new_AGEMA_signal_6647 ;
    wire new_AGEMA_signal_6648 ;
    wire new_AGEMA_signal_6649 ;
    wire new_AGEMA_signal_6650 ;
    wire new_AGEMA_signal_6651 ;
    wire new_AGEMA_signal_6652 ;
    wire new_AGEMA_signal_6653 ;
    wire new_AGEMA_signal_6654 ;
    wire new_AGEMA_signal_6655 ;
    wire new_AGEMA_signal_6656 ;
    wire new_AGEMA_signal_6657 ;
    wire new_AGEMA_signal_6658 ;
    wire new_AGEMA_signal_6659 ;
    wire new_AGEMA_signal_6660 ;
    wire new_AGEMA_signal_6661 ;
    wire new_AGEMA_signal_6662 ;
    wire new_AGEMA_signal_6663 ;
    wire new_AGEMA_signal_6664 ;
    wire new_AGEMA_signal_6665 ;
    wire new_AGEMA_signal_6666 ;
    wire new_AGEMA_signal_6667 ;
    wire new_AGEMA_signal_6668 ;
    wire new_AGEMA_signal_6669 ;
    wire new_AGEMA_signal_6670 ;
    wire new_AGEMA_signal_6671 ;
    wire new_AGEMA_signal_6672 ;
    wire new_AGEMA_signal_6673 ;
    wire new_AGEMA_signal_6674 ;
    wire new_AGEMA_signal_6675 ;
    wire new_AGEMA_signal_6676 ;
    wire new_AGEMA_signal_6677 ;
    wire new_AGEMA_signal_6678 ;
    wire new_AGEMA_signal_6679 ;
    wire new_AGEMA_signal_6680 ;
    wire new_AGEMA_signal_6681 ;
    wire new_AGEMA_signal_6682 ;
    wire new_AGEMA_signal_6683 ;
    wire new_AGEMA_signal_6684 ;
    wire new_AGEMA_signal_6685 ;
    wire new_AGEMA_signal_6686 ;
    wire new_AGEMA_signal_6687 ;
    wire new_AGEMA_signal_6688 ;
    wire new_AGEMA_signal_6689 ;
    wire new_AGEMA_signal_6690 ;
    wire new_AGEMA_signal_6691 ;
    wire new_AGEMA_signal_6692 ;
    wire new_AGEMA_signal_6693 ;
    wire new_AGEMA_signal_6694 ;
    wire new_AGEMA_signal_6695 ;
    wire new_AGEMA_signal_6696 ;
    wire new_AGEMA_signal_6697 ;
    wire new_AGEMA_signal_6698 ;
    wire new_AGEMA_signal_6699 ;
    wire new_AGEMA_signal_6700 ;
    wire new_AGEMA_signal_6701 ;
    wire new_AGEMA_signal_6702 ;
    wire new_AGEMA_signal_6703 ;
    wire new_AGEMA_signal_6704 ;
    wire new_AGEMA_signal_6705 ;
    wire new_AGEMA_signal_6706 ;
    wire new_AGEMA_signal_6707 ;
    wire new_AGEMA_signal_6708 ;
    wire new_AGEMA_signal_6709 ;
    wire new_AGEMA_signal_6710 ;
    wire new_AGEMA_signal_6711 ;
    wire new_AGEMA_signal_6712 ;
    wire new_AGEMA_signal_6713 ;
    wire new_AGEMA_signal_6714 ;
    wire new_AGEMA_signal_6715 ;
    wire new_AGEMA_signal_6716 ;
    wire new_AGEMA_signal_6717 ;
    wire new_AGEMA_signal_6718 ;
    wire new_AGEMA_signal_6719 ;
    wire new_AGEMA_signal_6720 ;
    wire new_AGEMA_signal_6721 ;
    wire new_AGEMA_signal_6722 ;
    wire new_AGEMA_signal_6723 ;
    wire new_AGEMA_signal_6724 ;
    wire new_AGEMA_signal_6725 ;
    wire new_AGEMA_signal_6726 ;
    wire new_AGEMA_signal_6727 ;
    wire new_AGEMA_signal_6728 ;
    wire new_AGEMA_signal_6729 ;
    wire new_AGEMA_signal_6730 ;
    wire new_AGEMA_signal_6731 ;
    wire new_AGEMA_signal_6732 ;
    wire new_AGEMA_signal_6733 ;
    wire new_AGEMA_signal_6734 ;
    wire new_AGEMA_signal_6735 ;
    wire new_AGEMA_signal_6736 ;
    wire new_AGEMA_signal_6737 ;
    wire new_AGEMA_signal_6738 ;
    wire new_AGEMA_signal_6739 ;
    wire new_AGEMA_signal_6740 ;
    wire new_AGEMA_signal_6741 ;
    wire new_AGEMA_signal_6742 ;
    wire new_AGEMA_signal_6743 ;
    wire new_AGEMA_signal_6744 ;
    wire new_AGEMA_signal_6745 ;
    wire new_AGEMA_signal_6746 ;
    wire new_AGEMA_signal_6747 ;
    wire new_AGEMA_signal_6748 ;
    wire new_AGEMA_signal_6749 ;
    wire new_AGEMA_signal_6750 ;
    wire new_AGEMA_signal_6751 ;
    wire new_AGEMA_signal_6752 ;
    wire new_AGEMA_signal_6753 ;
    wire new_AGEMA_signal_6754 ;
    wire new_AGEMA_signal_6755 ;
    wire new_AGEMA_signal_6756 ;
    wire new_AGEMA_signal_6757 ;
    wire new_AGEMA_signal_6758 ;
    wire new_AGEMA_signal_6759 ;
    wire new_AGEMA_signal_6760 ;
    wire new_AGEMA_signal_6761 ;
    wire new_AGEMA_signal_6762 ;
    wire new_AGEMA_signal_6763 ;
    wire new_AGEMA_signal_6764 ;
    wire new_AGEMA_signal_6765 ;
    wire new_AGEMA_signal_6766 ;
    wire new_AGEMA_signal_6767 ;
    wire new_AGEMA_signal_6768 ;
    wire new_AGEMA_signal_6769 ;
    wire new_AGEMA_signal_6770 ;
    wire new_AGEMA_signal_6771 ;
    wire new_AGEMA_signal_6772 ;
    wire new_AGEMA_signal_6773 ;
    wire new_AGEMA_signal_6774 ;
    wire new_AGEMA_signal_6775 ;
    wire new_AGEMA_signal_6776 ;
    wire new_AGEMA_signal_6777 ;
    wire new_AGEMA_signal_6778 ;
    wire new_AGEMA_signal_6779 ;
    wire new_AGEMA_signal_6780 ;
    wire new_AGEMA_signal_6781 ;
    wire new_AGEMA_signal_6782 ;
    wire new_AGEMA_signal_6783 ;
    wire new_AGEMA_signal_6784 ;
    wire new_AGEMA_signal_6785 ;
    wire new_AGEMA_signal_6786 ;
    wire new_AGEMA_signal_6787 ;
    wire new_AGEMA_signal_6788 ;
    wire new_AGEMA_signal_6789 ;
    wire new_AGEMA_signal_6790 ;
    wire new_AGEMA_signal_6791 ;
    wire new_AGEMA_signal_6792 ;
    wire new_AGEMA_signal_6793 ;
    wire new_AGEMA_signal_6794 ;
    wire new_AGEMA_signal_6795 ;
    wire new_AGEMA_signal_6796 ;
    wire new_AGEMA_signal_6797 ;
    wire new_AGEMA_signal_6798 ;
    wire new_AGEMA_signal_6799 ;
    wire new_AGEMA_signal_6800 ;
    wire new_AGEMA_signal_6801 ;
    wire new_AGEMA_signal_6802 ;
    wire new_AGEMA_signal_6803 ;
    wire new_AGEMA_signal_6804 ;
    wire new_AGEMA_signal_6805 ;
    wire new_AGEMA_signal_6806 ;
    wire new_AGEMA_signal_6807 ;
    wire new_AGEMA_signal_6808 ;
    wire new_AGEMA_signal_6809 ;
    wire new_AGEMA_signal_6810 ;
    wire new_AGEMA_signal_6811 ;
    wire new_AGEMA_signal_6812 ;
    wire new_AGEMA_signal_6813 ;
    wire new_AGEMA_signal_6814 ;
    wire new_AGEMA_signal_6815 ;
    wire new_AGEMA_signal_6816 ;
    wire new_AGEMA_signal_6817 ;
    wire new_AGEMA_signal_6818 ;
    wire new_AGEMA_signal_6819 ;
    wire new_AGEMA_signal_6820 ;
    wire new_AGEMA_signal_6821 ;
    wire new_AGEMA_signal_6822 ;
    wire new_AGEMA_signal_6823 ;
    wire new_AGEMA_signal_6824 ;
    wire new_AGEMA_signal_6825 ;
    wire new_AGEMA_signal_6826 ;
    wire new_AGEMA_signal_6827 ;
    wire new_AGEMA_signal_6828 ;
    wire new_AGEMA_signal_6829 ;
    wire new_AGEMA_signal_6830 ;
    wire new_AGEMA_signal_6831 ;
    wire new_AGEMA_signal_6832 ;
    wire new_AGEMA_signal_6833 ;
    wire new_AGEMA_signal_6834 ;
    wire new_AGEMA_signal_6835 ;
    wire new_AGEMA_signal_6836 ;
    wire new_AGEMA_signal_6837 ;
    wire new_AGEMA_signal_6838 ;
    wire new_AGEMA_signal_6839 ;
    wire new_AGEMA_signal_6840 ;
    wire new_AGEMA_signal_6841 ;
    wire new_AGEMA_signal_6842 ;
    wire new_AGEMA_signal_6843 ;
    wire new_AGEMA_signal_6844 ;
    wire new_AGEMA_signal_6845 ;
    wire new_AGEMA_signal_6846 ;
    wire new_AGEMA_signal_6847 ;
    wire new_AGEMA_signal_6848 ;
    wire new_AGEMA_signal_6849 ;
    wire new_AGEMA_signal_6850 ;
    wire new_AGEMA_signal_6851 ;
    wire new_AGEMA_signal_6852 ;
    wire new_AGEMA_signal_6853 ;
    wire new_AGEMA_signal_6854 ;
    wire new_AGEMA_signal_6855 ;
    wire new_AGEMA_signal_6856 ;
    wire new_AGEMA_signal_6857 ;
    wire new_AGEMA_signal_6858 ;
    wire new_AGEMA_signal_6859 ;
    wire new_AGEMA_signal_6860 ;
    wire new_AGEMA_signal_6861 ;
    wire new_AGEMA_signal_6862 ;
    wire new_AGEMA_signal_6863 ;
    wire new_AGEMA_signal_6864 ;
    wire new_AGEMA_signal_6865 ;
    wire new_AGEMA_signal_6866 ;
    wire new_AGEMA_signal_6867 ;
    wire new_AGEMA_signal_6868 ;
    wire new_AGEMA_signal_6869 ;
    wire new_AGEMA_signal_6870 ;
    wire new_AGEMA_signal_6871 ;
    wire new_AGEMA_signal_6872 ;
    wire new_AGEMA_signal_6873 ;
    wire new_AGEMA_signal_6874 ;
    wire new_AGEMA_signal_6875 ;
    wire new_AGEMA_signal_6876 ;
    wire new_AGEMA_signal_6877 ;
    wire new_AGEMA_signal_6878 ;
    wire new_AGEMA_signal_6879 ;
    wire new_AGEMA_signal_6880 ;
    wire new_AGEMA_signal_6881 ;
    wire new_AGEMA_signal_6882 ;
    wire new_AGEMA_signal_6883 ;
    wire new_AGEMA_signal_6884 ;
    wire new_AGEMA_signal_6885 ;
    wire new_AGEMA_signal_6886 ;
    wire new_AGEMA_signal_6887 ;
    wire new_AGEMA_signal_6888 ;
    wire new_AGEMA_signal_6889 ;
    wire new_AGEMA_signal_6890 ;
    wire new_AGEMA_signal_6891 ;
    wire new_AGEMA_signal_6892 ;
    wire new_AGEMA_signal_6893 ;
    wire new_AGEMA_signal_6894 ;
    wire new_AGEMA_signal_6895 ;
    wire new_AGEMA_signal_6896 ;
    wire new_AGEMA_signal_6897 ;
    wire new_AGEMA_signal_6898 ;
    wire new_AGEMA_signal_6899 ;
    wire new_AGEMA_signal_6900 ;
    wire new_AGEMA_signal_6901 ;
    wire new_AGEMA_signal_6902 ;
    wire new_AGEMA_signal_6903 ;
    wire new_AGEMA_signal_6904 ;
    wire new_AGEMA_signal_6905 ;
    wire new_AGEMA_signal_6906 ;
    wire new_AGEMA_signal_6907 ;
    wire new_AGEMA_signal_6908 ;
    wire new_AGEMA_signal_6909 ;
    wire new_AGEMA_signal_6910 ;
    wire new_AGEMA_signal_6911 ;
    wire new_AGEMA_signal_6912 ;
    wire new_AGEMA_signal_6913 ;
    wire new_AGEMA_signal_6914 ;
    wire new_AGEMA_signal_6915 ;
    wire new_AGEMA_signal_6916 ;
    wire new_AGEMA_signal_6917 ;
    wire new_AGEMA_signal_6918 ;
    wire new_AGEMA_signal_6919 ;
    wire new_AGEMA_signal_6920 ;
    wire new_AGEMA_signal_6921 ;
    wire new_AGEMA_signal_6922 ;
    wire new_AGEMA_signal_6923 ;
    wire new_AGEMA_signal_6924 ;
    wire new_AGEMA_signal_6925 ;
    wire new_AGEMA_signal_6926 ;
    wire new_AGEMA_signal_6927 ;
    wire new_AGEMA_signal_6928 ;
    wire new_AGEMA_signal_6929 ;
    wire new_AGEMA_signal_6930 ;
    wire new_AGEMA_signal_6931 ;
    wire new_AGEMA_signal_6932 ;
    wire new_AGEMA_signal_6933 ;
    wire new_AGEMA_signal_6934 ;
    wire new_AGEMA_signal_6935 ;
    wire new_AGEMA_signal_6936 ;
    wire new_AGEMA_signal_6937 ;
    wire new_AGEMA_signal_6938 ;
    wire new_AGEMA_signal_6939 ;
    wire new_AGEMA_signal_6940 ;
    wire new_AGEMA_signal_6941 ;
    wire new_AGEMA_signal_6942 ;
    wire new_AGEMA_signal_6943 ;
    wire new_AGEMA_signal_6944 ;
    wire new_AGEMA_signal_6945 ;
    wire new_AGEMA_signal_6946 ;
    wire new_AGEMA_signal_6947 ;
    wire new_AGEMA_signal_6948 ;
    wire new_AGEMA_signal_6949 ;
    wire new_AGEMA_signal_6950 ;
    wire new_AGEMA_signal_6951 ;
    wire new_AGEMA_signal_6952 ;
    wire new_AGEMA_signal_6953 ;
    wire new_AGEMA_signal_6954 ;
    wire new_AGEMA_signal_6955 ;
    wire new_AGEMA_signal_6956 ;
    wire new_AGEMA_signal_6957 ;
    wire new_AGEMA_signal_6958 ;
    wire new_AGEMA_signal_6959 ;
    wire new_AGEMA_signal_6960 ;
    wire new_AGEMA_signal_6961 ;
    wire new_AGEMA_signal_6962 ;
    wire new_AGEMA_signal_6963 ;
    wire new_AGEMA_signal_6964 ;
    wire new_AGEMA_signal_6965 ;
    wire new_AGEMA_signal_6966 ;
    wire new_AGEMA_signal_6967 ;
    wire new_AGEMA_signal_6968 ;
    wire new_AGEMA_signal_6969 ;
    wire new_AGEMA_signal_6970 ;
    wire new_AGEMA_signal_6971 ;
    wire new_AGEMA_signal_6972 ;
    wire new_AGEMA_signal_6973 ;
    wire new_AGEMA_signal_6974 ;
    wire new_AGEMA_signal_6975 ;
    wire new_AGEMA_signal_6976 ;
    wire new_AGEMA_signal_6977 ;
    wire new_AGEMA_signal_6978 ;
    wire new_AGEMA_signal_6979 ;
    wire new_AGEMA_signal_6980 ;
    wire new_AGEMA_signal_6981 ;
    wire new_AGEMA_signal_6982 ;
    wire new_AGEMA_signal_6983 ;
    wire new_AGEMA_signal_6984 ;
    wire new_AGEMA_signal_6985 ;
    wire new_AGEMA_signal_6986 ;
    wire new_AGEMA_signal_6987 ;
    wire new_AGEMA_signal_6988 ;
    wire new_AGEMA_signal_6989 ;
    wire new_AGEMA_signal_6990 ;
    wire new_AGEMA_signal_6991 ;
    wire new_AGEMA_signal_6992 ;
    wire new_AGEMA_signal_6993 ;
    wire new_AGEMA_signal_6994 ;
    wire new_AGEMA_signal_6995 ;
    wire new_AGEMA_signal_6996 ;
    wire new_AGEMA_signal_6997 ;
    wire new_AGEMA_signal_6998 ;
    wire new_AGEMA_signal_6999 ;
    wire new_AGEMA_signal_7000 ;
    wire new_AGEMA_signal_7001 ;
    wire new_AGEMA_signal_7002 ;
    wire new_AGEMA_signal_7003 ;
    wire new_AGEMA_signal_7004 ;
    wire new_AGEMA_signal_7005 ;
    wire new_AGEMA_signal_7006 ;
    wire new_AGEMA_signal_7007 ;
    wire new_AGEMA_signal_7008 ;
    wire new_AGEMA_signal_7009 ;
    wire new_AGEMA_signal_7010 ;
    wire new_AGEMA_signal_7011 ;
    wire new_AGEMA_signal_7012 ;
    wire new_AGEMA_signal_7013 ;
    wire new_AGEMA_signal_7014 ;
    wire new_AGEMA_signal_7015 ;
    wire new_AGEMA_signal_7016 ;
    wire new_AGEMA_signal_7017 ;
    wire new_AGEMA_signal_7018 ;
    wire new_AGEMA_signal_7019 ;
    wire new_AGEMA_signal_7020 ;
    wire new_AGEMA_signal_7021 ;
    wire new_AGEMA_signal_7022 ;
    wire new_AGEMA_signal_7023 ;
    wire new_AGEMA_signal_7024 ;
    wire new_AGEMA_signal_7025 ;
    wire new_AGEMA_signal_7026 ;
    wire new_AGEMA_signal_7027 ;
    wire new_AGEMA_signal_7028 ;
    wire new_AGEMA_signal_7029 ;
    wire new_AGEMA_signal_7030 ;
    wire new_AGEMA_signal_7031 ;
    wire new_AGEMA_signal_7032 ;
    wire new_AGEMA_signal_7033 ;
    wire new_AGEMA_signal_7034 ;
    wire new_AGEMA_signal_7035 ;
    wire new_AGEMA_signal_7036 ;
    wire new_AGEMA_signal_7037 ;
    wire new_AGEMA_signal_7038 ;
    wire new_AGEMA_signal_7039 ;
    wire new_AGEMA_signal_7040 ;
    wire new_AGEMA_signal_7041 ;
    wire new_AGEMA_signal_7042 ;
    wire new_AGEMA_signal_7043 ;
    wire new_AGEMA_signal_7044 ;
    wire new_AGEMA_signal_7045 ;
    wire new_AGEMA_signal_7046 ;
    wire new_AGEMA_signal_7047 ;
    wire new_AGEMA_signal_7048 ;
    wire new_AGEMA_signal_7049 ;
    wire new_AGEMA_signal_7050 ;
    wire new_AGEMA_signal_7051 ;
    wire new_AGEMA_signal_7052 ;
    wire new_AGEMA_signal_7053 ;
    wire new_AGEMA_signal_7054 ;
    wire new_AGEMA_signal_7055 ;
    wire new_AGEMA_signal_7056 ;
    wire new_AGEMA_signal_7057 ;
    wire new_AGEMA_signal_7058 ;
    wire new_AGEMA_signal_7059 ;
    wire new_AGEMA_signal_7060 ;
    wire new_AGEMA_signal_7061 ;
    wire new_AGEMA_signal_7062 ;
    wire new_AGEMA_signal_7063 ;
    wire new_AGEMA_signal_7064 ;
    wire new_AGEMA_signal_7065 ;
    wire new_AGEMA_signal_7066 ;
    wire new_AGEMA_signal_7067 ;
    wire new_AGEMA_signal_7068 ;
    wire new_AGEMA_signal_7069 ;
    wire new_AGEMA_signal_7070 ;
    wire new_AGEMA_signal_7071 ;
    wire new_AGEMA_signal_7072 ;
    wire new_AGEMA_signal_7073 ;
    wire new_AGEMA_signal_7074 ;
    wire new_AGEMA_signal_7075 ;
    wire new_AGEMA_signal_7076 ;
    wire new_AGEMA_signal_7077 ;
    wire new_AGEMA_signal_7078 ;
    wire new_AGEMA_signal_7079 ;
    wire new_AGEMA_signal_7080 ;
    wire new_AGEMA_signal_7081 ;
    wire new_AGEMA_signal_7082 ;
    wire new_AGEMA_signal_7083 ;
    wire new_AGEMA_signal_7084 ;
    wire new_AGEMA_signal_7085 ;
    wire new_AGEMA_signal_7086 ;
    wire new_AGEMA_signal_7087 ;
    wire new_AGEMA_signal_7088 ;
    wire new_AGEMA_signal_7089 ;
    wire new_AGEMA_signal_7090 ;
    wire new_AGEMA_signal_7091 ;
    wire new_AGEMA_signal_7092 ;
    wire new_AGEMA_signal_7093 ;
    wire new_AGEMA_signal_7094 ;
    wire new_AGEMA_signal_7095 ;
    wire new_AGEMA_signal_7096 ;
    wire new_AGEMA_signal_7097 ;
    wire new_AGEMA_signal_7098 ;
    wire new_AGEMA_signal_7099 ;
    wire new_AGEMA_signal_7100 ;
    wire new_AGEMA_signal_7101 ;
    wire new_AGEMA_signal_7102 ;
    wire new_AGEMA_signal_7103 ;
    wire new_AGEMA_signal_7104 ;
    wire new_AGEMA_signal_7105 ;
    wire new_AGEMA_signal_7106 ;
    wire new_AGEMA_signal_7107 ;
    wire new_AGEMA_signal_7108 ;
    wire new_AGEMA_signal_7109 ;
    wire new_AGEMA_signal_7110 ;
    wire new_AGEMA_signal_7111 ;
    wire new_AGEMA_signal_7112 ;
    wire new_AGEMA_signal_7113 ;
    wire new_AGEMA_signal_7114 ;
    wire new_AGEMA_signal_7115 ;
    wire new_AGEMA_signal_7116 ;
    wire new_AGEMA_signal_7117 ;
    wire new_AGEMA_signal_7118 ;
    wire new_AGEMA_signal_7119 ;
    wire new_AGEMA_signal_7120 ;
    wire new_AGEMA_signal_7121 ;
    wire new_AGEMA_signal_7122 ;
    wire new_AGEMA_signal_7123 ;
    wire new_AGEMA_signal_7124 ;
    wire new_AGEMA_signal_7125 ;
    wire new_AGEMA_signal_7126 ;
    wire new_AGEMA_signal_7127 ;
    wire new_AGEMA_signal_7128 ;
    wire new_AGEMA_signal_7129 ;
    wire new_AGEMA_signal_7130 ;
    wire new_AGEMA_signal_7131 ;
    wire new_AGEMA_signal_7132 ;
    wire new_AGEMA_signal_7133 ;
    wire new_AGEMA_signal_7134 ;
    wire new_AGEMA_signal_7135 ;
    wire new_AGEMA_signal_7136 ;
    wire new_AGEMA_signal_7137 ;
    wire new_AGEMA_signal_7138 ;
    wire new_AGEMA_signal_7139 ;
    wire new_AGEMA_signal_7140 ;
    wire new_AGEMA_signal_7141 ;
    wire new_AGEMA_signal_7142 ;
    wire new_AGEMA_signal_7143 ;
    wire new_AGEMA_signal_7144 ;
    wire new_AGEMA_signal_7145 ;
    wire new_AGEMA_signal_7146 ;
    wire new_AGEMA_signal_7147 ;
    wire new_AGEMA_signal_7148 ;
    wire new_AGEMA_signal_7149 ;
    wire new_AGEMA_signal_7150 ;
    wire new_AGEMA_signal_7151 ;
    wire new_AGEMA_signal_7152 ;
    wire new_AGEMA_signal_7153 ;
    wire new_AGEMA_signal_7154 ;
    wire new_AGEMA_signal_7155 ;
    wire new_AGEMA_signal_7156 ;
    wire new_AGEMA_signal_7157 ;
    wire new_AGEMA_signal_7158 ;
    wire new_AGEMA_signal_7159 ;
    wire new_AGEMA_signal_7160 ;
    wire new_AGEMA_signal_7161 ;
    wire new_AGEMA_signal_7162 ;
    wire new_AGEMA_signal_7163 ;
    wire new_AGEMA_signal_7164 ;
    wire new_AGEMA_signal_7165 ;
    wire new_AGEMA_signal_7166 ;
    wire new_AGEMA_signal_7167 ;
    wire new_AGEMA_signal_7168 ;
    wire new_AGEMA_signal_7169 ;
    wire new_AGEMA_signal_7170 ;
    wire new_AGEMA_signal_7171 ;
    wire new_AGEMA_signal_7172 ;
    wire new_AGEMA_signal_7173 ;
    wire new_AGEMA_signal_7174 ;
    wire new_AGEMA_signal_7175 ;
    wire new_AGEMA_signal_7176 ;
    wire new_AGEMA_signal_7177 ;
    wire new_AGEMA_signal_7178 ;
    wire new_AGEMA_signal_7179 ;
    wire new_AGEMA_signal_7180 ;
    wire new_AGEMA_signal_7181 ;
    wire new_AGEMA_signal_7182 ;
    wire new_AGEMA_signal_7183 ;
    wire new_AGEMA_signal_7184 ;
    wire new_AGEMA_signal_7185 ;
    wire new_AGEMA_signal_7186 ;
    wire new_AGEMA_signal_7187 ;
    wire new_AGEMA_signal_7188 ;
    wire new_AGEMA_signal_7189 ;
    wire new_AGEMA_signal_7190 ;
    wire new_AGEMA_signal_7191 ;
    wire new_AGEMA_signal_7192 ;
    wire new_AGEMA_signal_7193 ;
    wire new_AGEMA_signal_7194 ;
    wire new_AGEMA_signal_7195 ;
    wire new_AGEMA_signal_7196 ;
    wire new_AGEMA_signal_7197 ;
    wire new_AGEMA_signal_7198 ;
    wire new_AGEMA_signal_7199 ;
    wire new_AGEMA_signal_7200 ;
    wire new_AGEMA_signal_7201 ;
    wire new_AGEMA_signal_7202 ;
    wire new_AGEMA_signal_7203 ;
    wire new_AGEMA_signal_7204 ;
    wire new_AGEMA_signal_7205 ;
    wire new_AGEMA_signal_7206 ;
    wire new_AGEMA_signal_7207 ;
    wire new_AGEMA_signal_7208 ;
    wire new_AGEMA_signal_7209 ;
    wire new_AGEMA_signal_7210 ;
    wire new_AGEMA_signal_7211 ;
    wire new_AGEMA_signal_7212 ;
    wire new_AGEMA_signal_7213 ;
    wire new_AGEMA_signal_7214 ;
    wire new_AGEMA_signal_7215 ;
    wire new_AGEMA_signal_7216 ;
    wire new_AGEMA_signal_7217 ;
    wire new_AGEMA_signal_7218 ;
    wire new_AGEMA_signal_7219 ;
    wire new_AGEMA_signal_7220 ;
    wire new_AGEMA_signal_7221 ;
    wire new_AGEMA_signal_7222 ;
    wire new_AGEMA_signal_7223 ;
    wire new_AGEMA_signal_7224 ;
    wire new_AGEMA_signal_7225 ;
    wire new_AGEMA_signal_7226 ;
    wire new_AGEMA_signal_7227 ;
    wire new_AGEMA_signal_7228 ;
    wire new_AGEMA_signal_7229 ;
    wire new_AGEMA_signal_7230 ;
    wire new_AGEMA_signal_7231 ;
    wire new_AGEMA_signal_7232 ;
    wire new_AGEMA_signal_7233 ;
    wire new_AGEMA_signal_7234 ;
    wire new_AGEMA_signal_7235 ;
    wire new_AGEMA_signal_7236 ;
    wire new_AGEMA_signal_7237 ;
    wire new_AGEMA_signal_7238 ;
    wire new_AGEMA_signal_7239 ;
    wire new_AGEMA_signal_7240 ;
    wire new_AGEMA_signal_7241 ;
    wire new_AGEMA_signal_7242 ;
    wire new_AGEMA_signal_7243 ;
    wire new_AGEMA_signal_7244 ;
    wire new_AGEMA_signal_7245 ;
    wire new_AGEMA_signal_7246 ;
    wire new_AGEMA_signal_7247 ;
    wire new_AGEMA_signal_7248 ;
    wire new_AGEMA_signal_7249 ;
    wire new_AGEMA_signal_7250 ;
    wire new_AGEMA_signal_7251 ;
    wire new_AGEMA_signal_7252 ;
    wire new_AGEMA_signal_7253 ;
    wire new_AGEMA_signal_7254 ;
    wire new_AGEMA_signal_7255 ;
    wire new_AGEMA_signal_7256 ;
    wire new_AGEMA_signal_7257 ;
    wire new_AGEMA_signal_7258 ;
    wire new_AGEMA_signal_7259 ;
    wire new_AGEMA_signal_7260 ;
    wire new_AGEMA_signal_7261 ;
    wire new_AGEMA_signal_7262 ;
    wire new_AGEMA_signal_7263 ;
    wire new_AGEMA_signal_7264 ;
    wire new_AGEMA_signal_7265 ;
    wire new_AGEMA_signal_7266 ;
    wire new_AGEMA_signal_7267 ;
    wire new_AGEMA_signal_7268 ;
    wire new_AGEMA_signal_7269 ;
    wire new_AGEMA_signal_7270 ;
    wire new_AGEMA_signal_7271 ;
    wire new_AGEMA_signal_7272 ;
    wire new_AGEMA_signal_7273 ;
    wire new_AGEMA_signal_7274 ;
    wire new_AGEMA_signal_7275 ;
    wire new_AGEMA_signal_7276 ;
    wire new_AGEMA_signal_7277 ;
    wire new_AGEMA_signal_7278 ;
    wire new_AGEMA_signal_7279 ;
    wire new_AGEMA_signal_7280 ;
    wire new_AGEMA_signal_7281 ;
    wire new_AGEMA_signal_7282 ;
    wire new_AGEMA_signal_7283 ;
    wire new_AGEMA_signal_7284 ;
    wire new_AGEMA_signal_7285 ;
    wire new_AGEMA_signal_7286 ;
    wire new_AGEMA_signal_7287 ;
    wire new_AGEMA_signal_7288 ;
    wire new_AGEMA_signal_7289 ;
    wire new_AGEMA_signal_7290 ;
    wire new_AGEMA_signal_7291 ;
    wire new_AGEMA_signal_7292 ;
    wire new_AGEMA_signal_7293 ;
    wire new_AGEMA_signal_7294 ;
    wire new_AGEMA_signal_7295 ;
    wire new_AGEMA_signal_7296 ;
    wire new_AGEMA_signal_7297 ;
    wire new_AGEMA_signal_7298 ;
    wire new_AGEMA_signal_7299 ;
    wire new_AGEMA_signal_7300 ;
    wire new_AGEMA_signal_7301 ;
    wire new_AGEMA_signal_7302 ;
    wire new_AGEMA_signal_7303 ;
    wire new_AGEMA_signal_7304 ;
    wire new_AGEMA_signal_7305 ;
    wire new_AGEMA_signal_7306 ;
    wire new_AGEMA_signal_7307 ;
    wire new_AGEMA_signal_7308 ;
    wire new_AGEMA_signal_7309 ;
    wire new_AGEMA_signal_7310 ;
    wire new_AGEMA_signal_7311 ;
    wire new_AGEMA_signal_7312 ;
    wire new_AGEMA_signal_7313 ;
    wire new_AGEMA_signal_7314 ;
    wire new_AGEMA_signal_7315 ;
    wire new_AGEMA_signal_7316 ;
    wire new_AGEMA_signal_7317 ;
    wire new_AGEMA_signal_7318 ;
    wire new_AGEMA_signal_7319 ;
    wire new_AGEMA_signal_7320 ;
    wire new_AGEMA_signal_7321 ;
    wire new_AGEMA_signal_7322 ;
    wire new_AGEMA_signal_7323 ;
    wire new_AGEMA_signal_7324 ;
    wire new_AGEMA_signal_7325 ;
    wire new_AGEMA_signal_7326 ;
    wire new_AGEMA_signal_7327 ;
    wire new_AGEMA_signal_7328 ;
    wire new_AGEMA_signal_7329 ;
    wire new_AGEMA_signal_7330 ;
    wire new_AGEMA_signal_7331 ;
    wire new_AGEMA_signal_7332 ;
    wire new_AGEMA_signal_7333 ;
    wire new_AGEMA_signal_7334 ;
    wire new_AGEMA_signal_7335 ;
    wire new_AGEMA_signal_7336 ;
    wire new_AGEMA_signal_7337 ;
    wire new_AGEMA_signal_7338 ;
    wire new_AGEMA_signal_7339 ;
    wire new_AGEMA_signal_7340 ;
    wire new_AGEMA_signal_7341 ;
    wire new_AGEMA_signal_7342 ;
    wire new_AGEMA_signal_7343 ;
    wire new_AGEMA_signal_7344 ;
    wire new_AGEMA_signal_7345 ;
    wire new_AGEMA_signal_7346 ;
    wire new_AGEMA_signal_7347 ;
    wire new_AGEMA_signal_7348 ;
    wire new_AGEMA_signal_7349 ;
    wire new_AGEMA_signal_7350 ;
    wire new_AGEMA_signal_7351 ;
    wire new_AGEMA_signal_7352 ;
    wire new_AGEMA_signal_7353 ;
    wire new_AGEMA_signal_7354 ;
    wire new_AGEMA_signal_7355 ;
    wire new_AGEMA_signal_7356 ;
    wire new_AGEMA_signal_7357 ;
    wire new_AGEMA_signal_7358 ;
    wire new_AGEMA_signal_7359 ;
    wire new_AGEMA_signal_7360 ;
    wire new_AGEMA_signal_7361 ;
    wire new_AGEMA_signal_7362 ;
    wire new_AGEMA_signal_7363 ;
    wire new_AGEMA_signal_7364 ;
    wire new_AGEMA_signal_7365 ;
    wire new_AGEMA_signal_7366 ;
    wire new_AGEMA_signal_7367 ;
    wire new_AGEMA_signal_7368 ;
    wire new_AGEMA_signal_7369 ;
    wire new_AGEMA_signal_7370 ;
    wire new_AGEMA_signal_7371 ;
    wire new_AGEMA_signal_7372 ;
    wire new_AGEMA_signal_7373 ;
    wire new_AGEMA_signal_7374 ;
    wire new_AGEMA_signal_7375 ;
    wire new_AGEMA_signal_7376 ;
    wire new_AGEMA_signal_7377 ;
    wire new_AGEMA_signal_7378 ;
    wire new_AGEMA_signal_7379 ;
    wire new_AGEMA_signal_7380 ;
    wire new_AGEMA_signal_7381 ;
    wire new_AGEMA_signal_7382 ;
    wire new_AGEMA_signal_7383 ;
    wire new_AGEMA_signal_7384 ;
    wire new_AGEMA_signal_7385 ;
    wire new_AGEMA_signal_7386 ;
    wire new_AGEMA_signal_7387 ;
    wire new_AGEMA_signal_7388 ;
    wire new_AGEMA_signal_7389 ;
    wire new_AGEMA_signal_7390 ;
    wire new_AGEMA_signal_7391 ;
    wire new_AGEMA_signal_7392 ;
    wire new_AGEMA_signal_7393 ;
    wire new_AGEMA_signal_7394 ;
    wire new_AGEMA_signal_7395 ;
    wire new_AGEMA_signal_7396 ;
    wire new_AGEMA_signal_7397 ;
    wire new_AGEMA_signal_7398 ;
    wire new_AGEMA_signal_7399 ;
    wire new_AGEMA_signal_7400 ;
    wire new_AGEMA_signal_7401 ;
    wire new_AGEMA_signal_7402 ;
    wire new_AGEMA_signal_7403 ;
    wire new_AGEMA_signal_7404 ;
    wire new_AGEMA_signal_7405 ;
    wire new_AGEMA_signal_7406 ;
    wire new_AGEMA_signal_7407 ;
    wire new_AGEMA_signal_7408 ;
    wire new_AGEMA_signal_7409 ;
    wire new_AGEMA_signal_7410 ;
    wire new_AGEMA_signal_7411 ;
    wire new_AGEMA_signal_7412 ;
    wire new_AGEMA_signal_7413 ;
    wire new_AGEMA_signal_7414 ;
    wire new_AGEMA_signal_7415 ;
    wire new_AGEMA_signal_7416 ;
    wire new_AGEMA_signal_7417 ;
    wire new_AGEMA_signal_7418 ;
    wire new_AGEMA_signal_7419 ;
    wire new_AGEMA_signal_7420 ;
    wire new_AGEMA_signal_7421 ;
    wire new_AGEMA_signal_7422 ;
    wire new_AGEMA_signal_7423 ;
    wire new_AGEMA_signal_7424 ;
    wire new_AGEMA_signal_7425 ;
    wire new_AGEMA_signal_7426 ;
    wire new_AGEMA_signal_7427 ;
    wire new_AGEMA_signal_7428 ;
    wire new_AGEMA_signal_7429 ;
    wire new_AGEMA_signal_7430 ;
    wire new_AGEMA_signal_7431 ;
    wire new_AGEMA_signal_7432 ;
    wire new_AGEMA_signal_7433 ;
    wire new_AGEMA_signal_7434 ;
    wire new_AGEMA_signal_7435 ;
    wire new_AGEMA_signal_7436 ;
    wire new_AGEMA_signal_7437 ;
    wire new_AGEMA_signal_7438 ;
    wire new_AGEMA_signal_7439 ;
    wire new_AGEMA_signal_7440 ;
    wire new_AGEMA_signal_7441 ;
    wire new_AGEMA_signal_7442 ;
    wire new_AGEMA_signal_7443 ;
    wire new_AGEMA_signal_7444 ;
    wire new_AGEMA_signal_7445 ;
    wire new_AGEMA_signal_7446 ;
    wire new_AGEMA_signal_7447 ;
    wire new_AGEMA_signal_7448 ;
    wire new_AGEMA_signal_7449 ;
    wire new_AGEMA_signal_7450 ;
    wire new_AGEMA_signal_7451 ;
    wire new_AGEMA_signal_7452 ;
    wire new_AGEMA_signal_7453 ;
    wire new_AGEMA_signal_7454 ;
    wire new_AGEMA_signal_7455 ;
    wire new_AGEMA_signal_7456 ;
    wire new_AGEMA_signal_7457 ;
    wire new_AGEMA_signal_7458 ;
    wire new_AGEMA_signal_7459 ;
    wire new_AGEMA_signal_7460 ;
    wire new_AGEMA_signal_7461 ;
    wire new_AGEMA_signal_7462 ;
    wire new_AGEMA_signal_7463 ;
    wire new_AGEMA_signal_7464 ;
    wire new_AGEMA_signal_7465 ;
    wire new_AGEMA_signal_7466 ;
    wire new_AGEMA_signal_7467 ;
    wire new_AGEMA_signal_7468 ;
    wire new_AGEMA_signal_7469 ;
    wire new_AGEMA_signal_7470 ;
    wire new_AGEMA_signal_7471 ;
    wire new_AGEMA_signal_7472 ;
    wire new_AGEMA_signal_7473 ;
    wire new_AGEMA_signal_7474 ;
    wire new_AGEMA_signal_7475 ;
    wire new_AGEMA_signal_7476 ;
    wire new_AGEMA_signal_7477 ;
    wire new_AGEMA_signal_7478 ;
    wire new_AGEMA_signal_7479 ;
    wire new_AGEMA_signal_7480 ;
    wire new_AGEMA_signal_7481 ;
    wire new_AGEMA_signal_7482 ;
    wire new_AGEMA_signal_7483 ;
    wire new_AGEMA_signal_7484 ;
    wire new_AGEMA_signal_7485 ;
    wire new_AGEMA_signal_7486 ;
    wire new_AGEMA_signal_7487 ;
    wire new_AGEMA_signal_7488 ;
    wire new_AGEMA_signal_7489 ;
    wire new_AGEMA_signal_7490 ;
    wire new_AGEMA_signal_7491 ;
    wire new_AGEMA_signal_7492 ;
    wire new_AGEMA_signal_7493 ;
    wire new_AGEMA_signal_7494 ;
    wire new_AGEMA_signal_7495 ;
    wire new_AGEMA_signal_7496 ;
    wire new_AGEMA_signal_7498 ;
    wire new_AGEMA_signal_7500 ;
    wire new_AGEMA_signal_7502 ;
    wire new_AGEMA_signal_7503 ;
    wire new_AGEMA_signal_7504 ;
    wire new_AGEMA_signal_7505 ;
    wire new_AGEMA_signal_7506 ;
    wire new_AGEMA_signal_7507 ;
    wire new_AGEMA_signal_7508 ;
    wire new_AGEMA_signal_7509 ;
    wire new_AGEMA_signal_7510 ;
    wire new_AGEMA_signal_7511 ;
    wire new_AGEMA_signal_7512 ;
    wire new_AGEMA_signal_7513 ;
    wire new_AGEMA_signal_7514 ;
    wire new_AGEMA_signal_7515 ;
    wire new_AGEMA_signal_7516 ;
    wire new_AGEMA_signal_7517 ;
    wire new_AGEMA_signal_7518 ;
    wire new_AGEMA_signal_7519 ;
    wire new_AGEMA_signal_7520 ;
    wire new_AGEMA_signal_7521 ;
    wire new_AGEMA_signal_7522 ;
    wire new_AGEMA_signal_7523 ;
    wire new_AGEMA_signal_7524 ;
    wire new_AGEMA_signal_7525 ;
    wire new_AGEMA_signal_7526 ;
    wire new_AGEMA_signal_7527 ;
    wire new_AGEMA_signal_7528 ;
    wire new_AGEMA_signal_7529 ;
    wire new_AGEMA_signal_7530 ;
    wire new_AGEMA_signal_7531 ;
    wire new_AGEMA_signal_7532 ;
    wire new_AGEMA_signal_7533 ;
    wire new_AGEMA_signal_7534 ;
    wire new_AGEMA_signal_7535 ;
    wire new_AGEMA_signal_7536 ;
    wire new_AGEMA_signal_7537 ;
    wire new_AGEMA_signal_7538 ;
    wire new_AGEMA_signal_7539 ;
    wire new_AGEMA_signal_7540 ;
    wire new_AGEMA_signal_7541 ;
    wire new_AGEMA_signal_7542 ;
    wire new_AGEMA_signal_7543 ;
    wire new_AGEMA_signal_7544 ;
    wire new_AGEMA_signal_7545 ;
    wire new_AGEMA_signal_7546 ;
    wire new_AGEMA_signal_7547 ;
    wire new_AGEMA_signal_7548 ;
    wire new_AGEMA_signal_7549 ;
    wire new_AGEMA_signal_7550 ;
    wire new_AGEMA_signal_7551 ;
    wire new_AGEMA_signal_7552 ;
    wire new_AGEMA_signal_7553 ;
    wire new_AGEMA_signal_7554 ;
    wire new_AGEMA_signal_7555 ;
    wire new_AGEMA_signal_7556 ;
    wire new_AGEMA_signal_7557 ;
    wire new_AGEMA_signal_7558 ;
    wire new_AGEMA_signal_7559 ;
    wire new_AGEMA_signal_7560 ;
    wire new_AGEMA_signal_7561 ;
    wire new_AGEMA_signal_7562 ;
    wire new_AGEMA_signal_7563 ;
    wire new_AGEMA_signal_7564 ;
    wire new_AGEMA_signal_7565 ;
    wire new_AGEMA_signal_7566 ;
    wire new_AGEMA_signal_7567 ;
    wire new_AGEMA_signal_7568 ;
    wire new_AGEMA_signal_7569 ;
    wire new_AGEMA_signal_7570 ;
    wire new_AGEMA_signal_7571 ;
    wire new_AGEMA_signal_7572 ;
    wire new_AGEMA_signal_7573 ;
    wire new_AGEMA_signal_7574 ;
    wire new_AGEMA_signal_7575 ;
    wire new_AGEMA_signal_7576 ;
    wire new_AGEMA_signal_7577 ;
    wire new_AGEMA_signal_7578 ;
    wire new_AGEMA_signal_7579 ;
    wire new_AGEMA_signal_7580 ;
    wire new_AGEMA_signal_7581 ;
    wire new_AGEMA_signal_7582 ;
    wire new_AGEMA_signal_7583 ;
    wire new_AGEMA_signal_7584 ;
    wire new_AGEMA_signal_7585 ;
    wire new_AGEMA_signal_7586 ;
    wire new_AGEMA_signal_7587 ;
    wire new_AGEMA_signal_7588 ;
    wire new_AGEMA_signal_7589 ;
    wire new_AGEMA_signal_7590 ;
    wire new_AGEMA_signal_7591 ;
    wire new_AGEMA_signal_7592 ;
    wire new_AGEMA_signal_7593 ;
    wire new_AGEMA_signal_7594 ;
    wire new_AGEMA_signal_7595 ;
    wire new_AGEMA_signal_7596 ;
    wire new_AGEMA_signal_7597 ;
    wire new_AGEMA_signal_7598 ;
    wire new_AGEMA_signal_7599 ;
    wire new_AGEMA_signal_7600 ;
    wire new_AGEMA_signal_7601 ;
    wire new_AGEMA_signal_7602 ;
    wire new_AGEMA_signal_7603 ;
    wire new_AGEMA_signal_7604 ;
    wire new_AGEMA_signal_7605 ;
    wire new_AGEMA_signal_7606 ;
    wire new_AGEMA_signal_7607 ;
    wire new_AGEMA_signal_7608 ;
    wire new_AGEMA_signal_7609 ;
    wire new_AGEMA_signal_7610 ;
    wire new_AGEMA_signal_7611 ;
    wire new_AGEMA_signal_7612 ;
    wire new_AGEMA_signal_7613 ;
    wire new_AGEMA_signal_7614 ;
    wire new_AGEMA_signal_7615 ;
    wire new_AGEMA_signal_7616 ;
    wire new_AGEMA_signal_7617 ;
    wire new_AGEMA_signal_7618 ;
    wire new_AGEMA_signal_7619 ;
    wire new_AGEMA_signal_7620 ;
    wire new_AGEMA_signal_7621 ;
    wire new_AGEMA_signal_7622 ;
    wire new_AGEMA_signal_7623 ;
    wire new_AGEMA_signal_7624 ;
    wire new_AGEMA_signal_7625 ;
    wire new_AGEMA_signal_7626 ;
    wire new_AGEMA_signal_7627 ;
    wire new_AGEMA_signal_7628 ;
    wire new_AGEMA_signal_7629 ;
    wire new_AGEMA_signal_7630 ;
    wire new_AGEMA_signal_7631 ;
    wire new_AGEMA_signal_7632 ;
    wire new_AGEMA_signal_7633 ;
    wire new_AGEMA_signal_7634 ;
    wire new_AGEMA_signal_7635 ;
    wire new_AGEMA_signal_7636 ;
    wire new_AGEMA_signal_7637 ;
    wire new_AGEMA_signal_7638 ;
    wire new_AGEMA_signal_7639 ;
    wire new_AGEMA_signal_7640 ;
    wire new_AGEMA_signal_7641 ;
    wire new_AGEMA_signal_7642 ;
    wire new_AGEMA_signal_7643 ;
    wire new_AGEMA_signal_7644 ;
    wire new_AGEMA_signal_7645 ;
    wire new_AGEMA_signal_7646 ;
    wire new_AGEMA_signal_7647 ;
    wire new_AGEMA_signal_7648 ;
    wire new_AGEMA_signal_7649 ;
    wire new_AGEMA_signal_7650 ;
    wire new_AGEMA_signal_7651 ;
    wire new_AGEMA_signal_7652 ;
    wire new_AGEMA_signal_7653 ;
    wire new_AGEMA_signal_7654 ;
    wire new_AGEMA_signal_7655 ;
    wire new_AGEMA_signal_7656 ;
    wire new_AGEMA_signal_7657 ;
    wire new_AGEMA_signal_7658 ;
    wire new_AGEMA_signal_7659 ;
    wire new_AGEMA_signal_7660 ;
    wire new_AGEMA_signal_7661 ;
    wire new_AGEMA_signal_7662 ;
    wire new_AGEMA_signal_7664 ;
    wire new_AGEMA_signal_7666 ;
    wire new_AGEMA_signal_7668 ;
    wire new_AGEMA_signal_7670 ;
    wire new_AGEMA_signal_7672 ;
    wire new_AGEMA_signal_7674 ;
    wire new_AGEMA_signal_7676 ;
    wire new_AGEMA_signal_7678 ;
    wire new_AGEMA_signal_7680 ;
    wire new_AGEMA_signal_7682 ;
    wire new_AGEMA_signal_7684 ;
    wire new_AGEMA_signal_7686 ;
    wire new_AGEMA_signal_7688 ;
    wire new_AGEMA_signal_7690 ;
    wire new_AGEMA_signal_7692 ;
    wire new_AGEMA_signal_7694 ;
    wire new_AGEMA_signal_7696 ;
    wire new_AGEMA_signal_7698 ;
    wire new_AGEMA_signal_7700 ;
    wire new_AGEMA_signal_7702 ;
    wire new_AGEMA_signal_7704 ;
    wire new_AGEMA_signal_7706 ;
    wire new_AGEMA_signal_7708 ;
    wire new_AGEMA_signal_7710 ;
    wire new_AGEMA_signal_7712 ;
    wire new_AGEMA_signal_7713 ;
    wire new_AGEMA_signal_7714 ;
    wire new_AGEMA_signal_7715 ;
    wire new_AGEMA_signal_7716 ;
    wire new_AGEMA_signal_7717 ;
    wire new_AGEMA_signal_7718 ;
    wire new_AGEMA_signal_7719 ;
    wire new_AGEMA_signal_7720 ;
    wire new_AGEMA_signal_7721 ;
    wire new_AGEMA_signal_7722 ;
    wire new_AGEMA_signal_7723 ;
    wire new_AGEMA_signal_7724 ;
    wire new_AGEMA_signal_7725 ;
    wire new_AGEMA_signal_7726 ;
    wire new_AGEMA_signal_7727 ;
    wire new_AGEMA_signal_7728 ;
    wire new_AGEMA_signal_7729 ;
    wire new_AGEMA_signal_7730 ;
    wire new_AGEMA_signal_7731 ;
    wire new_AGEMA_signal_7732 ;
    wire new_AGEMA_signal_7733 ;
    wire new_AGEMA_signal_7734 ;
    wire new_AGEMA_signal_7735 ;
    wire new_AGEMA_signal_7736 ;
    wire new_AGEMA_signal_7737 ;
    wire new_AGEMA_signal_7738 ;
    wire new_AGEMA_signal_7739 ;
    wire new_AGEMA_signal_7740 ;
    wire new_AGEMA_signal_7741 ;
    wire new_AGEMA_signal_7742 ;
    wire new_AGEMA_signal_7743 ;
    wire new_AGEMA_signal_7744 ;
    wire new_AGEMA_signal_7745 ;
    wire new_AGEMA_signal_7746 ;
    wire new_AGEMA_signal_7747 ;
    wire new_AGEMA_signal_7748 ;
    wire new_AGEMA_signal_7749 ;
    wire new_AGEMA_signal_7750 ;
    wire new_AGEMA_signal_7751 ;
    wire new_AGEMA_signal_7752 ;
    wire new_AGEMA_signal_7753 ;
    wire new_AGEMA_signal_7754 ;
    wire new_AGEMA_signal_7755 ;
    wire new_AGEMA_signal_7756 ;
    wire new_AGEMA_signal_7757 ;
    wire new_AGEMA_signal_7758 ;
    wire new_AGEMA_signal_7759 ;
    wire new_AGEMA_signal_7760 ;
    wire new_AGEMA_signal_7761 ;
    wire new_AGEMA_signal_7762 ;
    wire new_AGEMA_signal_7763 ;
    wire new_AGEMA_signal_7764 ;
    wire new_AGEMA_signal_7765 ;
    wire new_AGEMA_signal_7766 ;
    wire new_AGEMA_signal_7767 ;
    wire new_AGEMA_signal_7768 ;
    wire new_AGEMA_signal_7769 ;
    wire new_AGEMA_signal_7770 ;
    wire new_AGEMA_signal_7771 ;
    wire new_AGEMA_signal_7772 ;
    wire new_AGEMA_signal_7773 ;
    wire new_AGEMA_signal_7774 ;
    wire new_AGEMA_signal_7775 ;
    wire new_AGEMA_signal_7776 ;
    wire new_AGEMA_signal_7777 ;
    wire new_AGEMA_signal_7778 ;
    wire new_AGEMA_signal_7779 ;
    wire new_AGEMA_signal_7780 ;
    wire new_AGEMA_signal_7781 ;
    wire new_AGEMA_signal_7782 ;
    wire new_AGEMA_signal_7783 ;
    wire new_AGEMA_signal_7784 ;
    wire new_AGEMA_signal_7785 ;
    wire new_AGEMA_signal_7786 ;
    wire new_AGEMA_signal_7787 ;
    wire new_AGEMA_signal_7788 ;
    wire new_AGEMA_signal_7789 ;
    wire new_AGEMA_signal_7790 ;
    wire new_AGEMA_signal_7791 ;
    wire new_AGEMA_signal_7792 ;
    wire new_AGEMA_signal_7793 ;
    wire new_AGEMA_signal_7794 ;
    wire new_AGEMA_signal_7795 ;
    wire new_AGEMA_signal_7796 ;
    wire new_AGEMA_signal_7797 ;
    wire new_AGEMA_signal_7798 ;
    wire new_AGEMA_signal_7799 ;
    wire new_AGEMA_signal_7800 ;
    wire new_AGEMA_signal_7801 ;
    wire new_AGEMA_signal_7802 ;
    wire new_AGEMA_signal_7803 ;
    wire new_AGEMA_signal_7804 ;
    wire new_AGEMA_signal_7805 ;
    wire new_AGEMA_signal_7806 ;
    wire new_AGEMA_signal_7807 ;
    wire new_AGEMA_signal_7808 ;
    wire new_AGEMA_signal_7809 ;
    wire new_AGEMA_signal_7810 ;
    wire new_AGEMA_signal_7811 ;
    wire new_AGEMA_signal_7812 ;
    wire new_AGEMA_signal_7813 ;
    wire new_AGEMA_signal_7814 ;
    wire new_AGEMA_signal_7815 ;
    wire new_AGEMA_signal_7816 ;
    wire new_AGEMA_signal_7817 ;
    wire new_AGEMA_signal_7818 ;
    wire new_AGEMA_signal_7819 ;
    wire new_AGEMA_signal_7820 ;
    wire new_AGEMA_signal_7821 ;
    wire new_AGEMA_signal_7822 ;
    wire new_AGEMA_signal_7823 ;
    wire new_AGEMA_signal_7824 ;
    wire new_AGEMA_signal_7825 ;
    wire new_AGEMA_signal_7826 ;
    wire new_AGEMA_signal_7827 ;
    wire new_AGEMA_signal_7828 ;
    wire new_AGEMA_signal_7829 ;
    wire new_AGEMA_signal_7830 ;
    wire new_AGEMA_signal_7831 ;
    wire new_AGEMA_signal_7832 ;
    wire new_AGEMA_signal_7833 ;
    wire new_AGEMA_signal_7834 ;
    wire new_AGEMA_signal_7835 ;
    wire new_AGEMA_signal_7836 ;
    wire new_AGEMA_signal_7837 ;
    wire new_AGEMA_signal_7838 ;
    wire new_AGEMA_signal_7839 ;
    wire new_AGEMA_signal_7840 ;
    wire new_AGEMA_signal_7841 ;
    wire new_AGEMA_signal_7842 ;
    wire new_AGEMA_signal_7843 ;
    wire new_AGEMA_signal_7844 ;
    wire new_AGEMA_signal_7845 ;
    wire new_AGEMA_signal_7846 ;
    wire new_AGEMA_signal_7847 ;
    wire new_AGEMA_signal_7848 ;
    wire new_AGEMA_signal_7849 ;
    wire new_AGEMA_signal_7850 ;
    wire new_AGEMA_signal_7851 ;
    wire new_AGEMA_signal_7852 ;
    wire new_AGEMA_signal_7853 ;
    wire new_AGEMA_signal_7854 ;
    wire new_AGEMA_signal_7855 ;
    wire new_AGEMA_signal_7856 ;
    wire new_AGEMA_signal_7857 ;
    wire new_AGEMA_signal_7858 ;
    wire new_AGEMA_signal_7859 ;
    wire new_AGEMA_signal_7860 ;
    wire new_AGEMA_signal_7861 ;
    wire new_AGEMA_signal_7862 ;
    wire new_AGEMA_signal_7863 ;
    wire new_AGEMA_signal_7864 ;
    wire new_AGEMA_signal_7865 ;
    wire new_AGEMA_signal_7866 ;
    wire new_AGEMA_signal_7867 ;
    wire new_AGEMA_signal_7868 ;
    wire new_AGEMA_signal_7869 ;
    wire new_AGEMA_signal_7870 ;
    wire new_AGEMA_signal_7871 ;
    wire new_AGEMA_signal_7872 ;
    wire new_AGEMA_signal_7874 ;
    wire new_AGEMA_signal_7876 ;
    wire new_AGEMA_signal_7878 ;
    wire new_AGEMA_signal_7880 ;
    wire new_AGEMA_signal_7882 ;
    wire new_AGEMA_signal_7884 ;
    wire new_AGEMA_signal_7886 ;
    wire new_AGEMA_signal_7888 ;
    wire new_AGEMA_signal_7890 ;
    wire new_AGEMA_signal_7892 ;
    wire new_AGEMA_signal_7894 ;
    wire new_AGEMA_signal_7896 ;
    wire new_AGEMA_signal_7898 ;
    wire new_AGEMA_signal_7900 ;
    wire new_AGEMA_signal_7902 ;
    wire new_AGEMA_signal_7904 ;
    wire new_AGEMA_signal_7906 ;
    wire new_AGEMA_signal_7908 ;
    wire new_AGEMA_signal_7910 ;
    wire new_AGEMA_signal_7912 ;
    wire new_AGEMA_signal_7914 ;
    wire new_AGEMA_signal_7916 ;
    wire new_AGEMA_signal_7918 ;
    wire new_AGEMA_signal_7920 ;
    wire new_AGEMA_signal_7922 ;
    wire new_AGEMA_signal_7924 ;
    wire new_AGEMA_signal_7926 ;
    wire new_AGEMA_signal_7928 ;
    wire new_AGEMA_signal_7930 ;
    wire new_AGEMA_signal_7932 ;
    wire new_AGEMA_signal_7934 ;
    wire new_AGEMA_signal_7936 ;
    wire new_AGEMA_signal_7937 ;
    wire new_AGEMA_signal_7938 ;
    wire new_AGEMA_signal_7939 ;
    wire new_AGEMA_signal_7940 ;
    wire new_AGEMA_signal_7941 ;
    wire new_AGEMA_signal_7942 ;
    wire new_AGEMA_signal_7943 ;
    wire new_AGEMA_signal_7944 ;
    wire new_AGEMA_signal_7945 ;
    wire new_AGEMA_signal_7946 ;
    wire new_AGEMA_signal_7947 ;
    wire new_AGEMA_signal_7948 ;
    wire new_AGEMA_signal_7949 ;
    wire new_AGEMA_signal_7950 ;
    wire new_AGEMA_signal_7951 ;
    wire new_AGEMA_signal_7952 ;
    wire new_AGEMA_signal_7953 ;
    wire new_AGEMA_signal_7954 ;
    wire new_AGEMA_signal_7955 ;
    wire new_AGEMA_signal_7956 ;
    wire new_AGEMA_signal_7957 ;
    wire new_AGEMA_signal_7958 ;
    wire new_AGEMA_signal_7959 ;
    wire new_AGEMA_signal_7960 ;
    wire new_AGEMA_signal_7961 ;
    wire new_AGEMA_signal_7962 ;
    wire new_AGEMA_signal_7963 ;
    wire new_AGEMA_signal_7964 ;
    wire new_AGEMA_signal_7965 ;
    wire new_AGEMA_signal_7966 ;
    wire new_AGEMA_signal_7967 ;
    wire new_AGEMA_signal_7968 ;
    wire new_AGEMA_signal_7969 ;
    wire new_AGEMA_signal_7970 ;
    wire new_AGEMA_signal_7971 ;
    wire new_AGEMA_signal_7972 ;
    wire new_AGEMA_signal_7973 ;
    wire new_AGEMA_signal_7974 ;
    wire new_AGEMA_signal_7975 ;
    wire new_AGEMA_signal_7976 ;
    wire new_AGEMA_signal_7977 ;
    wire new_AGEMA_signal_7978 ;
    wire new_AGEMA_signal_7979 ;
    wire new_AGEMA_signal_7980 ;
    wire new_AGEMA_signal_7981 ;
    wire new_AGEMA_signal_7982 ;
    wire new_AGEMA_signal_7983 ;
    wire new_AGEMA_signal_7984 ;
    wire new_AGEMA_signal_7985 ;
    wire new_AGEMA_signal_7986 ;
    wire new_AGEMA_signal_7987 ;
    wire new_AGEMA_signal_7988 ;
    wire new_AGEMA_signal_7989 ;
    wire new_AGEMA_signal_7990 ;
    wire new_AGEMA_signal_7991 ;
    wire new_AGEMA_signal_7992 ;
    wire new_AGEMA_signal_7993 ;
    wire new_AGEMA_signal_7994 ;
    wire new_AGEMA_signal_7995 ;
    wire new_AGEMA_signal_7996 ;
    wire new_AGEMA_signal_7997 ;
    wire new_AGEMA_signal_7998 ;
    wire new_AGEMA_signal_7999 ;
    wire new_AGEMA_signal_8000 ;
    wire new_AGEMA_signal_8001 ;
    wire new_AGEMA_signal_8002 ;
    wire new_AGEMA_signal_8003 ;
    wire new_AGEMA_signal_8004 ;
    wire new_AGEMA_signal_8005 ;
    wire new_AGEMA_signal_8006 ;
    wire new_AGEMA_signal_8007 ;
    wire new_AGEMA_signal_8008 ;
    wire new_AGEMA_signal_8009 ;
    wire new_AGEMA_signal_8010 ;
    wire new_AGEMA_signal_8011 ;
    wire new_AGEMA_signal_8012 ;
    wire new_AGEMA_signal_8013 ;
    wire new_AGEMA_signal_8014 ;
    wire new_AGEMA_signal_8015 ;
    wire new_AGEMA_signal_8016 ;
    wire new_AGEMA_signal_8017 ;
    wire new_AGEMA_signal_8018 ;
    wire new_AGEMA_signal_8019 ;
    wire new_AGEMA_signal_8020 ;
    wire new_AGEMA_signal_8021 ;
    wire new_AGEMA_signal_8022 ;
    wire new_AGEMA_signal_8023 ;
    wire new_AGEMA_signal_8024 ;
    wire new_AGEMA_signal_8025 ;
    wire new_AGEMA_signal_8026 ;
    wire new_AGEMA_signal_8027 ;
    wire new_AGEMA_signal_8028 ;
    wire new_AGEMA_signal_8029 ;
    wire new_AGEMA_signal_8030 ;
    wire new_AGEMA_signal_8031 ;
    wire new_AGEMA_signal_8032 ;
    wire new_AGEMA_signal_8033 ;
    wire new_AGEMA_signal_8034 ;
    wire new_AGEMA_signal_8035 ;
    wire new_AGEMA_signal_8036 ;
    wire new_AGEMA_signal_8037 ;
    wire new_AGEMA_signal_8038 ;
    wire new_AGEMA_signal_8039 ;
    wire new_AGEMA_signal_8040 ;
    wire new_AGEMA_signal_8041 ;
    wire new_AGEMA_signal_8042 ;
    wire new_AGEMA_signal_8043 ;
    wire new_AGEMA_signal_8044 ;
    wire new_AGEMA_signal_8045 ;
    wire new_AGEMA_signal_8046 ;
    wire new_AGEMA_signal_8047 ;
    wire new_AGEMA_signal_8048 ;
    wire new_AGEMA_signal_8049 ;
    wire new_AGEMA_signal_8050 ;
    wire new_AGEMA_signal_8051 ;
    wire new_AGEMA_signal_8052 ;
    wire new_AGEMA_signal_8053 ;
    wire new_AGEMA_signal_8054 ;
    wire new_AGEMA_signal_8055 ;
    wire new_AGEMA_signal_8056 ;
    wire new_AGEMA_signal_8057 ;
    wire new_AGEMA_signal_8058 ;
    wire new_AGEMA_signal_8059 ;
    wire new_AGEMA_signal_8060 ;
    wire new_AGEMA_signal_8061 ;
    wire new_AGEMA_signal_8062 ;
    wire new_AGEMA_signal_8063 ;
    wire new_AGEMA_signal_8064 ;
    wire new_AGEMA_signal_8065 ;
    wire new_AGEMA_signal_8066 ;
    wire new_AGEMA_signal_8067 ;
    wire new_AGEMA_signal_8068 ;
    wire new_AGEMA_signal_8069 ;
    wire new_AGEMA_signal_8070 ;
    wire new_AGEMA_signal_8071 ;
    wire new_AGEMA_signal_8072 ;
    wire new_AGEMA_signal_8073 ;
    wire new_AGEMA_signal_8074 ;
    wire new_AGEMA_signal_8075 ;
    wire new_AGEMA_signal_8076 ;
    wire new_AGEMA_signal_8077 ;
    wire new_AGEMA_signal_8078 ;
    wire new_AGEMA_signal_8079 ;
    wire new_AGEMA_signal_8080 ;
    wire new_AGEMA_signal_8081 ;
    wire new_AGEMA_signal_8082 ;
    wire new_AGEMA_signal_8083 ;
    wire new_AGEMA_signal_8084 ;
    wire new_AGEMA_signal_8085 ;
    wire new_AGEMA_signal_8086 ;
    wire new_AGEMA_signal_8087 ;
    wire new_AGEMA_signal_8088 ;
    wire new_AGEMA_signal_8089 ;
    wire new_AGEMA_signal_8090 ;
    wire new_AGEMA_signal_8091 ;
    wire new_AGEMA_signal_8092 ;
    wire new_AGEMA_signal_8093 ;
    wire new_AGEMA_signal_8094 ;
    wire new_AGEMA_signal_8095 ;
    wire new_AGEMA_signal_8096 ;
    wire new_AGEMA_signal_8098 ;
    wire new_AGEMA_signal_8100 ;
    wire new_AGEMA_signal_8102 ;
    wire new_AGEMA_signal_8104 ;
    wire new_AGEMA_signal_8106 ;
    wire new_AGEMA_signal_8108 ;
    wire new_AGEMA_signal_8110 ;
    wire new_AGEMA_signal_8112 ;
    wire new_AGEMA_signal_8114 ;
    wire new_AGEMA_signal_8116 ;
    wire new_AGEMA_signal_8118 ;
    wire new_AGEMA_signal_8120 ;
    wire new_AGEMA_signal_8122 ;
    wire new_AGEMA_signal_8124 ;
    wire new_AGEMA_signal_8126 ;
    wire new_AGEMA_signal_8128 ;
    wire new_AGEMA_signal_8130 ;
    wire new_AGEMA_signal_8132 ;
    wire new_AGEMA_signal_8134 ;
    wire new_AGEMA_signal_8136 ;
    wire new_AGEMA_signal_8138 ;
    wire new_AGEMA_signal_8140 ;
    wire new_AGEMA_signal_8142 ;
    wire new_AGEMA_signal_8144 ;
    wire new_AGEMA_signal_8146 ;
    wire new_AGEMA_signal_8148 ;
    wire new_AGEMA_signal_8150 ;
    wire new_AGEMA_signal_8152 ;
    wire new_AGEMA_signal_8154 ;
    wire new_AGEMA_signal_8156 ;
    wire new_AGEMA_signal_8158 ;
    wire new_AGEMA_signal_8160 ;
    wire new_AGEMA_signal_8161 ;
    wire new_AGEMA_signal_8162 ;
    wire new_AGEMA_signal_8163 ;
    wire new_AGEMA_signal_8164 ;
    wire new_AGEMA_signal_8165 ;
    wire new_AGEMA_signal_8166 ;
    wire new_AGEMA_signal_8167 ;
    wire new_AGEMA_signal_8168 ;
    wire new_AGEMA_signal_8169 ;
    wire new_AGEMA_signal_8170 ;
    wire new_AGEMA_signal_8171 ;
    wire new_AGEMA_signal_8172 ;
    wire new_AGEMA_signal_8173 ;
    wire new_AGEMA_signal_8174 ;
    wire new_AGEMA_signal_8175 ;
    wire new_AGEMA_signal_8176 ;
    wire new_AGEMA_signal_8177 ;
    wire new_AGEMA_signal_8178 ;
    wire new_AGEMA_signal_8179 ;
    wire new_AGEMA_signal_8180 ;
    wire new_AGEMA_signal_8181 ;
    wire new_AGEMA_signal_8182 ;
    wire new_AGEMA_signal_8183 ;
    wire new_AGEMA_signal_8184 ;
    wire new_AGEMA_signal_8185 ;
    wire new_AGEMA_signal_8186 ;
    wire new_AGEMA_signal_8187 ;
    wire new_AGEMA_signal_8188 ;
    wire new_AGEMA_signal_8189 ;
    wire new_AGEMA_signal_8190 ;
    wire new_AGEMA_signal_8191 ;
    wire new_AGEMA_signal_8192 ;
    wire new_AGEMA_signal_8193 ;
    wire new_AGEMA_signal_8194 ;
    wire new_AGEMA_signal_8195 ;
    wire new_AGEMA_signal_8196 ;
    wire new_AGEMA_signal_8197 ;
    wire new_AGEMA_signal_8198 ;
    wire new_AGEMA_signal_8199 ;
    wire new_AGEMA_signal_8200 ;
    wire new_AGEMA_signal_8201 ;
    wire new_AGEMA_signal_8202 ;
    wire new_AGEMA_signal_8203 ;
    wire new_AGEMA_signal_8204 ;
    wire new_AGEMA_signal_8205 ;
    wire new_AGEMA_signal_8206 ;
    wire new_AGEMA_signal_8207 ;
    wire new_AGEMA_signal_8208 ;
    wire new_AGEMA_signal_8209 ;
    wire new_AGEMA_signal_8210 ;
    wire new_AGEMA_signal_8211 ;
    wire new_AGEMA_signal_8212 ;
    wire new_AGEMA_signal_8213 ;
    wire new_AGEMA_signal_8214 ;
    wire new_AGEMA_signal_8215 ;
    wire new_AGEMA_signal_8216 ;
    wire new_AGEMA_signal_8217 ;
    wire new_AGEMA_signal_8218 ;
    wire new_AGEMA_signal_8219 ;
    wire new_AGEMA_signal_8220 ;
    wire new_AGEMA_signal_8221 ;
    wire new_AGEMA_signal_8222 ;
    wire new_AGEMA_signal_8223 ;
    wire new_AGEMA_signal_8224 ;
    wire new_AGEMA_signal_8225 ;
    wire new_AGEMA_signal_8226 ;
    wire new_AGEMA_signal_8227 ;
    wire new_AGEMA_signal_8228 ;
    wire new_AGEMA_signal_8229 ;
    wire new_AGEMA_signal_8230 ;
    wire new_AGEMA_signal_8231 ;
    wire new_AGEMA_signal_8232 ;
    wire new_AGEMA_signal_8233 ;
    wire new_AGEMA_signal_8234 ;
    wire new_AGEMA_signal_8235 ;
    wire new_AGEMA_signal_8236 ;
    wire new_AGEMA_signal_8237 ;
    wire new_AGEMA_signal_8238 ;
    wire new_AGEMA_signal_8239 ;
    wire new_AGEMA_signal_8240 ;
    wire new_AGEMA_signal_8241 ;
    wire new_AGEMA_signal_8242 ;
    wire new_AGEMA_signal_8243 ;
    wire new_AGEMA_signal_8244 ;
    wire new_AGEMA_signal_8245 ;
    wire new_AGEMA_signal_8246 ;
    wire new_AGEMA_signal_8247 ;
    wire new_AGEMA_signal_8248 ;
    wire new_AGEMA_signal_8249 ;
    wire new_AGEMA_signal_8250 ;
    wire new_AGEMA_signal_8251 ;
    wire new_AGEMA_signal_8252 ;
    wire new_AGEMA_signal_8253 ;
    wire new_AGEMA_signal_8254 ;
    wire new_AGEMA_signal_8255 ;
    wire new_AGEMA_signal_8256 ;
    wire new_AGEMA_signal_8257 ;
    wire new_AGEMA_signal_8258 ;
    wire new_AGEMA_signal_8259 ;
    wire new_AGEMA_signal_8260 ;
    wire new_AGEMA_signal_8261 ;
    wire new_AGEMA_signal_8262 ;
    wire new_AGEMA_signal_8263 ;
    wire new_AGEMA_signal_8264 ;
    wire new_AGEMA_signal_8265 ;
    wire new_AGEMA_signal_8266 ;
    wire new_AGEMA_signal_8267 ;
    wire new_AGEMA_signal_8268 ;
    wire new_AGEMA_signal_8269 ;
    wire new_AGEMA_signal_8270 ;
    wire new_AGEMA_signal_8271 ;
    wire new_AGEMA_signal_8272 ;
    wire new_AGEMA_signal_8273 ;
    wire new_AGEMA_signal_8274 ;
    wire new_AGEMA_signal_8275 ;
    wire new_AGEMA_signal_8276 ;
    wire new_AGEMA_signal_8277 ;
    wire new_AGEMA_signal_8278 ;
    wire new_AGEMA_signal_8279 ;
    wire new_AGEMA_signal_8280 ;
    wire new_AGEMA_signal_8281 ;
    wire new_AGEMA_signal_8282 ;
    wire new_AGEMA_signal_8283 ;
    wire new_AGEMA_signal_8284 ;
    wire new_AGEMA_signal_8285 ;
    wire new_AGEMA_signal_8286 ;
    wire new_AGEMA_signal_8287 ;
    wire new_AGEMA_signal_8288 ;
    wire new_AGEMA_signal_8289 ;
    wire new_AGEMA_signal_8290 ;
    wire new_AGEMA_signal_8291 ;
    wire new_AGEMA_signal_8292 ;
    wire new_AGEMA_signal_8293 ;
    wire new_AGEMA_signal_8294 ;
    wire new_AGEMA_signal_8295 ;
    wire new_AGEMA_signal_8296 ;
    wire new_AGEMA_signal_8297 ;
    wire new_AGEMA_signal_8298 ;
    wire new_AGEMA_signal_8299 ;
    wire new_AGEMA_signal_8300 ;
    wire new_AGEMA_signal_8301 ;
    wire new_AGEMA_signal_8302 ;
    wire new_AGEMA_signal_8303 ;
    wire new_AGEMA_signal_8304 ;
    wire new_AGEMA_signal_8305 ;
    wire new_AGEMA_signal_8306 ;
    wire new_AGEMA_signal_8307 ;
    wire new_AGEMA_signal_8308 ;
    wire new_AGEMA_signal_8309 ;
    wire new_AGEMA_signal_8310 ;
    wire new_AGEMA_signal_8311 ;
    wire new_AGEMA_signal_8312 ;
    wire new_AGEMA_signal_8313 ;
    wire new_AGEMA_signal_8314 ;
    wire new_AGEMA_signal_8315 ;
    wire new_AGEMA_signal_8316 ;
    wire new_AGEMA_signal_8317 ;
    wire new_AGEMA_signal_8319 ;
    wire new_AGEMA_signal_8321 ;
    wire new_AGEMA_signal_8323 ;
    wire new_AGEMA_signal_8325 ;
    wire new_AGEMA_signal_8327 ;
    wire new_AGEMA_signal_8329 ;
    wire new_AGEMA_signal_8331 ;
    wire new_AGEMA_signal_8333 ;
    wire new_AGEMA_signal_8335 ;
    wire new_AGEMA_signal_8337 ;
    wire new_AGEMA_signal_8339 ;
    wire new_AGEMA_signal_8341 ;
    wire new_AGEMA_signal_8343 ;
    wire new_AGEMA_signal_8345 ;
    wire new_AGEMA_signal_8347 ;
    wire new_AGEMA_signal_8349 ;
    wire new_AGEMA_signal_8351 ;
    wire new_AGEMA_signal_8353 ;
    wire new_AGEMA_signal_8355 ;
    wire new_AGEMA_signal_8357 ;
    wire new_AGEMA_signal_8359 ;
    wire new_AGEMA_signal_8361 ;
    wire new_AGEMA_signal_8363 ;
    wire new_AGEMA_signal_8365 ;
    wire new_AGEMA_signal_8367 ;
    wire new_AGEMA_signal_8369 ;
    wire new_AGEMA_signal_8371 ;
    wire new_AGEMA_signal_8373 ;
    wire new_AGEMA_signal_8375 ;
    wire new_AGEMA_signal_8376 ;
    wire new_AGEMA_signal_8377 ;
    wire new_AGEMA_signal_8378 ;
    wire new_AGEMA_signal_8379 ;
    wire new_AGEMA_signal_8380 ;
    wire new_AGEMA_signal_8381 ;
    wire new_AGEMA_signal_8382 ;
    wire new_AGEMA_signal_8383 ;
    wire new_AGEMA_signal_8384 ;
    wire new_AGEMA_signal_8385 ;
    wire new_AGEMA_signal_8386 ;
    wire new_AGEMA_signal_8387 ;
    wire new_AGEMA_signal_8388 ;
    wire new_AGEMA_signal_8389 ;
    wire new_AGEMA_signal_8390 ;
    wire new_AGEMA_signal_8391 ;
    wire new_AGEMA_signal_8392 ;
    wire new_AGEMA_signal_8393 ;
    wire new_AGEMA_signal_8394 ;
    wire new_AGEMA_signal_8395 ;
    wire new_AGEMA_signal_8396 ;
    wire new_AGEMA_signal_8397 ;
    wire new_AGEMA_signal_8398 ;
    wire new_AGEMA_signal_8399 ;
    wire new_AGEMA_signal_8400 ;
    wire new_AGEMA_signal_8401 ;
    wire new_AGEMA_signal_8402 ;
    wire new_AGEMA_signal_8403 ;
    wire new_AGEMA_signal_8404 ;
    wire new_AGEMA_signal_8405 ;
    wire new_AGEMA_signal_8406 ;
    wire new_AGEMA_signal_8407 ;
    wire new_AGEMA_signal_8408 ;
    wire new_AGEMA_signal_8409 ;
    wire new_AGEMA_signal_8410 ;
    wire new_AGEMA_signal_8411 ;
    wire new_AGEMA_signal_8412 ;
    wire new_AGEMA_signal_8413 ;
    wire new_AGEMA_signal_8414 ;
    wire new_AGEMA_signal_8415 ;
    wire new_AGEMA_signal_8416 ;
    wire new_AGEMA_signal_8417 ;
    wire new_AGEMA_signal_8418 ;
    wire new_AGEMA_signal_8419 ;
    wire new_AGEMA_signal_8420 ;
    wire new_AGEMA_signal_8421 ;
    wire new_AGEMA_signal_8422 ;
    wire new_AGEMA_signal_8423 ;
    wire new_AGEMA_signal_8424 ;
    wire new_AGEMA_signal_8425 ;
    wire new_AGEMA_signal_8426 ;
    wire new_AGEMA_signal_8427 ;
    wire new_AGEMA_signal_8428 ;
    wire new_AGEMA_signal_8429 ;
    wire new_AGEMA_signal_8430 ;
    wire new_AGEMA_signal_8432 ;
    wire new_AGEMA_signal_8434 ;
    wire new_AGEMA_signal_8436 ;
    wire new_AGEMA_signal_8438 ;
    wire new_AGEMA_signal_8440 ;
    wire new_AGEMA_signal_8442 ;
    wire new_AGEMA_signal_8444 ;
    wire new_AGEMA_signal_8446 ;
    wire new_AGEMA_signal_8448 ;
    wire new_AGEMA_signal_8450 ;
    wire new_AGEMA_signal_8452 ;
    wire new_AGEMA_signal_8454 ;
    wire new_AGEMA_signal_8456 ;
    wire new_AGEMA_signal_8458 ;
    wire new_AGEMA_signal_8460 ;
    wire new_AGEMA_signal_8462 ;
    wire new_AGEMA_signal_8464 ;
    wire new_AGEMA_signal_8466 ;
    wire new_AGEMA_signal_8468 ;
    wire new_AGEMA_signal_8470 ;
    wire new_AGEMA_signal_8472 ;
    wire new_AGEMA_signal_8474 ;
    wire new_AGEMA_signal_8476 ;
    wire new_AGEMA_signal_8478 ;
    wire new_AGEMA_signal_8480 ;
    wire new_AGEMA_signal_8482 ;
    wire new_AGEMA_signal_8484 ;
    wire new_AGEMA_signal_8486 ;
    wire new_AGEMA_signal_8488 ;
    wire new_AGEMA_signal_8490 ;
    wire new_AGEMA_signal_8492 ;
    wire new_AGEMA_signal_8494 ;
    wire new_AGEMA_signal_8496 ;
    wire new_AGEMA_signal_8498 ;
    wire new_AGEMA_signal_8500 ;
    wire new_AGEMA_signal_8502 ;
    wire new_AGEMA_signal_8504 ;
    wire new_AGEMA_signal_8506 ;
    wire new_AGEMA_signal_8508 ;
    wire new_AGEMA_signal_8510 ;
    wire new_AGEMA_signal_8512 ;
    wire new_AGEMA_signal_8514 ;
    wire new_AGEMA_signal_8516 ;
    wire new_AGEMA_signal_8518 ;
    wire new_AGEMA_signal_8520 ;
    wire new_AGEMA_signal_8522 ;
    wire new_AGEMA_signal_8524 ;
    wire new_AGEMA_signal_8526 ;
    wire new_AGEMA_signal_8528 ;
    wire new_AGEMA_signal_8530 ;
    wire new_AGEMA_signal_8532 ;
    wire new_AGEMA_signal_8534 ;
    wire new_AGEMA_signal_8536 ;
    wire new_AGEMA_signal_8538 ;
    wire new_AGEMA_signal_8540 ;
    wire new_AGEMA_signal_8542 ;
    wire new_AGEMA_signal_8544 ;
    wire new_AGEMA_signal_8546 ;
    wire new_AGEMA_signal_8548 ;
    wire new_AGEMA_signal_8550 ;
    wire new_AGEMA_signal_8552 ;
    wire new_AGEMA_signal_8554 ;
    wire new_AGEMA_signal_8556 ;
    wire new_AGEMA_signal_8558 ;
    wire new_AGEMA_signal_8560 ;
    wire new_AGEMA_signal_8562 ;
    wire new_AGEMA_signal_8564 ;
    wire new_AGEMA_signal_8566 ;
    wire new_AGEMA_signal_8568 ;
    wire new_AGEMA_signal_8570 ;
    wire new_AGEMA_signal_8572 ;
    wire new_AGEMA_signal_8574 ;
    wire new_AGEMA_signal_8576 ;
    wire new_AGEMA_signal_8578 ;
    wire new_AGEMA_signal_8580 ;
    wire new_AGEMA_signal_8582 ;
    wire new_AGEMA_signal_8584 ;
    wire new_AGEMA_signal_8586 ;
    wire new_AGEMA_signal_8588 ;
    wire new_AGEMA_signal_8590 ;
    wire new_AGEMA_signal_8592 ;
    wire new_AGEMA_signal_8594 ;
    wire new_AGEMA_signal_8596 ;
    wire new_AGEMA_signal_8598 ;
    wire new_AGEMA_signal_8600 ;
    wire new_AGEMA_signal_8602 ;
    wire new_AGEMA_signal_8604 ;
    wire new_AGEMA_signal_8606 ;
    wire new_AGEMA_signal_8608 ;
    wire new_AGEMA_signal_8610 ;
    wire new_AGEMA_signal_8612 ;
    wire new_AGEMA_signal_8614 ;
    wire new_AGEMA_signal_8616 ;
    wire new_AGEMA_signal_8618 ;
    wire new_AGEMA_signal_8620 ;
    wire new_AGEMA_signal_8622 ;
    wire new_AGEMA_signal_8624 ;
    wire new_AGEMA_signal_8626 ;
    wire new_AGEMA_signal_8628 ;
    wire new_AGEMA_signal_8630 ;
    wire new_AGEMA_signal_8632 ;
    wire new_AGEMA_signal_8634 ;
    wire new_AGEMA_signal_8636 ;
    wire new_AGEMA_signal_8638 ;
    wire new_AGEMA_signal_8640 ;
    wire new_AGEMA_signal_8642 ;
    wire new_AGEMA_signal_8644 ;
    wire new_AGEMA_signal_8646 ;
    wire new_AGEMA_signal_8648 ;
    wire new_AGEMA_signal_8650 ;
    wire new_AGEMA_signal_8652 ;
    wire new_AGEMA_signal_8654 ;
    wire new_AGEMA_signal_8656 ;
    wire new_AGEMA_signal_8658 ;
    wire new_AGEMA_signal_8660 ;
    wire new_AGEMA_signal_8662 ;
    wire new_AGEMA_signal_8664 ;
    wire new_AGEMA_signal_8666 ;
    wire new_AGEMA_signal_8668 ;
    wire new_AGEMA_signal_8670 ;
    wire new_AGEMA_signal_8672 ;
    wire new_AGEMA_signal_8674 ;
    wire new_AGEMA_signal_8676 ;
    wire new_AGEMA_signal_8678 ;
    wire new_AGEMA_signal_8680 ;
    wire new_AGEMA_signal_8682 ;
    wire new_AGEMA_signal_8684 ;
    wire new_AGEMA_signal_8686 ;
    wire new_AGEMA_signal_8688 ;
    wire new_AGEMA_signal_8690 ;
    wire new_AGEMA_signal_8692 ;
    wire new_AGEMA_signal_8694 ;
    wire new_AGEMA_signal_8696 ;
    wire new_AGEMA_signal_8698 ;
    wire new_AGEMA_signal_8700 ;
    wire new_AGEMA_signal_10061 ;
    wire new_AGEMA_signal_10062 ;
    wire new_AGEMA_signal_10063 ;
    wire new_AGEMA_signal_10064 ;
    wire new_AGEMA_signal_10065 ;
    wire new_AGEMA_signal_10066 ;
    wire new_AGEMA_signal_10067 ;
    wire new_AGEMA_signal_10068 ;
    wire new_AGEMA_signal_10069 ;
    wire new_AGEMA_signal_10070 ;
    wire new_AGEMA_signal_10071 ;
    wire new_AGEMA_signal_10072 ;
    wire new_AGEMA_signal_10073 ;
    wire new_AGEMA_signal_10074 ;
    wire new_AGEMA_signal_10075 ;
    wire new_AGEMA_signal_10076 ;
    wire new_AGEMA_signal_10077 ;
    wire new_AGEMA_signal_10078 ;
    wire new_AGEMA_signal_10079 ;
    wire new_AGEMA_signal_10080 ;
    wire new_AGEMA_signal_10081 ;
    wire new_AGEMA_signal_10082 ;
    wire new_AGEMA_signal_10083 ;
    wire new_AGEMA_signal_10084 ;
    wire new_AGEMA_signal_10085 ;
    wire new_AGEMA_signal_10086 ;
    wire new_AGEMA_signal_10087 ;
    wire new_AGEMA_signal_10088 ;
    wire new_AGEMA_signal_10089 ;
    wire new_AGEMA_signal_10090 ;
    wire new_AGEMA_signal_10091 ;
    wire new_AGEMA_signal_10092 ;
    wire new_AGEMA_signal_10093 ;
    wire new_AGEMA_signal_10094 ;
    wire new_AGEMA_signal_10095 ;
    wire new_AGEMA_signal_10096 ;
    wire new_AGEMA_signal_10097 ;
    wire new_AGEMA_signal_10098 ;
    wire new_AGEMA_signal_10099 ;
    wire new_AGEMA_signal_10100 ;
    wire new_AGEMA_signal_10101 ;
    wire new_AGEMA_signal_10102 ;
    wire new_AGEMA_signal_10103 ;
    wire new_AGEMA_signal_10104 ;
    wire new_AGEMA_signal_10105 ;
    wire new_AGEMA_signal_10106 ;
    wire new_AGEMA_signal_10107 ;
    wire new_AGEMA_signal_10108 ;
    wire new_AGEMA_signal_10109 ;
    wire new_AGEMA_signal_10110 ;
    wire new_AGEMA_signal_10111 ;
    wire new_AGEMA_signal_10112 ;
    wire new_AGEMA_signal_10113 ;
    wire new_AGEMA_signal_10114 ;
    wire new_AGEMA_signal_10115 ;
    wire new_AGEMA_signal_10116 ;
    wire new_AGEMA_signal_10117 ;
    wire new_AGEMA_signal_10118 ;
    wire new_AGEMA_signal_10119 ;
    wire new_AGEMA_signal_10120 ;
    wire new_AGEMA_signal_10121 ;
    wire new_AGEMA_signal_10122 ;
    wire new_AGEMA_signal_10123 ;
    wire new_AGEMA_signal_10124 ;
    wire new_AGEMA_signal_10125 ;
    wire new_AGEMA_signal_10126 ;
    wire new_AGEMA_signal_10127 ;
    wire new_AGEMA_signal_10128 ;
    wire new_AGEMA_signal_10129 ;
    wire new_AGEMA_signal_10130 ;
    wire new_AGEMA_signal_10131 ;
    wire new_AGEMA_signal_10132 ;
    wire new_AGEMA_signal_10133 ;
    wire new_AGEMA_signal_10134 ;
    wire new_AGEMA_signal_10135 ;
    wire new_AGEMA_signal_10136 ;
    wire new_AGEMA_signal_10137 ;
    wire new_AGEMA_signal_10138 ;
    wire new_AGEMA_signal_10139 ;
    wire new_AGEMA_signal_10140 ;
    wire new_AGEMA_signal_10141 ;
    wire new_AGEMA_signal_10142 ;
    wire new_AGEMA_signal_10143 ;
    wire new_AGEMA_signal_10144 ;
    wire new_AGEMA_signal_10145 ;
    wire new_AGEMA_signal_10146 ;
    wire new_AGEMA_signal_10147 ;
    wire new_AGEMA_signal_10148 ;
    wire new_AGEMA_signal_10149 ;
    wire new_AGEMA_signal_10150 ;
    wire new_AGEMA_signal_10151 ;
    wire new_AGEMA_signal_10152 ;
    wire new_AGEMA_signal_10153 ;
    wire new_AGEMA_signal_10154 ;
    wire new_AGEMA_signal_10155 ;
    wire new_AGEMA_signal_10156 ;
    wire new_AGEMA_signal_10157 ;
    wire new_AGEMA_signal_10158 ;
    wire new_AGEMA_signal_10159 ;
    wire new_AGEMA_signal_10160 ;
    wire new_AGEMA_signal_10161 ;
    wire new_AGEMA_signal_10162 ;
    wire new_AGEMA_signal_10163 ;
    wire new_AGEMA_signal_10164 ;
    wire new_AGEMA_signal_10165 ;
    wire new_AGEMA_signal_10166 ;
    wire new_AGEMA_signal_10167 ;
    wire new_AGEMA_signal_10168 ;
    wire new_AGEMA_signal_10169 ;
    wire new_AGEMA_signal_10170 ;
    wire new_AGEMA_signal_10171 ;
    wire new_AGEMA_signal_10172 ;
    wire new_AGEMA_signal_10173 ;
    wire new_AGEMA_signal_10174 ;
    wire new_AGEMA_signal_10175 ;
    wire new_AGEMA_signal_10176 ;
    wire new_AGEMA_signal_10177 ;
    wire new_AGEMA_signal_10178 ;
    wire new_AGEMA_signal_10179 ;
    wire new_AGEMA_signal_10180 ;
    wire new_AGEMA_signal_10181 ;
    wire new_AGEMA_signal_10182 ;
    wire new_AGEMA_signal_10183 ;
    wire new_AGEMA_signal_10184 ;
    wire new_AGEMA_signal_10185 ;
    wire new_AGEMA_signal_10186 ;
    wire new_AGEMA_signal_10187 ;
    wire new_AGEMA_signal_10188 ;
    wire new_AGEMA_signal_10189 ;
    wire new_AGEMA_signal_10190 ;
    wire new_AGEMA_signal_10191 ;
    wire new_AGEMA_signal_10192 ;
    wire new_AGEMA_signal_10193 ;
    wire new_AGEMA_signal_10194 ;
    wire new_AGEMA_signal_10195 ;
    wire new_AGEMA_signal_10196 ;
    wire new_AGEMA_signal_10197 ;
    wire new_AGEMA_signal_10198 ;
    wire new_AGEMA_signal_10199 ;
    wire new_AGEMA_signal_10200 ;
    wire new_AGEMA_signal_10201 ;
    wire new_AGEMA_signal_10202 ;
    wire new_AGEMA_signal_10203 ;
    wire new_AGEMA_signal_10204 ;
    wire new_AGEMA_signal_10205 ;
    wire new_AGEMA_signal_10206 ;
    wire new_AGEMA_signal_10207 ;
    wire new_AGEMA_signal_10208 ;
    wire new_AGEMA_signal_10209 ;
    wire new_AGEMA_signal_10210 ;
    wire new_AGEMA_signal_10211 ;
    wire new_AGEMA_signal_10212 ;
    wire new_AGEMA_signal_10213 ;
    wire new_AGEMA_signal_10214 ;
    wire new_AGEMA_signal_10215 ;
    wire new_AGEMA_signal_10216 ;
    wire new_AGEMA_signal_10217 ;
    wire new_AGEMA_signal_10218 ;
    wire new_AGEMA_signal_10219 ;
    wire new_AGEMA_signal_10220 ;
    wire new_AGEMA_signal_10221 ;
    wire new_AGEMA_signal_10222 ;
    wire new_AGEMA_signal_10223 ;
    wire new_AGEMA_signal_10224 ;
    wire new_AGEMA_signal_10225 ;
    wire new_AGEMA_signal_10226 ;
    wire new_AGEMA_signal_10227 ;
    wire new_AGEMA_signal_10228 ;
    wire new_AGEMA_signal_10229 ;
    wire new_AGEMA_signal_10230 ;
    wire new_AGEMA_signal_10231 ;
    wire new_AGEMA_signal_10232 ;
    wire new_AGEMA_signal_10233 ;
    wire new_AGEMA_signal_10234 ;
    wire new_AGEMA_signal_10235 ;
    wire new_AGEMA_signal_10236 ;
    wire new_AGEMA_signal_10237 ;
    wire new_AGEMA_signal_10238 ;
    wire new_AGEMA_signal_10239 ;
    wire new_AGEMA_signal_10240 ;
    wire new_AGEMA_signal_10241 ;
    wire new_AGEMA_signal_10242 ;
    wire new_AGEMA_signal_10243 ;
    wire new_AGEMA_signal_10244 ;
    wire new_AGEMA_signal_10245 ;
    wire new_AGEMA_signal_10246 ;
    wire new_AGEMA_signal_10247 ;
    wire new_AGEMA_signal_10248 ;
    wire new_AGEMA_signal_10249 ;
    wire new_AGEMA_signal_10250 ;
    wire new_AGEMA_signal_10251 ;
    wire new_AGEMA_signal_10252 ;
    wire new_AGEMA_signal_10253 ;
    wire new_AGEMA_signal_10254 ;
    wire new_AGEMA_signal_10255 ;
    wire new_AGEMA_signal_10256 ;
    wire new_AGEMA_signal_10257 ;
    wire new_AGEMA_signal_10258 ;
    wire new_AGEMA_signal_10259 ;
    wire new_AGEMA_signal_10260 ;
    wire new_AGEMA_signal_10261 ;
    wire new_AGEMA_signal_10262 ;
    wire new_AGEMA_signal_10263 ;
    wire new_AGEMA_signal_10264 ;
    wire new_AGEMA_signal_10265 ;
    wire new_AGEMA_signal_10266 ;
    wire new_AGEMA_signal_10267 ;
    wire new_AGEMA_signal_10268 ;
    wire new_AGEMA_signal_10269 ;
    wire new_AGEMA_signal_10270 ;
    wire new_AGEMA_signal_10271 ;
    wire new_AGEMA_signal_10272 ;
    wire new_AGEMA_signal_10273 ;
    wire new_AGEMA_signal_10274 ;
    wire new_AGEMA_signal_10275 ;
    wire new_AGEMA_signal_10276 ;
    wire new_AGEMA_signal_10277 ;
    wire new_AGEMA_signal_10278 ;
    wire new_AGEMA_signal_10279 ;
    wire new_AGEMA_signal_10280 ;
    wire new_AGEMA_signal_10281 ;
    wire new_AGEMA_signal_10282 ;
    wire new_AGEMA_signal_10283 ;
    wire new_AGEMA_signal_10284 ;
    wire new_AGEMA_signal_10285 ;
    wire new_AGEMA_signal_10286 ;
    wire new_AGEMA_signal_10287 ;
    wire new_AGEMA_signal_10288 ;
    wire new_AGEMA_signal_10289 ;
    wire new_AGEMA_signal_10290 ;
    wire new_AGEMA_signal_10291 ;
    wire new_AGEMA_signal_10292 ;
    wire new_AGEMA_signal_10293 ;
    wire new_AGEMA_signal_10294 ;
    wire new_AGEMA_signal_10295 ;
    wire new_AGEMA_signal_10296 ;
    wire new_AGEMA_signal_10297 ;
    wire new_AGEMA_signal_10298 ;
    wire new_AGEMA_signal_10299 ;
    wire new_AGEMA_signal_10300 ;
    wire new_AGEMA_signal_10301 ;
    wire new_AGEMA_signal_10302 ;
    wire new_AGEMA_signal_10303 ;
    wire new_AGEMA_signal_10304 ;
    wire new_AGEMA_signal_10305 ;
    wire new_AGEMA_signal_10306 ;
    wire new_AGEMA_signal_10307 ;
    wire new_AGEMA_signal_10308 ;
    wire new_AGEMA_signal_10309 ;
    wire new_AGEMA_signal_10310 ;
    wire new_AGEMA_signal_10311 ;
    wire new_AGEMA_signal_10312 ;
    wire new_AGEMA_signal_10313 ;
    wire new_AGEMA_signal_10314 ;
    wire new_AGEMA_signal_10315 ;
    wire new_AGEMA_signal_10316 ;
    wire new_AGEMA_signal_10317 ;
    wire new_AGEMA_signal_10318 ;
    wire new_AGEMA_signal_10319 ;
    wire new_AGEMA_signal_10320 ;
    wire new_AGEMA_signal_10321 ;
    wire new_AGEMA_signal_10322 ;
    wire new_AGEMA_signal_10323 ;
    wire new_AGEMA_signal_10324 ;
    wire new_AGEMA_signal_10325 ;
    wire new_AGEMA_signal_10326 ;
    wire new_AGEMA_signal_10327 ;
    wire new_AGEMA_signal_10328 ;
    wire new_AGEMA_signal_10329 ;
    wire new_AGEMA_signal_10330 ;
    wire new_AGEMA_signal_10331 ;
    wire new_AGEMA_signal_10332 ;
    wire new_AGEMA_signal_10333 ;
    wire new_AGEMA_signal_10334 ;
    wire new_AGEMA_signal_10335 ;
    wire new_AGEMA_signal_10336 ;
    wire new_AGEMA_signal_10337 ;
    wire new_AGEMA_signal_10338 ;
    wire new_AGEMA_signal_10339 ;
    wire new_AGEMA_signal_10340 ;
    wire new_AGEMA_signal_10341 ;
    wire new_AGEMA_signal_10342 ;
    wire new_AGEMA_signal_10343 ;
    wire new_AGEMA_signal_10344 ;
    wire new_AGEMA_signal_10345 ;
    wire new_AGEMA_signal_10346 ;
    wire new_AGEMA_signal_10347 ;
    wire new_AGEMA_signal_10348 ;
    wire new_AGEMA_signal_10349 ;
    wire new_AGEMA_signal_10350 ;
    wire new_AGEMA_signal_10351 ;
    wire new_AGEMA_signal_10352 ;
    wire new_AGEMA_signal_10353 ;
    wire new_AGEMA_signal_10354 ;
    wire new_AGEMA_signal_10355 ;
    wire new_AGEMA_signal_10356 ;
    wire new_AGEMA_signal_10357 ;
    wire new_AGEMA_signal_10358 ;
    wire new_AGEMA_signal_10359 ;
    wire new_AGEMA_signal_10360 ;
    wire new_AGEMA_signal_10361 ;
    wire new_AGEMA_signal_10362 ;
    wire new_AGEMA_signal_10363 ;
    wire new_AGEMA_signal_10364 ;
    wire new_AGEMA_signal_10365 ;
    wire new_AGEMA_signal_10366 ;
    wire new_AGEMA_signal_10367 ;
    wire new_AGEMA_signal_10368 ;
    wire new_AGEMA_signal_10369 ;
    wire new_AGEMA_signal_10370 ;
    wire new_AGEMA_signal_10371 ;
    wire new_AGEMA_signal_10372 ;
    wire new_AGEMA_signal_10373 ;
    wire new_AGEMA_signal_10374 ;
    wire new_AGEMA_signal_10375 ;
    wire new_AGEMA_signal_10376 ;
    wire new_AGEMA_signal_10377 ;
    wire new_AGEMA_signal_10378 ;
    wire new_AGEMA_signal_10379 ;
    wire new_AGEMA_signal_10380 ;
    wire new_AGEMA_signal_10381 ;
    wire new_AGEMA_signal_10382 ;
    wire new_AGEMA_signal_10383 ;
    wire new_AGEMA_signal_10384 ;
    wire new_AGEMA_signal_10385 ;
    wire new_AGEMA_signal_10386 ;
    wire new_AGEMA_signal_10387 ;
    wire new_AGEMA_signal_10388 ;
    wire new_AGEMA_signal_10389 ;
    wire new_AGEMA_signal_10390 ;
    wire new_AGEMA_signal_10391 ;
    wire new_AGEMA_signal_10392 ;
    wire new_AGEMA_signal_10393 ;
    wire new_AGEMA_signal_10394 ;
    wire new_AGEMA_signal_10395 ;
    wire new_AGEMA_signal_10396 ;
    wire new_AGEMA_signal_10397 ;
    wire new_AGEMA_signal_10398 ;
    wire new_AGEMA_signal_10399 ;
    wire new_AGEMA_signal_10400 ;
    wire new_AGEMA_signal_10401 ;
    wire new_AGEMA_signal_10402 ;
    wire new_AGEMA_signal_10403 ;
    wire new_AGEMA_signal_10404 ;
    wire new_AGEMA_signal_10405 ;
    wire new_AGEMA_signal_10406 ;
    wire new_AGEMA_signal_10407 ;
    wire new_AGEMA_signal_10408 ;
    wire new_AGEMA_signal_10409 ;
    wire new_AGEMA_signal_10410 ;
    wire new_AGEMA_signal_10411 ;
    wire new_AGEMA_signal_10412 ;
    wire new_AGEMA_signal_10413 ;
    wire new_AGEMA_signal_10414 ;
    wire new_AGEMA_signal_10415 ;
    wire new_AGEMA_signal_10416 ;
    wire new_AGEMA_signal_10417 ;
    wire new_AGEMA_signal_10418 ;
    wire new_AGEMA_signal_10419 ;
    wire new_AGEMA_signal_10420 ;
    wire new_AGEMA_signal_10421 ;
    wire new_AGEMA_signal_10422 ;
    wire new_AGEMA_signal_10423 ;
    wire new_AGEMA_signal_10424 ;
    wire new_AGEMA_signal_10425 ;
    wire new_AGEMA_signal_10426 ;
    wire new_AGEMA_signal_10427 ;
    wire new_AGEMA_signal_10428 ;
    wire new_AGEMA_signal_10429 ;
    wire new_AGEMA_signal_10430 ;
    wire new_AGEMA_signal_10431 ;
    wire new_AGEMA_signal_10432 ;
    wire new_AGEMA_signal_10433 ;
    wire new_AGEMA_signal_10434 ;
    wire new_AGEMA_signal_10435 ;
    wire new_AGEMA_signal_10436 ;
    wire new_AGEMA_signal_10437 ;
    wire new_AGEMA_signal_10438 ;
    wire new_AGEMA_signal_10439 ;
    wire new_AGEMA_signal_10440 ;
    wire new_AGEMA_signal_10441 ;
    wire new_AGEMA_signal_10442 ;
    wire new_AGEMA_signal_10443 ;
    wire new_AGEMA_signal_10444 ;
    wire new_AGEMA_signal_10445 ;
    wire new_AGEMA_signal_10446 ;
    wire new_AGEMA_signal_10447 ;
    wire new_AGEMA_signal_10448 ;
    wire new_AGEMA_signal_10449 ;
    wire new_AGEMA_signal_10450 ;
    wire new_AGEMA_signal_10451 ;
    wire new_AGEMA_signal_10452 ;
    wire new_AGEMA_signal_10453 ;
    wire new_AGEMA_signal_10454 ;
    wire new_AGEMA_signal_10455 ;
    wire new_AGEMA_signal_10456 ;
    wire new_AGEMA_signal_10457 ;
    wire new_AGEMA_signal_10458 ;
    wire new_AGEMA_signal_10459 ;
    wire new_AGEMA_signal_10460 ;
    wire new_AGEMA_signal_10461 ;
    wire new_AGEMA_signal_10462 ;
    wire new_AGEMA_signal_10463 ;
    wire new_AGEMA_signal_10464 ;
    wire new_AGEMA_signal_10465 ;
    wire new_AGEMA_signal_10466 ;
    wire new_AGEMA_signal_10467 ;
    wire new_AGEMA_signal_10468 ;
    wire new_AGEMA_signal_10469 ;
    wire new_AGEMA_signal_10470 ;
    wire new_AGEMA_signal_10471 ;
    wire new_AGEMA_signal_10472 ;
    wire new_AGEMA_signal_10473 ;
    wire new_AGEMA_signal_10474 ;
    wire new_AGEMA_signal_10475 ;
    wire new_AGEMA_signal_10476 ;
    wire new_AGEMA_signal_10477 ;
    wire new_AGEMA_signal_10478 ;
    wire new_AGEMA_signal_10479 ;
    wire new_AGEMA_signal_10480 ;
    wire new_AGEMA_signal_10481 ;
    wire new_AGEMA_signal_10482 ;
    wire new_AGEMA_signal_10483 ;
    wire new_AGEMA_signal_10484 ;
    wire new_AGEMA_signal_10485 ;
    wire new_AGEMA_signal_10486 ;
    wire new_AGEMA_signal_10487 ;
    wire new_AGEMA_signal_10488 ;
    wire new_AGEMA_signal_10489 ;
    wire new_AGEMA_signal_10490 ;
    wire new_AGEMA_signal_10491 ;
    wire new_AGEMA_signal_10492 ;
    wire new_AGEMA_signal_10493 ;
    wire new_AGEMA_signal_10494 ;
    wire new_AGEMA_signal_10495 ;
    wire new_AGEMA_signal_10496 ;
    wire new_AGEMA_signal_10497 ;
    wire new_AGEMA_signal_10498 ;
    wire new_AGEMA_signal_10499 ;
    wire new_AGEMA_signal_10500 ;
    wire new_AGEMA_signal_10501 ;
    wire new_AGEMA_signal_10502 ;
    wire new_AGEMA_signal_10503 ;
    wire new_AGEMA_signal_10504 ;
    wire new_AGEMA_signal_10505 ;
    wire new_AGEMA_signal_10506 ;
    wire new_AGEMA_signal_10507 ;
    wire new_AGEMA_signal_10508 ;
    wire new_AGEMA_signal_10509 ;
    wire new_AGEMA_signal_10510 ;
    wire new_AGEMA_signal_10511 ;
    wire new_AGEMA_signal_10512 ;
    wire new_AGEMA_signal_10513 ;
    wire new_AGEMA_signal_10514 ;
    wire new_AGEMA_signal_10515 ;
    wire new_AGEMA_signal_10516 ;
    wire new_AGEMA_signal_10517 ;
    wire new_AGEMA_signal_10518 ;
    wire new_AGEMA_signal_10519 ;
    wire new_AGEMA_signal_10520 ;
    wire new_AGEMA_signal_10521 ;
    wire new_AGEMA_signal_10522 ;
    wire new_AGEMA_signal_10523 ;
    wire new_AGEMA_signal_10524 ;
    wire new_AGEMA_signal_10525 ;
    wire new_AGEMA_signal_10526 ;
    wire new_AGEMA_signal_10527 ;
    wire new_AGEMA_signal_10528 ;
    wire new_AGEMA_signal_10529 ;
    wire new_AGEMA_signal_10530 ;
    wire new_AGEMA_signal_10531 ;
    wire new_AGEMA_signal_10532 ;
    wire new_AGEMA_signal_10533 ;
    wire new_AGEMA_signal_10534 ;
    wire new_AGEMA_signal_10535 ;
    wire new_AGEMA_signal_10536 ;
    wire new_AGEMA_signal_10537 ;
    wire new_AGEMA_signal_10538 ;
    wire new_AGEMA_signal_10539 ;
    wire new_AGEMA_signal_10540 ;
    wire new_AGEMA_signal_10541 ;
    wire new_AGEMA_signal_10542 ;
    wire new_AGEMA_signal_10543 ;
    wire new_AGEMA_signal_10544 ;
    wire new_AGEMA_signal_10545 ;
    wire new_AGEMA_signal_10546 ;
    wire new_AGEMA_signal_10547 ;
    wire new_AGEMA_signal_10548 ;
    wire new_AGEMA_signal_10549 ;
    wire new_AGEMA_signal_10550 ;
    wire new_AGEMA_signal_10551 ;
    wire new_AGEMA_signal_10552 ;
    wire new_AGEMA_signal_10553 ;
    wire new_AGEMA_signal_10554 ;
    wire new_AGEMA_signal_10555 ;
    wire new_AGEMA_signal_10556 ;
    wire new_AGEMA_signal_10557 ;
    wire new_AGEMA_signal_10558 ;
    wire new_AGEMA_signal_10559 ;
    wire new_AGEMA_signal_10560 ;
    wire new_AGEMA_signal_10561 ;
    wire new_AGEMA_signal_10562 ;
    wire new_AGEMA_signal_10563 ;
    wire new_AGEMA_signal_10564 ;
    wire new_AGEMA_signal_10565 ;
    wire new_AGEMA_signal_10566 ;
    wire new_AGEMA_signal_10567 ;
    wire new_AGEMA_signal_10568 ;
    wire new_AGEMA_signal_10569 ;
    wire new_AGEMA_signal_10570 ;
    wire new_AGEMA_signal_10571 ;
    wire new_AGEMA_signal_10572 ;
    wire new_AGEMA_signal_10573 ;
    wire new_AGEMA_signal_10574 ;
    wire new_AGEMA_signal_10575 ;
    wire new_AGEMA_signal_10576 ;
    wire new_AGEMA_signal_10577 ;
    wire new_AGEMA_signal_10578 ;
    wire new_AGEMA_signal_10579 ;
    wire new_AGEMA_signal_10580 ;
    wire new_AGEMA_signal_10581 ;
    wire new_AGEMA_signal_10582 ;
    wire new_AGEMA_signal_10583 ;
    wire new_AGEMA_signal_10584 ;
    wire new_AGEMA_signal_10585 ;
    wire new_AGEMA_signal_10586 ;
    wire new_AGEMA_signal_10587 ;
    wire new_AGEMA_signal_10588 ;
    wire new_AGEMA_signal_10589 ;
    wire new_AGEMA_signal_10590 ;
    wire new_AGEMA_signal_10591 ;
    wire new_AGEMA_signal_10592 ;
    wire new_AGEMA_signal_10593 ;
    wire new_AGEMA_signal_10594 ;
    wire new_AGEMA_signal_10595 ;
    wire new_AGEMA_signal_10596 ;
    wire new_AGEMA_signal_10597 ;
    wire new_AGEMA_signal_10598 ;
    wire new_AGEMA_signal_10599 ;
    wire new_AGEMA_signal_10600 ;
    wire new_AGEMA_signal_10601 ;
    wire new_AGEMA_signal_10602 ;
    wire new_AGEMA_signal_10603 ;
    wire new_AGEMA_signal_10604 ;
    wire new_AGEMA_signal_10605 ;
    wire new_AGEMA_signal_10606 ;
    wire new_AGEMA_signal_10607 ;
    wire new_AGEMA_signal_10608 ;
    wire new_AGEMA_signal_10609 ;
    wire new_AGEMA_signal_10610 ;
    wire new_AGEMA_signal_10611 ;
    wire new_AGEMA_signal_10612 ;
    wire new_AGEMA_signal_10613 ;
    wire new_AGEMA_signal_10614 ;
    wire new_AGEMA_signal_10615 ;
    wire new_AGEMA_signal_10616 ;
    wire new_AGEMA_signal_10617 ;
    wire new_AGEMA_signal_10618 ;
    wire new_AGEMA_signal_10619 ;
    wire new_AGEMA_signal_10620 ;
    wire new_AGEMA_signal_10621 ;
    wire new_AGEMA_signal_10622 ;
    wire new_AGEMA_signal_10623 ;
    wire new_AGEMA_signal_10624 ;
    wire new_AGEMA_signal_10625 ;
    wire new_AGEMA_signal_10626 ;
    wire new_AGEMA_signal_10627 ;
    wire new_AGEMA_signal_10628 ;
    wire new_AGEMA_signal_10629 ;
    wire new_AGEMA_signal_10630 ;
    wire new_AGEMA_signal_10631 ;
    wire new_AGEMA_signal_10632 ;
    wire new_AGEMA_signal_10633 ;
    wire new_AGEMA_signal_10634 ;
    wire new_AGEMA_signal_10635 ;
    wire new_AGEMA_signal_10636 ;
    wire new_AGEMA_signal_10637 ;
    wire new_AGEMA_signal_10638 ;
    wire new_AGEMA_signal_10639 ;
    wire new_AGEMA_signal_10640 ;
    wire new_AGEMA_signal_10641 ;
    wire new_AGEMA_signal_10642 ;
    wire new_AGEMA_signal_10643 ;
    wire new_AGEMA_signal_10644 ;
    wire new_AGEMA_signal_10645 ;
    wire new_AGEMA_signal_10646 ;
    wire new_AGEMA_signal_10647 ;
    wire new_AGEMA_signal_10648 ;
    wire new_AGEMA_signal_10649 ;
    wire new_AGEMA_signal_10650 ;
    wire new_AGEMA_signal_10651 ;
    wire new_AGEMA_signal_10652 ;
    wire new_AGEMA_signal_10653 ;
    wire new_AGEMA_signal_10654 ;
    wire new_AGEMA_signal_10655 ;
    wire new_AGEMA_signal_10656 ;
    wire new_AGEMA_signal_10657 ;
    wire new_AGEMA_signal_10658 ;
    wire new_AGEMA_signal_10659 ;
    wire new_AGEMA_signal_10660 ;
    wire new_AGEMA_signal_10661 ;
    wire new_AGEMA_signal_10662 ;
    wire new_AGEMA_signal_10663 ;
    wire new_AGEMA_signal_10664 ;
    wire new_AGEMA_signal_10665 ;
    wire new_AGEMA_signal_10666 ;
    wire new_AGEMA_signal_10667 ;
    wire new_AGEMA_signal_10668 ;
    wire new_AGEMA_signal_10669 ;
    wire new_AGEMA_signal_10670 ;
    wire new_AGEMA_signal_10671 ;
    wire new_AGEMA_signal_10672 ;
    wire new_AGEMA_signal_10673 ;
    wire new_AGEMA_signal_10674 ;
    wire new_AGEMA_signal_10675 ;
    wire new_AGEMA_signal_10676 ;
    wire new_AGEMA_signal_10677 ;
    wire new_AGEMA_signal_10678 ;
    wire new_AGEMA_signal_10679 ;
    wire new_AGEMA_signal_10680 ;
    wire new_AGEMA_signal_10681 ;
    wire new_AGEMA_signal_10682 ;
    wire new_AGEMA_signal_10683 ;
    wire new_AGEMA_signal_10684 ;
    wire new_AGEMA_signal_10685 ;
    wire new_AGEMA_signal_10686 ;
    wire new_AGEMA_signal_10687 ;
    wire new_AGEMA_signal_10688 ;
    wire new_AGEMA_signal_10689 ;
    wire new_AGEMA_signal_10690 ;
    wire new_AGEMA_signal_10691 ;
    wire new_AGEMA_signal_10692 ;
    wire new_AGEMA_signal_10693 ;
    wire new_AGEMA_signal_10694 ;
    wire new_AGEMA_signal_10695 ;
    wire new_AGEMA_signal_10696 ;
    wire new_AGEMA_signal_10697 ;
    wire new_AGEMA_signal_10698 ;
    wire new_AGEMA_signal_10699 ;
    wire new_AGEMA_signal_10700 ;
    wire new_AGEMA_signal_10701 ;
    wire new_AGEMA_signal_10702 ;
    wire new_AGEMA_signal_10703 ;
    wire new_AGEMA_signal_10704 ;
    wire new_AGEMA_signal_10705 ;
    wire new_AGEMA_signal_10706 ;
    wire new_AGEMA_signal_10707 ;
    wire new_AGEMA_signal_10708 ;
    wire new_AGEMA_signal_10709 ;
    wire new_AGEMA_signal_10710 ;
    wire new_AGEMA_signal_10711 ;
    wire new_AGEMA_signal_10712 ;
    wire new_AGEMA_signal_10713 ;
    wire new_AGEMA_signal_10714 ;
    wire new_AGEMA_signal_10715 ;
    wire new_AGEMA_signal_10716 ;
    wire new_AGEMA_signal_10717 ;
    wire new_AGEMA_signal_10718 ;
    wire new_AGEMA_signal_10719 ;
    wire new_AGEMA_signal_10720 ;
    wire new_AGEMA_signal_10721 ;
    wire new_AGEMA_signal_10722 ;
    wire new_AGEMA_signal_10723 ;
    wire new_AGEMA_signal_10724 ;
    wire new_AGEMA_signal_10725 ;
    wire new_AGEMA_signal_10726 ;
    wire new_AGEMA_signal_10727 ;
    wire new_AGEMA_signal_10728 ;
    wire new_AGEMA_signal_10729 ;
    wire new_AGEMA_signal_10730 ;
    wire new_AGEMA_signal_10731 ;
    wire new_AGEMA_signal_10732 ;
    wire new_AGEMA_signal_10733 ;
    wire new_AGEMA_signal_10734 ;
    wire new_AGEMA_signal_10735 ;
    wire new_AGEMA_signal_10736 ;
    wire new_AGEMA_signal_10737 ;
    wire new_AGEMA_signal_10738 ;
    wire new_AGEMA_signal_10739 ;
    wire new_AGEMA_signal_10740 ;
    wire new_AGEMA_signal_10741 ;
    wire new_AGEMA_signal_10742 ;
    wire new_AGEMA_signal_10743 ;
    wire new_AGEMA_signal_10744 ;
    wire new_AGEMA_signal_10745 ;
    wire new_AGEMA_signal_10746 ;
    wire new_AGEMA_signal_10747 ;
    wire new_AGEMA_signal_10748 ;
    wire new_AGEMA_signal_10749 ;
    wire new_AGEMA_signal_10750 ;
    wire new_AGEMA_signal_10751 ;
    wire new_AGEMA_signal_10752 ;
    wire new_AGEMA_signal_10753 ;
    wire new_AGEMA_signal_10754 ;
    wire new_AGEMA_signal_10755 ;
    wire new_AGEMA_signal_10756 ;
    wire new_AGEMA_signal_10757 ;
    wire new_AGEMA_signal_10758 ;
    wire new_AGEMA_signal_10759 ;
    wire new_AGEMA_signal_10760 ;
    wire new_AGEMA_signal_10761 ;
    wire new_AGEMA_signal_10762 ;
    wire new_AGEMA_signal_10763 ;
    wire new_AGEMA_signal_10764 ;
    wire new_AGEMA_signal_10765 ;
    wire new_AGEMA_signal_10766 ;
    wire new_AGEMA_signal_10767 ;
    wire new_AGEMA_signal_10768 ;
    wire new_AGEMA_signal_10769 ;
    wire new_AGEMA_signal_10770 ;
    wire new_AGEMA_signal_10771 ;
    wire new_AGEMA_signal_10772 ;
    wire new_AGEMA_signal_10773 ;
    wire new_AGEMA_signal_10774 ;
    wire new_AGEMA_signal_10775 ;
    wire new_AGEMA_signal_10776 ;
    wire new_AGEMA_signal_10777 ;
    wire new_AGEMA_signal_10778 ;
    wire new_AGEMA_signal_10779 ;
    wire new_AGEMA_signal_10780 ;
    wire new_AGEMA_signal_10781 ;
    wire new_AGEMA_signal_10782 ;
    wire new_AGEMA_signal_10783 ;
    wire new_AGEMA_signal_10784 ;
    wire new_AGEMA_signal_10785 ;
    wire new_AGEMA_signal_10786 ;
    wire new_AGEMA_signal_10787 ;
    wire new_AGEMA_signal_10788 ;
    wire new_AGEMA_signal_10789 ;
    wire new_AGEMA_signal_10790 ;
    wire new_AGEMA_signal_10791 ;
    wire new_AGEMA_signal_10792 ;
    wire new_AGEMA_signal_10793 ;
    wire new_AGEMA_signal_10794 ;
    wire new_AGEMA_signal_10795 ;
    wire new_AGEMA_signal_10796 ;
    wire new_AGEMA_signal_10797 ;
    wire new_AGEMA_signal_10798 ;
    wire new_AGEMA_signal_10799 ;
    wire new_AGEMA_signal_10800 ;
    wire new_AGEMA_signal_10801 ;
    wire new_AGEMA_signal_10802 ;
    wire new_AGEMA_signal_10803 ;
    wire new_AGEMA_signal_10804 ;
    wire new_AGEMA_signal_10805 ;
    wire new_AGEMA_signal_10806 ;
    wire new_AGEMA_signal_10807 ;
    wire new_AGEMA_signal_10808 ;
    wire new_AGEMA_signal_10809 ;
    wire new_AGEMA_signal_10810 ;
    wire new_AGEMA_signal_10811 ;
    wire new_AGEMA_signal_10812 ;
    wire new_AGEMA_signal_10813 ;
    wire new_AGEMA_signal_10814 ;
    wire new_AGEMA_signal_10815 ;
    wire new_AGEMA_signal_10816 ;
    wire new_AGEMA_signal_10817 ;
    wire new_AGEMA_signal_10818 ;
    wire new_AGEMA_signal_10819 ;
    wire new_AGEMA_signal_10820 ;
    wire new_AGEMA_signal_10821 ;
    wire new_AGEMA_signal_10822 ;
    wire new_AGEMA_signal_10823 ;
    wire new_AGEMA_signal_10824 ;
    wire new_AGEMA_signal_10825 ;
    wire new_AGEMA_signal_10826 ;
    wire new_AGEMA_signal_10827 ;
    wire new_AGEMA_signal_10828 ;
    wire new_AGEMA_signal_10829 ;
    wire new_AGEMA_signal_10830 ;
    wire new_AGEMA_signal_10831 ;
    wire new_AGEMA_signal_10832 ;
    wire new_AGEMA_signal_10833 ;
    wire new_AGEMA_signal_10834 ;
    wire new_AGEMA_signal_10835 ;
    wire new_AGEMA_signal_10836 ;
    wire new_AGEMA_signal_10837 ;
    wire new_AGEMA_signal_10838 ;
    wire new_AGEMA_signal_10839 ;
    wire new_AGEMA_signal_10840 ;
    wire new_AGEMA_signal_10841 ;
    wire new_AGEMA_signal_10842 ;
    wire new_AGEMA_signal_10843 ;
    wire new_AGEMA_signal_10844 ;
    wire new_AGEMA_signal_10845 ;
    wire new_AGEMA_signal_10846 ;
    wire new_AGEMA_signal_10847 ;
    wire new_AGEMA_signal_10848 ;
    wire new_AGEMA_signal_10849 ;
    wire new_AGEMA_signal_10850 ;
    wire new_AGEMA_signal_10851 ;
    wire new_AGEMA_signal_10852 ;
    wire new_AGEMA_signal_10853 ;
    wire new_AGEMA_signal_10854 ;
    wire new_AGEMA_signal_10855 ;
    wire new_AGEMA_signal_10856 ;
    wire new_AGEMA_signal_10857 ;
    wire new_AGEMA_signal_10858 ;
    wire new_AGEMA_signal_10859 ;
    wire new_AGEMA_signal_10860 ;
    wire new_AGEMA_signal_10861 ;
    wire new_AGEMA_signal_10862 ;
    wire new_AGEMA_signal_10863 ;
    wire new_AGEMA_signal_10864 ;
    wire new_AGEMA_signal_10865 ;
    wire new_AGEMA_signal_10866 ;
    wire new_AGEMA_signal_10867 ;
    wire new_AGEMA_signal_10868 ;
    wire new_AGEMA_signal_10869 ;
    wire new_AGEMA_signal_10870 ;
    wire new_AGEMA_signal_10871 ;
    wire new_AGEMA_signal_10872 ;
    wire new_AGEMA_signal_10873 ;
    wire new_AGEMA_signal_10874 ;
    wire new_AGEMA_signal_10875 ;
    wire new_AGEMA_signal_10876 ;
    wire new_AGEMA_signal_10877 ;
    wire new_AGEMA_signal_10878 ;
    wire new_AGEMA_signal_10879 ;
    wire new_AGEMA_signal_10880 ;
    wire new_AGEMA_signal_10881 ;
    wire new_AGEMA_signal_10882 ;
    wire new_AGEMA_signal_10883 ;
    wire new_AGEMA_signal_10884 ;
    wire new_AGEMA_signal_10885 ;
    wire new_AGEMA_signal_10886 ;
    wire new_AGEMA_signal_10887 ;
    wire new_AGEMA_signal_10888 ;
    wire new_AGEMA_signal_10889 ;
    wire new_AGEMA_signal_10890 ;
    wire new_AGEMA_signal_10891 ;
    wire new_AGEMA_signal_10892 ;
    wire new_AGEMA_signal_10893 ;
    wire new_AGEMA_signal_10894 ;
    wire new_AGEMA_signal_10895 ;
    wire new_AGEMA_signal_10896 ;
    wire new_AGEMA_signal_10897 ;
    wire new_AGEMA_signal_10898 ;
    wire new_AGEMA_signal_10899 ;
    wire new_AGEMA_signal_10900 ;
    wire new_AGEMA_signal_10901 ;
    wire new_AGEMA_signal_10902 ;
    wire new_AGEMA_signal_10903 ;
    wire new_AGEMA_signal_10904 ;
    wire new_AGEMA_signal_10905 ;
    wire new_AGEMA_signal_10906 ;
    wire new_AGEMA_signal_10907 ;
    wire new_AGEMA_signal_10908 ;
    wire new_AGEMA_signal_10909 ;
    wire new_AGEMA_signal_10910 ;
    wire new_AGEMA_signal_10911 ;
    wire new_AGEMA_signal_10912 ;
    wire new_AGEMA_signal_10913 ;
    wire new_AGEMA_signal_10914 ;
    wire new_AGEMA_signal_10915 ;
    wire new_AGEMA_signal_10916 ;
    wire new_AGEMA_signal_10917 ;
    wire new_AGEMA_signal_10918 ;
    wire new_AGEMA_signal_10919 ;
    wire new_AGEMA_signal_10920 ;
    wire new_AGEMA_signal_10921 ;
    wire new_AGEMA_signal_10922 ;
    wire new_AGEMA_signal_10923 ;
    wire new_AGEMA_signal_10924 ;
    wire new_AGEMA_signal_10925 ;
    wire new_AGEMA_signal_10926 ;
    wire new_AGEMA_signal_10927 ;
    wire new_AGEMA_signal_10928 ;
    wire new_AGEMA_signal_10929 ;
    wire new_AGEMA_signal_10930 ;
    wire new_AGEMA_signal_10931 ;
    wire new_AGEMA_signal_10932 ;
    wire new_AGEMA_signal_10933 ;
    wire new_AGEMA_signal_10934 ;
    wire new_AGEMA_signal_10935 ;
    wire new_AGEMA_signal_10936 ;
    wire new_AGEMA_signal_10937 ;
    wire new_AGEMA_signal_10938 ;
    wire new_AGEMA_signal_10939 ;
    wire new_AGEMA_signal_10940 ;
    wire new_AGEMA_signal_10941 ;
    wire new_AGEMA_signal_10942 ;
    wire new_AGEMA_signal_10943 ;
    wire new_AGEMA_signal_10944 ;
    wire new_AGEMA_signal_10945 ;
    wire new_AGEMA_signal_10946 ;
    wire new_AGEMA_signal_10947 ;
    wire new_AGEMA_signal_10948 ;
    wire new_AGEMA_signal_10949 ;
    wire new_AGEMA_signal_10950 ;
    wire new_AGEMA_signal_10951 ;
    wire new_AGEMA_signal_10952 ;
    wire new_AGEMA_signal_10953 ;
    wire new_AGEMA_signal_10954 ;
    wire new_AGEMA_signal_10955 ;
    wire new_AGEMA_signal_10956 ;
    wire new_AGEMA_signal_10957 ;
    wire new_AGEMA_signal_10958 ;
    wire new_AGEMA_signal_10959 ;
    wire new_AGEMA_signal_10960 ;
    wire new_AGEMA_signal_10961 ;
    wire new_AGEMA_signal_10962 ;
    wire new_AGEMA_signal_10963 ;
    wire new_AGEMA_signal_10964 ;
    wire new_AGEMA_signal_10965 ;
    wire new_AGEMA_signal_10966 ;
    wire new_AGEMA_signal_10967 ;
    wire new_AGEMA_signal_10968 ;
    wire new_AGEMA_signal_10969 ;
    wire new_AGEMA_signal_10970 ;
    wire new_AGEMA_signal_10971 ;
    wire new_AGEMA_signal_10972 ;
    wire new_AGEMA_signal_10973 ;
    wire new_AGEMA_signal_10974 ;
    wire new_AGEMA_signal_10975 ;
    wire new_AGEMA_signal_10976 ;
    wire new_AGEMA_signal_10977 ;
    wire new_AGEMA_signal_10978 ;
    wire new_AGEMA_signal_10979 ;
    wire new_AGEMA_signal_10980 ;
    wire new_AGEMA_signal_10981 ;
    wire new_AGEMA_signal_10982 ;
    wire new_AGEMA_signal_10983 ;
    wire new_AGEMA_signal_10984 ;
    wire new_AGEMA_signal_10985 ;
    wire new_AGEMA_signal_10986 ;
    wire new_AGEMA_signal_10987 ;
    wire new_AGEMA_signal_10988 ;
    wire new_AGEMA_signal_10989 ;
    wire new_AGEMA_signal_10990 ;
    wire new_AGEMA_signal_10991 ;
    wire new_AGEMA_signal_10992 ;
    wire new_AGEMA_signal_10993 ;
    wire new_AGEMA_signal_10994 ;
    wire new_AGEMA_signal_10995 ;
    wire new_AGEMA_signal_10996 ;
    wire new_AGEMA_signal_10997 ;
    wire new_AGEMA_signal_10998 ;
    wire new_AGEMA_signal_10999 ;
    wire new_AGEMA_signal_11000 ;
    wire new_AGEMA_signal_11001 ;
    wire new_AGEMA_signal_11002 ;
    wire new_AGEMA_signal_11003 ;
    wire new_AGEMA_signal_11004 ;
    wire new_AGEMA_signal_11005 ;
    wire new_AGEMA_signal_11006 ;
    wire new_AGEMA_signal_11007 ;
    wire new_AGEMA_signal_11008 ;
    wire new_AGEMA_signal_11009 ;
    wire new_AGEMA_signal_11010 ;
    wire new_AGEMA_signal_11011 ;
    wire new_AGEMA_signal_11012 ;
    wire new_AGEMA_signal_11013 ;
    wire new_AGEMA_signal_11014 ;
    wire new_AGEMA_signal_11015 ;
    wire new_AGEMA_signal_11016 ;
    wire new_AGEMA_signal_11017 ;
    wire new_AGEMA_signal_11018 ;
    wire new_AGEMA_signal_11019 ;
    wire new_AGEMA_signal_11020 ;
    wire new_AGEMA_signal_11021 ;
    wire new_AGEMA_signal_11022 ;
    wire new_AGEMA_signal_11023 ;
    wire new_AGEMA_signal_11024 ;
    wire new_AGEMA_signal_11025 ;
    wire new_AGEMA_signal_11026 ;
    wire new_AGEMA_signal_11027 ;
    wire new_AGEMA_signal_11028 ;
    wire new_AGEMA_signal_11029 ;
    wire new_AGEMA_signal_11030 ;
    wire new_AGEMA_signal_11031 ;
    wire new_AGEMA_signal_11032 ;
    wire new_AGEMA_signal_11033 ;
    wire new_AGEMA_signal_11034 ;
    wire new_AGEMA_signal_11035 ;
    wire new_AGEMA_signal_11036 ;
    wire new_AGEMA_signal_11037 ;
    wire new_AGEMA_signal_11038 ;
    wire new_AGEMA_signal_11039 ;
    wire new_AGEMA_signal_11040 ;
    wire new_AGEMA_signal_11041 ;
    wire new_AGEMA_signal_11042 ;
    wire new_AGEMA_signal_11043 ;
    wire new_AGEMA_signal_11044 ;
    wire new_AGEMA_signal_11045 ;
    wire new_AGEMA_signal_11046 ;
    wire new_AGEMA_signal_11047 ;
    wire new_AGEMA_signal_11048 ;
    wire new_AGEMA_signal_11049 ;
    wire new_AGEMA_signal_11050 ;
    wire new_AGEMA_signal_11051 ;
    wire new_AGEMA_signal_11052 ;
    wire new_AGEMA_signal_11053 ;
    wire new_AGEMA_signal_11054 ;
    wire new_AGEMA_signal_11055 ;
    wire new_AGEMA_signal_11056 ;
    wire new_AGEMA_signal_11057 ;
    wire new_AGEMA_signal_11058 ;
    wire new_AGEMA_signal_11059 ;
    wire new_AGEMA_signal_11060 ;
    wire new_AGEMA_signal_11061 ;
    wire new_AGEMA_signal_11062 ;
    wire new_AGEMA_signal_11063 ;
    wire new_AGEMA_signal_11064 ;
    wire new_AGEMA_signal_11065 ;
    wire new_AGEMA_signal_11066 ;
    wire new_AGEMA_signal_11067 ;
    wire new_AGEMA_signal_11068 ;
    wire new_AGEMA_signal_11069 ;
    wire new_AGEMA_signal_11070 ;
    wire new_AGEMA_signal_11071 ;
    wire new_AGEMA_signal_11072 ;
    wire new_AGEMA_signal_11073 ;
    wire new_AGEMA_signal_11074 ;
    wire new_AGEMA_signal_11075 ;
    wire new_AGEMA_signal_11076 ;
    wire new_AGEMA_signal_11077 ;
    wire new_AGEMA_signal_11078 ;
    wire new_AGEMA_signal_11079 ;
    wire new_AGEMA_signal_11080 ;
    wire new_AGEMA_signal_11081 ;
    wire new_AGEMA_signal_11082 ;
    wire new_AGEMA_signal_11083 ;
    wire new_AGEMA_signal_11084 ;
    wire new_AGEMA_signal_11085 ;
    wire new_AGEMA_signal_11086 ;
    wire new_AGEMA_signal_11087 ;
    wire new_AGEMA_signal_11088 ;
    wire new_AGEMA_signal_11089 ;
    wire new_AGEMA_signal_11090 ;
    wire new_AGEMA_signal_11091 ;
    wire new_AGEMA_signal_11092 ;
    wire new_AGEMA_signal_11093 ;
    wire new_AGEMA_signal_11094 ;
    wire new_AGEMA_signal_11095 ;
    wire new_AGEMA_signal_11096 ;
    wire new_AGEMA_signal_11097 ;
    wire new_AGEMA_signal_11098 ;
    wire new_AGEMA_signal_11099 ;
    wire new_AGEMA_signal_11100 ;
    wire new_AGEMA_signal_11101 ;
    wire new_AGEMA_signal_11102 ;
    wire new_AGEMA_signal_11103 ;
    wire new_AGEMA_signal_11104 ;
    wire new_AGEMA_signal_11105 ;
    wire new_AGEMA_signal_11106 ;
    wire new_AGEMA_signal_11107 ;
    wire new_AGEMA_signal_11108 ;
    wire new_AGEMA_signal_11109 ;
    wire new_AGEMA_signal_11110 ;
    wire new_AGEMA_signal_11111 ;
    wire new_AGEMA_signal_11112 ;
    wire new_AGEMA_signal_11113 ;
    wire new_AGEMA_signal_11114 ;
    wire new_AGEMA_signal_11115 ;
    wire new_AGEMA_signal_11116 ;
    wire new_AGEMA_signal_11117 ;
    wire new_AGEMA_signal_11118 ;
    wire new_AGEMA_signal_11119 ;
    wire new_AGEMA_signal_11120 ;
    wire new_AGEMA_signal_11121 ;
    wire new_AGEMA_signal_11122 ;
    wire new_AGEMA_signal_11123 ;
    wire new_AGEMA_signal_11124 ;
    wire new_AGEMA_signal_11125 ;
    wire new_AGEMA_signal_11126 ;
    wire new_AGEMA_signal_11127 ;
    wire new_AGEMA_signal_11128 ;
    wire new_AGEMA_signal_11129 ;
    wire new_AGEMA_signal_11130 ;
    wire new_AGEMA_signal_11131 ;
    wire new_AGEMA_signal_11132 ;
    wire new_AGEMA_signal_11133 ;
    wire new_AGEMA_signal_11134 ;
    wire new_AGEMA_signal_11135 ;
    wire new_AGEMA_signal_11136 ;
    wire new_AGEMA_signal_11137 ;
    wire new_AGEMA_signal_11138 ;
    wire new_AGEMA_signal_11139 ;
    wire new_AGEMA_signal_11140 ;
    wire new_AGEMA_signal_11141 ;
    wire new_AGEMA_signal_11142 ;
    wire new_AGEMA_signal_11143 ;
    wire new_AGEMA_signal_11144 ;
    wire new_AGEMA_signal_11145 ;
    wire new_AGEMA_signal_11146 ;
    wire new_AGEMA_signal_11147 ;
    wire new_AGEMA_signal_11148 ;
    wire new_AGEMA_signal_11149 ;
    wire new_AGEMA_signal_11150 ;
    wire new_AGEMA_signal_11151 ;
    wire new_AGEMA_signal_11152 ;
    wire new_AGEMA_signal_11153 ;
    wire new_AGEMA_signal_11154 ;
    wire new_AGEMA_signal_11155 ;
    wire new_AGEMA_signal_11156 ;
    wire new_AGEMA_signal_11157 ;
    wire new_AGEMA_signal_11158 ;
    wire new_AGEMA_signal_11159 ;
    wire new_AGEMA_signal_11160 ;
    wire new_AGEMA_signal_11161 ;
    wire new_AGEMA_signal_11162 ;
    wire new_AGEMA_signal_11163 ;
    wire new_AGEMA_signal_11164 ;
    wire new_AGEMA_signal_11165 ;
    wire new_AGEMA_signal_11166 ;
    wire new_AGEMA_signal_11167 ;
    wire new_AGEMA_signal_11168 ;
    wire new_AGEMA_signal_11169 ;
    wire new_AGEMA_signal_11170 ;
    wire new_AGEMA_signal_11171 ;
    wire new_AGEMA_signal_11172 ;
    wire new_AGEMA_signal_11173 ;
    wire new_AGEMA_signal_11174 ;
    wire new_AGEMA_signal_11175 ;
    wire new_AGEMA_signal_11176 ;
    wire new_AGEMA_signal_11177 ;
    wire new_AGEMA_signal_11178 ;
    wire new_AGEMA_signal_11179 ;
    wire new_AGEMA_signal_11180 ;
    wire new_AGEMA_signal_11181 ;
    wire new_AGEMA_signal_11182 ;
    wire new_AGEMA_signal_11183 ;
    wire new_AGEMA_signal_11184 ;
    wire new_AGEMA_signal_11185 ;
    wire new_AGEMA_signal_11186 ;
    wire new_AGEMA_signal_11187 ;
    wire new_AGEMA_signal_11188 ;
    wire new_AGEMA_signal_11189 ;
    wire new_AGEMA_signal_11190 ;
    wire new_AGEMA_signal_11191 ;
    wire new_AGEMA_signal_11192 ;
    wire new_AGEMA_signal_11193 ;
    wire new_AGEMA_signal_11194 ;
    wire new_AGEMA_signal_11195 ;
    wire new_AGEMA_signal_11196 ;
    wire new_AGEMA_signal_11197 ;
    wire new_AGEMA_signal_11198 ;
    wire new_AGEMA_signal_11199 ;
    wire new_AGEMA_signal_11200 ;
    wire new_AGEMA_signal_11201 ;
    wire new_AGEMA_signal_11202 ;
    wire new_AGEMA_signal_11203 ;
    wire new_AGEMA_signal_11204 ;
    wire new_AGEMA_signal_11205 ;
    wire new_AGEMA_signal_11206 ;
    wire new_AGEMA_signal_11207 ;
    wire new_AGEMA_signal_11208 ;
    wire new_AGEMA_signal_11209 ;
    wire new_AGEMA_signal_11210 ;
    wire new_AGEMA_signal_11211 ;
    wire new_AGEMA_signal_11212 ;
    wire new_AGEMA_signal_11213 ;
    wire new_AGEMA_signal_11214 ;
    wire new_AGEMA_signal_11215 ;
    wire new_AGEMA_signal_11216 ;
    wire new_AGEMA_signal_11217 ;
    wire new_AGEMA_signal_11218 ;
    wire new_AGEMA_signal_11219 ;
    wire new_AGEMA_signal_11220 ;
    wire new_AGEMA_signal_11221 ;
    wire new_AGEMA_signal_11222 ;
    wire new_AGEMA_signal_11223 ;
    wire new_AGEMA_signal_11224 ;
    wire new_AGEMA_signal_11225 ;
    wire new_AGEMA_signal_11226 ;
    wire new_AGEMA_signal_11227 ;
    wire new_AGEMA_signal_11228 ;
    wire new_AGEMA_signal_11229 ;
    wire new_AGEMA_signal_11230 ;
    wire new_AGEMA_signal_11231 ;
    wire new_AGEMA_signal_11232 ;
    wire new_AGEMA_signal_11233 ;
    wire new_AGEMA_signal_11234 ;
    wire new_AGEMA_signal_11235 ;
    wire new_AGEMA_signal_11236 ;
    wire new_AGEMA_signal_11237 ;
    wire new_AGEMA_signal_11238 ;
    wire new_AGEMA_signal_11239 ;
    wire new_AGEMA_signal_11240 ;
    wire new_AGEMA_signal_11241 ;
    wire new_AGEMA_signal_11242 ;
    wire new_AGEMA_signal_11243 ;
    wire new_AGEMA_signal_11244 ;
    wire new_AGEMA_signal_11245 ;
    wire new_AGEMA_signal_11246 ;
    wire new_AGEMA_signal_11247 ;
    wire new_AGEMA_signal_11248 ;
    wire new_AGEMA_signal_11249 ;
    wire new_AGEMA_signal_11250 ;
    wire new_AGEMA_signal_11251 ;
    wire new_AGEMA_signal_11252 ;
    wire new_AGEMA_signal_11253 ;
    wire new_AGEMA_signal_11254 ;
    wire new_AGEMA_signal_11255 ;
    wire new_AGEMA_signal_11256 ;
    wire new_AGEMA_signal_11257 ;
    wire new_AGEMA_signal_11258 ;
    wire new_AGEMA_signal_11259 ;
    wire new_AGEMA_signal_11260 ;
    wire new_AGEMA_signal_11261 ;
    wire new_AGEMA_signal_11262 ;
    wire new_AGEMA_signal_11263 ;
    wire new_AGEMA_signal_11264 ;
    wire new_AGEMA_signal_11265 ;
    wire new_AGEMA_signal_11266 ;
    wire new_AGEMA_signal_11267 ;
    wire new_AGEMA_signal_11268 ;
    wire new_AGEMA_signal_11269 ;
    wire new_AGEMA_signal_11270 ;
    wire new_AGEMA_signal_11271 ;
    wire new_AGEMA_signal_11272 ;
    wire new_AGEMA_signal_11273 ;
    wire new_AGEMA_signal_11274 ;
    wire new_AGEMA_signal_11275 ;
    wire new_AGEMA_signal_11276 ;
    wire new_AGEMA_signal_11277 ;
    wire new_AGEMA_signal_11278 ;
    wire new_AGEMA_signal_11279 ;
    wire new_AGEMA_signal_11280 ;
    wire new_AGEMA_signal_11281 ;
    wire new_AGEMA_signal_11282 ;
    wire new_AGEMA_signal_11283 ;
    wire new_AGEMA_signal_11284 ;
    wire new_AGEMA_signal_11285 ;
    wire new_AGEMA_signal_11286 ;
    wire new_AGEMA_signal_11287 ;
    wire new_AGEMA_signal_11288 ;
    wire new_AGEMA_signal_11289 ;
    wire new_AGEMA_signal_11290 ;
    wire new_AGEMA_signal_11291 ;
    wire new_AGEMA_signal_11292 ;
    wire new_AGEMA_signal_11293 ;
    wire new_AGEMA_signal_11294 ;
    wire new_AGEMA_signal_11295 ;
    wire new_AGEMA_signal_11296 ;
    wire new_AGEMA_signal_11297 ;
    wire new_AGEMA_signal_11298 ;
    wire new_AGEMA_signal_11299 ;
    wire new_AGEMA_signal_11300 ;
    wire new_AGEMA_signal_11301 ;
    wire new_AGEMA_signal_11302 ;
    wire new_AGEMA_signal_11303 ;
    wire new_AGEMA_signal_11304 ;
    wire new_AGEMA_signal_11305 ;
    wire new_AGEMA_signal_11306 ;
    wire new_AGEMA_signal_11307 ;
    wire new_AGEMA_signal_11308 ;
    wire new_AGEMA_signal_11309 ;
    wire new_AGEMA_signal_11310 ;
    wire new_AGEMA_signal_11311 ;
    wire new_AGEMA_signal_11312 ;
    wire new_AGEMA_signal_11313 ;
    wire new_AGEMA_signal_11314 ;
    wire new_AGEMA_signal_11315 ;
    wire new_AGEMA_signal_11316 ;
    wire new_AGEMA_signal_11317 ;
    wire new_AGEMA_signal_11318 ;
    wire new_AGEMA_signal_11319 ;
    wire new_AGEMA_signal_11320 ;
    wire new_AGEMA_signal_11321 ;
    wire new_AGEMA_signal_11322 ;
    wire new_AGEMA_signal_11323 ;
    wire new_AGEMA_signal_11324 ;
    wire new_AGEMA_signal_11325 ;
    wire new_AGEMA_signal_11326 ;
    wire new_AGEMA_signal_11327 ;
    wire new_AGEMA_signal_11328 ;
    wire new_AGEMA_signal_11329 ;
    wire new_AGEMA_signal_11330 ;
    wire new_AGEMA_signal_11331 ;
    wire new_AGEMA_signal_11332 ;
    wire new_AGEMA_signal_11333 ;
    wire new_AGEMA_signal_11334 ;
    wire new_AGEMA_signal_11335 ;
    wire new_AGEMA_signal_11336 ;
    wire new_AGEMA_signal_11337 ;
    wire new_AGEMA_signal_11338 ;
    wire new_AGEMA_signal_11339 ;
    wire new_AGEMA_signal_11340 ;
    wire new_AGEMA_signal_11341 ;
    wire new_AGEMA_signal_11342 ;
    wire new_AGEMA_signal_11343 ;
    wire new_AGEMA_signal_11344 ;
    wire new_AGEMA_signal_11345 ;
    wire new_AGEMA_signal_11346 ;
    wire new_AGEMA_signal_11347 ;
    wire new_AGEMA_signal_11348 ;
    wire new_AGEMA_signal_11349 ;
    wire new_AGEMA_signal_11350 ;
    wire new_AGEMA_signal_11351 ;
    wire new_AGEMA_signal_11352 ;
    wire new_AGEMA_signal_11353 ;
    wire new_AGEMA_signal_11354 ;
    wire new_AGEMA_signal_11355 ;
    wire new_AGEMA_signal_11356 ;
    wire new_AGEMA_signal_11357 ;
    wire new_AGEMA_signal_11358 ;
    wire new_AGEMA_signal_11359 ;
    wire new_AGEMA_signal_11360 ;
    wire new_AGEMA_signal_11361 ;
    wire new_AGEMA_signal_11362 ;
    wire new_AGEMA_signal_11363 ;
    wire new_AGEMA_signal_11364 ;
    wire new_AGEMA_signal_11365 ;
    wire new_AGEMA_signal_11366 ;
    wire new_AGEMA_signal_11367 ;
    wire new_AGEMA_signal_11368 ;
    wire new_AGEMA_signal_11369 ;
    wire new_AGEMA_signal_11370 ;
    wire new_AGEMA_signal_11371 ;
    wire new_AGEMA_signal_11372 ;
    wire new_AGEMA_signal_11373 ;
    wire new_AGEMA_signal_11374 ;
    wire new_AGEMA_signal_11375 ;
    wire new_AGEMA_signal_11376 ;
    wire new_AGEMA_signal_11377 ;
    wire new_AGEMA_signal_11378 ;
    wire new_AGEMA_signal_11379 ;
    wire new_AGEMA_signal_11380 ;
    wire new_AGEMA_signal_11381 ;
    wire new_AGEMA_signal_11382 ;
    wire new_AGEMA_signal_11383 ;
    wire new_AGEMA_signal_11384 ;
    wire new_AGEMA_signal_11385 ;
    wire new_AGEMA_signal_11386 ;
    wire new_AGEMA_signal_11387 ;
    wire new_AGEMA_signal_11388 ;
    wire new_AGEMA_signal_11389 ;
    wire new_AGEMA_signal_11390 ;
    wire new_AGEMA_signal_11391 ;
    wire new_AGEMA_signal_11392 ;
    wire new_AGEMA_signal_11393 ;
    wire new_AGEMA_signal_11394 ;
    wire new_AGEMA_signal_11395 ;
    wire new_AGEMA_signal_11396 ;
    wire new_AGEMA_signal_11397 ;
    wire new_AGEMA_signal_11398 ;
    wire new_AGEMA_signal_11399 ;
    wire new_AGEMA_signal_11400 ;
    wire new_AGEMA_signal_11401 ;
    wire new_AGEMA_signal_11402 ;
    wire new_AGEMA_signal_11403 ;
    wire new_AGEMA_signal_11404 ;
    wire new_AGEMA_signal_11405 ;
    wire new_AGEMA_signal_11406 ;
    wire new_AGEMA_signal_11407 ;
    wire new_AGEMA_signal_11408 ;
    wire new_AGEMA_signal_11409 ;
    wire new_AGEMA_signal_11410 ;
    wire new_AGEMA_signal_11411 ;
    wire new_AGEMA_signal_11412 ;
    wire new_AGEMA_signal_11413 ;
    wire new_AGEMA_signal_11414 ;
    wire new_AGEMA_signal_11415 ;
    wire new_AGEMA_signal_11416 ;
    wire new_AGEMA_signal_11417 ;
    wire new_AGEMA_signal_11418 ;
    wire new_AGEMA_signal_11419 ;
    wire new_AGEMA_signal_11420 ;
    wire new_AGEMA_signal_11421 ;
    wire new_AGEMA_signal_11422 ;
    wire new_AGEMA_signal_11423 ;
    wire new_AGEMA_signal_11424 ;
    wire new_AGEMA_signal_11425 ;
    wire new_AGEMA_signal_11426 ;
    wire new_AGEMA_signal_11427 ;
    wire new_AGEMA_signal_11428 ;
    wire new_AGEMA_signal_11429 ;
    wire new_AGEMA_signal_11430 ;
    wire new_AGEMA_signal_11431 ;
    wire new_AGEMA_signal_11432 ;
    wire new_AGEMA_signal_11433 ;
    wire new_AGEMA_signal_11434 ;
    wire new_AGEMA_signal_11435 ;
    wire new_AGEMA_signal_11436 ;
    wire new_AGEMA_signal_11437 ;
    wire new_AGEMA_signal_11438 ;
    wire new_AGEMA_signal_11439 ;
    wire new_AGEMA_signal_11440 ;
    wire new_AGEMA_signal_11441 ;
    wire new_AGEMA_signal_11442 ;
    wire new_AGEMA_signal_11443 ;
    wire new_AGEMA_signal_11444 ;
    wire new_AGEMA_signal_11445 ;
    wire new_AGEMA_signal_11446 ;
    wire new_AGEMA_signal_11447 ;
    wire new_AGEMA_signal_11448 ;
    wire new_AGEMA_signal_11449 ;
    wire new_AGEMA_signal_11450 ;
    wire new_AGEMA_signal_11451 ;
    wire new_AGEMA_signal_11452 ;
    wire new_AGEMA_signal_11453 ;
    wire new_AGEMA_signal_11454 ;
    wire new_AGEMA_signal_11455 ;
    wire new_AGEMA_signal_11456 ;
    wire new_AGEMA_signal_11457 ;
    wire new_AGEMA_signal_11458 ;
    wire new_AGEMA_signal_11459 ;
    wire new_AGEMA_signal_11460 ;
    wire new_AGEMA_signal_11461 ;
    wire new_AGEMA_signal_11462 ;
    wire new_AGEMA_signal_11463 ;
    wire new_AGEMA_signal_11464 ;
    wire new_AGEMA_signal_11465 ;
    wire new_AGEMA_signal_11466 ;
    wire new_AGEMA_signal_11467 ;
    wire new_AGEMA_signal_11468 ;
    wire new_AGEMA_signal_11469 ;
    wire new_AGEMA_signal_11470 ;
    wire new_AGEMA_signal_11471 ;
    wire new_AGEMA_signal_11472 ;
    wire new_AGEMA_signal_11473 ;
    wire new_AGEMA_signal_11474 ;
    wire new_AGEMA_signal_11475 ;
    wire new_AGEMA_signal_11476 ;
    wire new_AGEMA_signal_11477 ;
    wire new_AGEMA_signal_11478 ;
    wire new_AGEMA_signal_11479 ;
    wire new_AGEMA_signal_11480 ;
    wire new_AGEMA_signal_11481 ;
    wire new_AGEMA_signal_11482 ;
    wire new_AGEMA_signal_11483 ;
    wire new_AGEMA_signal_11484 ;
    wire new_AGEMA_signal_11485 ;
    wire new_AGEMA_signal_11486 ;
    wire new_AGEMA_signal_11487 ;
    wire new_AGEMA_signal_11488 ;
    wire new_AGEMA_signal_11489 ;
    wire new_AGEMA_signal_11490 ;
    wire new_AGEMA_signal_11491 ;
    wire new_AGEMA_signal_11492 ;
    wire new_AGEMA_signal_11493 ;
    wire new_AGEMA_signal_11494 ;
    wire new_AGEMA_signal_11495 ;
    wire new_AGEMA_signal_11496 ;
    wire new_AGEMA_signal_11497 ;
    wire new_AGEMA_signal_11498 ;
    wire new_AGEMA_signal_11499 ;
    wire new_AGEMA_signal_11500 ;
    wire new_AGEMA_signal_11501 ;
    wire new_AGEMA_signal_11502 ;
    wire new_AGEMA_signal_11503 ;
    wire new_AGEMA_signal_11504 ;
    wire new_AGEMA_signal_11505 ;
    wire new_AGEMA_signal_11506 ;
    wire new_AGEMA_signal_11507 ;
    wire new_AGEMA_signal_11508 ;
    wire new_AGEMA_signal_11509 ;
    wire new_AGEMA_signal_11510 ;
    wire new_AGEMA_signal_11511 ;
    wire new_AGEMA_signal_11512 ;
    wire new_AGEMA_signal_11513 ;
    wire new_AGEMA_signal_11514 ;
    wire new_AGEMA_signal_11515 ;
    wire new_AGEMA_signal_11516 ;
    wire new_AGEMA_signal_11517 ;
    wire new_AGEMA_signal_11518 ;
    wire new_AGEMA_signal_11519 ;
    wire new_AGEMA_signal_11520 ;
    wire new_AGEMA_signal_11521 ;
    wire new_AGEMA_signal_11522 ;
    wire new_AGEMA_signal_11523 ;
    wire new_AGEMA_signal_11524 ;
    wire new_AGEMA_signal_11525 ;
    wire new_AGEMA_signal_11526 ;
    wire new_AGEMA_signal_11527 ;
    wire new_AGEMA_signal_11528 ;
    wire new_AGEMA_signal_11529 ;
    wire new_AGEMA_signal_11530 ;
    wire new_AGEMA_signal_11531 ;
    wire new_AGEMA_signal_11532 ;
    wire new_AGEMA_signal_11533 ;
    wire new_AGEMA_signal_11534 ;
    wire new_AGEMA_signal_11535 ;
    wire new_AGEMA_signal_11536 ;
    wire new_AGEMA_signal_11537 ;
    wire new_AGEMA_signal_11538 ;
    wire new_AGEMA_signal_11539 ;
    wire new_AGEMA_signal_11540 ;
    wire new_AGEMA_signal_11541 ;
    wire new_AGEMA_signal_11542 ;
    wire new_AGEMA_signal_11543 ;
    wire new_AGEMA_signal_11544 ;
    wire new_AGEMA_signal_11545 ;
    wire new_AGEMA_signal_11546 ;
    wire new_AGEMA_signal_11547 ;
    wire new_AGEMA_signal_11548 ;
    wire new_AGEMA_signal_11549 ;
    wire new_AGEMA_signal_11550 ;
    wire new_AGEMA_signal_11551 ;
    wire new_AGEMA_signal_11552 ;
    wire new_AGEMA_signal_11553 ;
    wire new_AGEMA_signal_11554 ;
    wire new_AGEMA_signal_11555 ;
    wire new_AGEMA_signal_11556 ;
    wire new_AGEMA_signal_11557 ;
    wire new_AGEMA_signal_11558 ;
    wire new_AGEMA_signal_11559 ;
    wire new_AGEMA_signal_11560 ;
    wire new_AGEMA_signal_11561 ;
    wire new_AGEMA_signal_11562 ;
    wire new_AGEMA_signal_11563 ;
    wire new_AGEMA_signal_11564 ;
    wire new_AGEMA_signal_11565 ;
    wire new_AGEMA_signal_11566 ;
    wire new_AGEMA_signal_11567 ;
    wire new_AGEMA_signal_11568 ;
    wire new_AGEMA_signal_11569 ;
    wire new_AGEMA_signal_11570 ;
    wire new_AGEMA_signal_11571 ;
    wire new_AGEMA_signal_11572 ;
    wire new_AGEMA_signal_11573 ;
    wire new_AGEMA_signal_11574 ;
    wire new_AGEMA_signal_11575 ;
    wire new_AGEMA_signal_11576 ;
    wire new_AGEMA_signal_11577 ;
    wire new_AGEMA_signal_11578 ;
    wire new_AGEMA_signal_11579 ;
    wire new_AGEMA_signal_11580 ;
    wire new_AGEMA_signal_11581 ;
    wire new_AGEMA_signal_11582 ;
    wire new_AGEMA_signal_11583 ;
    wire new_AGEMA_signal_11584 ;
    wire new_AGEMA_signal_11585 ;
    wire new_AGEMA_signal_11586 ;
    wire new_AGEMA_signal_11587 ;
    wire new_AGEMA_signal_11588 ;
    wire new_AGEMA_signal_11589 ;
    wire new_AGEMA_signal_11590 ;
    wire new_AGEMA_signal_11591 ;
    wire new_AGEMA_signal_11592 ;
    wire new_AGEMA_signal_11593 ;
    wire new_AGEMA_signal_11594 ;
    wire new_AGEMA_signal_11595 ;
    wire new_AGEMA_signal_11596 ;
    wire new_AGEMA_signal_11597 ;
    wire new_AGEMA_signal_11598 ;
    wire new_AGEMA_signal_11599 ;
    wire new_AGEMA_signal_11600 ;
    wire new_AGEMA_signal_11601 ;
    wire new_AGEMA_signal_11602 ;
    wire new_AGEMA_signal_11603 ;
    wire new_AGEMA_signal_11604 ;
    wire new_AGEMA_signal_11605 ;
    wire new_AGEMA_signal_11606 ;
    wire new_AGEMA_signal_11607 ;
    wire new_AGEMA_signal_11608 ;
    wire new_AGEMA_signal_11609 ;
    wire new_AGEMA_signal_11610 ;
    wire new_AGEMA_signal_11611 ;
    wire new_AGEMA_signal_11612 ;
    wire new_AGEMA_signal_11613 ;
    wire new_AGEMA_signal_11614 ;
    wire new_AGEMA_signal_11615 ;
    wire new_AGEMA_signal_11616 ;
    wire new_AGEMA_signal_11617 ;
    wire new_AGEMA_signal_11618 ;
    wire new_AGEMA_signal_11619 ;
    wire new_AGEMA_signal_11620 ;
    wire new_AGEMA_signal_11621 ;
    wire new_AGEMA_signal_11622 ;
    wire new_AGEMA_signal_11623 ;
    wire new_AGEMA_signal_11624 ;
    wire new_AGEMA_signal_11625 ;
    wire new_AGEMA_signal_11626 ;
    wire new_AGEMA_signal_11627 ;
    wire new_AGEMA_signal_11628 ;
    wire new_AGEMA_signal_11629 ;
    wire new_AGEMA_signal_11630 ;
    wire new_AGEMA_signal_11631 ;
    wire new_AGEMA_signal_11632 ;
    wire new_AGEMA_signal_11633 ;
    wire new_AGEMA_signal_11634 ;
    wire new_AGEMA_signal_11635 ;
    wire new_AGEMA_signal_11636 ;
    wire new_AGEMA_signal_11637 ;
    wire new_AGEMA_signal_11638 ;
    wire new_AGEMA_signal_11639 ;
    wire new_AGEMA_signal_11640 ;
    wire new_AGEMA_signal_11641 ;
    wire new_AGEMA_signal_11642 ;
    wire new_AGEMA_signal_11643 ;
    wire new_AGEMA_signal_11644 ;
    wire new_AGEMA_signal_11645 ;
    wire new_AGEMA_signal_11646 ;
    wire new_AGEMA_signal_11647 ;
    wire new_AGEMA_signal_11648 ;
    wire new_AGEMA_signal_11649 ;
    wire new_AGEMA_signal_11650 ;
    wire new_AGEMA_signal_11651 ;
    wire new_AGEMA_signal_11652 ;
    wire new_AGEMA_signal_11653 ;
    wire new_AGEMA_signal_11654 ;
    wire new_AGEMA_signal_11655 ;
    wire new_AGEMA_signal_11656 ;
    wire new_AGEMA_signal_11657 ;
    wire new_AGEMA_signal_11658 ;
    wire new_AGEMA_signal_11659 ;
    wire new_AGEMA_signal_11660 ;
    wire new_AGEMA_signal_11661 ;
    wire new_AGEMA_signal_11662 ;
    wire new_AGEMA_signal_11663 ;
    wire new_AGEMA_signal_11664 ;
    wire new_AGEMA_signal_11665 ;
    wire new_AGEMA_signal_11666 ;
    wire new_AGEMA_signal_11667 ;
    wire new_AGEMA_signal_11668 ;
    wire new_AGEMA_signal_11669 ;
    wire new_AGEMA_signal_11670 ;
    wire new_AGEMA_signal_11671 ;
    wire new_AGEMA_signal_11672 ;
    wire new_AGEMA_signal_11673 ;
    wire new_AGEMA_signal_11674 ;
    wire new_AGEMA_signal_11675 ;
    wire new_AGEMA_signal_11676 ;
    wire new_AGEMA_signal_11677 ;
    wire new_AGEMA_signal_11678 ;
    wire new_AGEMA_signal_11679 ;
    wire new_AGEMA_signal_11680 ;
    wire new_AGEMA_signal_11681 ;
    wire new_AGEMA_signal_11682 ;
    wire new_AGEMA_signal_11683 ;
    wire new_AGEMA_signal_11684 ;
    wire new_AGEMA_signal_11685 ;
    wire new_AGEMA_signal_11686 ;
    wire new_AGEMA_signal_11687 ;
    wire new_AGEMA_signal_11688 ;
    wire new_AGEMA_signal_11689 ;
    wire new_AGEMA_signal_11690 ;
    wire new_AGEMA_signal_11691 ;
    wire new_AGEMA_signal_11692 ;
    wire new_AGEMA_signal_11693 ;
    wire new_AGEMA_signal_11694 ;
    wire new_AGEMA_signal_11695 ;
    wire new_AGEMA_signal_11696 ;
    wire new_AGEMA_signal_11697 ;
    wire new_AGEMA_signal_11698 ;
    wire new_AGEMA_signal_11699 ;
    wire new_AGEMA_signal_11700 ;
    wire new_AGEMA_signal_11701 ;
    wire new_AGEMA_signal_11702 ;
    wire new_AGEMA_signal_11703 ;
    wire new_AGEMA_signal_11704 ;
    wire new_AGEMA_signal_11705 ;
    wire new_AGEMA_signal_11706 ;
    wire new_AGEMA_signal_11707 ;
    wire new_AGEMA_signal_11708 ;
    wire new_AGEMA_signal_11709 ;
    wire new_AGEMA_signal_11710 ;
    wire new_AGEMA_signal_11711 ;
    wire new_AGEMA_signal_11712 ;
    wire new_AGEMA_signal_11713 ;
    wire new_AGEMA_signal_11714 ;
    wire new_AGEMA_signal_11715 ;
    wire new_AGEMA_signal_11716 ;
    wire new_AGEMA_signal_11717 ;
    wire new_AGEMA_signal_11718 ;
    wire new_AGEMA_signal_11719 ;
    wire new_AGEMA_signal_11720 ;
    wire new_AGEMA_signal_11721 ;
    wire new_AGEMA_signal_11722 ;
    wire new_AGEMA_signal_11723 ;
    wire new_AGEMA_signal_11724 ;
    wire new_AGEMA_signal_11725 ;
    wire new_AGEMA_signal_11726 ;
    wire new_AGEMA_signal_11727 ;
    wire new_AGEMA_signal_11728 ;
    wire new_AGEMA_signal_11729 ;
    wire new_AGEMA_signal_11730 ;
    wire new_AGEMA_signal_11731 ;
    wire new_AGEMA_signal_11732 ;
    wire new_AGEMA_signal_11733 ;
    wire new_AGEMA_signal_11734 ;
    wire new_AGEMA_signal_11735 ;
    wire new_AGEMA_signal_11736 ;
    wire new_AGEMA_signal_11737 ;
    wire new_AGEMA_signal_11738 ;
    wire new_AGEMA_signal_11739 ;
    wire new_AGEMA_signal_11740 ;
    wire new_AGEMA_signal_11741 ;
    wire new_AGEMA_signal_11742 ;
    wire new_AGEMA_signal_11743 ;
    wire new_AGEMA_signal_11744 ;
    wire new_AGEMA_signal_11745 ;
    wire new_AGEMA_signal_11746 ;
    wire new_AGEMA_signal_11747 ;
    wire new_AGEMA_signal_11748 ;
    wire new_AGEMA_signal_11749 ;
    wire new_AGEMA_signal_11750 ;
    wire new_AGEMA_signal_11751 ;
    wire new_AGEMA_signal_11752 ;
    wire new_AGEMA_signal_11753 ;
    wire new_AGEMA_signal_11754 ;
    wire new_AGEMA_signal_11755 ;
    wire new_AGEMA_signal_11756 ;
    wire new_AGEMA_signal_11757 ;
    wire new_AGEMA_signal_11758 ;
    wire new_AGEMA_signal_11759 ;
    wire new_AGEMA_signal_11760 ;
    wire new_AGEMA_signal_11761 ;
    wire new_AGEMA_signal_11762 ;
    wire new_AGEMA_signal_11763 ;
    wire new_AGEMA_signal_11764 ;
    wire new_AGEMA_signal_11765 ;
    wire new_AGEMA_signal_11766 ;
    wire new_AGEMA_signal_11767 ;
    wire new_AGEMA_signal_11768 ;
    wire new_AGEMA_signal_11769 ;
    wire new_AGEMA_signal_11770 ;
    wire new_AGEMA_signal_11771 ;
    wire new_AGEMA_signal_11772 ;
    wire new_AGEMA_signal_11773 ;
    wire new_AGEMA_signal_11774 ;
    wire new_AGEMA_signal_11775 ;
    wire new_AGEMA_signal_11776 ;
    wire new_AGEMA_signal_11777 ;
    wire new_AGEMA_signal_11778 ;
    wire new_AGEMA_signal_11779 ;
    wire new_AGEMA_signal_11780 ;
    wire new_AGEMA_signal_11781 ;
    wire new_AGEMA_signal_11782 ;
    wire new_AGEMA_signal_11783 ;
    wire new_AGEMA_signal_11784 ;
    wire new_AGEMA_signal_11785 ;
    wire new_AGEMA_signal_11786 ;
    wire new_AGEMA_signal_11787 ;
    wire new_AGEMA_signal_11788 ;
    wire new_AGEMA_signal_11789 ;
    wire new_AGEMA_signal_11790 ;
    wire new_AGEMA_signal_11791 ;
    wire new_AGEMA_signal_11792 ;
    wire new_AGEMA_signal_11793 ;
    wire new_AGEMA_signal_11794 ;
    wire new_AGEMA_signal_11795 ;
    wire new_AGEMA_signal_11796 ;
    wire new_AGEMA_signal_11797 ;
    wire new_AGEMA_signal_11798 ;
    wire new_AGEMA_signal_11799 ;
    wire new_AGEMA_signal_11800 ;
    wire new_AGEMA_signal_11801 ;
    wire new_AGEMA_signal_11802 ;
    wire new_AGEMA_signal_11803 ;
    wire new_AGEMA_signal_11804 ;
    wire new_AGEMA_signal_11805 ;
    wire new_AGEMA_signal_11806 ;
    wire new_AGEMA_signal_11807 ;
    wire new_AGEMA_signal_11808 ;
    wire new_AGEMA_signal_11809 ;
    wire new_AGEMA_signal_11810 ;
    wire new_AGEMA_signal_11811 ;
    wire new_AGEMA_signal_11812 ;
    wire new_AGEMA_signal_11813 ;
    wire new_AGEMA_signal_11814 ;
    wire new_AGEMA_signal_11815 ;
    wire new_AGEMA_signal_11816 ;
    wire new_AGEMA_signal_11817 ;
    wire new_AGEMA_signal_11818 ;
    wire new_AGEMA_signal_11819 ;
    wire new_AGEMA_signal_11820 ;
    wire new_AGEMA_signal_11821 ;
    wire new_AGEMA_signal_11822 ;
    wire new_AGEMA_signal_11823 ;
    wire new_AGEMA_signal_11824 ;
    wire new_AGEMA_signal_11825 ;
    wire new_AGEMA_signal_11826 ;
    wire new_AGEMA_signal_11827 ;
    wire new_AGEMA_signal_11828 ;
    wire new_AGEMA_signal_11829 ;
    wire new_AGEMA_signal_11830 ;
    wire new_AGEMA_signal_11831 ;
    wire new_AGEMA_signal_11832 ;
    wire new_AGEMA_signal_11833 ;
    wire new_AGEMA_signal_11834 ;
    wire new_AGEMA_signal_11835 ;
    wire new_AGEMA_signal_11836 ;
    wire new_AGEMA_signal_11837 ;
    wire new_AGEMA_signal_11838 ;
    wire new_AGEMA_signal_11839 ;
    wire new_AGEMA_signal_11840 ;
    wire new_AGEMA_signal_11841 ;
    wire new_AGEMA_signal_11842 ;
    wire new_AGEMA_signal_11843 ;
    wire new_AGEMA_signal_11844 ;
    wire new_AGEMA_signal_11845 ;
    wire new_AGEMA_signal_11846 ;
    wire new_AGEMA_signal_11847 ;
    wire new_AGEMA_signal_11848 ;
    wire new_AGEMA_signal_11849 ;
    wire new_AGEMA_signal_11850 ;
    wire new_AGEMA_signal_11851 ;
    wire new_AGEMA_signal_11852 ;
    wire new_AGEMA_signal_11853 ;
    wire new_AGEMA_signal_11854 ;
    wire new_AGEMA_signal_11855 ;
    wire new_AGEMA_signal_11856 ;
    wire new_AGEMA_signal_11857 ;
    wire new_AGEMA_signal_11858 ;
    wire new_AGEMA_signal_11859 ;
    wire new_AGEMA_signal_11860 ;
    wire new_AGEMA_signal_11861 ;
    wire new_AGEMA_signal_11862 ;
    wire new_AGEMA_signal_11863 ;
    wire new_AGEMA_signal_11864 ;
    wire new_AGEMA_signal_11865 ;
    wire new_AGEMA_signal_11866 ;
    wire new_AGEMA_signal_11867 ;
    wire new_AGEMA_signal_11868 ;
    wire new_AGEMA_signal_11869 ;
    wire new_AGEMA_signal_11870 ;
    wire new_AGEMA_signal_11871 ;
    wire new_AGEMA_signal_11872 ;
    wire new_AGEMA_signal_11873 ;
    wire new_AGEMA_signal_11874 ;
    wire new_AGEMA_signal_11875 ;
    wire new_AGEMA_signal_11876 ;
    wire new_AGEMA_signal_11877 ;
    wire new_AGEMA_signal_11878 ;
    wire new_AGEMA_signal_11879 ;
    wire new_AGEMA_signal_11880 ;
    wire new_AGEMA_signal_11881 ;
    wire new_AGEMA_signal_11882 ;
    wire new_AGEMA_signal_11883 ;
    wire new_AGEMA_signal_11884 ;
    wire new_AGEMA_signal_11885 ;
    wire new_AGEMA_signal_11886 ;
    wire new_AGEMA_signal_11887 ;
    wire new_AGEMA_signal_11888 ;
    wire new_AGEMA_signal_11889 ;
    wire new_AGEMA_signal_11890 ;
    wire new_AGEMA_signal_11891 ;
    wire new_AGEMA_signal_11892 ;
    wire new_AGEMA_signal_11893 ;
    wire new_AGEMA_signal_11894 ;
    wire new_AGEMA_signal_11895 ;
    wire new_AGEMA_signal_11896 ;
    wire new_AGEMA_signal_11897 ;
    wire new_AGEMA_signal_11898 ;
    wire new_AGEMA_signal_11899 ;
    wire new_AGEMA_signal_11900 ;
    wire new_AGEMA_signal_11901 ;
    wire new_AGEMA_signal_11902 ;
    wire new_AGEMA_signal_11903 ;
    wire new_AGEMA_signal_11904 ;
    wire new_AGEMA_signal_11905 ;
    wire new_AGEMA_signal_11906 ;
    wire new_AGEMA_signal_11907 ;
    wire new_AGEMA_signal_11908 ;
    wire new_AGEMA_signal_11909 ;
    wire new_AGEMA_signal_11910 ;
    wire new_AGEMA_signal_11911 ;
    wire new_AGEMA_signal_11912 ;
    wire new_AGEMA_signal_11913 ;
    wire new_AGEMA_signal_11914 ;
    wire new_AGEMA_signal_11915 ;
    wire new_AGEMA_signal_11916 ;
    wire new_AGEMA_signal_11917 ;
    wire new_AGEMA_signal_11918 ;
    wire new_AGEMA_signal_11919 ;
    wire new_AGEMA_signal_11920 ;
    wire new_AGEMA_signal_11921 ;
    wire new_AGEMA_signal_11922 ;
    wire new_AGEMA_signal_11923 ;
    wire new_AGEMA_signal_11924 ;
    wire new_AGEMA_signal_11925 ;
    wire new_AGEMA_signal_11926 ;
    wire new_AGEMA_signal_11927 ;
    wire new_AGEMA_signal_11928 ;
    wire new_AGEMA_signal_11929 ;
    wire new_AGEMA_signal_11930 ;
    wire new_AGEMA_signal_11931 ;
    wire new_AGEMA_signal_11932 ;
    wire new_AGEMA_signal_11933 ;
    wire new_AGEMA_signal_11934 ;
    wire new_AGEMA_signal_11935 ;
    wire new_AGEMA_signal_11936 ;
    wire new_AGEMA_signal_11937 ;
    wire new_AGEMA_signal_11938 ;
    wire new_AGEMA_signal_11939 ;
    wire new_AGEMA_signal_11940 ;
    wire new_AGEMA_signal_11941 ;
    wire new_AGEMA_signal_11942 ;
    wire new_AGEMA_signal_11943 ;
    wire new_AGEMA_signal_11944 ;
    wire new_AGEMA_signal_11945 ;
    wire new_AGEMA_signal_11946 ;
    wire new_AGEMA_signal_11947 ;
    wire new_AGEMA_signal_11948 ;
    wire new_AGEMA_signal_11949 ;
    wire new_AGEMA_signal_11950 ;
    wire new_AGEMA_signal_11951 ;
    wire new_AGEMA_signal_11952 ;
    wire new_AGEMA_signal_11953 ;
    wire new_AGEMA_signal_11954 ;
    wire new_AGEMA_signal_11955 ;
    wire new_AGEMA_signal_11956 ;
    wire new_AGEMA_signal_11957 ;
    wire new_AGEMA_signal_11958 ;
    wire new_AGEMA_signal_11959 ;
    wire new_AGEMA_signal_11960 ;
    wire new_AGEMA_signal_11961 ;
    wire new_AGEMA_signal_11962 ;
    wire new_AGEMA_signal_11963 ;
    wire new_AGEMA_signal_11964 ;
    wire new_AGEMA_signal_11965 ;
    wire new_AGEMA_signal_11966 ;
    wire new_AGEMA_signal_11967 ;
    wire new_AGEMA_signal_11968 ;
    wire new_AGEMA_signal_11969 ;
    wire new_AGEMA_signal_11970 ;
    wire new_AGEMA_signal_11971 ;
    wire new_AGEMA_signal_11972 ;
    wire new_AGEMA_signal_11973 ;
    wire new_AGEMA_signal_11974 ;
    wire new_AGEMA_signal_11975 ;
    wire new_AGEMA_signal_11976 ;
    wire new_AGEMA_signal_11977 ;
    wire new_AGEMA_signal_11978 ;
    wire new_AGEMA_signal_11979 ;
    wire new_AGEMA_signal_11980 ;
    wire new_AGEMA_signal_11981 ;
    wire new_AGEMA_signal_11982 ;
    wire new_AGEMA_signal_11983 ;
    wire new_AGEMA_signal_11984 ;
    wire new_AGEMA_signal_11985 ;
    wire new_AGEMA_signal_11986 ;
    wire new_AGEMA_signal_11987 ;
    wire new_AGEMA_signal_11988 ;
    wire new_AGEMA_signal_11989 ;
    wire new_AGEMA_signal_11990 ;
    wire new_AGEMA_signal_11991 ;
    wire new_AGEMA_signal_11992 ;
    wire new_AGEMA_signal_11993 ;
    wire new_AGEMA_signal_11994 ;
    wire new_AGEMA_signal_11995 ;
    wire new_AGEMA_signal_11996 ;
    wire new_AGEMA_signal_11997 ;
    wire new_AGEMA_signal_11998 ;
    wire new_AGEMA_signal_11999 ;
    wire new_AGEMA_signal_12000 ;
    wire new_AGEMA_signal_12001 ;
    wire new_AGEMA_signal_12002 ;
    wire new_AGEMA_signal_12003 ;
    wire new_AGEMA_signal_12004 ;
    wire new_AGEMA_signal_12005 ;
    wire new_AGEMA_signal_12006 ;
    wire new_AGEMA_signal_12007 ;
    wire new_AGEMA_signal_12008 ;
    wire new_AGEMA_signal_12009 ;
    wire new_AGEMA_signal_12010 ;
    wire new_AGEMA_signal_12011 ;
    wire new_AGEMA_signal_12012 ;
    wire new_AGEMA_signal_12013 ;
    wire new_AGEMA_signal_12014 ;
    wire new_AGEMA_signal_12015 ;
    wire new_AGEMA_signal_12016 ;
    wire new_AGEMA_signal_12017 ;
    wire new_AGEMA_signal_12018 ;
    wire new_AGEMA_signal_12019 ;
    wire new_AGEMA_signal_12020 ;
    wire new_AGEMA_signal_12021 ;
    wire new_AGEMA_signal_12022 ;
    wire new_AGEMA_signal_12023 ;
    wire new_AGEMA_signal_12024 ;
    wire new_AGEMA_signal_12025 ;
    wire new_AGEMA_signal_12026 ;
    wire new_AGEMA_signal_12027 ;
    wire new_AGEMA_signal_12028 ;
    wire new_AGEMA_signal_12029 ;
    wire new_AGEMA_signal_12030 ;
    wire new_AGEMA_signal_12031 ;
    wire new_AGEMA_signal_12032 ;
    wire new_AGEMA_signal_12033 ;
    wire new_AGEMA_signal_12034 ;
    wire new_AGEMA_signal_12035 ;
    wire new_AGEMA_signal_12036 ;
    wire new_AGEMA_signal_12037 ;
    wire new_AGEMA_signal_12038 ;
    wire new_AGEMA_signal_12039 ;
    wire new_AGEMA_signal_12040 ;
    wire new_AGEMA_signal_12041 ;
    wire new_AGEMA_signal_12042 ;
    wire new_AGEMA_signal_12043 ;
    wire new_AGEMA_signal_12044 ;
    wire new_AGEMA_signal_12045 ;
    wire new_AGEMA_signal_12046 ;
    wire new_AGEMA_signal_12047 ;
    wire new_AGEMA_signal_12048 ;
    wire new_AGEMA_signal_12049 ;
    wire new_AGEMA_signal_12050 ;
    wire new_AGEMA_signal_12051 ;
    wire new_AGEMA_signal_12052 ;
    wire new_AGEMA_signal_12053 ;
    wire new_AGEMA_signal_12054 ;
    wire new_AGEMA_signal_12055 ;
    wire new_AGEMA_signal_12056 ;
    wire new_AGEMA_signal_12057 ;
    wire new_AGEMA_signal_12058 ;
    wire new_AGEMA_signal_12059 ;
    wire new_AGEMA_signal_12060 ;
    wire new_AGEMA_signal_12061 ;
    wire new_AGEMA_signal_12062 ;
    wire new_AGEMA_signal_12063 ;
    wire new_AGEMA_signal_12064 ;
    wire new_AGEMA_signal_12065 ;
    wire new_AGEMA_signal_12066 ;
    wire new_AGEMA_signal_12067 ;
    wire new_AGEMA_signal_12068 ;
    wire new_AGEMA_signal_12069 ;
    wire new_AGEMA_signal_12070 ;
    wire new_AGEMA_signal_12071 ;
    wire new_AGEMA_signal_12072 ;
    wire new_AGEMA_signal_12073 ;
    wire new_AGEMA_signal_12074 ;
    wire new_AGEMA_signal_12075 ;
    wire new_AGEMA_signal_12076 ;
    wire new_AGEMA_signal_12077 ;
    wire new_AGEMA_signal_12078 ;
    wire new_AGEMA_signal_12079 ;
    wire new_AGEMA_signal_12080 ;
    wire new_AGEMA_signal_12081 ;
    wire new_AGEMA_signal_12082 ;
    wire new_AGEMA_signal_12083 ;
    wire new_AGEMA_signal_12084 ;
    wire new_AGEMA_signal_12085 ;
    wire new_AGEMA_signal_12086 ;
    wire new_AGEMA_signal_12087 ;
    wire new_AGEMA_signal_12088 ;
    wire new_AGEMA_signal_12089 ;
    wire new_AGEMA_signal_12090 ;
    wire new_AGEMA_signal_12091 ;
    wire new_AGEMA_signal_12092 ;
    wire new_AGEMA_signal_12093 ;
    wire new_AGEMA_signal_12094 ;
    wire new_AGEMA_signal_12095 ;
    wire new_AGEMA_signal_12096 ;
    wire new_AGEMA_signal_12097 ;
    wire new_AGEMA_signal_12098 ;
    wire new_AGEMA_signal_12099 ;
    wire new_AGEMA_signal_12100 ;
    wire new_AGEMA_signal_12101 ;
    wire new_AGEMA_signal_12102 ;
    wire new_AGEMA_signal_12103 ;
    wire new_AGEMA_signal_12104 ;
    wire new_AGEMA_signal_12105 ;
    wire new_AGEMA_signal_12106 ;
    wire new_AGEMA_signal_12107 ;
    wire new_AGEMA_signal_12108 ;
    wire new_AGEMA_signal_12109 ;
    wire new_AGEMA_signal_12110 ;
    wire new_AGEMA_signal_12111 ;
    wire new_AGEMA_signal_12112 ;
    wire new_AGEMA_signal_12113 ;
    wire new_AGEMA_signal_12114 ;
    wire new_AGEMA_signal_12115 ;
    wire new_AGEMA_signal_12116 ;
    wire new_AGEMA_signal_12117 ;
    wire new_AGEMA_signal_12118 ;
    wire new_AGEMA_signal_12119 ;
    wire new_AGEMA_signal_12120 ;
    wire new_AGEMA_signal_12121 ;
    wire new_AGEMA_signal_12122 ;
    wire new_AGEMA_signal_12123 ;
    wire new_AGEMA_signal_12124 ;
    wire new_AGEMA_signal_12125 ;
    wire new_AGEMA_signal_12126 ;
    wire new_AGEMA_signal_12127 ;
    wire new_AGEMA_signal_12128 ;
    wire new_AGEMA_signal_12129 ;
    wire new_AGEMA_signal_12130 ;
    wire new_AGEMA_signal_12131 ;
    wire new_AGEMA_signal_12132 ;
    wire new_AGEMA_signal_12133 ;
    wire new_AGEMA_signal_12134 ;
    wire new_AGEMA_signal_12135 ;
    wire new_AGEMA_signal_12136 ;
    wire new_AGEMA_signal_12137 ;
    wire new_AGEMA_signal_12138 ;
    wire new_AGEMA_signal_12139 ;
    wire new_AGEMA_signal_12140 ;
    wire new_AGEMA_signal_12141 ;
    wire new_AGEMA_signal_12142 ;
    wire new_AGEMA_signal_12143 ;
    wire new_AGEMA_signal_12144 ;
    wire new_AGEMA_signal_12145 ;
    wire new_AGEMA_signal_12146 ;
    wire new_AGEMA_signal_12147 ;
    wire new_AGEMA_signal_12148 ;
    wire new_AGEMA_signal_12149 ;
    wire new_AGEMA_signal_12150 ;
    wire new_AGEMA_signal_12151 ;
    wire new_AGEMA_signal_12152 ;
    wire new_AGEMA_signal_12153 ;
    wire new_AGEMA_signal_12154 ;
    wire new_AGEMA_signal_12155 ;
    wire new_AGEMA_signal_12156 ;
    wire new_AGEMA_signal_12157 ;
    wire new_AGEMA_signal_12158 ;
    wire new_AGEMA_signal_12159 ;
    wire new_AGEMA_signal_12160 ;
    wire new_AGEMA_signal_12161 ;
    wire new_AGEMA_signal_12162 ;
    wire new_AGEMA_signal_12163 ;
    wire new_AGEMA_signal_12164 ;
    wire new_AGEMA_signal_12165 ;
    wire new_AGEMA_signal_12166 ;
    wire new_AGEMA_signal_12167 ;
    wire new_AGEMA_signal_12168 ;
    wire new_AGEMA_signal_12169 ;
    wire new_AGEMA_signal_12170 ;
    wire new_AGEMA_signal_12171 ;
    wire new_AGEMA_signal_12172 ;
    wire new_AGEMA_signal_12173 ;
    wire new_AGEMA_signal_12174 ;
    wire new_AGEMA_signal_12175 ;
    wire new_AGEMA_signal_12176 ;
    wire new_AGEMA_signal_12177 ;
    wire new_AGEMA_signal_12178 ;
    wire new_AGEMA_signal_12179 ;
    wire new_AGEMA_signal_12180 ;
    wire new_AGEMA_signal_12181 ;
    wire new_AGEMA_signal_12182 ;
    wire new_AGEMA_signal_12183 ;
    wire new_AGEMA_signal_12184 ;
    wire new_AGEMA_signal_12185 ;
    wire new_AGEMA_signal_12186 ;
    wire new_AGEMA_signal_12187 ;
    wire new_AGEMA_signal_12188 ;
    wire new_AGEMA_signal_12189 ;
    wire new_AGEMA_signal_12190 ;
    wire new_AGEMA_signal_12191 ;
    wire new_AGEMA_signal_12192 ;
    wire new_AGEMA_signal_12193 ;
    wire new_AGEMA_signal_12194 ;
    wire new_AGEMA_signal_12195 ;
    wire new_AGEMA_signal_12196 ;
    wire new_AGEMA_signal_12197 ;
    wire new_AGEMA_signal_12198 ;
    wire new_AGEMA_signal_12199 ;
    wire new_AGEMA_signal_12200 ;
    wire new_AGEMA_signal_12201 ;
    wire new_AGEMA_signal_12202 ;
    wire new_AGEMA_signal_12203 ;
    wire new_AGEMA_signal_12204 ;
    wire new_AGEMA_signal_12205 ;
    wire new_AGEMA_signal_12206 ;
    wire new_AGEMA_signal_12207 ;
    wire new_AGEMA_signal_12208 ;
    wire new_AGEMA_signal_12209 ;
    wire new_AGEMA_signal_12210 ;
    wire new_AGEMA_signal_12211 ;
    wire new_AGEMA_signal_12212 ;
    wire new_AGEMA_signal_12213 ;
    wire new_AGEMA_signal_12214 ;
    wire new_AGEMA_signal_12215 ;
    wire new_AGEMA_signal_12216 ;
    wire new_AGEMA_signal_12217 ;
    wire new_AGEMA_signal_12218 ;
    wire new_AGEMA_signal_12219 ;
    wire new_AGEMA_signal_12220 ;
    wire new_AGEMA_signal_12221 ;
    wire new_AGEMA_signal_12222 ;
    wire new_AGEMA_signal_12223 ;
    wire new_AGEMA_signal_12224 ;
    wire new_AGEMA_signal_12225 ;
    wire new_AGEMA_signal_12226 ;
    wire new_AGEMA_signal_12227 ;
    wire new_AGEMA_signal_12228 ;
    wire new_AGEMA_signal_12229 ;
    wire new_AGEMA_signal_12230 ;
    wire new_AGEMA_signal_12231 ;
    wire new_AGEMA_signal_12232 ;
    wire new_AGEMA_signal_12233 ;
    wire new_AGEMA_signal_12234 ;
    wire new_AGEMA_signal_12235 ;
    wire new_AGEMA_signal_12236 ;
    wire new_AGEMA_signal_12237 ;
    wire new_AGEMA_signal_12238 ;
    wire new_AGEMA_signal_12239 ;
    wire new_AGEMA_signal_12240 ;
    wire new_AGEMA_signal_12241 ;
    wire new_AGEMA_signal_12242 ;
    wire new_AGEMA_signal_12243 ;
    wire new_AGEMA_signal_12244 ;
    wire new_AGEMA_signal_12245 ;
    wire new_AGEMA_signal_12246 ;
    wire new_AGEMA_signal_12247 ;
    wire new_AGEMA_signal_12248 ;
    wire new_AGEMA_signal_12249 ;
    wire new_AGEMA_signal_12250 ;
    wire new_AGEMA_signal_12251 ;
    wire new_AGEMA_signal_12252 ;
    wire new_AGEMA_signal_12253 ;
    wire new_AGEMA_signal_12254 ;
    wire new_AGEMA_signal_12255 ;
    wire new_AGEMA_signal_12256 ;
    wire new_AGEMA_signal_12257 ;
    wire new_AGEMA_signal_12258 ;
    wire new_AGEMA_signal_12259 ;
    wire new_AGEMA_signal_12260 ;
    wire new_AGEMA_signal_12261 ;
    wire new_AGEMA_signal_12262 ;
    wire new_AGEMA_signal_12263 ;
    wire new_AGEMA_signal_12264 ;
    wire new_AGEMA_signal_12265 ;
    wire new_AGEMA_signal_12266 ;
    wire new_AGEMA_signal_12267 ;
    wire new_AGEMA_signal_12268 ;
    wire new_AGEMA_signal_12269 ;
    wire new_AGEMA_signal_12270 ;
    wire new_AGEMA_signal_12271 ;
    wire new_AGEMA_signal_12272 ;
    wire new_AGEMA_signal_12273 ;
    wire new_AGEMA_signal_12274 ;
    wire new_AGEMA_signal_12275 ;
    wire new_AGEMA_signal_12276 ;
    wire new_AGEMA_signal_12277 ;
    wire new_AGEMA_signal_12278 ;
    wire new_AGEMA_signal_12279 ;
    wire new_AGEMA_signal_12280 ;
    wire new_AGEMA_signal_12281 ;
    wire new_AGEMA_signal_12282 ;
    wire new_AGEMA_signal_12283 ;
    wire new_AGEMA_signal_12284 ;
    wire new_AGEMA_signal_12285 ;
    wire new_AGEMA_signal_12286 ;
    wire new_AGEMA_signal_12287 ;
    wire new_AGEMA_signal_12288 ;
    wire new_AGEMA_signal_12289 ;
    wire new_AGEMA_signal_12290 ;
    wire new_AGEMA_signal_12291 ;
    wire new_AGEMA_signal_12292 ;
    wire new_AGEMA_signal_12293 ;
    wire new_AGEMA_signal_12294 ;
    wire new_AGEMA_signal_12295 ;
    wire new_AGEMA_signal_12296 ;
    wire new_AGEMA_signal_12297 ;
    wire new_AGEMA_signal_12298 ;
    wire new_AGEMA_signal_12299 ;
    wire new_AGEMA_signal_12300 ;
    wire new_AGEMA_signal_12301 ;
    wire new_AGEMA_signal_12302 ;
    wire new_AGEMA_signal_12303 ;
    wire new_AGEMA_signal_12304 ;
    wire new_AGEMA_signal_12305 ;
    wire new_AGEMA_signal_12306 ;
    wire new_AGEMA_signal_12307 ;
    wire new_AGEMA_signal_12308 ;
    wire new_AGEMA_signal_12309 ;
    wire new_AGEMA_signal_12310 ;
    wire new_AGEMA_signal_12311 ;
    wire new_AGEMA_signal_12312 ;
    wire new_AGEMA_signal_12313 ;
    wire new_AGEMA_signal_12314 ;
    wire new_AGEMA_signal_12315 ;
    wire new_AGEMA_signal_12316 ;
    wire new_AGEMA_signal_12317 ;
    wire new_AGEMA_signal_12318 ;
    wire new_AGEMA_signal_12319 ;
    wire new_AGEMA_signal_12320 ;
    wire new_AGEMA_signal_12321 ;
    wire new_AGEMA_signal_12322 ;
    wire new_AGEMA_signal_12323 ;
    wire new_AGEMA_signal_12324 ;
    wire new_AGEMA_signal_12325 ;
    wire new_AGEMA_signal_12326 ;
    wire new_AGEMA_signal_12327 ;
    wire new_AGEMA_signal_12328 ;
    wire new_AGEMA_signal_12329 ;
    wire new_AGEMA_signal_12330 ;
    wire new_AGEMA_signal_12331 ;
    wire new_AGEMA_signal_12332 ;
    wire new_AGEMA_signal_12333 ;
    wire new_AGEMA_signal_12334 ;
    wire new_AGEMA_signal_12335 ;
    wire new_AGEMA_signal_12336 ;
    wire new_AGEMA_signal_12337 ;
    wire new_AGEMA_signal_12338 ;
    wire new_AGEMA_signal_12339 ;
    wire new_AGEMA_signal_12340 ;
    wire new_AGEMA_signal_12341 ;
    wire new_AGEMA_signal_12342 ;
    wire new_AGEMA_signal_12343 ;
    wire new_AGEMA_signal_12344 ;
    wire new_AGEMA_signal_12345 ;
    wire new_AGEMA_signal_12346 ;
    wire new_AGEMA_signal_12347 ;
    wire new_AGEMA_signal_12348 ;
    wire new_AGEMA_signal_12349 ;
    wire new_AGEMA_signal_12350 ;
    wire new_AGEMA_signal_12351 ;
    wire new_AGEMA_signal_12352 ;
    wire new_AGEMA_signal_12353 ;
    wire new_AGEMA_signal_12354 ;
    wire new_AGEMA_signal_12355 ;
    wire new_AGEMA_signal_12356 ;
    wire new_AGEMA_signal_12357 ;
    wire new_AGEMA_signal_12358 ;
    wire new_AGEMA_signal_12359 ;
    wire new_AGEMA_signal_12360 ;
    wire new_AGEMA_signal_12361 ;
    wire new_AGEMA_signal_12362 ;
    wire new_AGEMA_signal_12363 ;
    wire new_AGEMA_signal_12364 ;
    wire new_AGEMA_signal_12365 ;
    wire new_AGEMA_signal_12366 ;
    wire new_AGEMA_signal_12367 ;
    wire new_AGEMA_signal_12368 ;
    wire new_AGEMA_signal_12369 ;
    wire new_AGEMA_signal_12370 ;
    wire new_AGEMA_signal_12371 ;
    wire new_AGEMA_signal_12372 ;
    wire new_AGEMA_signal_12373 ;
    wire new_AGEMA_signal_12374 ;
    wire new_AGEMA_signal_12375 ;
    wire new_AGEMA_signal_12376 ;
    wire new_AGEMA_signal_12377 ;
    wire new_AGEMA_signal_12378 ;
    wire new_AGEMA_signal_12379 ;
    wire new_AGEMA_signal_12380 ;
    wire new_AGEMA_signal_12381 ;
    wire new_AGEMA_signal_12382 ;
    wire new_AGEMA_signal_12383 ;
    wire new_AGEMA_signal_12384 ;
    wire new_AGEMA_signal_12385 ;
    wire new_AGEMA_signal_12386 ;
    wire new_AGEMA_signal_12387 ;
    wire new_AGEMA_signal_12388 ;
    wire new_AGEMA_signal_12389 ;
    wire new_AGEMA_signal_12390 ;
    wire new_AGEMA_signal_12391 ;
    wire new_AGEMA_signal_12392 ;
    wire new_AGEMA_signal_12393 ;
    wire new_AGEMA_signal_12394 ;
    wire new_AGEMA_signal_12395 ;
    wire new_AGEMA_signal_12396 ;
    wire new_AGEMA_signal_12397 ;
    wire new_AGEMA_signal_12398 ;
    wire new_AGEMA_signal_12399 ;
    wire new_AGEMA_signal_12400 ;
    wire new_AGEMA_signal_12401 ;
    wire new_AGEMA_signal_12402 ;
    wire new_AGEMA_signal_12403 ;
    wire new_AGEMA_signal_12404 ;
    wire new_AGEMA_signal_12405 ;
    wire new_AGEMA_signal_12406 ;
    wire new_AGEMA_signal_12407 ;
    wire new_AGEMA_signal_12408 ;
    wire new_AGEMA_signal_12409 ;
    wire new_AGEMA_signal_12410 ;
    wire new_AGEMA_signal_12411 ;
    wire new_AGEMA_signal_12412 ;
    wire new_AGEMA_signal_12413 ;
    wire new_AGEMA_signal_12414 ;
    wire new_AGEMA_signal_12415 ;
    wire new_AGEMA_signal_12416 ;
    wire new_AGEMA_signal_12417 ;
    wire new_AGEMA_signal_12418 ;
    wire new_AGEMA_signal_12419 ;
    wire new_AGEMA_signal_12420 ;
    wire new_AGEMA_signal_12421 ;
    wire new_AGEMA_signal_12422 ;
    wire new_AGEMA_signal_12423 ;
    wire new_AGEMA_signal_12424 ;
    wire new_AGEMA_signal_12425 ;
    wire new_AGEMA_signal_12426 ;
    wire new_AGEMA_signal_12427 ;
    wire new_AGEMA_signal_12428 ;
    wire new_AGEMA_signal_12429 ;
    wire new_AGEMA_signal_12430 ;
    wire new_AGEMA_signal_12431 ;
    wire new_AGEMA_signal_12432 ;
    wire new_AGEMA_signal_12433 ;
    wire new_AGEMA_signal_12434 ;
    wire new_AGEMA_signal_12435 ;
    wire new_AGEMA_signal_12436 ;
    wire new_AGEMA_signal_12437 ;
    wire new_AGEMA_signal_12438 ;
    wire new_AGEMA_signal_12439 ;
    wire new_AGEMA_signal_12440 ;
    wire new_AGEMA_signal_12441 ;
    wire new_AGEMA_signal_12442 ;
    wire new_AGEMA_signal_12443 ;
    wire new_AGEMA_signal_12444 ;
    wire new_AGEMA_signal_12445 ;
    wire new_AGEMA_signal_12446 ;
    wire new_AGEMA_signal_12447 ;
    wire new_AGEMA_signal_12448 ;
    wire new_AGEMA_signal_12449 ;
    wire new_AGEMA_signal_12450 ;
    wire new_AGEMA_signal_12451 ;
    wire new_AGEMA_signal_12452 ;
    wire new_AGEMA_signal_12453 ;
    wire new_AGEMA_signal_12454 ;
    wire new_AGEMA_signal_12455 ;
    wire new_AGEMA_signal_12456 ;
    wire new_AGEMA_signal_12457 ;
    wire new_AGEMA_signal_12458 ;
    wire new_AGEMA_signal_12459 ;
    wire new_AGEMA_signal_12460 ;
    wire new_AGEMA_signal_12461 ;
    wire new_AGEMA_signal_12462 ;
    wire new_AGEMA_signal_12463 ;
    wire new_AGEMA_signal_12464 ;
    wire new_AGEMA_signal_12465 ;
    wire new_AGEMA_signal_12466 ;
    wire new_AGEMA_signal_12467 ;
    wire new_AGEMA_signal_12468 ;
    wire new_AGEMA_signal_12469 ;
    wire new_AGEMA_signal_12470 ;
    wire new_AGEMA_signal_12471 ;
    wire new_AGEMA_signal_12472 ;
    wire new_AGEMA_signal_12473 ;
    wire new_AGEMA_signal_12474 ;
    wire new_AGEMA_signal_12475 ;
    wire new_AGEMA_signal_12476 ;
    wire new_AGEMA_signal_12477 ;
    wire new_AGEMA_signal_12478 ;
    wire new_AGEMA_signal_12479 ;
    wire new_AGEMA_signal_12480 ;
    wire new_AGEMA_signal_12481 ;
    wire new_AGEMA_signal_12482 ;
    wire new_AGEMA_signal_12483 ;
    wire new_AGEMA_signal_12484 ;
    wire new_AGEMA_signal_12485 ;
    wire new_AGEMA_signal_12486 ;
    wire new_AGEMA_signal_12487 ;
    wire new_AGEMA_signal_12488 ;
    wire new_AGEMA_signal_12489 ;
    wire new_AGEMA_signal_12490 ;
    wire new_AGEMA_signal_12491 ;
    wire new_AGEMA_signal_12492 ;
    wire new_AGEMA_signal_12493 ;
    wire new_AGEMA_signal_12494 ;
    wire new_AGEMA_signal_12495 ;
    wire new_AGEMA_signal_12496 ;
    wire new_AGEMA_signal_12497 ;
    wire new_AGEMA_signal_12498 ;
    wire new_AGEMA_signal_12499 ;
    wire new_AGEMA_signal_12500 ;
    wire new_AGEMA_signal_12501 ;
    wire new_AGEMA_signal_12502 ;
    wire new_AGEMA_signal_12503 ;
    wire new_AGEMA_signal_12504 ;
    wire new_AGEMA_signal_12505 ;
    wire new_AGEMA_signal_12506 ;
    wire new_AGEMA_signal_12507 ;
    wire new_AGEMA_signal_12508 ;
    wire new_AGEMA_signal_12509 ;
    wire new_AGEMA_signal_12510 ;
    wire new_AGEMA_signal_12511 ;
    wire new_AGEMA_signal_12512 ;
    wire new_AGEMA_signal_12513 ;
    wire new_AGEMA_signal_12514 ;
    wire new_AGEMA_signal_12515 ;
    wire new_AGEMA_signal_12516 ;
    wire new_AGEMA_signal_12517 ;
    wire new_AGEMA_signal_12518 ;
    wire new_AGEMA_signal_12519 ;
    wire new_AGEMA_signal_12520 ;
    wire new_AGEMA_signal_12521 ;
    wire new_AGEMA_signal_12522 ;
    wire new_AGEMA_signal_12523 ;
    wire new_AGEMA_signal_12524 ;
    wire new_AGEMA_signal_12525 ;
    wire new_AGEMA_signal_12526 ;
    wire new_AGEMA_signal_12527 ;
    wire new_AGEMA_signal_12528 ;
    wire new_AGEMA_signal_12529 ;
    wire new_AGEMA_signal_12530 ;
    wire new_AGEMA_signal_12531 ;
    wire new_AGEMA_signal_12532 ;
    wire new_AGEMA_signal_12533 ;
    wire new_AGEMA_signal_12534 ;
    wire new_AGEMA_signal_12535 ;
    wire new_AGEMA_signal_12536 ;
    wire new_AGEMA_signal_12537 ;
    wire new_AGEMA_signal_12538 ;
    wire new_AGEMA_signal_12539 ;
    wire new_AGEMA_signal_12540 ;
    wire new_AGEMA_signal_12541 ;
    wire new_AGEMA_signal_12542 ;
    wire new_AGEMA_signal_12543 ;
    wire new_AGEMA_signal_12544 ;
    wire new_AGEMA_signal_12545 ;
    wire new_AGEMA_signal_12546 ;
    wire new_AGEMA_signal_12547 ;
    wire new_AGEMA_signal_12548 ;
    wire new_AGEMA_signal_12549 ;
    wire new_AGEMA_signal_12550 ;
    wire new_AGEMA_signal_12551 ;
    wire new_AGEMA_signal_12552 ;
    wire new_AGEMA_signal_12553 ;
    wire new_AGEMA_signal_12554 ;
    wire new_AGEMA_signal_12555 ;
    wire new_AGEMA_signal_12556 ;
    wire new_AGEMA_signal_12557 ;
    wire new_AGEMA_signal_12558 ;
    wire new_AGEMA_signal_12559 ;
    wire new_AGEMA_signal_12560 ;
    wire new_AGEMA_signal_12561 ;
    wire new_AGEMA_signal_12562 ;
    wire new_AGEMA_signal_12563 ;
    wire new_AGEMA_signal_12564 ;
    wire new_AGEMA_signal_12565 ;
    wire new_AGEMA_signal_12566 ;
    wire new_AGEMA_signal_12567 ;
    wire new_AGEMA_signal_12568 ;
    wire new_AGEMA_signal_12569 ;
    wire new_AGEMA_signal_12570 ;
    wire new_AGEMA_signal_12571 ;
    wire new_AGEMA_signal_12572 ;
    wire new_AGEMA_signal_12573 ;
    wire new_AGEMA_signal_12574 ;
    wire new_AGEMA_signal_12575 ;
    wire new_AGEMA_signal_12576 ;
    wire new_AGEMA_signal_12577 ;
    wire new_AGEMA_signal_12578 ;
    wire new_AGEMA_signal_12579 ;
    wire new_AGEMA_signal_12580 ;
    wire new_AGEMA_signal_12581 ;
    wire new_AGEMA_signal_12582 ;
    wire new_AGEMA_signal_12583 ;
    wire new_AGEMA_signal_12584 ;
    wire new_AGEMA_signal_12585 ;
    wire new_AGEMA_signal_12586 ;
    wire new_AGEMA_signal_12587 ;
    wire new_AGEMA_signal_12588 ;
    wire new_AGEMA_signal_12589 ;
    wire new_AGEMA_signal_12590 ;
    wire new_AGEMA_signal_12591 ;
    wire new_AGEMA_signal_12592 ;
    wire new_AGEMA_signal_12593 ;
    wire new_AGEMA_signal_12594 ;
    wire new_AGEMA_signal_12595 ;
    wire new_AGEMA_signal_12596 ;
    wire new_AGEMA_signal_12597 ;
    wire new_AGEMA_signal_12598 ;
    wire new_AGEMA_signal_12599 ;
    wire new_AGEMA_signal_12600 ;
    wire new_AGEMA_signal_12601 ;
    wire new_AGEMA_signal_12602 ;
    wire new_AGEMA_signal_12603 ;
    wire new_AGEMA_signal_12604 ;
    wire new_AGEMA_signal_12605 ;
    wire new_AGEMA_signal_12606 ;
    wire new_AGEMA_signal_12607 ;
    wire new_AGEMA_signal_12608 ;
    wire new_AGEMA_signal_12609 ;
    wire new_AGEMA_signal_12610 ;
    wire new_AGEMA_signal_12611 ;
    wire new_AGEMA_signal_12612 ;
    wire new_AGEMA_signal_12613 ;
    wire new_AGEMA_signal_12614 ;
    wire new_AGEMA_signal_12615 ;
    wire new_AGEMA_signal_12616 ;
    wire new_AGEMA_signal_12617 ;
    wire new_AGEMA_signal_12618 ;
    wire new_AGEMA_signal_12619 ;
    wire new_AGEMA_signal_12620 ;
    wire new_AGEMA_signal_12621 ;
    wire new_AGEMA_signal_12622 ;
    wire new_AGEMA_signal_12623 ;
    wire new_AGEMA_signal_12624 ;
    wire new_AGEMA_signal_12625 ;
    wire new_AGEMA_signal_12626 ;
    wire new_AGEMA_signal_12627 ;
    wire new_AGEMA_signal_12628 ;
    wire new_AGEMA_signal_12629 ;
    wire new_AGEMA_signal_12630 ;
    wire new_AGEMA_signal_12631 ;
    wire new_AGEMA_signal_12632 ;
    wire new_AGEMA_signal_12633 ;
    wire new_AGEMA_signal_12634 ;
    wire new_AGEMA_signal_12635 ;
    wire new_AGEMA_signal_12636 ;
    wire new_AGEMA_signal_12637 ;
    wire new_AGEMA_signal_12638 ;
    wire new_AGEMA_signal_12639 ;
    wire new_AGEMA_signal_12640 ;
    wire new_AGEMA_signal_12641 ;
    wire new_AGEMA_signal_12642 ;
    wire new_AGEMA_signal_12643 ;
    wire new_AGEMA_signal_12644 ;
    wire new_AGEMA_signal_12645 ;
    wire new_AGEMA_signal_12646 ;
    wire new_AGEMA_signal_12647 ;
    wire new_AGEMA_signal_12648 ;
    wire new_AGEMA_signal_12649 ;
    wire new_AGEMA_signal_12650 ;
    wire new_AGEMA_signal_12651 ;
    wire new_AGEMA_signal_12652 ;
    wire new_AGEMA_signal_12653 ;
    wire new_AGEMA_signal_12654 ;
    wire new_AGEMA_signal_12655 ;
    wire new_AGEMA_signal_12656 ;
    wire new_AGEMA_signal_12657 ;
    wire new_AGEMA_signal_12658 ;
    wire new_AGEMA_signal_12659 ;
    wire new_AGEMA_signal_12660 ;
    wire new_AGEMA_signal_12661 ;
    wire new_AGEMA_signal_12662 ;
    wire new_AGEMA_signal_12663 ;
    wire new_AGEMA_signal_12664 ;
    wire new_AGEMA_signal_12665 ;
    wire new_AGEMA_signal_12666 ;
    wire new_AGEMA_signal_12667 ;
    wire new_AGEMA_signal_12668 ;
    wire new_AGEMA_signal_12669 ;
    wire new_AGEMA_signal_12670 ;
    wire new_AGEMA_signal_12671 ;
    wire new_AGEMA_signal_12672 ;
    wire new_AGEMA_signal_12673 ;
    wire new_AGEMA_signal_12674 ;
    wire new_AGEMA_signal_12675 ;
    wire new_AGEMA_signal_12676 ;
    wire new_AGEMA_signal_12677 ;
    wire new_AGEMA_signal_12678 ;
    wire new_AGEMA_signal_12679 ;
    wire new_AGEMA_signal_12680 ;
    wire new_AGEMA_signal_12681 ;
    wire new_AGEMA_signal_12682 ;
    wire new_AGEMA_signal_12683 ;
    wire new_AGEMA_signal_12684 ;
    wire new_AGEMA_signal_12685 ;
    wire new_AGEMA_signal_12686 ;
    wire new_AGEMA_signal_12687 ;
    wire new_AGEMA_signal_12688 ;
    wire new_AGEMA_signal_12689 ;
    wire new_AGEMA_signal_12690 ;
    wire new_AGEMA_signal_12691 ;
    wire new_AGEMA_signal_12692 ;
    wire new_AGEMA_signal_12693 ;
    wire new_AGEMA_signal_12694 ;
    wire new_AGEMA_signal_12695 ;
    wire new_AGEMA_signal_12696 ;
    wire new_AGEMA_signal_12697 ;
    wire new_AGEMA_signal_12698 ;
    wire new_AGEMA_signal_12699 ;
    wire new_AGEMA_signal_12700 ;
    wire new_AGEMA_signal_12701 ;
    wire new_AGEMA_signal_12702 ;
    wire new_AGEMA_signal_12703 ;
    wire new_AGEMA_signal_12704 ;
    wire new_AGEMA_signal_12705 ;
    wire new_AGEMA_signal_12706 ;
    wire new_AGEMA_signal_12707 ;
    wire new_AGEMA_signal_12708 ;
    wire new_AGEMA_signal_12709 ;
    wire new_AGEMA_signal_12710 ;
    wire new_AGEMA_signal_12711 ;
    wire new_AGEMA_signal_12712 ;
    wire new_AGEMA_signal_12713 ;
    wire new_AGEMA_signal_12714 ;
    wire new_AGEMA_signal_12715 ;
    wire new_AGEMA_signal_12716 ;
    wire new_AGEMA_signal_12717 ;
    wire new_AGEMA_signal_12718 ;
    wire new_AGEMA_signal_12719 ;
    wire new_AGEMA_signal_12720 ;
    wire new_AGEMA_signal_12721 ;
    wire new_AGEMA_signal_12722 ;
    wire new_AGEMA_signal_12723 ;
    wire new_AGEMA_signal_12724 ;
    wire new_AGEMA_signal_12725 ;
    wire new_AGEMA_signal_12726 ;
    wire new_AGEMA_signal_12727 ;
    wire new_AGEMA_signal_12728 ;
    wire new_AGEMA_signal_12729 ;
    wire new_AGEMA_signal_12730 ;
    wire new_AGEMA_signal_12731 ;
    wire new_AGEMA_signal_12732 ;
    wire new_AGEMA_signal_12733 ;
    wire new_AGEMA_signal_12734 ;
    wire new_AGEMA_signal_12735 ;
    wire new_AGEMA_signal_12736 ;
    wire new_AGEMA_signal_12737 ;
    wire new_AGEMA_signal_12738 ;
    wire new_AGEMA_signal_12739 ;
    wire new_AGEMA_signal_12740 ;
    wire new_AGEMA_signal_12741 ;
    wire new_AGEMA_signal_12742 ;
    wire new_AGEMA_signal_12743 ;
    wire new_AGEMA_signal_12744 ;
    wire new_AGEMA_signal_12745 ;
    wire new_AGEMA_signal_12746 ;
    wire new_AGEMA_signal_12747 ;
    wire new_AGEMA_signal_12748 ;
    wire new_AGEMA_signal_12749 ;
    wire new_AGEMA_signal_12750 ;
    wire new_AGEMA_signal_12751 ;
    wire new_AGEMA_signal_12752 ;
    wire new_AGEMA_signal_12753 ;
    wire new_AGEMA_signal_12754 ;
    wire new_AGEMA_signal_12755 ;
    wire new_AGEMA_signal_12756 ;
    wire new_AGEMA_signal_12757 ;
    wire new_AGEMA_signal_12758 ;
    wire new_AGEMA_signal_12759 ;
    wire new_AGEMA_signal_12760 ;
    wire new_AGEMA_signal_12761 ;
    wire new_AGEMA_signal_12762 ;
    wire new_AGEMA_signal_12763 ;
    wire new_AGEMA_signal_12764 ;
    wire new_AGEMA_signal_12765 ;
    wire new_AGEMA_signal_12766 ;
    wire new_AGEMA_signal_12767 ;
    wire new_AGEMA_signal_12768 ;
    wire new_AGEMA_signal_12769 ;
    wire new_AGEMA_signal_12770 ;
    wire new_AGEMA_signal_12771 ;
    wire new_AGEMA_signal_12772 ;
    wire new_AGEMA_signal_12773 ;
    wire new_AGEMA_signal_12774 ;
    wire new_AGEMA_signal_12775 ;
    wire new_AGEMA_signal_12776 ;
    wire new_AGEMA_signal_12777 ;
    wire new_AGEMA_signal_12778 ;
    wire new_AGEMA_signal_12779 ;
    wire new_AGEMA_signal_12780 ;
    wire new_AGEMA_signal_12781 ;
    wire new_AGEMA_signal_12782 ;
    wire new_AGEMA_signal_12783 ;
    wire new_AGEMA_signal_12784 ;
    wire new_AGEMA_signal_12785 ;
    wire new_AGEMA_signal_12786 ;
    wire new_AGEMA_signal_12787 ;
    wire new_AGEMA_signal_12788 ;
    wire new_AGEMA_signal_12789 ;
    wire new_AGEMA_signal_12790 ;
    wire new_AGEMA_signal_12791 ;
    wire new_AGEMA_signal_12792 ;
    wire new_AGEMA_signal_12793 ;
    wire new_AGEMA_signal_12794 ;
    wire new_AGEMA_signal_12795 ;
    wire new_AGEMA_signal_12796 ;
    wire new_AGEMA_signal_12797 ;
    wire new_AGEMA_signal_12798 ;
    wire new_AGEMA_signal_12799 ;
    wire new_AGEMA_signal_12800 ;
    wire new_AGEMA_signal_12801 ;
    wire new_AGEMA_signal_12802 ;
    wire new_AGEMA_signal_12803 ;
    wire new_AGEMA_signal_12804 ;
    wire new_AGEMA_signal_12805 ;
    wire new_AGEMA_signal_12806 ;
    wire new_AGEMA_signal_12807 ;
    wire new_AGEMA_signal_12808 ;
    wire new_AGEMA_signal_12809 ;
    wire new_AGEMA_signal_12810 ;
    wire new_AGEMA_signal_12811 ;
    wire new_AGEMA_signal_12812 ;
    wire new_AGEMA_signal_12813 ;
    wire new_AGEMA_signal_12814 ;
    wire new_AGEMA_signal_12815 ;
    wire new_AGEMA_signal_12816 ;
    wire new_AGEMA_signal_12817 ;
    wire new_AGEMA_signal_12818 ;
    wire new_AGEMA_signal_12819 ;
    wire new_AGEMA_signal_12820 ;
    wire new_AGEMA_signal_12821 ;
    wire new_AGEMA_signal_12822 ;
    wire new_AGEMA_signal_12823 ;
    wire new_AGEMA_signal_12824 ;
    wire new_AGEMA_signal_12825 ;
    wire new_AGEMA_signal_12826 ;
    wire new_AGEMA_signal_12827 ;
    wire new_AGEMA_signal_12828 ;
    wire new_AGEMA_signal_12829 ;
    wire new_AGEMA_signal_12830 ;
    wire new_AGEMA_signal_12831 ;
    wire new_AGEMA_signal_12832 ;
    wire new_AGEMA_signal_12833 ;
    wire new_AGEMA_signal_12834 ;
    wire new_AGEMA_signal_12835 ;
    wire new_AGEMA_signal_12836 ;
    wire new_AGEMA_signal_12837 ;
    wire new_AGEMA_signal_12838 ;
    wire new_AGEMA_signal_12839 ;
    wire new_AGEMA_signal_12840 ;
    wire new_AGEMA_signal_12841 ;
    wire new_AGEMA_signal_12842 ;
    wire new_AGEMA_signal_12843 ;
    wire new_AGEMA_signal_12844 ;
    wire new_AGEMA_signal_12845 ;
    wire new_AGEMA_signal_12846 ;
    wire new_AGEMA_signal_12847 ;
    wire new_AGEMA_signal_12848 ;
    wire new_AGEMA_signal_12849 ;
    wire new_AGEMA_signal_12850 ;
    wire new_AGEMA_signal_12851 ;
    wire new_AGEMA_signal_12852 ;
    wire new_AGEMA_signal_12853 ;
    wire new_AGEMA_signal_12854 ;
    wire new_AGEMA_signal_12855 ;
    wire new_AGEMA_signal_12856 ;
    wire new_AGEMA_signal_12857 ;
    wire new_AGEMA_signal_12858 ;
    wire new_AGEMA_signal_12859 ;
    wire new_AGEMA_signal_12860 ;
    wire new_AGEMA_signal_12861 ;
    wire new_AGEMA_signal_12862 ;
    wire new_AGEMA_signal_12863 ;
    wire new_AGEMA_signal_12864 ;
    wire new_AGEMA_signal_12865 ;
    wire new_AGEMA_signal_12866 ;
    wire new_AGEMA_signal_12867 ;
    wire new_AGEMA_signal_12868 ;
    wire new_AGEMA_signal_12869 ;
    wire new_AGEMA_signal_12870 ;
    wire new_AGEMA_signal_12871 ;
    wire new_AGEMA_signal_12872 ;
    wire new_AGEMA_signal_12873 ;
    wire new_AGEMA_signal_12874 ;
    wire new_AGEMA_signal_12875 ;
    wire new_AGEMA_signal_12876 ;
    wire new_AGEMA_signal_12877 ;
    wire new_AGEMA_signal_12878 ;
    wire new_AGEMA_signal_12879 ;
    wire new_AGEMA_signal_12880 ;
    wire new_AGEMA_signal_12881 ;
    wire new_AGEMA_signal_12882 ;
    wire new_AGEMA_signal_12883 ;
    wire new_AGEMA_signal_12884 ;
    wire new_AGEMA_signal_12885 ;
    wire new_AGEMA_signal_12886 ;
    wire new_AGEMA_signal_12887 ;
    wire new_AGEMA_signal_12888 ;
    wire new_AGEMA_signal_12889 ;
    wire new_AGEMA_signal_12890 ;
    wire new_AGEMA_signal_12891 ;
    wire new_AGEMA_signal_12892 ;
    wire new_AGEMA_signal_12893 ;
    wire new_AGEMA_signal_12894 ;
    wire new_AGEMA_signal_12895 ;
    wire new_AGEMA_signal_12896 ;
    wire new_AGEMA_signal_12897 ;
    wire new_AGEMA_signal_12898 ;
    wire new_AGEMA_signal_12899 ;
    wire new_AGEMA_signal_12900 ;
    wire new_AGEMA_signal_12901 ;
    wire new_AGEMA_signal_12902 ;
    wire new_AGEMA_signal_12903 ;
    wire new_AGEMA_signal_12904 ;
    wire new_AGEMA_signal_12905 ;
    wire new_AGEMA_signal_12906 ;
    wire new_AGEMA_signal_12907 ;
    wire new_AGEMA_signal_12908 ;
    wire new_AGEMA_signal_12909 ;
    wire new_AGEMA_signal_12910 ;
    wire new_AGEMA_signal_12911 ;
    wire new_AGEMA_signal_12912 ;
    wire new_AGEMA_signal_12913 ;
    wire new_AGEMA_signal_12914 ;
    wire new_AGEMA_signal_12915 ;
    wire new_AGEMA_signal_12916 ;
    wire new_AGEMA_signal_12917 ;
    wire new_AGEMA_signal_12918 ;
    wire new_AGEMA_signal_12919 ;
    wire new_AGEMA_signal_12920 ;
    wire new_AGEMA_signal_12921 ;
    wire new_AGEMA_signal_12922 ;
    wire new_AGEMA_signal_12923 ;
    wire new_AGEMA_signal_12924 ;
    wire new_AGEMA_signal_12925 ;
    wire new_AGEMA_signal_12926 ;
    wire new_AGEMA_signal_12927 ;
    wire new_AGEMA_signal_12928 ;
    wire new_AGEMA_signal_12929 ;
    wire new_AGEMA_signal_12930 ;
    wire new_AGEMA_signal_12931 ;
    wire new_AGEMA_signal_12932 ;
    wire new_AGEMA_signal_12933 ;
    wire new_AGEMA_signal_12934 ;
    wire new_AGEMA_signal_12935 ;
    wire new_AGEMA_signal_12936 ;
    wire new_AGEMA_signal_12937 ;
    wire new_AGEMA_signal_12938 ;
    wire new_AGEMA_signal_12939 ;
    wire new_AGEMA_signal_12940 ;
    wire new_AGEMA_signal_12941 ;
    wire new_AGEMA_signal_12942 ;
    wire new_AGEMA_signal_12943 ;
    wire new_AGEMA_signal_12944 ;
    wire new_AGEMA_signal_12945 ;
    wire new_AGEMA_signal_12946 ;
    wire new_AGEMA_signal_12947 ;
    wire new_AGEMA_signal_12948 ;
    wire new_AGEMA_signal_12949 ;
    wire new_AGEMA_signal_12950 ;
    wire new_AGEMA_signal_12951 ;
    wire new_AGEMA_signal_12952 ;
    wire new_AGEMA_signal_12953 ;
    wire new_AGEMA_signal_12954 ;
    wire new_AGEMA_signal_12955 ;
    wire new_AGEMA_signal_12956 ;
    wire new_AGEMA_signal_12957 ;
    wire new_AGEMA_signal_12958 ;
    wire new_AGEMA_signal_12959 ;
    wire new_AGEMA_signal_12960 ;
    wire new_AGEMA_signal_12961 ;
    wire new_AGEMA_signal_12962 ;
    wire new_AGEMA_signal_12963 ;
    wire new_AGEMA_signal_12964 ;
    wire new_AGEMA_signal_12965 ;
    wire new_AGEMA_signal_12966 ;
    wire new_AGEMA_signal_12967 ;
    wire new_AGEMA_signal_12968 ;
    wire new_AGEMA_signal_12969 ;
    wire new_AGEMA_signal_12970 ;
    wire new_AGEMA_signal_12971 ;
    wire new_AGEMA_signal_12972 ;
    wire new_AGEMA_signal_12973 ;
    wire new_AGEMA_signal_12974 ;
    wire new_AGEMA_signal_12975 ;
    wire new_AGEMA_signal_12976 ;
    wire new_AGEMA_signal_12977 ;
    wire new_AGEMA_signal_12978 ;
    wire new_AGEMA_signal_12979 ;
    wire new_AGEMA_signal_12980 ;
    wire new_AGEMA_signal_12981 ;
    wire new_AGEMA_signal_12982 ;
    wire new_AGEMA_signal_12983 ;
    wire new_AGEMA_signal_12984 ;
    wire new_AGEMA_signal_12985 ;
    wire new_AGEMA_signal_12986 ;
    wire new_AGEMA_signal_12987 ;
    wire new_AGEMA_signal_12988 ;
    wire new_AGEMA_signal_12989 ;
    wire new_AGEMA_signal_12990 ;
    wire new_AGEMA_signal_12991 ;
    wire new_AGEMA_signal_12992 ;
    wire new_AGEMA_signal_12993 ;
    wire new_AGEMA_signal_12994 ;
    wire new_AGEMA_signal_12995 ;
    wire new_AGEMA_signal_12996 ;
    wire new_AGEMA_signal_12997 ;
    wire new_AGEMA_signal_12998 ;
    wire new_AGEMA_signal_12999 ;
    wire new_AGEMA_signal_13000 ;
    wire new_AGEMA_signal_13001 ;
    wire new_AGEMA_signal_13002 ;
    wire new_AGEMA_signal_13003 ;
    wire new_AGEMA_signal_13004 ;
    wire new_AGEMA_signal_13005 ;
    wire new_AGEMA_signal_13006 ;
    wire new_AGEMA_signal_13007 ;
    wire new_AGEMA_signal_13008 ;
    wire new_AGEMA_signal_13009 ;
    wire new_AGEMA_signal_13010 ;
    wire new_AGEMA_signal_13011 ;
    wire new_AGEMA_signal_13012 ;
    wire new_AGEMA_signal_13013 ;
    wire new_AGEMA_signal_13014 ;
    wire new_AGEMA_signal_13015 ;
    wire new_AGEMA_signal_13016 ;
    wire new_AGEMA_signal_13017 ;
    wire new_AGEMA_signal_13018 ;
    wire new_AGEMA_signal_13019 ;
    wire new_AGEMA_signal_13020 ;
    wire new_AGEMA_signal_13021 ;
    wire new_AGEMA_signal_13022 ;
    wire new_AGEMA_signal_13023 ;
    wire new_AGEMA_signal_13024 ;
    wire new_AGEMA_signal_13025 ;
    wire new_AGEMA_signal_13026 ;
    wire new_AGEMA_signal_13027 ;
    wire new_AGEMA_signal_13028 ;
    wire new_AGEMA_signal_13029 ;
    wire new_AGEMA_signal_13030 ;
    wire new_AGEMA_signal_13031 ;
    wire new_AGEMA_signal_13032 ;
    wire new_AGEMA_signal_13033 ;
    wire new_AGEMA_signal_13034 ;
    wire new_AGEMA_signal_13035 ;
    wire new_AGEMA_signal_13036 ;
    wire new_AGEMA_signal_13037 ;
    wire new_AGEMA_signal_13038 ;
    wire new_AGEMA_signal_13039 ;
    wire new_AGEMA_signal_13040 ;
    wire new_AGEMA_signal_13041 ;
    wire new_AGEMA_signal_13042 ;
    wire new_AGEMA_signal_13043 ;
    wire new_AGEMA_signal_13044 ;
    wire new_AGEMA_signal_13045 ;
    wire new_AGEMA_signal_13046 ;
    wire new_AGEMA_signal_13047 ;
    wire new_AGEMA_signal_13048 ;
    wire new_AGEMA_signal_13049 ;
    wire new_AGEMA_signal_13050 ;
    wire new_AGEMA_signal_13051 ;
    wire new_AGEMA_signal_13052 ;
    wire new_AGEMA_signal_13053 ;
    wire new_AGEMA_signal_13054 ;
    wire new_AGEMA_signal_13055 ;
    wire new_AGEMA_signal_13056 ;
    wire new_AGEMA_signal_13057 ;
    wire new_AGEMA_signal_13058 ;
    wire new_AGEMA_signal_13059 ;
    wire new_AGEMA_signal_13060 ;
    wire new_AGEMA_signal_13061 ;
    wire new_AGEMA_signal_13062 ;
    wire new_AGEMA_signal_13063 ;
    wire new_AGEMA_signal_13064 ;
    wire new_AGEMA_signal_13065 ;
    wire new_AGEMA_signal_13066 ;
    wire new_AGEMA_signal_13067 ;
    wire new_AGEMA_signal_13068 ;
    wire new_AGEMA_signal_13069 ;
    wire new_AGEMA_signal_13070 ;
    wire new_AGEMA_signal_13071 ;
    wire new_AGEMA_signal_13072 ;
    wire new_AGEMA_signal_13073 ;
    wire new_AGEMA_signal_13074 ;
    wire new_AGEMA_signal_13075 ;
    wire new_AGEMA_signal_13076 ;
    wire new_AGEMA_signal_13077 ;
    wire new_AGEMA_signal_13078 ;
    wire new_AGEMA_signal_13079 ;
    wire new_AGEMA_signal_13080 ;
    wire new_AGEMA_signal_13081 ;
    wire new_AGEMA_signal_13082 ;
    wire new_AGEMA_signal_13083 ;
    wire new_AGEMA_signal_13084 ;
    wire new_AGEMA_signal_13085 ;
    wire new_AGEMA_signal_13086 ;
    wire new_AGEMA_signal_13087 ;
    wire new_AGEMA_signal_13088 ;
    wire new_AGEMA_signal_13089 ;
    wire new_AGEMA_signal_13090 ;
    wire new_AGEMA_signal_13091 ;
    wire new_AGEMA_signal_13092 ;
    wire new_AGEMA_signal_13093 ;
    wire new_AGEMA_signal_13094 ;
    wire new_AGEMA_signal_13095 ;
    wire new_AGEMA_signal_13096 ;
    wire new_AGEMA_signal_13097 ;
    wire new_AGEMA_signal_13098 ;
    wire new_AGEMA_signal_13099 ;
    wire new_AGEMA_signal_13100 ;
    wire new_AGEMA_signal_13101 ;
    wire new_AGEMA_signal_13102 ;
    wire new_AGEMA_signal_13103 ;
    wire new_AGEMA_signal_13104 ;
    wire new_AGEMA_signal_13105 ;
    wire new_AGEMA_signal_13106 ;
    wire new_AGEMA_signal_13107 ;
    wire new_AGEMA_signal_13108 ;
    wire new_AGEMA_signal_13109 ;
    wire new_AGEMA_signal_13110 ;
    wire new_AGEMA_signal_13111 ;
    wire new_AGEMA_signal_13112 ;
    wire new_AGEMA_signal_13113 ;
    wire new_AGEMA_signal_13114 ;
    wire new_AGEMA_signal_13115 ;
    wire new_AGEMA_signal_13116 ;
    wire new_AGEMA_signal_13117 ;
    wire new_AGEMA_signal_13118 ;
    wire new_AGEMA_signal_13119 ;
    wire new_AGEMA_signal_13120 ;
    wire new_AGEMA_signal_13121 ;
    wire new_AGEMA_signal_13122 ;
    wire new_AGEMA_signal_13123 ;
    wire new_AGEMA_signal_13124 ;
    wire new_AGEMA_signal_13125 ;
    wire new_AGEMA_signal_13126 ;
    wire new_AGEMA_signal_13127 ;
    wire new_AGEMA_signal_13128 ;
    wire new_AGEMA_signal_13129 ;
    wire new_AGEMA_signal_13130 ;
    wire new_AGEMA_signal_13131 ;
    wire new_AGEMA_signal_13132 ;
    wire new_AGEMA_signal_13133 ;
    wire new_AGEMA_signal_13134 ;
    wire new_AGEMA_signal_13135 ;
    wire new_AGEMA_signal_13136 ;
    wire new_AGEMA_signal_13137 ;
    wire new_AGEMA_signal_13138 ;
    wire new_AGEMA_signal_13139 ;
    wire new_AGEMA_signal_13140 ;
    wire new_AGEMA_signal_13141 ;
    wire new_AGEMA_signal_13142 ;
    wire new_AGEMA_signal_13143 ;
    wire new_AGEMA_signal_13144 ;
    wire new_AGEMA_signal_13145 ;
    wire new_AGEMA_signal_13146 ;
    wire new_AGEMA_signal_13147 ;
    wire new_AGEMA_signal_13148 ;
    wire new_AGEMA_signal_13149 ;
    wire new_AGEMA_signal_13150 ;
    wire new_AGEMA_signal_13151 ;
    wire new_AGEMA_signal_13152 ;
    wire new_AGEMA_signal_13153 ;
    wire new_AGEMA_signal_13154 ;
    wire new_AGEMA_signal_13155 ;
    wire new_AGEMA_signal_13156 ;
    wire new_AGEMA_signal_13157 ;
    wire new_AGEMA_signal_13158 ;
    wire new_AGEMA_signal_13159 ;
    wire new_AGEMA_signal_13160 ;
    wire new_AGEMA_signal_13161 ;
    wire new_AGEMA_signal_13162 ;
    wire new_AGEMA_signal_13163 ;
    wire new_AGEMA_signal_13164 ;
    wire new_AGEMA_signal_13165 ;
    wire new_AGEMA_signal_13166 ;
    wire new_AGEMA_signal_13167 ;
    wire new_AGEMA_signal_13168 ;
    wire new_AGEMA_signal_13169 ;
    wire new_AGEMA_signal_13170 ;
    wire new_AGEMA_signal_13171 ;
    wire new_AGEMA_signal_13172 ;
    wire new_AGEMA_signal_13173 ;
    wire new_AGEMA_signal_13174 ;
    wire new_AGEMA_signal_13175 ;
    wire new_AGEMA_signal_13176 ;
    wire new_AGEMA_signal_13177 ;
    wire new_AGEMA_signal_13178 ;
    wire new_AGEMA_signal_13179 ;
    wire new_AGEMA_signal_13180 ;
    wire new_AGEMA_signal_13181 ;
    wire new_AGEMA_signal_13182 ;
    wire new_AGEMA_signal_13183 ;
    wire new_AGEMA_signal_13184 ;
    wire new_AGEMA_signal_13185 ;
    wire new_AGEMA_signal_13186 ;
    wire new_AGEMA_signal_13187 ;
    wire new_AGEMA_signal_13188 ;
    wire new_AGEMA_signal_13189 ;
    wire new_AGEMA_signal_13190 ;
    wire new_AGEMA_signal_13191 ;
    wire new_AGEMA_signal_13192 ;
    wire new_AGEMA_signal_13193 ;
    wire new_AGEMA_signal_13194 ;
    wire new_AGEMA_signal_13195 ;
    wire new_AGEMA_signal_13196 ;
    wire new_AGEMA_signal_13197 ;
    wire new_AGEMA_signal_13198 ;
    wire new_AGEMA_signal_13199 ;
    wire new_AGEMA_signal_13200 ;
    wire new_AGEMA_signal_13201 ;
    wire new_AGEMA_signal_13202 ;
    wire new_AGEMA_signal_13203 ;
    wire new_AGEMA_signal_13204 ;
    wire new_AGEMA_signal_13205 ;
    wire new_AGEMA_signal_13206 ;
    wire new_AGEMA_signal_13207 ;
    wire new_AGEMA_signal_13208 ;
    wire new_AGEMA_signal_13209 ;
    wire new_AGEMA_signal_13210 ;
    wire new_AGEMA_signal_13211 ;
    wire new_AGEMA_signal_13212 ;
    wire new_AGEMA_signal_13213 ;
    wire new_AGEMA_signal_13214 ;
    wire new_AGEMA_signal_13215 ;
    wire new_AGEMA_signal_13216 ;
    wire new_AGEMA_signal_13217 ;
    wire new_AGEMA_signal_13218 ;
    wire new_AGEMA_signal_13219 ;
    wire new_AGEMA_signal_13220 ;
    wire new_AGEMA_signal_13221 ;
    wire new_AGEMA_signal_13222 ;
    wire new_AGEMA_signal_13223 ;
    wire new_AGEMA_signal_13224 ;
    wire new_AGEMA_signal_13225 ;
    wire new_AGEMA_signal_13226 ;
    wire new_AGEMA_signal_13227 ;
    wire new_AGEMA_signal_13228 ;
    wire new_AGEMA_signal_13229 ;
    wire new_AGEMA_signal_13230 ;
    wire new_AGEMA_signal_13231 ;
    wire new_AGEMA_signal_13232 ;
    wire new_AGEMA_signal_13233 ;
    wire new_AGEMA_signal_13234 ;
    wire new_AGEMA_signal_13235 ;
    wire new_AGEMA_signal_13236 ;
    wire new_AGEMA_signal_13237 ;
    wire new_AGEMA_signal_13238 ;
    wire new_AGEMA_signal_13239 ;
    wire new_AGEMA_signal_13240 ;
    wire new_AGEMA_signal_13241 ;
    wire new_AGEMA_signal_13242 ;
    wire new_AGEMA_signal_13243 ;
    wire new_AGEMA_signal_13244 ;
    wire new_AGEMA_signal_13245 ;
    wire new_AGEMA_signal_13246 ;
    wire new_AGEMA_signal_13247 ;
    wire new_AGEMA_signal_13248 ;
    wire new_AGEMA_signal_13249 ;
    wire new_AGEMA_signal_13250 ;
    wire new_AGEMA_signal_13251 ;
    wire new_AGEMA_signal_13252 ;
    wire new_AGEMA_signal_13253 ;
    wire new_AGEMA_signal_13254 ;
    wire new_AGEMA_signal_13255 ;
    wire new_AGEMA_signal_13256 ;
    wire new_AGEMA_signal_13257 ;
    wire new_AGEMA_signal_13258 ;
    wire new_AGEMA_signal_13259 ;
    wire new_AGEMA_signal_13260 ;
    wire new_AGEMA_signal_13261 ;
    wire new_AGEMA_signal_13262 ;
    wire new_AGEMA_signal_13263 ;
    wire new_AGEMA_signal_13264 ;
    wire new_AGEMA_signal_13265 ;
    wire new_AGEMA_signal_13266 ;
    wire new_AGEMA_signal_13267 ;
    wire new_AGEMA_signal_13268 ;
    wire new_AGEMA_signal_13269 ;
    wire new_AGEMA_signal_13270 ;
    wire new_AGEMA_signal_13271 ;
    wire new_AGEMA_signal_13272 ;
    wire new_AGEMA_signal_13273 ;
    wire new_AGEMA_signal_13274 ;
    wire new_AGEMA_signal_13275 ;
    wire new_AGEMA_signal_13276 ;
    wire new_AGEMA_signal_13277 ;
    wire new_AGEMA_signal_13278 ;
    wire new_AGEMA_signal_13279 ;
    wire new_AGEMA_signal_13280 ;
    wire new_AGEMA_signal_13281 ;
    wire new_AGEMA_signal_13282 ;
    wire new_AGEMA_signal_13283 ;
    wire new_AGEMA_signal_13284 ;
    wire new_AGEMA_signal_13285 ;
    wire new_AGEMA_signal_13286 ;
    wire new_AGEMA_signal_13287 ;
    wire new_AGEMA_signal_13288 ;
    wire new_AGEMA_signal_13289 ;
    wire new_AGEMA_signal_13290 ;
    wire new_AGEMA_signal_13291 ;
    wire new_AGEMA_signal_13292 ;
    wire new_AGEMA_signal_13293 ;
    wire new_AGEMA_signal_13294 ;
    wire new_AGEMA_signal_13295 ;
    wire new_AGEMA_signal_13296 ;
    wire new_AGEMA_signal_13297 ;
    wire new_AGEMA_signal_13298 ;
    wire new_AGEMA_signal_13299 ;
    wire new_AGEMA_signal_13300 ;
    wire new_AGEMA_signal_13301 ;
    wire new_AGEMA_signal_13302 ;
    wire new_AGEMA_signal_13303 ;
    wire new_AGEMA_signal_13304 ;
    wire new_AGEMA_signal_13305 ;
    wire new_AGEMA_signal_13306 ;
    wire new_AGEMA_signal_13307 ;
    wire new_AGEMA_signal_13308 ;
    wire new_AGEMA_signal_13309 ;
    wire new_AGEMA_signal_13310 ;
    wire new_AGEMA_signal_13311 ;
    wire new_AGEMA_signal_13312 ;
    wire new_AGEMA_signal_13313 ;
    wire new_AGEMA_signal_13314 ;
    wire new_AGEMA_signal_13315 ;
    wire new_AGEMA_signal_13316 ;
    wire new_AGEMA_signal_13317 ;
    wire new_AGEMA_signal_13318 ;
    wire new_AGEMA_signal_13319 ;
    wire new_AGEMA_signal_13320 ;
    wire new_AGEMA_signal_13321 ;
    wire new_AGEMA_signal_13322 ;
    wire new_AGEMA_signal_13323 ;
    wire new_AGEMA_signal_13324 ;
    wire new_AGEMA_signal_13325 ;
    wire new_AGEMA_signal_13326 ;
    wire new_AGEMA_signal_13327 ;
    wire new_AGEMA_signal_13328 ;
    wire new_AGEMA_signal_13329 ;
    wire new_AGEMA_signal_13330 ;
    wire new_AGEMA_signal_13331 ;
    wire new_AGEMA_signal_13332 ;
    wire new_AGEMA_signal_13333 ;
    wire new_AGEMA_signal_13334 ;
    wire new_AGEMA_signal_13335 ;
    wire new_AGEMA_signal_13336 ;
    wire new_AGEMA_signal_13337 ;
    wire new_AGEMA_signal_13338 ;
    wire new_AGEMA_signal_13339 ;
    wire new_AGEMA_signal_13340 ;
    wire new_AGEMA_signal_13341 ;
    wire new_AGEMA_signal_13342 ;
    wire new_AGEMA_signal_13343 ;
    wire new_AGEMA_signal_13344 ;
    wire new_AGEMA_signal_13345 ;
    wire new_AGEMA_signal_13346 ;
    wire new_AGEMA_signal_13347 ;
    wire new_AGEMA_signal_13348 ;
    wire new_AGEMA_signal_13349 ;
    wire new_AGEMA_signal_13350 ;
    wire new_AGEMA_signal_13351 ;
    wire new_AGEMA_signal_13352 ;
    wire new_AGEMA_signal_13353 ;
    wire new_AGEMA_signal_13354 ;
    wire new_AGEMA_signal_13355 ;
    wire new_AGEMA_signal_13356 ;
    wire new_AGEMA_signal_13357 ;
    wire new_AGEMA_signal_13358 ;
    wire new_AGEMA_signal_13359 ;
    wire new_AGEMA_signal_13360 ;
    wire new_AGEMA_signal_13361 ;
    wire new_AGEMA_signal_13362 ;
    wire new_AGEMA_signal_13363 ;
    wire new_AGEMA_signal_13364 ;
    wire new_AGEMA_signal_13365 ;
    wire new_AGEMA_signal_13366 ;
    wire new_AGEMA_signal_13367 ;
    wire new_AGEMA_signal_13368 ;
    wire new_AGEMA_signal_13369 ;
    wire new_AGEMA_signal_13370 ;
    wire new_AGEMA_signal_13371 ;
    wire new_AGEMA_signal_13372 ;
    wire new_AGEMA_signal_13373 ;
    wire new_AGEMA_signal_13374 ;
    wire new_AGEMA_signal_13375 ;
    wire new_AGEMA_signal_13376 ;
    wire new_AGEMA_signal_13377 ;
    wire new_AGEMA_signal_13378 ;
    wire new_AGEMA_signal_13379 ;
    wire new_AGEMA_signal_13380 ;
    wire new_AGEMA_signal_13381 ;
    wire new_AGEMA_signal_13382 ;
    wire new_AGEMA_signal_13383 ;
    wire new_AGEMA_signal_13384 ;
    wire new_AGEMA_signal_13385 ;
    wire new_AGEMA_signal_13386 ;
    wire new_AGEMA_signal_13387 ;
    wire new_AGEMA_signal_13388 ;
    wire new_AGEMA_signal_13389 ;
    wire new_AGEMA_signal_13390 ;
    wire new_AGEMA_signal_13391 ;
    wire new_AGEMA_signal_13392 ;
    wire new_AGEMA_signal_13393 ;
    wire new_AGEMA_signal_13394 ;
    wire new_AGEMA_signal_13395 ;
    wire new_AGEMA_signal_13396 ;
    wire new_AGEMA_signal_13397 ;
    wire new_AGEMA_signal_13398 ;
    wire new_AGEMA_signal_13399 ;
    wire new_AGEMA_signal_13400 ;
    wire new_AGEMA_signal_13401 ;
    wire new_AGEMA_signal_13402 ;
    wire new_AGEMA_signal_13403 ;
    wire new_AGEMA_signal_13404 ;
    wire new_AGEMA_signal_13405 ;
    wire new_AGEMA_signal_13406 ;
    wire new_AGEMA_signal_13407 ;
    wire new_AGEMA_signal_13408 ;
    wire new_AGEMA_signal_13409 ;
    wire new_AGEMA_signal_13410 ;
    wire new_AGEMA_signal_13411 ;
    wire new_AGEMA_signal_13412 ;
    wire new_AGEMA_signal_13413 ;
    wire new_AGEMA_signal_13414 ;
    wire new_AGEMA_signal_13415 ;
    wire new_AGEMA_signal_13416 ;
    wire new_AGEMA_signal_13417 ;
    wire new_AGEMA_signal_13418 ;
    wire new_AGEMA_signal_13419 ;
    wire new_AGEMA_signal_13420 ;
    wire new_AGEMA_signal_13421 ;
    wire new_AGEMA_signal_13422 ;
    wire new_AGEMA_signal_13423 ;
    wire new_AGEMA_signal_13424 ;
    wire new_AGEMA_signal_13425 ;
    wire new_AGEMA_signal_13426 ;
    wire new_AGEMA_signal_13427 ;
    wire new_AGEMA_signal_13428 ;
    wire new_AGEMA_signal_13429 ;
    wire new_AGEMA_signal_13430 ;
    wire new_AGEMA_signal_13431 ;
    wire new_AGEMA_signal_13432 ;
    wire new_AGEMA_signal_13433 ;
    wire new_AGEMA_signal_13434 ;
    wire new_AGEMA_signal_13435 ;
    wire new_AGEMA_signal_13436 ;
    wire new_AGEMA_signal_13437 ;
    wire new_AGEMA_signal_13438 ;
    wire new_AGEMA_signal_13439 ;
    wire new_AGEMA_signal_13440 ;
    wire new_AGEMA_signal_13441 ;
    wire new_AGEMA_signal_13442 ;
    wire new_AGEMA_signal_13443 ;
    wire new_AGEMA_signal_13444 ;
    wire new_AGEMA_signal_13445 ;
    wire new_AGEMA_signal_13446 ;
    wire new_AGEMA_signal_13447 ;
    wire new_AGEMA_signal_13448 ;
    wire new_AGEMA_signal_13449 ;
    wire new_AGEMA_signal_13450 ;
    wire new_AGEMA_signal_13451 ;
    wire new_AGEMA_signal_13452 ;
    wire new_AGEMA_signal_13453 ;
    wire new_AGEMA_signal_13454 ;
    wire new_AGEMA_signal_13455 ;
    wire new_AGEMA_signal_13456 ;
    wire new_AGEMA_signal_13457 ;
    wire new_AGEMA_signal_13458 ;
    wire new_AGEMA_signal_13459 ;
    wire new_AGEMA_signal_13460 ;
    wire new_AGEMA_signal_13461 ;
    wire new_AGEMA_signal_13462 ;
    wire new_AGEMA_signal_13463 ;
    wire new_AGEMA_signal_13464 ;
    wire new_AGEMA_signal_13465 ;
    wire new_AGEMA_signal_13466 ;
    wire new_AGEMA_signal_13467 ;
    wire new_AGEMA_signal_13468 ;
    wire new_AGEMA_signal_13469 ;
    wire new_AGEMA_signal_13470 ;
    wire new_AGEMA_signal_13471 ;
    wire new_AGEMA_signal_13472 ;
    wire new_AGEMA_signal_13473 ;
    wire new_AGEMA_signal_13474 ;
    wire new_AGEMA_signal_13475 ;
    wire new_AGEMA_signal_13476 ;
    wire new_AGEMA_signal_13477 ;
    wire new_AGEMA_signal_13478 ;
    wire new_AGEMA_signal_13479 ;
    wire new_AGEMA_signal_13480 ;
    wire new_AGEMA_signal_13481 ;
    wire new_AGEMA_signal_13482 ;
    wire new_AGEMA_signal_13483 ;
    wire new_AGEMA_signal_13484 ;
    wire new_AGEMA_signal_13485 ;
    wire new_AGEMA_signal_13486 ;
    wire new_AGEMA_signal_13487 ;
    wire new_AGEMA_signal_13488 ;
    wire new_AGEMA_signal_13489 ;
    wire new_AGEMA_signal_13490 ;
    wire new_AGEMA_signal_13491 ;
    wire new_AGEMA_signal_13492 ;
    wire new_AGEMA_signal_13493 ;
    wire new_AGEMA_signal_13494 ;
    wire new_AGEMA_signal_13495 ;
    wire new_AGEMA_signal_13496 ;
    wire new_AGEMA_signal_13497 ;
    wire new_AGEMA_signal_13498 ;
    wire new_AGEMA_signal_13499 ;
    wire new_AGEMA_signal_13500 ;
    wire new_AGEMA_signal_13501 ;
    wire new_AGEMA_signal_13502 ;
    wire new_AGEMA_signal_13503 ;
    wire new_AGEMA_signal_13504 ;
    wire new_AGEMA_signal_13505 ;
    wire new_AGEMA_signal_13506 ;
    wire new_AGEMA_signal_13507 ;
    wire new_AGEMA_signal_13508 ;
    wire new_AGEMA_signal_13509 ;
    wire new_AGEMA_signal_13510 ;
    wire new_AGEMA_signal_13511 ;
    wire new_AGEMA_signal_13512 ;
    wire new_AGEMA_signal_13513 ;
    wire new_AGEMA_signal_13514 ;
    wire new_AGEMA_signal_13515 ;
    wire new_AGEMA_signal_13516 ;
    wire new_AGEMA_signal_13517 ;
    wire new_AGEMA_signal_13518 ;
    wire new_AGEMA_signal_13519 ;
    wire new_AGEMA_signal_13520 ;
    wire new_AGEMA_signal_13521 ;
    wire new_AGEMA_signal_13522 ;
    wire new_AGEMA_signal_13523 ;
    wire new_AGEMA_signal_13524 ;
    wire new_AGEMA_signal_13525 ;
    wire new_AGEMA_signal_13526 ;
    wire new_AGEMA_signal_13527 ;
    wire new_AGEMA_signal_13528 ;
    wire new_AGEMA_signal_13529 ;
    wire new_AGEMA_signal_13530 ;
    wire new_AGEMA_signal_13531 ;
    wire new_AGEMA_signal_13532 ;
    wire new_AGEMA_signal_13533 ;
    wire new_AGEMA_signal_13534 ;
    wire new_AGEMA_signal_13535 ;
    wire new_AGEMA_signal_13536 ;
    wire new_AGEMA_signal_13537 ;
    wire new_AGEMA_signal_13538 ;
    wire new_AGEMA_signal_13539 ;
    wire new_AGEMA_signal_13540 ;
    wire new_AGEMA_signal_13541 ;
    wire new_AGEMA_signal_13542 ;
    wire new_AGEMA_signal_13543 ;
    wire new_AGEMA_signal_13544 ;
    wire new_AGEMA_signal_13545 ;
    wire new_AGEMA_signal_13546 ;
    wire new_AGEMA_signal_13547 ;
    wire new_AGEMA_signal_13548 ;
    wire new_AGEMA_signal_13549 ;
    wire new_AGEMA_signal_13550 ;
    wire new_AGEMA_signal_13551 ;
    wire new_AGEMA_signal_13552 ;
    wire new_AGEMA_signal_13553 ;
    wire new_AGEMA_signal_13554 ;
    wire new_AGEMA_signal_13555 ;
    wire new_AGEMA_signal_13556 ;
    wire new_AGEMA_signal_13557 ;
    wire new_AGEMA_signal_13558 ;
    wire new_AGEMA_signal_13559 ;
    wire new_AGEMA_signal_13560 ;
    wire new_AGEMA_signal_13561 ;
    wire new_AGEMA_signal_13562 ;
    wire new_AGEMA_signal_13563 ;
    wire new_AGEMA_signal_13564 ;
    wire new_AGEMA_signal_13565 ;
    wire new_AGEMA_signal_13566 ;
    wire new_AGEMA_signal_13567 ;
    wire new_AGEMA_signal_13568 ;
    wire new_AGEMA_signal_13569 ;
    wire new_AGEMA_signal_13570 ;
    wire new_AGEMA_signal_13571 ;
    wire new_AGEMA_signal_13572 ;
    wire new_AGEMA_signal_13573 ;
    wire new_AGEMA_signal_13574 ;
    wire new_AGEMA_signal_13575 ;
    wire new_AGEMA_signal_13576 ;
    wire new_AGEMA_signal_13577 ;
    wire new_AGEMA_signal_13578 ;
    wire new_AGEMA_signal_13579 ;
    wire new_AGEMA_signal_13580 ;
    wire new_AGEMA_signal_13581 ;
    wire new_AGEMA_signal_13582 ;
    wire new_AGEMA_signal_13583 ;
    wire new_AGEMA_signal_13584 ;
    wire new_AGEMA_signal_13585 ;
    wire new_AGEMA_signal_13586 ;
    wire new_AGEMA_signal_13587 ;
    wire new_AGEMA_signal_13588 ;
    wire new_AGEMA_signal_13589 ;
    wire new_AGEMA_signal_13590 ;
    wire new_AGEMA_signal_13591 ;
    wire new_AGEMA_signal_13592 ;
    wire new_AGEMA_signal_13593 ;
    wire new_AGEMA_signal_13594 ;
    wire new_AGEMA_signal_13595 ;
    wire new_AGEMA_signal_13596 ;
    wire new_AGEMA_signal_13597 ;
    wire new_AGEMA_signal_13598 ;
    wire new_AGEMA_signal_13599 ;
    wire new_AGEMA_signal_13600 ;
    wire new_AGEMA_signal_13601 ;
    wire new_AGEMA_signal_13602 ;
    wire new_AGEMA_signal_13603 ;
    wire new_AGEMA_signal_13604 ;
    wire new_AGEMA_signal_13605 ;
    wire new_AGEMA_signal_13606 ;
    wire new_AGEMA_signal_13607 ;
    wire new_AGEMA_signal_13608 ;
    wire new_AGEMA_signal_13609 ;
    wire new_AGEMA_signal_13610 ;
    wire new_AGEMA_signal_13611 ;
    wire new_AGEMA_signal_13612 ;
    wire new_AGEMA_signal_13613 ;
    wire new_AGEMA_signal_13614 ;
    wire new_AGEMA_signal_13615 ;
    wire new_AGEMA_signal_13616 ;
    wire new_AGEMA_signal_13617 ;
    wire new_AGEMA_signal_13618 ;
    wire new_AGEMA_signal_13619 ;
    wire new_AGEMA_signal_13620 ;
    wire new_AGEMA_signal_13621 ;
    wire new_AGEMA_signal_13622 ;
    wire new_AGEMA_signal_13623 ;
    wire new_AGEMA_signal_13624 ;
    wire new_AGEMA_signal_13625 ;
    wire new_AGEMA_signal_13626 ;
    wire new_AGEMA_signal_13627 ;
    wire new_AGEMA_signal_13628 ;
    wire new_AGEMA_signal_13629 ;
    wire new_AGEMA_signal_13630 ;
    wire new_AGEMA_signal_13631 ;
    wire new_AGEMA_signal_13632 ;
    wire new_AGEMA_signal_13633 ;
    wire new_AGEMA_signal_13634 ;
    wire new_AGEMA_signal_13635 ;
    wire new_AGEMA_signal_13636 ;
    wire new_AGEMA_signal_13637 ;
    wire new_AGEMA_signal_13638 ;
    wire new_AGEMA_signal_13639 ;
    wire new_AGEMA_signal_13640 ;
    wire new_AGEMA_signal_13641 ;
    wire new_AGEMA_signal_13642 ;
    wire new_AGEMA_signal_13643 ;
    wire new_AGEMA_signal_13644 ;
    wire new_AGEMA_signal_13645 ;
    wire new_AGEMA_signal_13646 ;
    wire new_AGEMA_signal_13647 ;
    wire new_AGEMA_signal_13648 ;
    wire new_AGEMA_signal_13649 ;
    wire new_AGEMA_signal_13650 ;
    wire new_AGEMA_signal_13651 ;
    wire new_AGEMA_signal_13652 ;
    wire new_AGEMA_signal_13653 ;
    wire new_AGEMA_signal_13654 ;
    wire new_AGEMA_signal_13655 ;
    wire new_AGEMA_signal_13656 ;
    wire new_AGEMA_signal_13657 ;
    wire new_AGEMA_signal_13658 ;
    wire new_AGEMA_signal_13659 ;
    wire new_AGEMA_signal_13660 ;
    wire new_AGEMA_signal_13661 ;
    wire new_AGEMA_signal_13662 ;
    wire new_AGEMA_signal_13663 ;
    wire new_AGEMA_signal_13664 ;
    wire new_AGEMA_signal_13665 ;
    wire new_AGEMA_signal_13666 ;
    wire new_AGEMA_signal_13667 ;
    wire new_AGEMA_signal_13668 ;
    wire new_AGEMA_signal_13669 ;
    wire new_AGEMA_signal_13670 ;
    wire new_AGEMA_signal_13671 ;
    wire new_AGEMA_signal_13672 ;
    wire new_AGEMA_signal_13673 ;
    wire new_AGEMA_signal_13674 ;
    wire new_AGEMA_signal_13675 ;
    wire new_AGEMA_signal_13676 ;
    wire new_AGEMA_signal_13677 ;
    wire new_AGEMA_signal_13678 ;
    wire new_AGEMA_signal_13679 ;
    wire new_AGEMA_signal_13680 ;
    wire new_AGEMA_signal_13681 ;
    wire new_AGEMA_signal_13682 ;
    wire new_AGEMA_signal_13683 ;
    wire new_AGEMA_signal_13684 ;
    wire new_AGEMA_signal_13685 ;
    wire new_AGEMA_signal_13686 ;
    wire new_AGEMA_signal_13687 ;
    wire new_AGEMA_signal_13688 ;
    wire new_AGEMA_signal_13689 ;
    wire new_AGEMA_signal_13690 ;
    wire new_AGEMA_signal_13691 ;
    wire new_AGEMA_signal_13692 ;
    wire new_AGEMA_signal_13693 ;
    wire new_AGEMA_signal_13694 ;
    wire new_AGEMA_signal_13695 ;
    wire new_AGEMA_signal_13696 ;
    wire new_AGEMA_signal_13697 ;
    wire new_AGEMA_signal_13698 ;
    wire new_AGEMA_signal_13699 ;
    wire new_AGEMA_signal_13700 ;
    wire new_AGEMA_signal_13701 ;
    wire new_AGEMA_signal_13702 ;
    wire new_AGEMA_signal_13703 ;
    wire new_AGEMA_signal_13704 ;
    wire new_AGEMA_signal_13705 ;
    wire new_AGEMA_signal_13706 ;
    wire new_AGEMA_signal_13707 ;
    wire new_AGEMA_signal_13708 ;
    wire new_AGEMA_signal_13709 ;
    wire new_AGEMA_signal_13710 ;
    wire new_AGEMA_signal_13711 ;
    wire new_AGEMA_signal_13712 ;
    wire new_AGEMA_signal_13713 ;
    wire new_AGEMA_signal_13714 ;
    wire new_AGEMA_signal_13715 ;
    wire new_AGEMA_signal_13716 ;
    wire new_AGEMA_signal_13717 ;
    wire new_AGEMA_signal_13718 ;
    wire new_AGEMA_signal_13719 ;
    wire new_AGEMA_signal_13720 ;
    wire new_AGEMA_signal_13721 ;
    wire new_AGEMA_signal_13722 ;
    wire new_AGEMA_signal_13723 ;
    wire new_AGEMA_signal_13724 ;
    wire new_AGEMA_signal_13725 ;
    wire new_AGEMA_signal_13726 ;
    wire new_AGEMA_signal_13727 ;
    wire new_AGEMA_signal_13728 ;
    wire new_AGEMA_signal_13729 ;
    wire new_AGEMA_signal_13730 ;
    wire new_AGEMA_signal_13731 ;
    wire new_AGEMA_signal_13732 ;
    wire new_AGEMA_signal_13733 ;
    wire new_AGEMA_signal_13734 ;
    wire new_AGEMA_signal_13735 ;
    wire new_AGEMA_signal_13736 ;
    wire new_AGEMA_signal_13737 ;
    wire new_AGEMA_signal_13738 ;
    wire new_AGEMA_signal_13739 ;
    wire new_AGEMA_signal_13740 ;
    wire new_AGEMA_signal_13741 ;
    wire new_AGEMA_signal_13742 ;
    wire new_AGEMA_signal_13743 ;
    wire new_AGEMA_signal_13744 ;
    wire new_AGEMA_signal_13745 ;
    wire new_AGEMA_signal_13746 ;
    wire new_AGEMA_signal_13747 ;
    wire new_AGEMA_signal_13748 ;
    wire new_AGEMA_signal_13749 ;
    wire new_AGEMA_signal_13750 ;
    wire new_AGEMA_signal_13751 ;
    wire new_AGEMA_signal_13752 ;
    wire new_AGEMA_signal_13753 ;
    wire new_AGEMA_signal_13754 ;
    wire new_AGEMA_signal_13755 ;
    wire new_AGEMA_signal_13756 ;
    wire new_AGEMA_signal_13757 ;
    wire new_AGEMA_signal_13758 ;
    wire new_AGEMA_signal_13759 ;
    wire new_AGEMA_signal_13760 ;
    wire new_AGEMA_signal_13761 ;
    wire new_AGEMA_signal_13762 ;
    wire new_AGEMA_signal_13763 ;
    wire new_AGEMA_signal_13764 ;
    wire new_AGEMA_signal_13765 ;
    wire new_AGEMA_signal_13766 ;
    wire new_AGEMA_signal_13767 ;
    wire new_AGEMA_signal_13768 ;
    wire new_AGEMA_signal_13769 ;
    wire new_AGEMA_signal_13770 ;
    wire new_AGEMA_signal_13771 ;
    wire new_AGEMA_signal_13772 ;
    wire new_AGEMA_signal_13773 ;
    wire new_AGEMA_signal_13774 ;
    wire new_AGEMA_signal_13775 ;
    wire new_AGEMA_signal_13776 ;
    wire new_AGEMA_signal_13777 ;
    wire new_AGEMA_signal_13778 ;
    wire new_AGEMA_signal_13779 ;
    wire new_AGEMA_signal_13780 ;
    wire new_AGEMA_signal_13781 ;
    wire new_AGEMA_signal_13782 ;
    wire new_AGEMA_signal_13783 ;
    wire new_AGEMA_signal_13784 ;
    wire new_AGEMA_signal_13785 ;
    wire new_AGEMA_signal_13786 ;
    wire new_AGEMA_signal_13787 ;
    wire new_AGEMA_signal_13788 ;
    wire new_AGEMA_signal_13789 ;
    wire new_AGEMA_signal_13790 ;
    wire new_AGEMA_signal_13791 ;
    wire new_AGEMA_signal_13792 ;
    wire new_AGEMA_signal_13793 ;
    wire new_AGEMA_signal_13794 ;
    wire new_AGEMA_signal_13795 ;
    wire new_AGEMA_signal_13796 ;
    wire new_AGEMA_signal_13797 ;
    wire new_AGEMA_signal_13798 ;
    wire new_AGEMA_signal_13799 ;
    wire new_AGEMA_signal_13800 ;
    wire new_AGEMA_signal_13801 ;
    wire new_AGEMA_signal_13802 ;
    wire new_AGEMA_signal_13803 ;
    wire new_AGEMA_signal_13804 ;
    wire new_AGEMA_signal_13805 ;
    wire new_AGEMA_signal_13806 ;
    wire new_AGEMA_signal_13807 ;
    wire new_AGEMA_signal_13808 ;
    wire new_AGEMA_signal_13809 ;
    wire new_AGEMA_signal_13810 ;
    wire new_AGEMA_signal_13811 ;
    wire new_AGEMA_signal_13812 ;
    wire new_AGEMA_signal_13813 ;
    wire new_AGEMA_signal_13814 ;
    wire new_AGEMA_signal_13815 ;
    wire new_AGEMA_signal_13816 ;
    wire new_AGEMA_signal_13817 ;
    wire new_AGEMA_signal_13818 ;
    wire new_AGEMA_signal_13819 ;
    wire new_AGEMA_signal_13820 ;
    wire new_AGEMA_signal_13821 ;
    wire new_AGEMA_signal_13822 ;
    wire new_AGEMA_signal_13823 ;
    wire new_AGEMA_signal_13824 ;
    wire new_AGEMA_signal_13825 ;
    wire new_AGEMA_signal_13826 ;
    wire new_AGEMA_signal_13827 ;
    wire new_AGEMA_signal_13828 ;
    wire new_AGEMA_signal_13829 ;
    wire new_AGEMA_signal_13830 ;
    wire new_AGEMA_signal_13831 ;
    wire new_AGEMA_signal_13832 ;
    wire new_AGEMA_signal_13833 ;
    wire new_AGEMA_signal_13834 ;
    wire new_AGEMA_signal_13835 ;
    wire new_AGEMA_signal_13836 ;
    wire new_AGEMA_signal_13837 ;
    wire new_AGEMA_signal_13838 ;
    wire new_AGEMA_signal_13839 ;
    wire new_AGEMA_signal_13840 ;
    wire new_AGEMA_signal_13841 ;
    wire new_AGEMA_signal_13842 ;
    wire new_AGEMA_signal_13843 ;
    wire new_AGEMA_signal_13844 ;
    wire new_AGEMA_signal_13845 ;
    wire new_AGEMA_signal_13846 ;
    wire new_AGEMA_signal_13847 ;
    wire new_AGEMA_signal_13848 ;
    wire new_AGEMA_signal_13849 ;
    wire new_AGEMA_signal_13850 ;
    wire new_AGEMA_signal_13851 ;
    wire new_AGEMA_signal_13852 ;
    wire new_AGEMA_signal_13853 ;
    wire new_AGEMA_signal_13854 ;
    wire new_AGEMA_signal_13855 ;
    wire new_AGEMA_signal_13856 ;
    wire new_AGEMA_signal_13857 ;
    wire new_AGEMA_signal_13858 ;
    wire new_AGEMA_signal_13859 ;
    wire new_AGEMA_signal_13860 ;
    wire new_AGEMA_signal_13861 ;
    wire new_AGEMA_signal_13862 ;
    wire new_AGEMA_signal_13863 ;
    wire new_AGEMA_signal_13864 ;
    wire new_AGEMA_signal_13865 ;
    wire new_AGEMA_signal_13866 ;
    wire new_AGEMA_signal_13867 ;
    wire new_AGEMA_signal_13868 ;
    wire new_AGEMA_signal_13869 ;
    wire new_AGEMA_signal_13870 ;
    wire new_AGEMA_signal_13871 ;
    wire new_AGEMA_signal_13872 ;
    wire new_AGEMA_signal_13873 ;
    wire new_AGEMA_signal_13874 ;
    wire new_AGEMA_signal_13875 ;
    wire new_AGEMA_signal_13876 ;
    wire new_AGEMA_signal_13877 ;
    wire new_AGEMA_signal_13878 ;
    wire new_AGEMA_signal_13879 ;
    wire new_AGEMA_signal_13880 ;
    wire new_AGEMA_signal_13881 ;
    wire new_AGEMA_signal_13882 ;
    wire new_AGEMA_signal_13883 ;
    wire new_AGEMA_signal_13884 ;
    wire new_AGEMA_signal_13885 ;
    wire new_AGEMA_signal_13886 ;
    wire new_AGEMA_signal_13887 ;
    wire new_AGEMA_signal_13888 ;
    wire new_AGEMA_signal_13889 ;
    wire new_AGEMA_signal_13890 ;
    wire new_AGEMA_signal_13891 ;
    wire new_AGEMA_signal_13892 ;
    wire new_AGEMA_signal_13893 ;
    wire new_AGEMA_signal_13894 ;
    wire new_AGEMA_signal_13895 ;
    wire new_AGEMA_signal_13896 ;
    wire new_AGEMA_signal_13897 ;
    wire new_AGEMA_signal_13898 ;
    wire new_AGEMA_signal_13899 ;
    wire new_AGEMA_signal_13900 ;
    wire new_AGEMA_signal_13901 ;
    wire new_AGEMA_signal_13902 ;
    wire new_AGEMA_signal_13903 ;
    wire new_AGEMA_signal_13904 ;
    wire new_AGEMA_signal_13905 ;
    wire new_AGEMA_signal_13906 ;
    wire new_AGEMA_signal_13907 ;
    wire new_AGEMA_signal_13908 ;
    wire new_AGEMA_signal_13909 ;
    wire new_AGEMA_signal_13910 ;
    wire new_AGEMA_signal_13911 ;
    wire new_AGEMA_signal_13912 ;
    wire new_AGEMA_signal_13913 ;
    wire new_AGEMA_signal_13914 ;
    wire new_AGEMA_signal_13915 ;
    wire new_AGEMA_signal_13916 ;
    wire new_AGEMA_signal_13917 ;
    wire new_AGEMA_signal_13918 ;
    wire new_AGEMA_signal_13919 ;
    wire new_AGEMA_signal_13920 ;
    wire new_AGEMA_signal_13921 ;
    wire new_AGEMA_signal_13922 ;
    wire new_AGEMA_signal_13923 ;
    wire new_AGEMA_signal_13924 ;
    wire new_AGEMA_signal_13925 ;
    wire new_AGEMA_signal_13926 ;
    wire new_AGEMA_signal_13927 ;
    wire new_AGEMA_signal_13928 ;
    wire new_AGEMA_signal_13929 ;
    wire new_AGEMA_signal_13930 ;
    wire new_AGEMA_signal_13931 ;
    wire new_AGEMA_signal_13932 ;
    wire new_AGEMA_signal_13933 ;
    wire new_AGEMA_signal_13934 ;
    wire new_AGEMA_signal_13935 ;
    wire new_AGEMA_signal_13936 ;
    wire new_AGEMA_signal_13937 ;
    wire new_AGEMA_signal_13938 ;
    wire new_AGEMA_signal_13939 ;
    wire new_AGEMA_signal_13940 ;
    wire new_AGEMA_signal_13941 ;
    wire new_AGEMA_signal_13942 ;
    wire new_AGEMA_signal_13943 ;
    wire new_AGEMA_signal_13944 ;
    wire new_AGEMA_signal_13945 ;
    wire new_AGEMA_signal_13946 ;
    wire new_AGEMA_signal_13947 ;
    wire new_AGEMA_signal_13948 ;
    wire new_AGEMA_signal_13949 ;
    wire new_AGEMA_signal_13950 ;
    wire new_AGEMA_signal_13951 ;
    wire new_AGEMA_signal_13952 ;
    wire new_AGEMA_signal_13953 ;
    wire new_AGEMA_signal_13954 ;
    wire new_AGEMA_signal_13955 ;
    wire new_AGEMA_signal_13956 ;
    wire new_AGEMA_signal_13957 ;
    wire new_AGEMA_signal_13958 ;
    wire new_AGEMA_signal_13959 ;
    wire new_AGEMA_signal_13960 ;
    wire new_AGEMA_signal_13961 ;
    wire new_AGEMA_signal_13962 ;
    wire new_AGEMA_signal_13963 ;
    wire new_AGEMA_signal_13964 ;
    wire new_AGEMA_signal_13965 ;
    wire new_AGEMA_signal_13966 ;
    wire new_AGEMA_signal_13967 ;
    wire new_AGEMA_signal_13968 ;
    wire new_AGEMA_signal_13969 ;
    wire new_AGEMA_signal_13970 ;
    wire new_AGEMA_signal_13971 ;
    wire new_AGEMA_signal_13972 ;
    wire new_AGEMA_signal_13973 ;
    wire new_AGEMA_signal_13974 ;
    wire new_AGEMA_signal_13975 ;
    wire new_AGEMA_signal_13976 ;
    wire new_AGEMA_signal_13977 ;
    wire new_AGEMA_signal_13978 ;
    wire new_AGEMA_signal_13979 ;
    wire new_AGEMA_signal_13980 ;
    wire new_AGEMA_signal_13981 ;
    wire new_AGEMA_signal_13982 ;
    wire new_AGEMA_signal_13983 ;
    wire new_AGEMA_signal_13984 ;
    wire new_AGEMA_signal_13985 ;
    wire new_AGEMA_signal_13986 ;
    wire new_AGEMA_signal_13987 ;
    wire new_AGEMA_signal_13988 ;
    wire new_AGEMA_signal_13989 ;
    wire new_AGEMA_signal_13990 ;
    wire new_AGEMA_signal_13991 ;
    wire new_AGEMA_signal_13992 ;
    wire new_AGEMA_signal_13993 ;
    wire new_AGEMA_signal_13994 ;
    wire new_AGEMA_signal_13995 ;
    wire new_AGEMA_signal_13996 ;
    wire new_AGEMA_signal_13997 ;
    wire new_AGEMA_signal_13998 ;
    wire new_AGEMA_signal_13999 ;
    wire new_AGEMA_signal_14000 ;
    wire new_AGEMA_signal_14001 ;
    wire new_AGEMA_signal_14002 ;
    wire new_AGEMA_signal_14003 ;
    wire new_AGEMA_signal_14004 ;
    wire new_AGEMA_signal_14005 ;
    wire new_AGEMA_signal_14006 ;
    wire new_AGEMA_signal_14007 ;
    wire new_AGEMA_signal_14008 ;
    wire new_AGEMA_signal_14009 ;
    wire new_AGEMA_signal_14010 ;
    wire new_AGEMA_signal_14011 ;
    wire new_AGEMA_signal_14012 ;
    wire new_AGEMA_signal_14013 ;
    wire new_AGEMA_signal_14014 ;
    wire new_AGEMA_signal_14015 ;
    wire new_AGEMA_signal_14016 ;
    wire new_AGEMA_signal_14017 ;
    wire new_AGEMA_signal_14018 ;
    wire new_AGEMA_signal_14019 ;
    wire new_AGEMA_signal_14020 ;
    wire new_AGEMA_signal_14021 ;
    wire new_AGEMA_signal_14022 ;
    wire new_AGEMA_signal_14023 ;
    wire new_AGEMA_signal_14024 ;
    wire new_AGEMA_signal_14025 ;
    wire new_AGEMA_signal_14026 ;
    wire new_AGEMA_signal_14027 ;
    wire new_AGEMA_signal_14028 ;
    wire new_AGEMA_signal_14029 ;
    wire new_AGEMA_signal_14030 ;
    wire new_AGEMA_signal_14031 ;
    wire new_AGEMA_signal_14032 ;
    wire new_AGEMA_signal_14033 ;
    wire new_AGEMA_signal_14034 ;
    wire new_AGEMA_signal_14035 ;
    wire new_AGEMA_signal_14036 ;
    wire new_AGEMA_signal_14037 ;
    wire new_AGEMA_signal_14038 ;
    wire new_AGEMA_signal_14039 ;
    wire new_AGEMA_signal_14040 ;
    wire new_AGEMA_signal_14041 ;
    wire new_AGEMA_signal_14042 ;
    wire new_AGEMA_signal_14043 ;
    wire new_AGEMA_signal_14044 ;
    wire new_AGEMA_signal_14045 ;
    wire new_AGEMA_signal_14046 ;
    wire new_AGEMA_signal_14047 ;
    wire new_AGEMA_signal_14048 ;
    wire new_AGEMA_signal_14049 ;
    wire new_AGEMA_signal_14050 ;
    wire new_AGEMA_signal_14051 ;
    wire new_AGEMA_signal_14052 ;
    wire new_AGEMA_signal_14053 ;
    wire new_AGEMA_signal_14054 ;
    wire new_AGEMA_signal_14055 ;
    wire new_AGEMA_signal_14056 ;
    wire new_AGEMA_signal_14057 ;
    wire new_AGEMA_signal_14058 ;
    wire new_AGEMA_signal_14059 ;
    wire new_AGEMA_signal_14060 ;
    wire new_AGEMA_signal_14061 ;
    wire new_AGEMA_signal_14062 ;
    wire new_AGEMA_signal_14063 ;
    wire new_AGEMA_signal_14064 ;
    wire new_AGEMA_signal_14065 ;
    wire new_AGEMA_signal_14066 ;
    wire new_AGEMA_signal_14067 ;
    wire new_AGEMA_signal_14068 ;
    wire new_AGEMA_signal_14069 ;
    wire new_AGEMA_signal_14070 ;
    wire new_AGEMA_signal_14071 ;
    wire new_AGEMA_signal_14072 ;
    wire new_AGEMA_signal_14073 ;
    wire new_AGEMA_signal_14074 ;
    wire new_AGEMA_signal_14075 ;
    wire new_AGEMA_signal_14076 ;
    wire new_AGEMA_signal_14077 ;
    wire new_AGEMA_signal_14078 ;
    wire new_AGEMA_signal_14079 ;
    wire new_AGEMA_signal_14080 ;
    wire new_AGEMA_signal_14081 ;
    wire new_AGEMA_signal_14082 ;
    wire new_AGEMA_signal_14083 ;
    wire new_AGEMA_signal_14084 ;
    wire new_AGEMA_signal_14085 ;
    wire new_AGEMA_signal_14086 ;
    wire new_AGEMA_signal_14087 ;
    wire new_AGEMA_signal_14088 ;
    wire new_AGEMA_signal_14089 ;
    wire new_AGEMA_signal_14090 ;
    wire new_AGEMA_signal_14091 ;
    wire new_AGEMA_signal_14092 ;
    wire new_AGEMA_signal_14093 ;
    wire new_AGEMA_signal_14094 ;
    wire new_AGEMA_signal_14095 ;
    wire new_AGEMA_signal_14096 ;
    wire new_AGEMA_signal_14097 ;
    wire new_AGEMA_signal_14098 ;
    wire new_AGEMA_signal_14099 ;
    wire new_AGEMA_signal_14100 ;
    wire new_AGEMA_signal_14101 ;
    wire new_AGEMA_signal_14102 ;
    wire new_AGEMA_signal_14103 ;
    wire new_AGEMA_signal_14104 ;
    wire new_AGEMA_signal_14105 ;
    wire new_AGEMA_signal_14106 ;
    wire new_AGEMA_signal_14107 ;
    wire new_AGEMA_signal_14108 ;
    wire new_AGEMA_signal_14109 ;
    wire new_AGEMA_signal_14110 ;
    wire new_AGEMA_signal_14111 ;
    wire new_AGEMA_signal_14112 ;
    wire new_AGEMA_signal_14113 ;
    wire new_AGEMA_signal_14114 ;
    wire new_AGEMA_signal_14115 ;
    wire new_AGEMA_signal_14116 ;
    wire new_AGEMA_signal_14117 ;
    wire new_AGEMA_signal_14118 ;
    wire new_AGEMA_signal_14119 ;
    wire new_AGEMA_signal_14120 ;
    wire new_AGEMA_signal_14121 ;
    wire new_AGEMA_signal_14122 ;
    wire new_AGEMA_signal_14123 ;
    wire new_AGEMA_signal_14124 ;
    wire new_AGEMA_signal_14125 ;
    wire new_AGEMA_signal_14126 ;
    wire new_AGEMA_signal_14127 ;
    wire new_AGEMA_signal_14128 ;
    wire new_AGEMA_signal_14129 ;
    wire new_AGEMA_signal_14130 ;
    wire new_AGEMA_signal_14131 ;
    wire new_AGEMA_signal_14132 ;
    wire new_AGEMA_signal_14133 ;
    wire new_AGEMA_signal_14134 ;
    wire new_AGEMA_signal_14135 ;
    wire new_AGEMA_signal_14136 ;
    wire new_AGEMA_signal_14137 ;
    wire new_AGEMA_signal_14138 ;
    wire new_AGEMA_signal_14139 ;
    wire new_AGEMA_signal_14140 ;
    wire new_AGEMA_signal_14141 ;
    wire new_AGEMA_signal_14142 ;
    wire new_AGEMA_signal_14143 ;
    wire new_AGEMA_signal_14144 ;
    wire new_AGEMA_signal_14145 ;
    wire new_AGEMA_signal_14146 ;
    wire new_AGEMA_signal_14147 ;
    wire new_AGEMA_signal_14148 ;
    wire new_AGEMA_signal_14149 ;
    wire new_AGEMA_signal_14150 ;
    wire new_AGEMA_signal_14151 ;
    wire new_AGEMA_signal_14152 ;
    wire new_AGEMA_signal_14153 ;
    wire new_AGEMA_signal_14154 ;
    wire new_AGEMA_signal_14155 ;
    wire new_AGEMA_signal_14156 ;
    wire new_AGEMA_signal_14157 ;
    wire new_AGEMA_signal_14158 ;
    wire new_AGEMA_signal_14159 ;
    wire new_AGEMA_signal_14160 ;
    wire new_AGEMA_signal_14161 ;
    wire new_AGEMA_signal_14162 ;
    wire new_AGEMA_signal_14163 ;
    wire new_AGEMA_signal_14164 ;
    wire new_AGEMA_signal_14165 ;
    wire new_AGEMA_signal_14166 ;
    wire new_AGEMA_signal_14167 ;
    wire new_AGEMA_signal_14168 ;
    wire new_AGEMA_signal_14169 ;
    wire new_AGEMA_signal_14170 ;
    wire new_AGEMA_signal_14171 ;
    wire new_AGEMA_signal_14172 ;
    wire new_AGEMA_signal_14173 ;
    wire new_AGEMA_signal_14174 ;
    wire new_AGEMA_signal_14175 ;
    wire new_AGEMA_signal_14176 ;
    wire new_AGEMA_signal_14177 ;
    wire new_AGEMA_signal_14178 ;
    wire new_AGEMA_signal_14179 ;
    wire new_AGEMA_signal_14180 ;
    wire new_AGEMA_signal_14181 ;
    wire new_AGEMA_signal_14182 ;
    wire new_AGEMA_signal_14183 ;
    wire new_AGEMA_signal_14184 ;
    wire new_AGEMA_signal_14185 ;
    wire new_AGEMA_signal_14186 ;
    wire new_AGEMA_signal_14187 ;
    wire new_AGEMA_signal_14188 ;
    wire new_AGEMA_signal_14189 ;
    wire new_AGEMA_signal_14190 ;
    wire new_AGEMA_signal_14191 ;
    wire new_AGEMA_signal_14192 ;
    wire new_AGEMA_signal_14193 ;
    wire new_AGEMA_signal_14194 ;
    wire new_AGEMA_signal_14195 ;
    wire new_AGEMA_signal_14196 ;
    wire new_AGEMA_signal_14197 ;
    wire new_AGEMA_signal_14198 ;
    wire new_AGEMA_signal_14199 ;
    wire new_AGEMA_signal_14200 ;
    wire new_AGEMA_signal_14201 ;
    wire new_AGEMA_signal_14202 ;
    wire new_AGEMA_signal_14203 ;
    wire new_AGEMA_signal_14204 ;
    wire new_AGEMA_signal_14205 ;
    wire new_AGEMA_signal_14206 ;
    wire new_AGEMA_signal_14207 ;
    wire new_AGEMA_signal_14208 ;
    wire new_AGEMA_signal_14209 ;
    wire new_AGEMA_signal_14210 ;
    wire new_AGEMA_signal_14211 ;
    wire new_AGEMA_signal_14212 ;
    wire new_AGEMA_signal_14213 ;
    wire new_AGEMA_signal_14214 ;
    wire new_AGEMA_signal_14215 ;
    wire new_AGEMA_signal_14216 ;
    wire new_AGEMA_signal_14217 ;
    wire new_AGEMA_signal_14218 ;
    wire new_AGEMA_signal_14219 ;
    wire new_AGEMA_signal_14220 ;
    wire new_AGEMA_signal_14221 ;
    wire new_AGEMA_signal_14222 ;
    wire new_AGEMA_signal_14223 ;
    wire new_AGEMA_signal_14224 ;
    wire new_AGEMA_signal_14225 ;
    wire new_AGEMA_signal_14226 ;
    wire new_AGEMA_signal_14227 ;
    wire new_AGEMA_signal_14228 ;
    wire new_AGEMA_signal_14229 ;
    wire new_AGEMA_signal_14230 ;
    wire new_AGEMA_signal_14231 ;
    wire new_AGEMA_signal_14232 ;
    wire new_AGEMA_signal_14233 ;
    wire new_AGEMA_signal_14234 ;
    wire new_AGEMA_signal_14235 ;
    wire new_AGEMA_signal_14236 ;
    wire new_AGEMA_signal_14237 ;
    wire new_AGEMA_signal_14238 ;
    wire new_AGEMA_signal_14239 ;
    wire new_AGEMA_signal_14240 ;
    wire new_AGEMA_signal_14241 ;
    wire new_AGEMA_signal_14242 ;
    wire new_AGEMA_signal_14243 ;
    wire new_AGEMA_signal_14244 ;
    wire new_AGEMA_signal_14245 ;
    wire new_AGEMA_signal_14246 ;
    wire new_AGEMA_signal_14247 ;
    wire new_AGEMA_signal_14248 ;
    wire new_AGEMA_signal_14249 ;
    wire new_AGEMA_signal_14250 ;
    wire new_AGEMA_signal_14251 ;
    wire new_AGEMA_signal_14252 ;
    wire new_AGEMA_signal_14253 ;
    wire new_AGEMA_signal_14254 ;
    wire new_AGEMA_signal_14255 ;
    wire new_AGEMA_signal_14256 ;
    wire new_AGEMA_signal_14257 ;
    wire new_AGEMA_signal_14258 ;
    wire new_AGEMA_signal_14259 ;
    wire new_AGEMA_signal_14260 ;
    wire new_AGEMA_signal_14261 ;
    wire new_AGEMA_signal_14262 ;
    wire new_AGEMA_signal_14263 ;
    wire new_AGEMA_signal_14264 ;
    wire new_AGEMA_signal_14265 ;
    wire new_AGEMA_signal_14266 ;
    wire new_AGEMA_signal_14267 ;
    wire new_AGEMA_signal_14268 ;
    wire new_AGEMA_signal_14269 ;
    wire new_AGEMA_signal_14270 ;
    wire new_AGEMA_signal_14271 ;
    wire new_AGEMA_signal_14272 ;
    wire new_AGEMA_signal_14273 ;
    wire new_AGEMA_signal_14274 ;
    wire new_AGEMA_signal_14275 ;
    wire new_AGEMA_signal_14276 ;
    wire new_AGEMA_signal_14277 ;
    wire new_AGEMA_signal_14278 ;
    wire new_AGEMA_signal_14279 ;
    wire new_AGEMA_signal_14280 ;
    wire new_AGEMA_signal_14281 ;
    wire new_AGEMA_signal_14282 ;
    wire new_AGEMA_signal_14283 ;
    wire new_AGEMA_signal_14284 ;
    wire new_AGEMA_signal_14285 ;
    wire new_AGEMA_signal_14286 ;
    wire new_AGEMA_signal_14287 ;
    wire new_AGEMA_signal_14288 ;
    wire new_AGEMA_signal_14289 ;
    wire new_AGEMA_signal_14290 ;
    wire new_AGEMA_signal_14291 ;
    wire new_AGEMA_signal_14292 ;
    wire new_AGEMA_signal_14293 ;
    wire new_AGEMA_signal_14294 ;
    wire new_AGEMA_signal_14295 ;
    wire new_AGEMA_signal_14296 ;
    wire new_AGEMA_signal_14297 ;
    wire new_AGEMA_signal_14298 ;
    wire new_AGEMA_signal_14299 ;
    wire new_AGEMA_signal_14300 ;
    wire new_AGEMA_signal_14301 ;
    wire new_AGEMA_signal_14302 ;
    wire new_AGEMA_signal_14303 ;
    wire new_AGEMA_signal_14304 ;
    wire new_AGEMA_signal_14305 ;
    wire new_AGEMA_signal_14306 ;
    wire new_AGEMA_signal_14307 ;
    wire new_AGEMA_signal_14308 ;
    wire new_AGEMA_signal_14309 ;
    wire new_AGEMA_signal_14310 ;
    wire new_AGEMA_signal_14311 ;
    wire new_AGEMA_signal_14312 ;
    wire new_AGEMA_signal_14313 ;
    wire new_AGEMA_signal_14314 ;
    wire new_AGEMA_signal_14315 ;
    wire new_AGEMA_signal_14316 ;
    wire new_AGEMA_signal_14317 ;
    wire new_AGEMA_signal_14318 ;
    wire new_AGEMA_signal_14319 ;
    wire new_AGEMA_signal_14320 ;
    wire new_AGEMA_signal_14321 ;
    wire new_AGEMA_signal_14322 ;
    wire new_AGEMA_signal_14323 ;
    wire new_AGEMA_signal_14324 ;
    wire new_AGEMA_signal_14325 ;
    wire new_AGEMA_signal_14326 ;
    wire new_AGEMA_signal_14327 ;
    wire new_AGEMA_signal_14328 ;
    wire new_AGEMA_signal_14329 ;
    wire new_AGEMA_signal_14330 ;
    wire new_AGEMA_signal_14331 ;
    wire new_AGEMA_signal_14332 ;
    wire new_AGEMA_signal_14333 ;
    wire new_AGEMA_signal_14334 ;
    wire new_AGEMA_signal_14335 ;
    wire new_AGEMA_signal_14336 ;
    wire new_AGEMA_signal_14337 ;
    wire new_AGEMA_signal_14338 ;
    wire new_AGEMA_signal_14339 ;
    wire new_AGEMA_signal_14340 ;
    wire new_AGEMA_signal_14341 ;
    wire new_AGEMA_signal_14342 ;
    wire new_AGEMA_signal_14343 ;
    wire new_AGEMA_signal_14344 ;
    wire new_AGEMA_signal_14345 ;
    wire new_AGEMA_signal_14346 ;
    wire new_AGEMA_signal_14347 ;
    wire new_AGEMA_signal_14348 ;
    wire new_AGEMA_signal_14349 ;
    wire new_AGEMA_signal_14350 ;
    wire new_AGEMA_signal_14351 ;
    wire new_AGEMA_signal_14352 ;
    wire new_AGEMA_signal_14353 ;
    wire new_AGEMA_signal_14354 ;
    wire new_AGEMA_signal_14355 ;
    wire new_AGEMA_signal_14356 ;
    wire new_AGEMA_signal_14357 ;
    wire new_AGEMA_signal_14358 ;
    wire new_AGEMA_signal_14359 ;
    wire new_AGEMA_signal_14360 ;
    wire new_AGEMA_signal_14361 ;
    wire new_AGEMA_signal_14362 ;
    wire new_AGEMA_signal_14363 ;
    wire new_AGEMA_signal_14364 ;
    wire new_AGEMA_signal_14365 ;
    wire new_AGEMA_signal_14366 ;
    wire new_AGEMA_signal_14367 ;
    wire new_AGEMA_signal_14368 ;
    wire new_AGEMA_signal_14369 ;
    wire new_AGEMA_signal_14370 ;
    wire new_AGEMA_signal_14371 ;
    wire new_AGEMA_signal_14372 ;
    wire new_AGEMA_signal_14373 ;
    wire new_AGEMA_signal_14374 ;
    wire new_AGEMA_signal_14375 ;
    wire new_AGEMA_signal_14376 ;
    wire new_AGEMA_signal_14377 ;
    wire new_AGEMA_signal_14378 ;
    wire new_AGEMA_signal_14379 ;
    wire new_AGEMA_signal_14380 ;
    wire new_AGEMA_signal_14381 ;
    wire new_AGEMA_signal_14382 ;
    wire new_AGEMA_signal_14383 ;
    wire new_AGEMA_signal_14384 ;
    wire new_AGEMA_signal_14385 ;
    wire new_AGEMA_signal_14386 ;
    wire new_AGEMA_signal_14387 ;
    wire new_AGEMA_signal_14388 ;
    wire new_AGEMA_signal_14389 ;
    wire new_AGEMA_signal_14390 ;
    wire new_AGEMA_signal_14391 ;
    wire new_AGEMA_signal_14392 ;
    wire new_AGEMA_signal_14393 ;
    wire new_AGEMA_signal_14394 ;
    wire new_AGEMA_signal_14395 ;
    wire new_AGEMA_signal_14396 ;
    wire new_AGEMA_signal_14397 ;
    wire new_AGEMA_signal_14398 ;
    wire new_AGEMA_signal_14399 ;
    wire new_AGEMA_signal_14400 ;
    wire new_AGEMA_signal_14401 ;
    wire new_AGEMA_signal_14402 ;
    wire new_AGEMA_signal_14403 ;
    wire new_AGEMA_signal_14404 ;
    wire new_AGEMA_signal_14405 ;
    wire new_AGEMA_signal_14406 ;
    wire new_AGEMA_signal_14407 ;
    wire new_AGEMA_signal_14408 ;
    wire new_AGEMA_signal_14409 ;
    wire new_AGEMA_signal_14410 ;
    wire new_AGEMA_signal_14411 ;
    wire new_AGEMA_signal_14412 ;
    wire new_AGEMA_signal_14413 ;
    wire new_AGEMA_signal_14414 ;
    wire new_AGEMA_signal_14415 ;
    wire new_AGEMA_signal_14416 ;
    wire new_AGEMA_signal_14417 ;
    wire new_AGEMA_signal_14418 ;
    wire new_AGEMA_signal_14419 ;
    wire new_AGEMA_signal_14420 ;
    wire new_AGEMA_signal_14421 ;
    wire new_AGEMA_signal_14422 ;
    wire new_AGEMA_signal_14423 ;
    wire new_AGEMA_signal_14424 ;
    wire new_AGEMA_signal_14425 ;
    wire new_AGEMA_signal_14426 ;
    wire new_AGEMA_signal_14427 ;
    wire new_AGEMA_signal_14428 ;
    wire new_AGEMA_signal_14429 ;
    wire new_AGEMA_signal_14430 ;
    wire new_AGEMA_signal_14431 ;
    wire new_AGEMA_signal_14432 ;
    wire new_AGEMA_signal_14433 ;
    wire new_AGEMA_signal_14434 ;
    wire new_AGEMA_signal_14435 ;
    wire new_AGEMA_signal_14436 ;
    wire new_AGEMA_signal_14437 ;
    wire new_AGEMA_signal_14438 ;
    wire new_AGEMA_signal_14439 ;
    wire new_AGEMA_signal_14440 ;
    wire new_AGEMA_signal_14441 ;
    wire new_AGEMA_signal_14442 ;
    wire new_AGEMA_signal_14443 ;
    wire new_AGEMA_signal_14444 ;
    wire new_AGEMA_signal_14445 ;
    wire new_AGEMA_signal_14446 ;
    wire new_AGEMA_signal_14447 ;
    wire new_AGEMA_signal_14448 ;
    wire new_AGEMA_signal_14449 ;
    wire new_AGEMA_signal_14450 ;
    wire new_AGEMA_signal_14451 ;
    wire new_AGEMA_signal_14452 ;
    wire new_AGEMA_signal_14453 ;
    wire new_AGEMA_signal_14454 ;
    wire new_AGEMA_signal_14455 ;
    wire new_AGEMA_signal_14456 ;
    wire new_AGEMA_signal_14457 ;
    wire new_AGEMA_signal_14458 ;
    wire new_AGEMA_signal_14459 ;
    wire new_AGEMA_signal_14460 ;
    wire new_AGEMA_signal_14461 ;
    wire new_AGEMA_signal_14462 ;
    wire new_AGEMA_signal_14463 ;
    wire new_AGEMA_signal_14464 ;
    wire new_AGEMA_signal_14465 ;
    wire new_AGEMA_signal_14466 ;
    wire new_AGEMA_signal_14467 ;
    wire new_AGEMA_signal_14468 ;
    wire new_AGEMA_signal_14469 ;
    wire new_AGEMA_signal_14470 ;
    wire new_AGEMA_signal_14471 ;
    wire new_AGEMA_signal_14472 ;
    wire new_AGEMA_signal_14473 ;
    wire new_AGEMA_signal_14474 ;
    wire new_AGEMA_signal_14475 ;
    wire new_AGEMA_signal_14476 ;
    wire new_AGEMA_signal_14477 ;
    wire new_AGEMA_signal_14478 ;
    wire new_AGEMA_signal_14479 ;
    wire new_AGEMA_signal_14480 ;
    wire new_AGEMA_signal_14481 ;
    wire new_AGEMA_signal_14482 ;
    wire new_AGEMA_signal_14483 ;
    wire new_AGEMA_signal_14484 ;
    wire new_AGEMA_signal_14485 ;
    wire new_AGEMA_signal_14486 ;
    wire new_AGEMA_signal_14487 ;
    wire new_AGEMA_signal_14488 ;
    wire new_AGEMA_signal_14489 ;
    wire new_AGEMA_signal_14490 ;
    wire new_AGEMA_signal_14491 ;
    wire new_AGEMA_signal_14492 ;
    wire new_AGEMA_signal_14493 ;
    wire new_AGEMA_signal_14494 ;
    wire new_AGEMA_signal_14495 ;
    wire new_AGEMA_signal_14496 ;
    wire new_AGEMA_signal_14497 ;
    wire new_AGEMA_signal_14498 ;
    wire new_AGEMA_signal_14499 ;
    wire new_AGEMA_signal_14500 ;
    wire new_AGEMA_signal_14501 ;
    wire new_AGEMA_signal_14502 ;
    wire new_AGEMA_signal_14503 ;
    wire new_AGEMA_signal_14504 ;
    wire new_AGEMA_signal_14505 ;
    wire new_AGEMA_signal_14506 ;
    wire new_AGEMA_signal_14507 ;
    wire new_AGEMA_signal_14508 ;
    wire new_AGEMA_signal_14509 ;
    wire new_AGEMA_signal_14510 ;
    wire new_AGEMA_signal_14511 ;
    wire new_AGEMA_signal_14512 ;
    wire new_AGEMA_signal_14513 ;
    wire new_AGEMA_signal_14514 ;
    wire new_AGEMA_signal_14515 ;
    wire new_AGEMA_signal_14516 ;
    wire new_AGEMA_signal_14517 ;
    wire new_AGEMA_signal_14518 ;
    wire new_AGEMA_signal_14519 ;
    wire new_AGEMA_signal_14520 ;
    wire new_AGEMA_signal_14521 ;
    wire new_AGEMA_signal_14522 ;
    wire new_AGEMA_signal_14523 ;
    wire new_AGEMA_signal_14524 ;
    wire new_AGEMA_signal_14525 ;
    wire new_AGEMA_signal_14526 ;
    wire new_AGEMA_signal_14527 ;
    wire new_AGEMA_signal_14528 ;
    wire new_AGEMA_signal_14529 ;
    wire new_AGEMA_signal_14530 ;
    wire new_AGEMA_signal_14531 ;
    wire new_AGEMA_signal_14532 ;
    wire new_AGEMA_signal_14533 ;
    wire new_AGEMA_signal_14534 ;
    wire new_AGEMA_signal_14535 ;
    wire new_AGEMA_signal_14536 ;
    wire new_AGEMA_signal_14537 ;
    wire new_AGEMA_signal_14538 ;
    wire new_AGEMA_signal_14539 ;
    wire new_AGEMA_signal_14540 ;
    wire new_AGEMA_signal_14541 ;
    wire new_AGEMA_signal_14542 ;
    wire new_AGEMA_signal_14543 ;
    wire new_AGEMA_signal_14544 ;
    wire new_AGEMA_signal_14545 ;
    wire new_AGEMA_signal_14546 ;
    wire new_AGEMA_signal_14547 ;
    wire new_AGEMA_signal_14548 ;
    wire new_AGEMA_signal_14549 ;
    wire new_AGEMA_signal_14550 ;
    wire new_AGEMA_signal_14551 ;
    wire new_AGEMA_signal_14552 ;
    wire new_AGEMA_signal_14553 ;
    wire new_AGEMA_signal_14554 ;
    wire new_AGEMA_signal_14555 ;
    wire new_AGEMA_signal_14556 ;
    wire new_AGEMA_signal_14557 ;
    wire new_AGEMA_signal_14558 ;
    wire new_AGEMA_signal_14559 ;
    wire new_AGEMA_signal_14560 ;
    wire new_AGEMA_signal_14561 ;
    wire new_AGEMA_signal_14562 ;
    wire new_AGEMA_signal_14563 ;
    wire new_AGEMA_signal_14564 ;
    wire new_AGEMA_signal_14565 ;
    wire new_AGEMA_signal_14566 ;
    wire new_AGEMA_signal_14567 ;
    wire new_AGEMA_signal_14568 ;
    wire new_AGEMA_signal_14569 ;
    wire new_AGEMA_signal_14570 ;
    wire new_AGEMA_signal_14571 ;
    wire new_AGEMA_signal_14572 ;
    wire new_AGEMA_signal_14573 ;
    wire new_AGEMA_signal_14574 ;
    wire new_AGEMA_signal_14575 ;
    wire new_AGEMA_signal_14576 ;
    wire new_AGEMA_signal_14577 ;
    wire new_AGEMA_signal_14578 ;
    wire new_AGEMA_signal_14579 ;
    wire new_AGEMA_signal_14580 ;
    wire new_AGEMA_signal_14581 ;
    wire new_AGEMA_signal_14582 ;
    wire new_AGEMA_signal_14583 ;
    wire new_AGEMA_signal_14584 ;
    wire new_AGEMA_signal_14585 ;
    wire new_AGEMA_signal_14586 ;
    wire new_AGEMA_signal_14587 ;
    wire new_AGEMA_signal_14588 ;
    wire new_AGEMA_signal_14589 ;
    wire new_AGEMA_signal_14590 ;
    wire new_AGEMA_signal_14591 ;
    wire new_AGEMA_signal_14592 ;
    wire new_AGEMA_signal_14593 ;
    wire new_AGEMA_signal_14594 ;
    wire new_AGEMA_signal_14595 ;
    wire new_AGEMA_signal_14596 ;
    wire new_AGEMA_signal_14597 ;
    wire new_AGEMA_signal_14598 ;
    wire new_AGEMA_signal_14599 ;
    wire new_AGEMA_signal_14600 ;
    wire new_AGEMA_signal_14601 ;
    wire new_AGEMA_signal_14602 ;
    wire new_AGEMA_signal_14603 ;
    wire new_AGEMA_signal_14604 ;
    wire new_AGEMA_signal_14605 ;
    wire new_AGEMA_signal_14606 ;
    wire new_AGEMA_signal_14607 ;
    wire new_AGEMA_signal_14608 ;
    wire new_AGEMA_signal_14609 ;
    wire new_AGEMA_signal_14610 ;
    wire new_AGEMA_signal_14611 ;
    wire new_AGEMA_signal_14612 ;
    wire new_AGEMA_signal_14613 ;
    wire new_AGEMA_signal_14614 ;
    wire new_AGEMA_signal_14615 ;
    wire new_AGEMA_signal_14616 ;
    wire new_AGEMA_signal_14617 ;
    wire new_AGEMA_signal_14618 ;
    wire new_AGEMA_signal_14619 ;
    wire new_AGEMA_signal_14620 ;
    wire new_AGEMA_signal_14621 ;
    wire new_AGEMA_signal_14622 ;
    wire new_AGEMA_signal_14623 ;
    wire new_AGEMA_signal_14624 ;
    wire new_AGEMA_signal_14625 ;
    wire new_AGEMA_signal_14626 ;
    wire new_AGEMA_signal_14627 ;
    wire new_AGEMA_signal_14628 ;
    wire new_AGEMA_signal_14629 ;
    wire new_AGEMA_signal_14630 ;
    wire new_AGEMA_signal_14631 ;
    wire new_AGEMA_signal_14632 ;
    wire new_AGEMA_signal_14633 ;
    wire new_AGEMA_signal_14634 ;
    wire new_AGEMA_signal_14635 ;
    wire new_AGEMA_signal_14636 ;
    wire new_AGEMA_signal_14637 ;
    wire new_AGEMA_signal_14638 ;
    wire new_AGEMA_signal_14639 ;
    wire new_AGEMA_signal_14640 ;
    wire new_AGEMA_signal_14641 ;
    wire new_AGEMA_signal_14642 ;
    wire new_AGEMA_signal_14643 ;
    wire new_AGEMA_signal_14644 ;
    wire new_AGEMA_signal_14645 ;
    wire new_AGEMA_signal_14646 ;
    wire new_AGEMA_signal_14647 ;
    wire new_AGEMA_signal_14648 ;
    wire new_AGEMA_signal_14649 ;
    wire new_AGEMA_signal_14650 ;
    wire new_AGEMA_signal_14651 ;
    wire new_AGEMA_signal_14652 ;
    wire new_AGEMA_signal_14653 ;
    wire new_AGEMA_signal_14654 ;
    wire new_AGEMA_signal_14655 ;
    wire new_AGEMA_signal_14656 ;
    wire new_AGEMA_signal_14657 ;
    wire new_AGEMA_signal_14658 ;
    wire new_AGEMA_signal_14659 ;
    wire new_AGEMA_signal_14660 ;
    wire new_AGEMA_signal_14661 ;
    wire new_AGEMA_signal_14662 ;
    wire new_AGEMA_signal_14663 ;
    wire new_AGEMA_signal_14664 ;
    wire new_AGEMA_signal_14665 ;
    wire new_AGEMA_signal_14666 ;
    wire new_AGEMA_signal_14667 ;
    wire new_AGEMA_signal_14668 ;
    wire new_AGEMA_signal_14669 ;
    wire new_AGEMA_signal_14670 ;
    wire new_AGEMA_signal_14671 ;
    wire new_AGEMA_signal_14672 ;
    wire new_AGEMA_signal_14673 ;
    wire new_AGEMA_signal_14674 ;
    wire new_AGEMA_signal_14675 ;
    wire new_AGEMA_signal_14676 ;
    wire new_AGEMA_signal_14677 ;
    wire new_AGEMA_signal_14678 ;
    wire new_AGEMA_signal_14679 ;
    wire new_AGEMA_signal_14680 ;
    wire new_AGEMA_signal_14681 ;
    wire new_AGEMA_signal_14682 ;
    wire new_AGEMA_signal_14683 ;
    wire new_AGEMA_signal_14684 ;
    wire new_AGEMA_signal_14685 ;
    wire new_AGEMA_signal_14686 ;
    wire new_AGEMA_signal_14687 ;
    wire new_AGEMA_signal_14688 ;
    wire new_AGEMA_signal_14689 ;
    wire new_AGEMA_signal_14690 ;
    wire new_AGEMA_signal_14691 ;
    wire new_AGEMA_signal_14692 ;
    wire new_AGEMA_signal_14693 ;
    wire new_AGEMA_signal_14694 ;
    wire new_AGEMA_signal_14695 ;
    wire new_AGEMA_signal_14696 ;
    wire new_AGEMA_signal_14697 ;
    wire new_AGEMA_signal_14698 ;
    wire new_AGEMA_signal_14699 ;
    wire new_AGEMA_signal_14700 ;
    wire new_AGEMA_signal_14701 ;
    wire new_AGEMA_signal_14702 ;
    wire new_AGEMA_signal_14703 ;
    wire new_AGEMA_signal_14704 ;
    wire new_AGEMA_signal_14705 ;
    wire new_AGEMA_signal_14706 ;
    wire new_AGEMA_signal_14707 ;
    wire new_AGEMA_signal_14708 ;
    wire new_AGEMA_signal_14709 ;
    wire new_AGEMA_signal_14710 ;
    wire new_AGEMA_signal_14711 ;
    wire new_AGEMA_signal_14712 ;
    wire new_AGEMA_signal_14713 ;
    wire new_AGEMA_signal_14714 ;
    wire new_AGEMA_signal_14715 ;
    wire new_AGEMA_signal_14716 ;
    wire new_AGEMA_signal_14717 ;
    wire new_AGEMA_signal_14718 ;
    wire new_AGEMA_signal_14719 ;
    wire new_AGEMA_signal_14720 ;
    wire new_AGEMA_signal_14721 ;
    wire new_AGEMA_signal_14722 ;
    wire new_AGEMA_signal_14723 ;
    wire new_AGEMA_signal_14724 ;
    wire new_AGEMA_signal_14725 ;
    wire new_AGEMA_signal_14726 ;
    wire new_AGEMA_signal_14727 ;
    wire new_AGEMA_signal_14728 ;
    wire new_AGEMA_signal_14729 ;
    wire new_AGEMA_signal_14730 ;
    wire new_AGEMA_signal_14731 ;
    wire new_AGEMA_signal_14732 ;
    wire new_AGEMA_signal_14733 ;
    wire new_AGEMA_signal_14734 ;
    wire new_AGEMA_signal_14735 ;
    wire new_AGEMA_signal_14736 ;
    wire new_AGEMA_signal_14737 ;
    wire new_AGEMA_signal_14738 ;
    wire new_AGEMA_signal_14739 ;
    wire new_AGEMA_signal_14740 ;
    wire new_AGEMA_signal_14741 ;
    wire new_AGEMA_signal_14742 ;
    wire new_AGEMA_signal_14743 ;
    wire new_AGEMA_signal_14744 ;
    wire new_AGEMA_signal_14745 ;
    wire new_AGEMA_signal_14746 ;
    wire new_AGEMA_signal_14747 ;
    wire new_AGEMA_signal_14748 ;
    wire new_AGEMA_signal_14749 ;
    wire new_AGEMA_signal_14750 ;
    wire new_AGEMA_signal_14751 ;
    wire new_AGEMA_signal_14752 ;
    wire new_AGEMA_signal_14753 ;
    wire new_AGEMA_signal_14754 ;
    wire new_AGEMA_signal_14755 ;
    wire new_AGEMA_signal_14756 ;
    wire new_AGEMA_signal_14757 ;
    wire new_AGEMA_signal_14758 ;
    wire new_AGEMA_signal_14759 ;
    wire new_AGEMA_signal_14760 ;
    wire new_AGEMA_signal_14761 ;
    wire new_AGEMA_signal_14762 ;
    wire new_AGEMA_signal_14763 ;
    wire new_AGEMA_signal_14764 ;
    wire new_AGEMA_signal_14765 ;
    wire new_AGEMA_signal_14766 ;
    wire new_AGEMA_signal_14767 ;
    wire new_AGEMA_signal_14768 ;
    wire new_AGEMA_signal_14769 ;
    wire new_AGEMA_signal_14770 ;
    wire new_AGEMA_signal_14771 ;
    wire new_AGEMA_signal_14772 ;
    wire new_AGEMA_signal_14773 ;
    wire new_AGEMA_signal_14774 ;
    wire new_AGEMA_signal_14775 ;
    wire new_AGEMA_signal_14776 ;
    wire new_AGEMA_signal_14777 ;
    wire new_AGEMA_signal_14778 ;
    wire new_AGEMA_signal_14779 ;
    wire new_AGEMA_signal_14780 ;
    wire new_AGEMA_signal_14781 ;
    wire new_AGEMA_signal_14782 ;
    wire new_AGEMA_signal_14783 ;
    wire new_AGEMA_signal_14784 ;
    wire new_AGEMA_signal_14785 ;
    wire new_AGEMA_signal_14786 ;
    wire new_AGEMA_signal_14787 ;
    wire new_AGEMA_signal_14788 ;
    wire new_AGEMA_signal_14789 ;
    wire new_AGEMA_signal_14790 ;
    wire new_AGEMA_signal_14791 ;
    wire new_AGEMA_signal_14792 ;
    wire new_AGEMA_signal_14793 ;
    wire new_AGEMA_signal_14794 ;
    wire new_AGEMA_signal_14795 ;
    wire new_AGEMA_signal_14796 ;
    wire new_AGEMA_signal_14797 ;
    wire new_AGEMA_signal_14798 ;
    wire new_AGEMA_signal_14799 ;
    wire new_AGEMA_signal_14800 ;
    wire new_AGEMA_signal_14801 ;
    wire new_AGEMA_signal_14802 ;
    wire new_AGEMA_signal_14803 ;
    wire new_AGEMA_signal_14804 ;
    wire new_AGEMA_signal_14805 ;
    wire new_AGEMA_signal_14806 ;
    wire new_AGEMA_signal_14807 ;
    wire new_AGEMA_signal_14808 ;
    wire new_AGEMA_signal_14809 ;
    wire new_AGEMA_signal_14810 ;
    wire new_AGEMA_signal_14811 ;
    wire new_AGEMA_signal_14812 ;
    wire new_AGEMA_signal_14813 ;
    wire new_AGEMA_signal_14814 ;
    wire new_AGEMA_signal_14815 ;
    wire new_AGEMA_signal_14816 ;
    wire new_AGEMA_signal_14817 ;
    wire new_AGEMA_signal_14818 ;
    wire new_AGEMA_signal_14819 ;
    wire new_AGEMA_signal_14820 ;
    wire new_AGEMA_signal_14821 ;
    wire new_AGEMA_signal_14822 ;
    wire new_AGEMA_signal_14823 ;
    wire new_AGEMA_signal_14824 ;
    wire new_AGEMA_signal_14825 ;
    wire new_AGEMA_signal_14826 ;
    wire new_AGEMA_signal_14827 ;
    wire new_AGEMA_signal_14828 ;
    wire new_AGEMA_signal_14829 ;
    wire new_AGEMA_signal_14830 ;
    wire new_AGEMA_signal_14831 ;
    wire new_AGEMA_signal_14832 ;
    wire new_AGEMA_signal_14833 ;
    wire new_AGEMA_signal_14834 ;
    wire new_AGEMA_signal_14835 ;
    wire new_AGEMA_signal_14836 ;
    wire new_AGEMA_signal_14837 ;
    wire new_AGEMA_signal_14838 ;
    wire new_AGEMA_signal_14839 ;
    wire new_AGEMA_signal_14840 ;
    wire new_AGEMA_signal_14841 ;
    wire new_AGEMA_signal_14842 ;
    wire new_AGEMA_signal_14843 ;
    wire new_AGEMA_signal_14844 ;
    wire new_AGEMA_signal_14845 ;
    wire new_AGEMA_signal_14846 ;
    wire new_AGEMA_signal_14847 ;
    wire new_AGEMA_signal_14848 ;
    wire new_AGEMA_signal_14849 ;
    wire new_AGEMA_signal_14850 ;
    wire new_AGEMA_signal_14851 ;
    wire new_AGEMA_signal_14852 ;
    wire new_AGEMA_signal_14853 ;
    wire new_AGEMA_signal_14854 ;
    wire new_AGEMA_signal_14855 ;
    wire new_AGEMA_signal_14856 ;
    wire new_AGEMA_signal_14857 ;
    wire new_AGEMA_signal_14858 ;
    wire new_AGEMA_signal_14859 ;
    wire new_AGEMA_signal_14860 ;
    wire new_AGEMA_signal_14861 ;
    wire new_AGEMA_signal_14862 ;
    wire new_AGEMA_signal_14863 ;
    wire new_AGEMA_signal_14864 ;
    wire new_AGEMA_signal_14865 ;
    wire new_AGEMA_signal_14866 ;
    wire new_AGEMA_signal_14867 ;
    wire new_AGEMA_signal_14868 ;
    wire new_AGEMA_signal_14869 ;
    wire new_AGEMA_signal_14870 ;
    wire new_AGEMA_signal_14871 ;
    wire new_AGEMA_signal_14872 ;
    wire new_AGEMA_signal_14873 ;
    wire new_AGEMA_signal_14874 ;
    wire new_AGEMA_signal_14875 ;
    wire new_AGEMA_signal_14876 ;
    wire new_AGEMA_signal_14877 ;
    wire new_AGEMA_signal_14878 ;
    wire new_AGEMA_signal_14879 ;
    wire new_AGEMA_signal_14880 ;
    wire new_AGEMA_signal_14881 ;
    wire new_AGEMA_signal_14882 ;
    wire new_AGEMA_signal_14883 ;
    wire new_AGEMA_signal_14884 ;
    wire new_AGEMA_signal_14885 ;
    wire new_AGEMA_signal_14886 ;
    wire new_AGEMA_signal_14887 ;
    wire new_AGEMA_signal_14888 ;
    wire new_AGEMA_signal_14889 ;
    wire new_AGEMA_signal_14890 ;
    wire new_AGEMA_signal_14891 ;
    wire new_AGEMA_signal_14892 ;
    wire new_AGEMA_signal_14893 ;
    wire new_AGEMA_signal_14894 ;
    wire new_AGEMA_signal_14895 ;
    wire new_AGEMA_signal_14896 ;
    wire new_AGEMA_signal_14897 ;
    wire new_AGEMA_signal_14898 ;
    wire new_AGEMA_signal_14899 ;
    wire new_AGEMA_signal_14900 ;
    wire new_AGEMA_signal_14901 ;
    wire new_AGEMA_signal_14902 ;
    wire new_AGEMA_signal_14903 ;
    wire new_AGEMA_signal_14904 ;
    wire new_AGEMA_signal_14905 ;
    wire new_AGEMA_signal_14906 ;
    wire new_AGEMA_signal_14907 ;
    wire new_AGEMA_signal_14908 ;
    wire new_AGEMA_signal_14909 ;
    wire new_AGEMA_signal_14910 ;
    wire new_AGEMA_signal_14911 ;
    wire new_AGEMA_signal_14912 ;
    wire new_AGEMA_signal_14913 ;
    wire new_AGEMA_signal_14914 ;
    wire new_AGEMA_signal_14915 ;
    wire new_AGEMA_signal_14916 ;
    wire new_AGEMA_signal_14917 ;
    wire new_AGEMA_signal_14918 ;
    wire new_AGEMA_signal_14919 ;
    wire new_AGEMA_signal_14920 ;
    wire new_AGEMA_signal_14921 ;
    wire new_AGEMA_signal_14922 ;
    wire new_AGEMA_signal_14923 ;
    wire new_AGEMA_signal_14924 ;
    wire new_AGEMA_signal_14925 ;
    wire new_AGEMA_signal_14926 ;
    wire new_AGEMA_signal_14927 ;
    wire new_AGEMA_signal_14928 ;
    wire new_AGEMA_signal_14929 ;
    wire new_AGEMA_signal_14930 ;
    wire new_AGEMA_signal_14931 ;
    wire new_AGEMA_signal_14932 ;
    wire new_AGEMA_signal_14933 ;
    wire new_AGEMA_signal_14934 ;
    wire new_AGEMA_signal_14935 ;
    wire new_AGEMA_signal_14936 ;
    wire new_AGEMA_signal_14937 ;
    wire new_AGEMA_signal_14938 ;
    wire new_AGEMA_signal_14939 ;
    wire new_AGEMA_signal_14940 ;
    wire new_AGEMA_signal_14941 ;
    wire new_AGEMA_signal_14942 ;
    wire new_AGEMA_signal_14943 ;
    wire new_AGEMA_signal_14944 ;
    wire new_AGEMA_signal_14945 ;
    wire new_AGEMA_signal_14946 ;
    wire new_AGEMA_signal_14947 ;
    wire new_AGEMA_signal_14948 ;
    wire new_AGEMA_signal_14949 ;
    wire new_AGEMA_signal_14950 ;
    wire new_AGEMA_signal_14951 ;
    wire new_AGEMA_signal_14952 ;
    wire new_AGEMA_signal_14953 ;
    wire new_AGEMA_signal_14954 ;
    wire new_AGEMA_signal_14955 ;
    wire new_AGEMA_signal_14956 ;
    wire new_AGEMA_signal_14957 ;
    wire new_AGEMA_signal_14958 ;
    wire new_AGEMA_signal_14959 ;
    wire new_AGEMA_signal_14960 ;
    wire new_AGEMA_signal_14961 ;
    wire new_AGEMA_signal_14962 ;
    wire new_AGEMA_signal_14963 ;
    wire new_AGEMA_signal_14964 ;
    wire new_AGEMA_signal_14965 ;
    wire new_AGEMA_signal_14966 ;
    wire new_AGEMA_signal_14967 ;
    wire new_AGEMA_signal_14968 ;
    wire new_AGEMA_signal_14969 ;
    wire new_AGEMA_signal_14970 ;
    wire new_AGEMA_signal_14971 ;
    wire new_AGEMA_signal_14972 ;
    wire new_AGEMA_signal_14973 ;
    wire new_AGEMA_signal_14974 ;
    wire new_AGEMA_signal_14975 ;
    wire new_AGEMA_signal_14976 ;
    wire new_AGEMA_signal_14977 ;
    wire new_AGEMA_signal_14978 ;
    wire new_AGEMA_signal_14979 ;
    wire new_AGEMA_signal_14980 ;
    wire new_AGEMA_signal_14981 ;
    wire new_AGEMA_signal_14982 ;
    wire new_AGEMA_signal_14983 ;
    wire new_AGEMA_signal_14984 ;
    wire new_AGEMA_signal_14985 ;
    wire new_AGEMA_signal_14986 ;
    wire new_AGEMA_signal_14987 ;
    wire new_AGEMA_signal_14988 ;
    wire new_AGEMA_signal_14989 ;
    wire new_AGEMA_signal_14990 ;
    wire new_AGEMA_signal_14991 ;
    wire new_AGEMA_signal_14992 ;
    wire new_AGEMA_signal_14993 ;
    wire new_AGEMA_signal_14994 ;
    wire new_AGEMA_signal_14995 ;
    wire new_AGEMA_signal_14996 ;
    wire new_AGEMA_signal_14997 ;
    wire new_AGEMA_signal_14998 ;
    wire new_AGEMA_signal_14999 ;
    wire new_AGEMA_signal_15000 ;
    wire new_AGEMA_signal_15001 ;
    wire new_AGEMA_signal_15002 ;
    wire new_AGEMA_signal_15003 ;
    wire new_AGEMA_signal_15004 ;
    wire new_AGEMA_signal_15005 ;
    wire new_AGEMA_signal_15006 ;
    wire new_AGEMA_signal_15007 ;
    wire new_AGEMA_signal_15008 ;
    wire new_AGEMA_signal_15009 ;
    wire new_AGEMA_signal_15010 ;
    wire new_AGEMA_signal_15011 ;
    wire new_AGEMA_signal_15012 ;
    wire new_AGEMA_signal_15013 ;
    wire new_AGEMA_signal_15014 ;
    wire new_AGEMA_signal_15015 ;
    wire new_AGEMA_signal_15016 ;
    wire new_AGEMA_signal_15017 ;
    wire new_AGEMA_signal_15018 ;
    wire new_AGEMA_signal_15019 ;
    wire new_AGEMA_signal_15020 ;
    wire new_AGEMA_signal_15021 ;
    wire new_AGEMA_signal_15022 ;
    wire new_AGEMA_signal_15023 ;
    wire new_AGEMA_signal_15024 ;
    wire new_AGEMA_signal_15025 ;
    wire new_AGEMA_signal_15026 ;
    wire new_AGEMA_signal_15027 ;
    wire new_AGEMA_signal_15028 ;
    wire new_AGEMA_signal_15029 ;
    wire new_AGEMA_signal_15030 ;
    wire new_AGEMA_signal_15031 ;
    wire new_AGEMA_signal_15032 ;
    wire new_AGEMA_signal_15033 ;
    wire new_AGEMA_signal_15034 ;
    wire new_AGEMA_signal_15035 ;
    wire new_AGEMA_signal_15036 ;
    wire new_AGEMA_signal_15037 ;
    wire new_AGEMA_signal_15038 ;
    wire new_AGEMA_signal_15039 ;
    wire new_AGEMA_signal_15040 ;
    wire new_AGEMA_signal_15041 ;
    wire new_AGEMA_signal_15042 ;
    wire new_AGEMA_signal_15043 ;
    wire new_AGEMA_signal_15044 ;
    wire new_AGEMA_signal_15045 ;
    wire new_AGEMA_signal_15046 ;
    wire new_AGEMA_signal_15047 ;
    wire new_AGEMA_signal_15048 ;
    wire new_AGEMA_signal_15049 ;
    wire new_AGEMA_signal_15050 ;
    wire new_AGEMA_signal_15051 ;
    wire new_AGEMA_signal_15052 ;
    wire new_AGEMA_signal_15053 ;
    wire new_AGEMA_signal_15054 ;
    wire new_AGEMA_signal_15055 ;
    wire new_AGEMA_signal_15056 ;
    wire new_AGEMA_signal_15057 ;
    wire new_AGEMA_signal_15058 ;
    wire new_AGEMA_signal_15059 ;
    wire new_AGEMA_signal_15060 ;
    wire new_AGEMA_signal_15061 ;
    wire new_AGEMA_signal_15062 ;
    wire new_AGEMA_signal_15063 ;
    wire new_AGEMA_signal_15064 ;
    wire new_AGEMA_signal_15065 ;
    wire new_AGEMA_signal_15066 ;
    wire new_AGEMA_signal_15067 ;
    wire new_AGEMA_signal_15068 ;
    wire new_AGEMA_signal_15069 ;
    wire new_AGEMA_signal_15070 ;
    wire new_AGEMA_signal_15071 ;
    wire new_AGEMA_signal_15072 ;
    wire new_AGEMA_signal_15073 ;
    wire new_AGEMA_signal_15074 ;
    wire new_AGEMA_signal_15075 ;
    wire new_AGEMA_signal_15076 ;
    wire new_AGEMA_signal_15077 ;
    wire new_AGEMA_signal_15078 ;
    wire new_AGEMA_signal_15079 ;
    wire new_AGEMA_signal_15080 ;
    wire new_AGEMA_signal_15081 ;
    wire new_AGEMA_signal_15082 ;
    wire new_AGEMA_signal_15083 ;
    wire new_AGEMA_signal_15084 ;
    wire new_AGEMA_signal_15085 ;
    wire new_AGEMA_signal_15086 ;
    wire new_AGEMA_signal_15087 ;
    wire new_AGEMA_signal_15088 ;
    wire new_AGEMA_signal_15089 ;
    wire new_AGEMA_signal_15090 ;
    wire new_AGEMA_signal_15091 ;
    wire new_AGEMA_signal_15092 ;
    wire new_AGEMA_signal_15093 ;
    wire new_AGEMA_signal_15094 ;
    wire new_AGEMA_signal_15095 ;
    wire new_AGEMA_signal_15096 ;
    wire new_AGEMA_signal_15097 ;
    wire new_AGEMA_signal_15098 ;
    wire new_AGEMA_signal_15099 ;
    wire new_AGEMA_signal_15100 ;
    wire new_AGEMA_signal_15101 ;
    wire new_AGEMA_signal_15102 ;
    wire new_AGEMA_signal_15103 ;
    wire new_AGEMA_signal_15104 ;
    wire new_AGEMA_signal_15105 ;
    wire new_AGEMA_signal_15106 ;
    wire new_AGEMA_signal_15107 ;
    wire new_AGEMA_signal_15108 ;
    wire new_AGEMA_signal_15109 ;
    wire new_AGEMA_signal_15110 ;
    wire new_AGEMA_signal_15111 ;
    wire new_AGEMA_signal_15112 ;
    wire new_AGEMA_signal_15113 ;
    wire new_AGEMA_signal_15114 ;
    wire new_AGEMA_signal_15115 ;
    wire new_AGEMA_signal_15116 ;
    wire new_AGEMA_signal_15117 ;
    wire new_AGEMA_signal_15118 ;
    wire new_AGEMA_signal_15119 ;
    wire new_AGEMA_signal_15120 ;
    wire new_AGEMA_signal_15121 ;
    wire new_AGEMA_signal_15122 ;
    wire new_AGEMA_signal_15123 ;
    wire new_AGEMA_signal_15124 ;
    wire new_AGEMA_signal_15125 ;
    wire new_AGEMA_signal_15126 ;
    wire new_AGEMA_signal_15127 ;
    wire new_AGEMA_signal_15128 ;
    wire new_AGEMA_signal_15129 ;
    wire new_AGEMA_signal_15130 ;
    wire new_AGEMA_signal_15131 ;
    wire new_AGEMA_signal_15132 ;
    wire new_AGEMA_signal_15133 ;
    wire new_AGEMA_signal_15134 ;
    wire new_AGEMA_signal_15135 ;
    wire new_AGEMA_signal_15136 ;
    wire new_AGEMA_signal_15137 ;
    wire new_AGEMA_signal_15138 ;
    wire new_AGEMA_signal_15139 ;
    wire new_AGEMA_signal_15140 ;
    wire new_AGEMA_signal_15141 ;
    wire new_AGEMA_signal_15142 ;
    wire new_AGEMA_signal_15143 ;
    wire new_AGEMA_signal_15144 ;
    wire new_AGEMA_signal_15145 ;
    wire new_AGEMA_signal_15146 ;
    wire new_AGEMA_signal_15147 ;
    wire new_AGEMA_signal_15148 ;
    wire new_AGEMA_signal_15149 ;
    wire new_AGEMA_signal_15150 ;
    wire new_AGEMA_signal_15151 ;
    wire new_AGEMA_signal_15152 ;
    wire new_AGEMA_signal_15153 ;
    wire new_AGEMA_signal_15154 ;
    wire new_AGEMA_signal_15155 ;
    wire new_AGEMA_signal_15156 ;
    wire new_AGEMA_signal_15157 ;
    wire new_AGEMA_signal_15158 ;
    wire new_AGEMA_signal_15159 ;
    wire new_AGEMA_signal_15160 ;
    wire new_AGEMA_signal_15161 ;
    wire new_AGEMA_signal_15162 ;
    wire new_AGEMA_signal_15163 ;
    wire new_AGEMA_signal_15164 ;
    wire new_AGEMA_signal_15165 ;
    wire new_AGEMA_signal_15166 ;
    wire new_AGEMA_signal_15167 ;
    wire new_AGEMA_signal_15168 ;
    wire new_AGEMA_signal_15169 ;
    wire new_AGEMA_signal_15170 ;
    wire new_AGEMA_signal_15171 ;
    wire new_AGEMA_signal_15172 ;
    wire new_AGEMA_signal_15173 ;
    wire new_AGEMA_signal_15174 ;
    wire new_AGEMA_signal_15175 ;
    wire new_AGEMA_signal_15176 ;
    wire new_AGEMA_signal_15177 ;
    wire new_AGEMA_signal_15178 ;
    wire new_AGEMA_signal_15179 ;
    wire new_AGEMA_signal_15180 ;
    wire new_AGEMA_signal_15181 ;
    wire new_AGEMA_signal_15182 ;
    wire new_AGEMA_signal_15183 ;
    wire new_AGEMA_signal_15184 ;
    wire new_AGEMA_signal_15185 ;
    wire new_AGEMA_signal_15186 ;
    wire new_AGEMA_signal_15187 ;
    wire new_AGEMA_signal_15188 ;
    wire new_AGEMA_signal_15189 ;
    wire new_AGEMA_signal_15190 ;
    wire new_AGEMA_signal_15191 ;
    wire new_AGEMA_signal_15192 ;
    wire new_AGEMA_signal_15193 ;
    wire new_AGEMA_signal_15194 ;
    wire new_AGEMA_signal_15195 ;
    wire new_AGEMA_signal_15196 ;
    wire new_AGEMA_signal_15197 ;
    wire new_AGEMA_signal_15198 ;
    wire new_AGEMA_signal_15199 ;
    wire new_AGEMA_signal_15200 ;
    wire new_AGEMA_signal_15201 ;
    wire new_AGEMA_signal_15202 ;
    wire new_AGEMA_signal_15203 ;
    wire new_AGEMA_signal_15204 ;
    wire new_AGEMA_signal_15205 ;
    wire new_AGEMA_signal_15206 ;
    wire new_AGEMA_signal_15207 ;
    wire new_AGEMA_signal_15208 ;
    wire new_AGEMA_signal_15209 ;
    wire new_AGEMA_signal_15210 ;
    wire new_AGEMA_signal_15211 ;
    wire new_AGEMA_signal_15212 ;
    wire new_AGEMA_signal_15213 ;
    wire new_AGEMA_signal_15214 ;
    wire new_AGEMA_signal_15215 ;
    wire new_AGEMA_signal_15216 ;
    wire new_AGEMA_signal_15217 ;
    wire new_AGEMA_signal_15218 ;
    wire new_AGEMA_signal_15219 ;
    wire new_AGEMA_signal_15220 ;
    wire new_AGEMA_signal_15221 ;
    wire new_AGEMA_signal_15222 ;
    wire new_AGEMA_signal_15223 ;
    wire new_AGEMA_signal_15224 ;
    wire new_AGEMA_signal_15225 ;
    wire new_AGEMA_signal_15226 ;
    wire new_AGEMA_signal_15227 ;
    wire new_AGEMA_signal_15228 ;
    wire new_AGEMA_signal_15229 ;
    wire new_AGEMA_signal_15230 ;
    wire new_AGEMA_signal_15231 ;
    wire new_AGEMA_signal_15232 ;
    wire new_AGEMA_signal_15233 ;
    wire new_AGEMA_signal_15234 ;
    wire new_AGEMA_signal_15235 ;
    wire new_AGEMA_signal_15236 ;
    wire new_AGEMA_signal_15237 ;
    wire new_AGEMA_signal_15238 ;
    wire new_AGEMA_signal_15239 ;
    wire new_AGEMA_signal_15240 ;
    wire new_AGEMA_signal_15241 ;
    wire new_AGEMA_signal_15242 ;
    wire new_AGEMA_signal_15243 ;
    wire new_AGEMA_signal_15244 ;
    wire new_AGEMA_signal_15245 ;
    wire new_AGEMA_signal_15246 ;
    wire new_AGEMA_signal_15247 ;
    wire new_AGEMA_signal_15248 ;
    wire new_AGEMA_signal_15249 ;
    wire new_AGEMA_signal_15250 ;
    wire new_AGEMA_signal_15251 ;
    wire new_AGEMA_signal_15252 ;
    wire new_AGEMA_signal_15253 ;
    wire new_AGEMA_signal_15254 ;
    wire new_AGEMA_signal_15255 ;
    wire new_AGEMA_signal_15256 ;
    wire new_AGEMA_signal_15257 ;
    wire new_AGEMA_signal_15258 ;
    wire new_AGEMA_signal_15259 ;
    wire new_AGEMA_signal_15260 ;
    wire new_AGEMA_signal_15261 ;
    wire new_AGEMA_signal_15262 ;
    wire new_AGEMA_signal_15263 ;
    wire new_AGEMA_signal_15264 ;
    wire new_AGEMA_signal_15265 ;
    wire new_AGEMA_signal_15266 ;
    wire new_AGEMA_signal_15267 ;
    wire new_AGEMA_signal_15268 ;
    wire new_AGEMA_signal_15269 ;
    wire new_AGEMA_signal_15270 ;
    wire new_AGEMA_signal_15271 ;
    wire new_AGEMA_signal_15272 ;
    wire new_AGEMA_signal_15273 ;
    wire new_AGEMA_signal_15274 ;
    wire new_AGEMA_signal_15275 ;
    wire new_AGEMA_signal_15276 ;
    wire new_AGEMA_signal_15277 ;
    wire new_AGEMA_signal_15278 ;
    wire new_AGEMA_signal_15279 ;
    wire new_AGEMA_signal_15280 ;
    wire new_AGEMA_signal_15281 ;
    wire new_AGEMA_signal_15282 ;
    wire new_AGEMA_signal_15283 ;
    wire new_AGEMA_signal_15284 ;
    wire new_AGEMA_signal_15285 ;
    wire new_AGEMA_signal_15286 ;
    wire new_AGEMA_signal_15287 ;
    wire new_AGEMA_signal_15288 ;
    wire new_AGEMA_signal_15289 ;
    wire new_AGEMA_signal_15290 ;
    wire new_AGEMA_signal_15291 ;
    wire new_AGEMA_signal_15292 ;
    wire new_AGEMA_signal_15293 ;
    wire new_AGEMA_signal_15294 ;
    wire new_AGEMA_signal_15295 ;
    wire new_AGEMA_signal_15296 ;
    wire new_AGEMA_signal_15297 ;
    wire new_AGEMA_signal_15298 ;
    wire new_AGEMA_signal_15299 ;
    wire new_AGEMA_signal_15300 ;
    wire new_AGEMA_signal_15301 ;
    wire new_AGEMA_signal_15302 ;
    wire new_AGEMA_signal_15303 ;
    wire new_AGEMA_signal_15304 ;
    wire new_AGEMA_signal_15305 ;
    wire new_AGEMA_signal_15306 ;
    wire new_AGEMA_signal_15307 ;
    wire new_AGEMA_signal_15308 ;
    wire new_AGEMA_signal_15309 ;
    wire new_AGEMA_signal_15310 ;
    wire new_AGEMA_signal_15311 ;
    wire new_AGEMA_signal_15312 ;
    wire new_AGEMA_signal_15313 ;
    wire new_AGEMA_signal_15314 ;
    wire new_AGEMA_signal_15315 ;
    wire new_AGEMA_signal_15316 ;
    wire new_AGEMA_signal_15317 ;
    wire new_AGEMA_signal_15318 ;
    wire new_AGEMA_signal_15319 ;
    wire new_AGEMA_signal_15320 ;
    wire new_AGEMA_signal_15321 ;
    wire new_AGEMA_signal_15322 ;
    wire new_AGEMA_signal_15323 ;
    wire new_AGEMA_signal_15324 ;
    wire new_AGEMA_signal_15325 ;
    wire new_AGEMA_signal_15326 ;
    wire new_AGEMA_signal_15327 ;
    wire new_AGEMA_signal_15328 ;
    wire new_AGEMA_signal_15329 ;
    wire new_AGEMA_signal_15330 ;
    wire new_AGEMA_signal_15331 ;
    wire new_AGEMA_signal_15332 ;
    wire new_AGEMA_signal_15333 ;
    wire new_AGEMA_signal_15334 ;
    wire new_AGEMA_signal_15335 ;
    wire new_AGEMA_signal_15336 ;
    wire new_AGEMA_signal_15337 ;
    wire new_AGEMA_signal_15338 ;
    wire new_AGEMA_signal_15339 ;
    wire new_AGEMA_signal_15340 ;
    wire new_AGEMA_signal_15341 ;
    wire new_AGEMA_signal_15342 ;
    wire new_AGEMA_signal_15343 ;
    wire new_AGEMA_signal_15344 ;
    wire new_AGEMA_signal_15345 ;
    wire new_AGEMA_signal_15346 ;
    wire new_AGEMA_signal_15347 ;
    wire new_AGEMA_signal_15348 ;
    wire new_AGEMA_signal_15349 ;
    wire new_AGEMA_signal_15350 ;
    wire new_AGEMA_signal_15351 ;
    wire new_AGEMA_signal_15352 ;
    wire new_AGEMA_signal_15353 ;
    wire new_AGEMA_signal_15354 ;
    wire new_AGEMA_signal_15355 ;
    wire new_AGEMA_signal_15356 ;
    wire new_AGEMA_signal_15357 ;
    wire new_AGEMA_signal_15358 ;
    wire new_AGEMA_signal_15359 ;
    wire new_AGEMA_signal_15360 ;
    wire new_AGEMA_signal_15361 ;
    wire new_AGEMA_signal_15362 ;
    wire new_AGEMA_signal_15363 ;
    wire new_AGEMA_signal_15364 ;
    wire new_AGEMA_signal_15365 ;
    wire new_AGEMA_signal_15366 ;
    wire new_AGEMA_signal_15367 ;
    wire new_AGEMA_signal_15368 ;
    wire new_AGEMA_signal_15369 ;
    wire new_AGEMA_signal_15370 ;
    wire new_AGEMA_signal_15371 ;
    wire new_AGEMA_signal_15372 ;
    wire new_AGEMA_signal_15373 ;
    wire new_AGEMA_signal_15374 ;
    wire new_AGEMA_signal_15375 ;
    wire new_AGEMA_signal_15376 ;
    wire new_AGEMA_signal_15377 ;
    wire new_AGEMA_signal_15378 ;
    wire new_AGEMA_signal_15379 ;
    wire new_AGEMA_signal_15380 ;
    wire new_AGEMA_signal_15381 ;
    wire new_AGEMA_signal_15382 ;
    wire new_AGEMA_signal_15383 ;
    wire new_AGEMA_signal_15384 ;
    wire new_AGEMA_signal_15385 ;
    wire new_AGEMA_signal_15386 ;
    wire new_AGEMA_signal_15387 ;
    wire new_AGEMA_signal_15388 ;
    wire new_AGEMA_signal_15389 ;
    wire new_AGEMA_signal_15390 ;
    wire new_AGEMA_signal_15391 ;
    wire new_AGEMA_signal_15392 ;
    wire new_AGEMA_signal_15393 ;
    wire new_AGEMA_signal_15394 ;
    wire new_AGEMA_signal_15395 ;
    wire new_AGEMA_signal_15396 ;
    wire new_AGEMA_signal_15397 ;
    wire new_AGEMA_signal_15398 ;
    wire new_AGEMA_signal_15399 ;
    wire new_AGEMA_signal_15400 ;
    wire new_AGEMA_signal_15401 ;
    wire new_AGEMA_signal_15402 ;
    wire new_AGEMA_signal_15403 ;
    wire new_AGEMA_signal_15404 ;
    wire new_AGEMA_signal_15405 ;
    wire new_AGEMA_signal_15406 ;
    wire new_AGEMA_signal_15407 ;
    wire new_AGEMA_signal_15408 ;
    wire new_AGEMA_signal_15409 ;
    wire new_AGEMA_signal_15410 ;
    wire new_AGEMA_signal_15411 ;
    wire new_AGEMA_signal_15412 ;
    wire new_AGEMA_signal_15413 ;
    wire new_AGEMA_signal_15414 ;
    wire new_AGEMA_signal_15415 ;
    wire new_AGEMA_signal_15416 ;
    wire new_AGEMA_signal_15417 ;
    wire new_AGEMA_signal_15418 ;
    wire new_AGEMA_signal_15419 ;
    wire new_AGEMA_signal_15420 ;
    wire new_AGEMA_signal_15421 ;
    wire new_AGEMA_signal_15422 ;
    wire new_AGEMA_signal_15423 ;
    wire new_AGEMA_signal_15424 ;
    wire new_AGEMA_signal_15425 ;
    wire new_AGEMA_signal_15426 ;
    wire new_AGEMA_signal_15427 ;
    wire new_AGEMA_signal_15428 ;
    wire new_AGEMA_signal_15429 ;
    wire new_AGEMA_signal_15430 ;
    wire new_AGEMA_signal_15431 ;
    wire new_AGEMA_signal_15432 ;
    wire new_AGEMA_signal_15433 ;
    wire new_AGEMA_signal_15434 ;
    wire new_AGEMA_signal_15435 ;
    wire new_AGEMA_signal_15436 ;
    wire new_AGEMA_signal_15437 ;
    wire new_AGEMA_signal_15438 ;
    wire new_AGEMA_signal_15439 ;
    wire new_AGEMA_signal_15440 ;
    wire new_AGEMA_signal_15441 ;
    wire new_AGEMA_signal_15442 ;
    wire new_AGEMA_signal_15443 ;
    wire new_AGEMA_signal_15444 ;
    wire new_AGEMA_signal_15445 ;
    wire new_AGEMA_signal_15446 ;
    wire new_AGEMA_signal_15447 ;
    wire new_AGEMA_signal_15448 ;
    wire new_AGEMA_signal_15449 ;
    wire new_AGEMA_signal_15450 ;
    wire new_AGEMA_signal_15451 ;
    wire new_AGEMA_signal_15452 ;
    wire new_AGEMA_signal_15453 ;
    wire new_AGEMA_signal_15454 ;
    wire new_AGEMA_signal_15455 ;
    wire new_AGEMA_signal_15456 ;
    wire new_AGEMA_signal_15457 ;
    wire new_AGEMA_signal_15458 ;
    wire new_AGEMA_signal_15459 ;
    wire new_AGEMA_signal_15460 ;
    wire new_AGEMA_signal_15461 ;
    wire new_AGEMA_signal_15462 ;
    wire new_AGEMA_signal_15463 ;
    wire new_AGEMA_signal_15464 ;
    wire new_AGEMA_signal_15465 ;
    wire new_AGEMA_signal_15466 ;
    wire new_AGEMA_signal_15467 ;
    wire new_AGEMA_signal_15468 ;
    wire new_AGEMA_signal_15469 ;
    wire new_AGEMA_signal_15470 ;
    wire new_AGEMA_signal_15471 ;
    wire new_AGEMA_signal_15472 ;
    wire new_AGEMA_signal_15473 ;
    wire new_AGEMA_signal_15474 ;
    wire new_AGEMA_signal_15475 ;
    wire new_AGEMA_signal_15476 ;
    wire new_AGEMA_signal_15477 ;
    wire new_AGEMA_signal_15478 ;
    wire new_AGEMA_signal_15479 ;
    wire new_AGEMA_signal_15480 ;
    wire new_AGEMA_signal_15481 ;
    wire new_AGEMA_signal_15482 ;
    wire new_AGEMA_signal_15483 ;
    wire new_AGEMA_signal_15484 ;
    wire new_AGEMA_signal_15485 ;
    wire new_AGEMA_signal_15486 ;
    wire new_AGEMA_signal_15487 ;
    wire new_AGEMA_signal_15488 ;
    wire new_AGEMA_signal_15489 ;
    wire new_AGEMA_signal_15490 ;
    wire new_AGEMA_signal_15491 ;
    wire new_AGEMA_signal_15492 ;
    wire new_AGEMA_signal_15493 ;
    wire new_AGEMA_signal_15494 ;
    wire new_AGEMA_signal_15495 ;
    wire new_AGEMA_signal_15496 ;
    wire new_AGEMA_signal_15497 ;
    wire new_AGEMA_signal_15498 ;
    wire new_AGEMA_signal_15499 ;
    wire new_AGEMA_signal_15500 ;
    wire new_AGEMA_signal_15501 ;
    wire new_AGEMA_signal_15502 ;
    wire new_AGEMA_signal_15503 ;
    wire new_AGEMA_signal_15504 ;
    wire new_AGEMA_signal_15505 ;
    wire new_AGEMA_signal_15506 ;
    wire new_AGEMA_signal_15507 ;
    wire new_AGEMA_signal_15508 ;
    wire new_AGEMA_signal_15509 ;
    wire new_AGEMA_signal_15510 ;
    wire new_AGEMA_signal_15511 ;
    wire new_AGEMA_signal_15512 ;
    wire new_AGEMA_signal_15513 ;
    wire new_AGEMA_signal_15514 ;
    wire new_AGEMA_signal_15515 ;
    wire new_AGEMA_signal_15516 ;
    wire new_AGEMA_signal_15517 ;
    wire new_AGEMA_signal_15518 ;
    wire new_AGEMA_signal_15519 ;
    wire new_AGEMA_signal_15520 ;
    wire new_AGEMA_signal_15521 ;
    wire new_AGEMA_signal_15522 ;
    wire new_AGEMA_signal_15523 ;
    wire new_AGEMA_signal_15524 ;
    wire new_AGEMA_signal_15525 ;
    wire new_AGEMA_signal_15526 ;
    wire new_AGEMA_signal_15527 ;
    wire new_AGEMA_signal_15528 ;
    wire new_AGEMA_signal_15529 ;
    wire new_AGEMA_signal_15530 ;
    wire new_AGEMA_signal_15531 ;
    wire new_AGEMA_signal_15532 ;
    wire new_AGEMA_signal_15533 ;
    wire new_AGEMA_signal_15534 ;
    wire new_AGEMA_signal_15535 ;
    wire new_AGEMA_signal_15536 ;
    wire new_AGEMA_signal_15537 ;
    wire new_AGEMA_signal_15538 ;
    wire new_AGEMA_signal_15539 ;
    wire new_AGEMA_signal_15540 ;
    wire new_AGEMA_signal_15541 ;
    wire new_AGEMA_signal_15542 ;
    wire new_AGEMA_signal_15543 ;
    wire new_AGEMA_signal_15544 ;
    wire new_AGEMA_signal_15545 ;
    wire new_AGEMA_signal_15546 ;
    wire new_AGEMA_signal_15547 ;
    wire new_AGEMA_signal_15548 ;
    wire new_AGEMA_signal_15549 ;
    wire new_AGEMA_signal_15550 ;
    wire new_AGEMA_signal_15551 ;
    wire new_AGEMA_signal_15552 ;
    wire new_AGEMA_signal_15553 ;
    wire new_AGEMA_signal_15554 ;
    wire new_AGEMA_signal_15555 ;
    wire new_AGEMA_signal_15556 ;
    wire new_AGEMA_signal_15557 ;
    wire new_AGEMA_signal_15558 ;
    wire new_AGEMA_signal_15559 ;
    wire new_AGEMA_signal_15560 ;
    wire new_AGEMA_signal_15561 ;
    wire new_AGEMA_signal_15562 ;
    wire new_AGEMA_signal_15563 ;
    wire new_AGEMA_signal_15564 ;
    wire new_AGEMA_signal_15565 ;
    wire new_AGEMA_signal_15566 ;
    wire new_AGEMA_signal_15567 ;
    wire new_AGEMA_signal_15568 ;
    wire new_AGEMA_signal_15569 ;
    wire new_AGEMA_signal_15570 ;
    wire new_AGEMA_signal_15571 ;
    wire new_AGEMA_signal_15572 ;
    wire new_AGEMA_signal_15573 ;
    wire new_AGEMA_signal_15574 ;
    wire new_AGEMA_signal_15575 ;
    wire new_AGEMA_signal_15576 ;
    wire new_AGEMA_signal_15577 ;
    wire new_AGEMA_signal_15578 ;
    wire new_AGEMA_signal_15579 ;
    wire new_AGEMA_signal_15580 ;
    wire new_AGEMA_signal_15581 ;
    wire new_AGEMA_signal_15582 ;
    wire new_AGEMA_signal_15583 ;
    wire new_AGEMA_signal_15584 ;
    wire new_AGEMA_signal_15585 ;
    wire new_AGEMA_signal_15586 ;
    wire new_AGEMA_signal_15587 ;
    wire new_AGEMA_signal_15588 ;
    wire new_AGEMA_signal_15589 ;
    wire new_AGEMA_signal_15590 ;
    wire new_AGEMA_signal_15591 ;
    wire new_AGEMA_signal_15592 ;
    wire new_AGEMA_signal_15593 ;
    wire new_AGEMA_signal_15594 ;
    wire new_AGEMA_signal_15595 ;
    wire new_AGEMA_signal_15596 ;
    wire new_AGEMA_signal_15597 ;
    wire new_AGEMA_signal_15598 ;
    wire new_AGEMA_signal_15599 ;
    wire new_AGEMA_signal_15600 ;
    wire new_AGEMA_signal_15601 ;
    wire new_AGEMA_signal_15602 ;
    wire new_AGEMA_signal_15603 ;
    wire new_AGEMA_signal_15604 ;
    wire new_AGEMA_signal_15605 ;
    wire new_AGEMA_signal_15606 ;
    wire new_AGEMA_signal_15607 ;
    wire new_AGEMA_signal_15608 ;
    wire new_AGEMA_signal_15609 ;
    wire new_AGEMA_signal_15610 ;
    wire new_AGEMA_signal_15611 ;
    wire new_AGEMA_signal_15612 ;
    wire new_AGEMA_signal_15613 ;
    wire new_AGEMA_signal_15614 ;
    wire new_AGEMA_signal_15615 ;
    wire new_AGEMA_signal_15616 ;
    wire new_AGEMA_signal_15617 ;
    wire new_AGEMA_signal_15618 ;
    wire new_AGEMA_signal_15619 ;
    wire new_AGEMA_signal_15620 ;
    wire new_AGEMA_signal_15621 ;
    wire new_AGEMA_signal_15622 ;
    wire new_AGEMA_signal_15623 ;
    wire new_AGEMA_signal_15624 ;
    wire new_AGEMA_signal_15625 ;
    wire new_AGEMA_signal_15626 ;
    wire new_AGEMA_signal_15627 ;
    wire new_AGEMA_signal_15628 ;
    wire new_AGEMA_signal_15629 ;
    wire new_AGEMA_signal_15630 ;
    wire new_AGEMA_signal_15631 ;
    wire new_AGEMA_signal_15632 ;
    wire new_AGEMA_signal_15633 ;
    wire new_AGEMA_signal_15634 ;
    wire new_AGEMA_signal_15635 ;
    wire new_AGEMA_signal_15636 ;
    wire new_AGEMA_signal_15637 ;
    wire new_AGEMA_signal_15638 ;
    wire new_AGEMA_signal_15639 ;
    wire new_AGEMA_signal_15640 ;
    wire new_AGEMA_signal_15641 ;
    wire new_AGEMA_signal_15642 ;
    wire new_AGEMA_signal_15643 ;
    wire new_AGEMA_signal_15644 ;
    wire new_AGEMA_signal_15645 ;
    wire new_AGEMA_signal_15646 ;
    wire new_AGEMA_signal_15647 ;
    wire new_AGEMA_signal_15648 ;
    wire new_AGEMA_signal_15649 ;
    wire new_AGEMA_signal_15650 ;
    wire new_AGEMA_signal_15651 ;
    wire new_AGEMA_signal_15652 ;
    wire new_AGEMA_signal_15653 ;
    wire new_AGEMA_signal_15654 ;
    wire new_AGEMA_signal_15655 ;
    wire new_AGEMA_signal_15656 ;
    wire new_AGEMA_signal_15657 ;
    wire new_AGEMA_signal_15658 ;
    wire new_AGEMA_signal_15659 ;
    wire new_AGEMA_signal_15660 ;
    wire new_AGEMA_signal_15661 ;
    wire new_AGEMA_signal_15662 ;
    wire new_AGEMA_signal_15663 ;
    wire new_AGEMA_signal_15664 ;
    wire new_AGEMA_signal_15665 ;
    wire new_AGEMA_signal_15666 ;
    wire new_AGEMA_signal_15667 ;
    wire new_AGEMA_signal_15668 ;
    wire new_AGEMA_signal_15669 ;
    wire new_AGEMA_signal_15670 ;
    wire new_AGEMA_signal_15671 ;
    wire new_AGEMA_signal_15672 ;
    wire new_AGEMA_signal_15673 ;
    wire new_AGEMA_signal_15674 ;
    wire new_AGEMA_signal_15675 ;
    wire new_AGEMA_signal_15676 ;
    wire new_AGEMA_signal_15677 ;
    wire new_AGEMA_signal_15678 ;
    wire new_AGEMA_signal_15679 ;
    wire new_AGEMA_signal_15680 ;
    wire new_AGEMA_signal_15681 ;
    wire new_AGEMA_signal_15682 ;
    wire new_AGEMA_signal_15683 ;
    wire new_AGEMA_signal_15684 ;
    wire new_AGEMA_signal_15685 ;
    wire new_AGEMA_signal_15686 ;
    wire new_AGEMA_signal_15687 ;
    wire new_AGEMA_signal_15688 ;
    wire new_AGEMA_signal_15689 ;
    wire new_AGEMA_signal_15690 ;
    wire new_AGEMA_signal_15691 ;
    wire new_AGEMA_signal_15692 ;
    wire new_AGEMA_signal_15693 ;
    wire new_AGEMA_signal_15694 ;
    wire new_AGEMA_signal_15695 ;
    wire new_AGEMA_signal_15696 ;
    wire new_AGEMA_signal_15697 ;
    wire new_AGEMA_signal_15698 ;
    wire new_AGEMA_signal_15699 ;
    wire new_AGEMA_signal_15700 ;
    wire new_AGEMA_signal_15701 ;
    wire new_AGEMA_signal_15702 ;
    wire new_AGEMA_signal_15703 ;
    wire new_AGEMA_signal_15704 ;
    wire new_AGEMA_signal_15705 ;
    wire new_AGEMA_signal_15706 ;
    wire new_AGEMA_signal_15707 ;
    wire new_AGEMA_signal_15708 ;
    wire new_AGEMA_signal_15709 ;
    wire new_AGEMA_signal_15710 ;
    wire new_AGEMA_signal_15711 ;
    wire new_AGEMA_signal_15712 ;
    wire new_AGEMA_signal_15713 ;
    wire new_AGEMA_signal_15714 ;
    wire new_AGEMA_signal_15715 ;
    wire new_AGEMA_signal_15716 ;
    wire new_AGEMA_signal_15717 ;
    wire new_AGEMA_signal_15718 ;
    wire new_AGEMA_signal_15719 ;
    wire new_AGEMA_signal_15720 ;
    wire new_AGEMA_signal_15721 ;
    wire new_AGEMA_signal_15722 ;
    wire new_AGEMA_signal_15723 ;
    wire new_AGEMA_signal_15724 ;
    wire new_AGEMA_signal_15725 ;
    wire new_AGEMA_signal_15726 ;
    wire new_AGEMA_signal_15727 ;
    wire new_AGEMA_signal_15728 ;
    wire new_AGEMA_signal_15729 ;
    wire new_AGEMA_signal_15730 ;
    wire new_AGEMA_signal_15731 ;
    wire new_AGEMA_signal_15732 ;
    wire new_AGEMA_signal_15733 ;
    wire new_AGEMA_signal_15734 ;
    wire new_AGEMA_signal_15735 ;
    wire new_AGEMA_signal_15736 ;
    wire new_AGEMA_signal_15737 ;
    wire new_AGEMA_signal_15738 ;
    wire new_AGEMA_signal_15739 ;
    wire new_AGEMA_signal_15740 ;
    wire new_AGEMA_signal_15741 ;
    wire new_AGEMA_signal_15742 ;
    wire new_AGEMA_signal_15743 ;
    wire new_AGEMA_signal_15744 ;
    wire new_AGEMA_signal_15745 ;
    wire new_AGEMA_signal_15746 ;
    wire new_AGEMA_signal_15747 ;
    wire new_AGEMA_signal_15748 ;
    wire new_AGEMA_signal_15749 ;
    wire new_AGEMA_signal_15750 ;
    wire new_AGEMA_signal_15751 ;
    wire new_AGEMA_signal_15752 ;
    wire new_AGEMA_signal_15753 ;
    wire new_AGEMA_signal_15754 ;
    wire new_AGEMA_signal_15755 ;
    wire new_AGEMA_signal_15756 ;
    wire new_AGEMA_signal_15757 ;
    wire new_AGEMA_signal_15758 ;
    wire new_AGEMA_signal_15759 ;
    wire new_AGEMA_signal_15760 ;
    wire new_AGEMA_signal_15761 ;
    wire new_AGEMA_signal_15762 ;
    wire new_AGEMA_signal_15763 ;
    wire new_AGEMA_signal_15764 ;
    wire new_AGEMA_signal_15765 ;
    wire new_AGEMA_signal_15766 ;
    wire new_AGEMA_signal_15767 ;
    wire new_AGEMA_signal_15768 ;
    wire new_AGEMA_signal_15769 ;
    wire new_AGEMA_signal_15770 ;
    wire new_AGEMA_signal_15771 ;
    wire new_AGEMA_signal_15772 ;
    wire new_AGEMA_signal_15773 ;
    wire new_AGEMA_signal_15774 ;
    wire new_AGEMA_signal_15775 ;
    wire new_AGEMA_signal_15776 ;
    wire new_AGEMA_signal_15777 ;
    wire new_AGEMA_signal_15778 ;
    wire new_AGEMA_signal_15779 ;
    wire new_AGEMA_signal_15780 ;
    wire new_AGEMA_signal_15781 ;
    wire new_AGEMA_signal_15782 ;
    wire new_AGEMA_signal_15783 ;
    wire new_AGEMA_signal_15784 ;
    wire new_AGEMA_signal_15785 ;
    wire new_AGEMA_signal_15786 ;
    wire new_AGEMA_signal_15787 ;
    wire new_AGEMA_signal_15788 ;
    wire new_AGEMA_signal_15789 ;
    wire new_AGEMA_signal_15790 ;
    wire new_AGEMA_signal_15791 ;
    wire new_AGEMA_signal_15792 ;
    wire new_AGEMA_signal_15793 ;
    wire new_AGEMA_signal_15794 ;
    wire new_AGEMA_signal_15795 ;
    wire new_AGEMA_signal_15796 ;
    wire new_AGEMA_signal_15797 ;
    wire new_AGEMA_signal_15798 ;
    wire new_AGEMA_signal_15799 ;
    wire new_AGEMA_signal_15800 ;
    wire new_AGEMA_signal_15801 ;
    wire new_AGEMA_signal_15802 ;
    wire new_AGEMA_signal_15803 ;
    wire new_AGEMA_signal_15804 ;
    wire new_AGEMA_signal_15805 ;
    wire new_AGEMA_signal_15806 ;
    wire new_AGEMA_signal_15807 ;
    wire new_AGEMA_signal_15808 ;
    wire new_AGEMA_signal_15809 ;
    wire new_AGEMA_signal_15810 ;
    wire new_AGEMA_signal_15811 ;
    wire new_AGEMA_signal_15812 ;
    wire new_AGEMA_signal_15813 ;
    wire new_AGEMA_signal_15814 ;
    wire new_AGEMA_signal_15815 ;
    wire new_AGEMA_signal_15816 ;
    wire new_AGEMA_signal_15817 ;
    wire new_AGEMA_signal_15818 ;
    wire new_AGEMA_signal_15819 ;
    wire new_AGEMA_signal_15820 ;
    wire new_AGEMA_signal_15821 ;
    wire new_AGEMA_signal_15822 ;
    wire new_AGEMA_signal_15823 ;
    wire new_AGEMA_signal_15824 ;
    wire new_AGEMA_signal_15825 ;
    wire new_AGEMA_signal_15826 ;
    wire new_AGEMA_signal_15827 ;
    wire new_AGEMA_signal_15828 ;

    /* cells in depth 0 */
    INV_X1 U830 ( .A (n314), .ZN (n319) ) ;
    INV_X1 U831 ( .A (n314), .ZN (n320) ) ;
    INV_X1 U832 ( .A (n314), .ZN (n317) ) ;
    INV_X1 U833 ( .A (n314), .ZN (n315) ) ;
    INV_X1 U834 ( .A (n314), .ZN (n316) ) ;
    INV_X1 U835 ( .A (n314), .ZN (n318) ) ;
    NOR2_X1 U836 ( .A1 (n325), .A2 (n330), .ZN (n314) ) ;
    INV_X1 U837 ( .A (RoundCounter[0]), .ZN (n325) ) ;
    INV_X1 U838 ( .A (n314), .ZN (n321) ) ;
    NOR2_X1 U839 ( .A1 (RoundCounter[2]), .A2 (RoundCounter[1]), .ZN (n323) ) ;
    INV_X1 U840 ( .A (n323), .ZN (n322) ) ;
    NOR2_X1 U841 ( .A1 (RoundCounter[0]), .A2 (n322), .ZN (Rcon[0]) ) ;
    NOR2_X1 U842 ( .A1 (RoundCounter[0]), .A2 (RoundCounter[3]), .ZN (n337) ) ;
    NOR2_X1 U843 ( .A1 (n337), .A2 (n322), .ZN (Rcon[1]) ) ;
    NAND2_X1 U844 ( .A1 (RoundCounter[3]), .A2 (n323), .ZN (n330) ) ;
    INV_X1 U845 ( .A (RoundCounter[2]), .ZN (n328) ) ;
    AND2_X1 U846 ( .A1 (n328), .A2 (RoundCounter[1]), .ZN (n333) ) ;
    NAND2_X1 U847 ( .A1 (n337), .A2 (n333), .ZN (n324) ) ;
    NAND2_X1 U848 ( .A1 (n321), .A2 (n324), .ZN (Rcon[2]) ) ;
    NOR2_X1 U849 ( .A1 (RoundCounter[3]), .A2 (n325), .ZN (n335) ) ;
    NAND2_X1 U850 ( .A1 (n333), .A2 (n335), .ZN (n327) ) ;
    NAND2_X1 U851 ( .A1 (RoundCounter[3]), .A2 (Rcon[0]), .ZN (n326) ) ;
    NAND2_X1 U852 ( .A1 (n327), .A2 (n326), .ZN (Rcon[3]) ) ;
    NOR2_X1 U853 ( .A1 (RoundCounter[1]), .A2 (n328), .ZN (n331) ) ;
    NAND2_X1 U854 ( .A1 (n337), .A2 (n331), .ZN (n329) ) ;
    NAND2_X1 U855 ( .A1 (n330), .A2 (n329), .ZN (Rcon[4]) ) ;
    NAND2_X1 U856 ( .A1 (n335), .A2 (n331), .ZN (n332) ) ;
    NAND2_X1 U857 ( .A1 (n321), .A2 (n332), .ZN (Rcon[5]) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U986 ( .a ({new_AGEMA_signal_4549, RoundInput[0]}), .b ({new_AGEMA_signal_4550, RoundKey[0]}), .c ({ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U987 ( .a ({new_AGEMA_signal_4552, RoundInput[100]}), .b ({new_AGEMA_signal_4553, RoundKey[100]}), .c ({ciphertext_s1[100], ciphertext_s0[100]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U988 ( .a ({new_AGEMA_signal_4555, RoundInput[101]}), .b ({new_AGEMA_signal_4556, RoundKey[101]}), .c ({ciphertext_s1[101], ciphertext_s0[101]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U989 ( .a ({new_AGEMA_signal_4558, RoundInput[102]}), .b ({new_AGEMA_signal_4559, RoundKey[102]}), .c ({ciphertext_s1[102], ciphertext_s0[102]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U990 ( .a ({new_AGEMA_signal_4561, RoundInput[103]}), .b ({new_AGEMA_signal_4562, RoundKey[103]}), .c ({ciphertext_s1[103], ciphertext_s0[103]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U991 ( .a ({new_AGEMA_signal_4564, RoundInput[104]}), .b ({new_AGEMA_signal_4565, RoundKey[104]}), .c ({ciphertext_s1[104], ciphertext_s0[104]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U992 ( .a ({new_AGEMA_signal_4567, RoundInput[105]}), .b ({new_AGEMA_signal_4568, RoundKey[105]}), .c ({ciphertext_s1[105], ciphertext_s0[105]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U993 ( .a ({new_AGEMA_signal_4570, RoundInput[106]}), .b ({new_AGEMA_signal_4571, RoundKey[106]}), .c ({ciphertext_s1[106], ciphertext_s0[106]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U994 ( .a ({new_AGEMA_signal_4573, RoundInput[107]}), .b ({new_AGEMA_signal_4574, RoundKey[107]}), .c ({ciphertext_s1[107], ciphertext_s0[107]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U995 ( .a ({new_AGEMA_signal_4576, RoundInput[108]}), .b ({new_AGEMA_signal_4577, RoundKey[108]}), .c ({ciphertext_s1[108], ciphertext_s0[108]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U996 ( .a ({new_AGEMA_signal_4579, RoundInput[109]}), .b ({new_AGEMA_signal_4580, RoundKey[109]}), .c ({ciphertext_s1[109], ciphertext_s0[109]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U997 ( .a ({new_AGEMA_signal_4582, RoundInput[10]}), .b ({new_AGEMA_signal_4583, RoundKey[10]}), .c ({ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U998 ( .a ({new_AGEMA_signal_4585, RoundInput[110]}), .b ({new_AGEMA_signal_4586, RoundKey[110]}), .c ({ciphertext_s1[110], ciphertext_s0[110]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U999 ( .a ({new_AGEMA_signal_4588, RoundInput[111]}), .b ({new_AGEMA_signal_4589, RoundKey[111]}), .c ({ciphertext_s1[111], ciphertext_s0[111]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1000 ( .a ({new_AGEMA_signal_4591, RoundInput[112]}), .b ({new_AGEMA_signal_4592, RoundKey[112]}), .c ({ciphertext_s1[112], ciphertext_s0[112]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1001 ( .a ({new_AGEMA_signal_4594, RoundInput[113]}), .b ({new_AGEMA_signal_4595, RoundKey[113]}), .c ({ciphertext_s1[113], ciphertext_s0[113]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1002 ( .a ({new_AGEMA_signal_4597, RoundInput[114]}), .b ({new_AGEMA_signal_4598, RoundKey[114]}), .c ({ciphertext_s1[114], ciphertext_s0[114]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1003 ( .a ({new_AGEMA_signal_4600, RoundInput[115]}), .b ({new_AGEMA_signal_4601, RoundKey[115]}), .c ({ciphertext_s1[115], ciphertext_s0[115]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1004 ( .a ({new_AGEMA_signal_4603, RoundInput[116]}), .b ({new_AGEMA_signal_4604, RoundKey[116]}), .c ({ciphertext_s1[116], ciphertext_s0[116]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1005 ( .a ({new_AGEMA_signal_4606, RoundInput[117]}), .b ({new_AGEMA_signal_4607, RoundKey[117]}), .c ({ciphertext_s1[117], ciphertext_s0[117]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1006 ( .a ({new_AGEMA_signal_4609, RoundInput[118]}), .b ({new_AGEMA_signal_4610, RoundKey[118]}), .c ({ciphertext_s1[118], ciphertext_s0[118]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1007 ( .a ({new_AGEMA_signal_4612, RoundInput[119]}), .b ({new_AGEMA_signal_4613, RoundKey[119]}), .c ({ciphertext_s1[119], ciphertext_s0[119]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1008 ( .a ({new_AGEMA_signal_4615, RoundInput[11]}), .b ({new_AGEMA_signal_4616, RoundKey[11]}), .c ({ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1009 ( .a ({new_AGEMA_signal_4618, RoundInput[120]}), .b ({new_AGEMA_signal_4619, RoundKey[120]}), .c ({ciphertext_s1[120], ciphertext_s0[120]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1010 ( .a ({new_AGEMA_signal_4621, RoundInput[121]}), .b ({new_AGEMA_signal_4622, RoundKey[121]}), .c ({ciphertext_s1[121], ciphertext_s0[121]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1011 ( .a ({new_AGEMA_signal_4624, RoundInput[122]}), .b ({new_AGEMA_signal_4625, RoundKey[122]}), .c ({ciphertext_s1[122], ciphertext_s0[122]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1012 ( .a ({new_AGEMA_signal_4627, RoundInput[123]}), .b ({new_AGEMA_signal_4628, RoundKey[123]}), .c ({ciphertext_s1[123], ciphertext_s0[123]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1013 ( .a ({new_AGEMA_signal_4630, RoundInput[124]}), .b ({new_AGEMA_signal_4631, RoundKey[124]}), .c ({ciphertext_s1[124], ciphertext_s0[124]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1014 ( .a ({new_AGEMA_signal_4633, RoundInput[125]}), .b ({new_AGEMA_signal_4634, RoundKey[125]}), .c ({ciphertext_s1[125], ciphertext_s0[125]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1015 ( .a ({new_AGEMA_signal_4636, RoundInput[126]}), .b ({new_AGEMA_signal_4637, RoundKey[126]}), .c ({ciphertext_s1[126], ciphertext_s0[126]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1016 ( .a ({new_AGEMA_signal_4639, RoundInput[127]}), .b ({new_AGEMA_signal_4640, RoundKey[127]}), .c ({ciphertext_s1[127], ciphertext_s0[127]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1017 ( .a ({new_AGEMA_signal_4642, RoundInput[12]}), .b ({new_AGEMA_signal_4643, RoundKey[12]}), .c ({ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1018 ( .a ({new_AGEMA_signal_4645, RoundInput[13]}), .b ({new_AGEMA_signal_4646, RoundKey[13]}), .c ({ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1019 ( .a ({new_AGEMA_signal_4648, RoundInput[14]}), .b ({new_AGEMA_signal_4649, RoundKey[14]}), .c ({ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1020 ( .a ({new_AGEMA_signal_4651, RoundInput[15]}), .b ({new_AGEMA_signal_4652, RoundKey[15]}), .c ({ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1021 ( .a ({new_AGEMA_signal_4654, RoundInput[16]}), .b ({new_AGEMA_signal_4655, RoundKey[16]}), .c ({ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1022 ( .a ({new_AGEMA_signal_4657, RoundInput[17]}), .b ({new_AGEMA_signal_4658, RoundKey[17]}), .c ({ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1023 ( .a ({new_AGEMA_signal_4660, RoundInput[18]}), .b ({new_AGEMA_signal_4661, RoundKey[18]}), .c ({ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1024 ( .a ({new_AGEMA_signal_4663, RoundInput[19]}), .b ({new_AGEMA_signal_4664, RoundKey[19]}), .c ({ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1025 ( .a ({new_AGEMA_signal_4666, RoundInput[1]}), .b ({new_AGEMA_signal_4667, RoundKey[1]}), .c ({ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1026 ( .a ({new_AGEMA_signal_4669, RoundInput[20]}), .b ({new_AGEMA_signal_4670, RoundKey[20]}), .c ({ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1027 ( .a ({new_AGEMA_signal_4672, RoundInput[21]}), .b ({new_AGEMA_signal_4673, RoundKey[21]}), .c ({ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1028 ( .a ({new_AGEMA_signal_4675, RoundInput[22]}), .b ({new_AGEMA_signal_4676, RoundKey[22]}), .c ({ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1029 ( .a ({new_AGEMA_signal_4678, RoundInput[23]}), .b ({new_AGEMA_signal_4679, RoundKey[23]}), .c ({ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1030 ( .a ({new_AGEMA_signal_4681, RoundInput[24]}), .b ({new_AGEMA_signal_4682, RoundKey[24]}), .c ({ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1031 ( .a ({new_AGEMA_signal_4684, RoundInput[25]}), .b ({new_AGEMA_signal_4685, RoundKey[25]}), .c ({ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1032 ( .a ({new_AGEMA_signal_4687, RoundInput[26]}), .b ({new_AGEMA_signal_4688, RoundKey[26]}), .c ({ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1033 ( .a ({new_AGEMA_signal_4690, RoundInput[27]}), .b ({new_AGEMA_signal_4691, RoundKey[27]}), .c ({ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1034 ( .a ({new_AGEMA_signal_4693, RoundInput[28]}), .b ({new_AGEMA_signal_4694, RoundKey[28]}), .c ({ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1035 ( .a ({new_AGEMA_signal_4696, RoundInput[29]}), .b ({new_AGEMA_signal_4697, RoundKey[29]}), .c ({ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1036 ( .a ({new_AGEMA_signal_4699, RoundInput[2]}), .b ({new_AGEMA_signal_4700, RoundKey[2]}), .c ({ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1037 ( .a ({new_AGEMA_signal_4702, RoundInput[30]}), .b ({new_AGEMA_signal_4703, RoundKey[30]}), .c ({ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1038 ( .a ({new_AGEMA_signal_4705, RoundInput[31]}), .b ({new_AGEMA_signal_4706, RoundKey[31]}), .c ({ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1039 ( .a ({new_AGEMA_signal_4708, RoundInput[32]}), .b ({new_AGEMA_signal_4709, RoundKey[32]}), .c ({ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1040 ( .a ({new_AGEMA_signal_4711, RoundInput[33]}), .b ({new_AGEMA_signal_4712, RoundKey[33]}), .c ({ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1041 ( .a ({new_AGEMA_signal_4714, RoundInput[34]}), .b ({new_AGEMA_signal_4715, RoundKey[34]}), .c ({ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1042 ( .a ({new_AGEMA_signal_4717, RoundInput[35]}), .b ({new_AGEMA_signal_4718, RoundKey[35]}), .c ({ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1043 ( .a ({new_AGEMA_signal_4720, RoundInput[36]}), .b ({new_AGEMA_signal_4721, RoundKey[36]}), .c ({ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1044 ( .a ({new_AGEMA_signal_4723, RoundInput[37]}), .b ({new_AGEMA_signal_4724, RoundKey[37]}), .c ({ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1045 ( .a ({new_AGEMA_signal_4726, RoundInput[38]}), .b ({new_AGEMA_signal_4727, RoundKey[38]}), .c ({ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1046 ( .a ({new_AGEMA_signal_4729, RoundInput[39]}), .b ({new_AGEMA_signal_4730, RoundKey[39]}), .c ({ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1047 ( .a ({new_AGEMA_signal_4732, RoundInput[3]}), .b ({new_AGEMA_signal_4733, RoundKey[3]}), .c ({ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1048 ( .a ({new_AGEMA_signal_4735, RoundInput[40]}), .b ({new_AGEMA_signal_4736, RoundKey[40]}), .c ({ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1049 ( .a ({new_AGEMA_signal_4738, RoundInput[41]}), .b ({new_AGEMA_signal_4739, RoundKey[41]}), .c ({ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1050 ( .a ({new_AGEMA_signal_4741, RoundInput[42]}), .b ({new_AGEMA_signal_4742, RoundKey[42]}), .c ({ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1051 ( .a ({new_AGEMA_signal_4744, RoundInput[43]}), .b ({new_AGEMA_signal_4745, RoundKey[43]}), .c ({ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1052 ( .a ({new_AGEMA_signal_4747, RoundInput[44]}), .b ({new_AGEMA_signal_4748, RoundKey[44]}), .c ({ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1053 ( .a ({new_AGEMA_signal_4750, RoundInput[45]}), .b ({new_AGEMA_signal_4751, RoundKey[45]}), .c ({ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1054 ( .a ({new_AGEMA_signal_4753, RoundInput[46]}), .b ({new_AGEMA_signal_4754, RoundKey[46]}), .c ({ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1055 ( .a ({new_AGEMA_signal_4756, RoundInput[47]}), .b ({new_AGEMA_signal_4757, RoundKey[47]}), .c ({ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1056 ( .a ({new_AGEMA_signal_4759, RoundInput[48]}), .b ({new_AGEMA_signal_4760, RoundKey[48]}), .c ({ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1057 ( .a ({new_AGEMA_signal_4762, RoundInput[49]}), .b ({new_AGEMA_signal_4763, RoundKey[49]}), .c ({ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1058 ( .a ({new_AGEMA_signal_4765, RoundInput[4]}), .b ({new_AGEMA_signal_4766, RoundKey[4]}), .c ({ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1059 ( .a ({new_AGEMA_signal_4768, RoundInput[50]}), .b ({new_AGEMA_signal_4769, RoundKey[50]}), .c ({ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1060 ( .a ({new_AGEMA_signal_4771, RoundInput[51]}), .b ({new_AGEMA_signal_4772, RoundKey[51]}), .c ({ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1061 ( .a ({new_AGEMA_signal_4774, RoundInput[52]}), .b ({new_AGEMA_signal_4775, RoundKey[52]}), .c ({ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1062 ( .a ({new_AGEMA_signal_4777, RoundInput[53]}), .b ({new_AGEMA_signal_4778, RoundKey[53]}), .c ({ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1063 ( .a ({new_AGEMA_signal_4780, RoundInput[54]}), .b ({new_AGEMA_signal_4781, RoundKey[54]}), .c ({ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1064 ( .a ({new_AGEMA_signal_4783, RoundInput[55]}), .b ({new_AGEMA_signal_4784, RoundKey[55]}), .c ({ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1065 ( .a ({new_AGEMA_signal_4786, RoundInput[56]}), .b ({new_AGEMA_signal_4787, RoundKey[56]}), .c ({ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1066 ( .a ({new_AGEMA_signal_4789, RoundInput[57]}), .b ({new_AGEMA_signal_4790, RoundKey[57]}), .c ({ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1067 ( .a ({new_AGEMA_signal_4792, RoundInput[58]}), .b ({new_AGEMA_signal_4793, RoundKey[58]}), .c ({ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1068 ( .a ({new_AGEMA_signal_4795, RoundInput[59]}), .b ({new_AGEMA_signal_4796, RoundKey[59]}), .c ({ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1069 ( .a ({new_AGEMA_signal_4798, RoundInput[5]}), .b ({new_AGEMA_signal_4799, RoundKey[5]}), .c ({ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1070 ( .a ({new_AGEMA_signal_4801, RoundInput[60]}), .b ({new_AGEMA_signal_4802, RoundKey[60]}), .c ({ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1071 ( .a ({new_AGEMA_signal_4804, RoundInput[61]}), .b ({new_AGEMA_signal_4805, RoundKey[61]}), .c ({ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1072 ( .a ({new_AGEMA_signal_4807, RoundInput[62]}), .b ({new_AGEMA_signal_4808, RoundKey[62]}), .c ({ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1073 ( .a ({new_AGEMA_signal_4810, RoundInput[63]}), .b ({new_AGEMA_signal_4811, RoundKey[63]}), .c ({ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1074 ( .a ({new_AGEMA_signal_4813, RoundInput[64]}), .b ({new_AGEMA_signal_4814, RoundKey[64]}), .c ({ciphertext_s1[64], ciphertext_s0[64]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1075 ( .a ({new_AGEMA_signal_4816, RoundInput[65]}), .b ({new_AGEMA_signal_4817, RoundKey[65]}), .c ({ciphertext_s1[65], ciphertext_s0[65]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1076 ( .a ({new_AGEMA_signal_4819, RoundInput[66]}), .b ({new_AGEMA_signal_4820, RoundKey[66]}), .c ({ciphertext_s1[66], ciphertext_s0[66]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1077 ( .a ({new_AGEMA_signal_4822, RoundInput[67]}), .b ({new_AGEMA_signal_4823, RoundKey[67]}), .c ({ciphertext_s1[67], ciphertext_s0[67]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1078 ( .a ({new_AGEMA_signal_4825, RoundInput[68]}), .b ({new_AGEMA_signal_4826, RoundKey[68]}), .c ({ciphertext_s1[68], ciphertext_s0[68]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1079 ( .a ({new_AGEMA_signal_4828, RoundInput[69]}), .b ({new_AGEMA_signal_4829, RoundKey[69]}), .c ({ciphertext_s1[69], ciphertext_s0[69]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1080 ( .a ({new_AGEMA_signal_4831, RoundInput[6]}), .b ({new_AGEMA_signal_4832, RoundKey[6]}), .c ({ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1081 ( .a ({new_AGEMA_signal_4834, RoundInput[70]}), .b ({new_AGEMA_signal_4835, RoundKey[70]}), .c ({ciphertext_s1[70], ciphertext_s0[70]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1082 ( .a ({new_AGEMA_signal_4837, RoundInput[71]}), .b ({new_AGEMA_signal_4838, RoundKey[71]}), .c ({ciphertext_s1[71], ciphertext_s0[71]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1083 ( .a ({new_AGEMA_signal_4840, RoundInput[72]}), .b ({new_AGEMA_signal_4841, RoundKey[72]}), .c ({ciphertext_s1[72], ciphertext_s0[72]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1084 ( .a ({new_AGEMA_signal_4843, RoundInput[73]}), .b ({new_AGEMA_signal_4844, RoundKey[73]}), .c ({ciphertext_s1[73], ciphertext_s0[73]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1085 ( .a ({new_AGEMA_signal_4846, RoundInput[74]}), .b ({new_AGEMA_signal_4847, RoundKey[74]}), .c ({ciphertext_s1[74], ciphertext_s0[74]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1086 ( .a ({new_AGEMA_signal_4849, RoundInput[75]}), .b ({new_AGEMA_signal_4850, RoundKey[75]}), .c ({ciphertext_s1[75], ciphertext_s0[75]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1087 ( .a ({new_AGEMA_signal_4852, RoundInput[76]}), .b ({new_AGEMA_signal_4853, RoundKey[76]}), .c ({ciphertext_s1[76], ciphertext_s0[76]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1088 ( .a ({new_AGEMA_signal_4855, RoundInput[77]}), .b ({new_AGEMA_signal_4856, RoundKey[77]}), .c ({ciphertext_s1[77], ciphertext_s0[77]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1089 ( .a ({new_AGEMA_signal_4858, RoundInput[78]}), .b ({new_AGEMA_signal_4859, RoundKey[78]}), .c ({ciphertext_s1[78], ciphertext_s0[78]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1090 ( .a ({new_AGEMA_signal_4861, RoundInput[79]}), .b ({new_AGEMA_signal_4862, RoundKey[79]}), .c ({ciphertext_s1[79], ciphertext_s0[79]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1091 ( .a ({new_AGEMA_signal_4864, RoundInput[7]}), .b ({new_AGEMA_signal_4865, RoundKey[7]}), .c ({ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1092 ( .a ({new_AGEMA_signal_4867, RoundInput[80]}), .b ({new_AGEMA_signal_4868, RoundKey[80]}), .c ({ciphertext_s1[80], ciphertext_s0[80]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1093 ( .a ({new_AGEMA_signal_4870, RoundInput[81]}), .b ({new_AGEMA_signal_4871, RoundKey[81]}), .c ({ciphertext_s1[81], ciphertext_s0[81]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1094 ( .a ({new_AGEMA_signal_4873, RoundInput[82]}), .b ({new_AGEMA_signal_4874, RoundKey[82]}), .c ({ciphertext_s1[82], ciphertext_s0[82]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1095 ( .a ({new_AGEMA_signal_4876, RoundInput[83]}), .b ({new_AGEMA_signal_4877, RoundKey[83]}), .c ({ciphertext_s1[83], ciphertext_s0[83]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1096 ( .a ({new_AGEMA_signal_4879, RoundInput[84]}), .b ({new_AGEMA_signal_4880, RoundKey[84]}), .c ({ciphertext_s1[84], ciphertext_s0[84]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1097 ( .a ({new_AGEMA_signal_4882, RoundInput[85]}), .b ({new_AGEMA_signal_4883, RoundKey[85]}), .c ({ciphertext_s1[85], ciphertext_s0[85]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1098 ( .a ({new_AGEMA_signal_4885, RoundInput[86]}), .b ({new_AGEMA_signal_4886, RoundKey[86]}), .c ({ciphertext_s1[86], ciphertext_s0[86]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1099 ( .a ({new_AGEMA_signal_4888, RoundInput[87]}), .b ({new_AGEMA_signal_4889, RoundKey[87]}), .c ({ciphertext_s1[87], ciphertext_s0[87]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1100 ( .a ({new_AGEMA_signal_4891, RoundInput[88]}), .b ({new_AGEMA_signal_4892, RoundKey[88]}), .c ({ciphertext_s1[88], ciphertext_s0[88]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1101 ( .a ({new_AGEMA_signal_4894, RoundInput[89]}), .b ({new_AGEMA_signal_4895, RoundKey[89]}), .c ({ciphertext_s1[89], ciphertext_s0[89]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1102 ( .a ({new_AGEMA_signal_4897, RoundInput[8]}), .b ({new_AGEMA_signal_4898, RoundKey[8]}), .c ({ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1103 ( .a ({new_AGEMA_signal_4900, RoundInput[90]}), .b ({new_AGEMA_signal_4901, RoundKey[90]}), .c ({ciphertext_s1[90], ciphertext_s0[90]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1104 ( .a ({new_AGEMA_signal_4903, RoundInput[91]}), .b ({new_AGEMA_signal_4904, RoundKey[91]}), .c ({ciphertext_s1[91], ciphertext_s0[91]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1105 ( .a ({new_AGEMA_signal_4906, RoundInput[92]}), .b ({new_AGEMA_signal_4907, RoundKey[92]}), .c ({ciphertext_s1[92], ciphertext_s0[92]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1106 ( .a ({new_AGEMA_signal_4909, RoundInput[93]}), .b ({new_AGEMA_signal_4910, RoundKey[93]}), .c ({ciphertext_s1[93], ciphertext_s0[93]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1107 ( .a ({new_AGEMA_signal_4912, RoundInput[94]}), .b ({new_AGEMA_signal_4913, RoundKey[94]}), .c ({ciphertext_s1[94], ciphertext_s0[94]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1108 ( .a ({new_AGEMA_signal_4915, RoundInput[95]}), .b ({new_AGEMA_signal_4916, RoundKey[95]}), .c ({ciphertext_s1[95], ciphertext_s0[95]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1109 ( .a ({new_AGEMA_signal_4918, RoundInput[96]}), .b ({new_AGEMA_signal_4919, RoundKey[96]}), .c ({ciphertext_s1[96], ciphertext_s0[96]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1110 ( .a ({new_AGEMA_signal_4921, RoundInput[97]}), .b ({new_AGEMA_signal_4922, RoundKey[97]}), .c ({ciphertext_s1[97], ciphertext_s0[97]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1111 ( .a ({new_AGEMA_signal_4924, RoundInput[98]}), .b ({new_AGEMA_signal_4925, RoundKey[98]}), .c ({ciphertext_s1[98], ciphertext_s0[98]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1112 ( .a ({new_AGEMA_signal_4927, RoundInput[99]}), .b ({new_AGEMA_signal_4928, RoundKey[99]}), .c ({ciphertext_s1[99], ciphertext_s0[99]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U1113 ( .a ({new_AGEMA_signal_4930, RoundInput[9]}), .b ({new_AGEMA_signal_4931, RoundKey[9]}), .c ({ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    NAND2_X1 U1114 ( .A1 (RoundCounter[3]), .A2 (n333), .ZN (n334) ) ;
    NOR2_X1 U1115 ( .A1 (RoundCounter[0]), .A2 (n334), .ZN (done) ) ;
    INV_X1 U1116 ( .A (n335), .ZN (n336) ) ;
    NAND2_X1 U1117 ( .A1 (RoundCounter[2]), .A2 (RoundCounter[1]), .ZN (n338) ) ;
    NOR2_X1 U1118 ( .A1 (n336), .A2 (n338), .ZN (n283) ) ;
    INV_X1 U1119 ( .A (n337), .ZN (n339) ) ;
    NOR2_X1 U1120 ( .A1 (n339), .A2 (n338), .ZN (n285) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T1_U1 ( .a ({ciphertext_s1[7], ciphertext_s0[7]}), .b ({ciphertext_s1[4], ciphertext_s0[4]}), .c ({new_AGEMA_signal_4973, SubBytesIns_Inst_Sbox_0_T1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T2_U1 ( .a ({ciphertext_s1[7], ciphertext_s0[7]}), .b ({ciphertext_s1[2], ciphertext_s0[2]}), .c ({new_AGEMA_signal_4974, SubBytesIns_Inst_Sbox_0_T2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T3_U1 ( .a ({ciphertext_s1[7], ciphertext_s0[7]}), .b ({ciphertext_s1[1], ciphertext_s0[1]}), .c ({new_AGEMA_signal_4975, SubBytesIns_Inst_Sbox_0_T3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T4_U1 ( .a ({ciphertext_s1[4], ciphertext_s0[4]}), .b ({ciphertext_s1[2], ciphertext_s0[2]}), .c ({new_AGEMA_signal_4976, SubBytesIns_Inst_Sbox_0_T4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T5_U1 ( .a ({ciphertext_s1[3], ciphertext_s0[3]}), .b ({ciphertext_s1[1], ciphertext_s0[1]}), .c ({new_AGEMA_signal_4977, SubBytesIns_Inst_Sbox_0_T5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T6_U1 ( .a ({new_AGEMA_signal_4973, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_4977, SubBytesIns_Inst_Sbox_0_T5}), .c ({new_AGEMA_signal_5165, SubBytesIns_Inst_Sbox_0_T6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T7_U1 ( .a ({ciphertext_s1[6], ciphertext_s0[6]}), .b ({ciphertext_s1[5], ciphertext_s0[5]}), .c ({new_AGEMA_signal_4978, SubBytesIns_Inst_Sbox_0_T7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T8_U1 ( .a ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({new_AGEMA_signal_5165, SubBytesIns_Inst_Sbox_0_T6}), .c ({new_AGEMA_signal_5345, SubBytesIns_Inst_Sbox_0_T8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T9_U1 ( .a ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({new_AGEMA_signal_4978, SubBytesIns_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_5166, SubBytesIns_Inst_Sbox_0_T9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T10_U1 ( .a ({new_AGEMA_signal_5165, SubBytesIns_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_4978, SubBytesIns_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_5346, SubBytesIns_Inst_Sbox_0_T10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T11_U1 ( .a ({ciphertext_s1[6], ciphertext_s0[6]}), .b ({ciphertext_s1[2], ciphertext_s0[2]}), .c ({new_AGEMA_signal_4979, SubBytesIns_Inst_Sbox_0_T11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T12_U1 ( .a ({ciphertext_s1[5], ciphertext_s0[5]}), .b ({ciphertext_s1[2], ciphertext_s0[2]}), .c ({new_AGEMA_signal_4980, SubBytesIns_Inst_Sbox_0_T12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T13_U1 ( .a ({new_AGEMA_signal_4975, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_4976, SubBytesIns_Inst_Sbox_0_T4}), .c ({new_AGEMA_signal_5167, SubBytesIns_Inst_Sbox_0_T13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T14_U1 ( .a ({new_AGEMA_signal_5165, SubBytesIns_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_4979, SubBytesIns_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_5347, SubBytesIns_Inst_Sbox_0_T14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T15_U1 ( .a ({new_AGEMA_signal_4977, SubBytesIns_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_4979, SubBytesIns_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_5168, SubBytesIns_Inst_Sbox_0_T15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T16_U1 ( .a ({new_AGEMA_signal_4977, SubBytesIns_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_4980, SubBytesIns_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_5169, SubBytesIns_Inst_Sbox_0_T16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T17_U1 ( .a ({new_AGEMA_signal_5166, SubBytesIns_Inst_Sbox_0_T9}), .b ({new_AGEMA_signal_5169, SubBytesIns_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_5348, SubBytesIns_Inst_Sbox_0_T17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T18_U1 ( .a ({ciphertext_s1[4], ciphertext_s0[4]}), .b ({ciphertext_s1[0], ciphertext_s0[0]}), .c ({new_AGEMA_signal_4981, SubBytesIns_Inst_Sbox_0_T18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T19_U1 ( .a ({new_AGEMA_signal_4978, SubBytesIns_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_4981, SubBytesIns_Inst_Sbox_0_T18}), .c ({new_AGEMA_signal_5170, SubBytesIns_Inst_Sbox_0_T19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T20_U1 ( .a ({new_AGEMA_signal_4973, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_5170, SubBytesIns_Inst_Sbox_0_T19}), .c ({new_AGEMA_signal_5349, SubBytesIns_Inst_Sbox_0_T20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T21_U1 ( .a ({ciphertext_s1[1], ciphertext_s0[1]}), .b ({ciphertext_s1[0], ciphertext_s0[0]}), .c ({new_AGEMA_signal_4982, SubBytesIns_Inst_Sbox_0_T21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T22_U1 ( .a ({new_AGEMA_signal_4978, SubBytesIns_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_4982, SubBytesIns_Inst_Sbox_0_T21}), .c ({new_AGEMA_signal_5171, SubBytesIns_Inst_Sbox_0_T22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T23_U1 ( .a ({new_AGEMA_signal_4974, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_5171, SubBytesIns_Inst_Sbox_0_T22}), .c ({new_AGEMA_signal_5350, SubBytesIns_Inst_Sbox_0_T23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T24_U1 ( .a ({new_AGEMA_signal_4974, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_5346, SubBytesIns_Inst_Sbox_0_T10}), .c ({new_AGEMA_signal_5589, SubBytesIns_Inst_Sbox_0_T24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T25_U1 ( .a ({new_AGEMA_signal_5349, SubBytesIns_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_5348, SubBytesIns_Inst_Sbox_0_T17}), .c ({new_AGEMA_signal_5590, SubBytesIns_Inst_Sbox_0_T25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T26_U1 ( .a ({new_AGEMA_signal_4975, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_5169, SubBytesIns_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_5351, SubBytesIns_Inst_Sbox_0_T26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T27_U1 ( .a ({new_AGEMA_signal_4973, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_4980, SubBytesIns_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_5172, SubBytesIns_Inst_Sbox_0_T27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T1_U1 ( .a ({ciphertext_s1[15], ciphertext_s0[15]}), .b ({ciphertext_s1[12], ciphertext_s0[12]}), .c ({new_AGEMA_signal_4983, SubBytesIns_Inst_Sbox_1_T1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T2_U1 ( .a ({ciphertext_s1[15], ciphertext_s0[15]}), .b ({ciphertext_s1[10], ciphertext_s0[10]}), .c ({new_AGEMA_signal_4984, SubBytesIns_Inst_Sbox_1_T2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T3_U1 ( .a ({ciphertext_s1[15], ciphertext_s0[15]}), .b ({ciphertext_s1[9], ciphertext_s0[9]}), .c ({new_AGEMA_signal_4985, SubBytesIns_Inst_Sbox_1_T3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T4_U1 ( .a ({ciphertext_s1[12], ciphertext_s0[12]}), .b ({ciphertext_s1[10], ciphertext_s0[10]}), .c ({new_AGEMA_signal_4986, SubBytesIns_Inst_Sbox_1_T4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T5_U1 ( .a ({ciphertext_s1[11], ciphertext_s0[11]}), .b ({ciphertext_s1[9], ciphertext_s0[9]}), .c ({new_AGEMA_signal_4987, SubBytesIns_Inst_Sbox_1_T5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T6_U1 ( .a ({new_AGEMA_signal_4983, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_4987, SubBytesIns_Inst_Sbox_1_T5}), .c ({new_AGEMA_signal_5173, SubBytesIns_Inst_Sbox_1_T6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T7_U1 ( .a ({ciphertext_s1[14], ciphertext_s0[14]}), .b ({ciphertext_s1[13], ciphertext_s0[13]}), .c ({new_AGEMA_signal_4988, SubBytesIns_Inst_Sbox_1_T7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T8_U1 ( .a ({ciphertext_s1[8], ciphertext_s0[8]}), .b ({new_AGEMA_signal_5173, SubBytesIns_Inst_Sbox_1_T6}), .c ({new_AGEMA_signal_5358, SubBytesIns_Inst_Sbox_1_T8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T9_U1 ( .a ({ciphertext_s1[8], ciphertext_s0[8]}), .b ({new_AGEMA_signal_4988, SubBytesIns_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_5174, SubBytesIns_Inst_Sbox_1_T9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T10_U1 ( .a ({new_AGEMA_signal_5173, SubBytesIns_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_4988, SubBytesIns_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_5359, SubBytesIns_Inst_Sbox_1_T10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T11_U1 ( .a ({ciphertext_s1[14], ciphertext_s0[14]}), .b ({ciphertext_s1[10], ciphertext_s0[10]}), .c ({new_AGEMA_signal_4989, SubBytesIns_Inst_Sbox_1_T11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T12_U1 ( .a ({ciphertext_s1[13], ciphertext_s0[13]}), .b ({ciphertext_s1[10], ciphertext_s0[10]}), .c ({new_AGEMA_signal_4990, SubBytesIns_Inst_Sbox_1_T12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T13_U1 ( .a ({new_AGEMA_signal_4985, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_4986, SubBytesIns_Inst_Sbox_1_T4}), .c ({new_AGEMA_signal_5175, SubBytesIns_Inst_Sbox_1_T13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T14_U1 ( .a ({new_AGEMA_signal_5173, SubBytesIns_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_4989, SubBytesIns_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_5360, SubBytesIns_Inst_Sbox_1_T14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T15_U1 ( .a ({new_AGEMA_signal_4987, SubBytesIns_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_4989, SubBytesIns_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_5176, SubBytesIns_Inst_Sbox_1_T15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T16_U1 ( .a ({new_AGEMA_signal_4987, SubBytesIns_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_4990, SubBytesIns_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_5177, SubBytesIns_Inst_Sbox_1_T16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T17_U1 ( .a ({new_AGEMA_signal_5174, SubBytesIns_Inst_Sbox_1_T9}), .b ({new_AGEMA_signal_5177, SubBytesIns_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_5361, SubBytesIns_Inst_Sbox_1_T17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T18_U1 ( .a ({ciphertext_s1[12], ciphertext_s0[12]}), .b ({ciphertext_s1[8], ciphertext_s0[8]}), .c ({new_AGEMA_signal_4991, SubBytesIns_Inst_Sbox_1_T18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T19_U1 ( .a ({new_AGEMA_signal_4988, SubBytesIns_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_4991, SubBytesIns_Inst_Sbox_1_T18}), .c ({new_AGEMA_signal_5178, SubBytesIns_Inst_Sbox_1_T19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T20_U1 ( .a ({new_AGEMA_signal_4983, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_5178, SubBytesIns_Inst_Sbox_1_T19}), .c ({new_AGEMA_signal_5362, SubBytesIns_Inst_Sbox_1_T20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T21_U1 ( .a ({ciphertext_s1[9], ciphertext_s0[9]}), .b ({ciphertext_s1[8], ciphertext_s0[8]}), .c ({new_AGEMA_signal_4992, SubBytesIns_Inst_Sbox_1_T21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T22_U1 ( .a ({new_AGEMA_signal_4988, SubBytesIns_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_4992, SubBytesIns_Inst_Sbox_1_T21}), .c ({new_AGEMA_signal_5179, SubBytesIns_Inst_Sbox_1_T22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T23_U1 ( .a ({new_AGEMA_signal_4984, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_5179, SubBytesIns_Inst_Sbox_1_T22}), .c ({new_AGEMA_signal_5363, SubBytesIns_Inst_Sbox_1_T23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T24_U1 ( .a ({new_AGEMA_signal_4984, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_5359, SubBytesIns_Inst_Sbox_1_T10}), .c ({new_AGEMA_signal_5598, SubBytesIns_Inst_Sbox_1_T24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T25_U1 ( .a ({new_AGEMA_signal_5362, SubBytesIns_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_5361, SubBytesIns_Inst_Sbox_1_T17}), .c ({new_AGEMA_signal_5599, SubBytesIns_Inst_Sbox_1_T25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T26_U1 ( .a ({new_AGEMA_signal_4985, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_5177, SubBytesIns_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_5364, SubBytesIns_Inst_Sbox_1_T26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T27_U1 ( .a ({new_AGEMA_signal_4983, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_4990, SubBytesIns_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_5180, SubBytesIns_Inst_Sbox_1_T27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T1_U1 ( .a ({ciphertext_s1[23], ciphertext_s0[23]}), .b ({ciphertext_s1[20], ciphertext_s0[20]}), .c ({new_AGEMA_signal_4993, SubBytesIns_Inst_Sbox_2_T1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T2_U1 ( .a ({ciphertext_s1[23], ciphertext_s0[23]}), .b ({ciphertext_s1[18], ciphertext_s0[18]}), .c ({new_AGEMA_signal_4994, SubBytesIns_Inst_Sbox_2_T2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T3_U1 ( .a ({ciphertext_s1[23], ciphertext_s0[23]}), .b ({ciphertext_s1[17], ciphertext_s0[17]}), .c ({new_AGEMA_signal_4995, SubBytesIns_Inst_Sbox_2_T3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T4_U1 ( .a ({ciphertext_s1[20], ciphertext_s0[20]}), .b ({ciphertext_s1[18], ciphertext_s0[18]}), .c ({new_AGEMA_signal_4996, SubBytesIns_Inst_Sbox_2_T4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T5_U1 ( .a ({ciphertext_s1[19], ciphertext_s0[19]}), .b ({ciphertext_s1[17], ciphertext_s0[17]}), .c ({new_AGEMA_signal_4997, SubBytesIns_Inst_Sbox_2_T5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T6_U1 ( .a ({new_AGEMA_signal_4993, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_4997, SubBytesIns_Inst_Sbox_2_T5}), .c ({new_AGEMA_signal_5181, SubBytesIns_Inst_Sbox_2_T6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T7_U1 ( .a ({ciphertext_s1[22], ciphertext_s0[22]}), .b ({ciphertext_s1[21], ciphertext_s0[21]}), .c ({new_AGEMA_signal_4998, SubBytesIns_Inst_Sbox_2_T7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T8_U1 ( .a ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({new_AGEMA_signal_5181, SubBytesIns_Inst_Sbox_2_T6}), .c ({new_AGEMA_signal_5371, SubBytesIns_Inst_Sbox_2_T8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T9_U1 ( .a ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({new_AGEMA_signal_4998, SubBytesIns_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_5182, SubBytesIns_Inst_Sbox_2_T9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T10_U1 ( .a ({new_AGEMA_signal_5181, SubBytesIns_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_4998, SubBytesIns_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_5372, SubBytesIns_Inst_Sbox_2_T10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T11_U1 ( .a ({ciphertext_s1[22], ciphertext_s0[22]}), .b ({ciphertext_s1[18], ciphertext_s0[18]}), .c ({new_AGEMA_signal_4999, SubBytesIns_Inst_Sbox_2_T11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T12_U1 ( .a ({ciphertext_s1[21], ciphertext_s0[21]}), .b ({ciphertext_s1[18], ciphertext_s0[18]}), .c ({new_AGEMA_signal_5000, SubBytesIns_Inst_Sbox_2_T12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T13_U1 ( .a ({new_AGEMA_signal_4995, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_4996, SubBytesIns_Inst_Sbox_2_T4}), .c ({new_AGEMA_signal_5183, SubBytesIns_Inst_Sbox_2_T13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T14_U1 ( .a ({new_AGEMA_signal_5181, SubBytesIns_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_4999, SubBytesIns_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_5373, SubBytesIns_Inst_Sbox_2_T14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T15_U1 ( .a ({new_AGEMA_signal_4997, SubBytesIns_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_4999, SubBytesIns_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_5184, SubBytesIns_Inst_Sbox_2_T15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T16_U1 ( .a ({new_AGEMA_signal_4997, SubBytesIns_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_5000, SubBytesIns_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_5185, SubBytesIns_Inst_Sbox_2_T16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T17_U1 ( .a ({new_AGEMA_signal_5182, SubBytesIns_Inst_Sbox_2_T9}), .b ({new_AGEMA_signal_5185, SubBytesIns_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_5374, SubBytesIns_Inst_Sbox_2_T17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T18_U1 ( .a ({ciphertext_s1[20], ciphertext_s0[20]}), .b ({ciphertext_s1[16], ciphertext_s0[16]}), .c ({new_AGEMA_signal_5001, SubBytesIns_Inst_Sbox_2_T18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T19_U1 ( .a ({new_AGEMA_signal_4998, SubBytesIns_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_5001, SubBytesIns_Inst_Sbox_2_T18}), .c ({new_AGEMA_signal_5186, SubBytesIns_Inst_Sbox_2_T19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T20_U1 ( .a ({new_AGEMA_signal_4993, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5186, SubBytesIns_Inst_Sbox_2_T19}), .c ({new_AGEMA_signal_5375, SubBytesIns_Inst_Sbox_2_T20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T21_U1 ( .a ({ciphertext_s1[17], ciphertext_s0[17]}), .b ({ciphertext_s1[16], ciphertext_s0[16]}), .c ({new_AGEMA_signal_5002, SubBytesIns_Inst_Sbox_2_T21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T22_U1 ( .a ({new_AGEMA_signal_4998, SubBytesIns_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_5002, SubBytesIns_Inst_Sbox_2_T21}), .c ({new_AGEMA_signal_5187, SubBytesIns_Inst_Sbox_2_T22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T23_U1 ( .a ({new_AGEMA_signal_4994, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_5187, SubBytesIns_Inst_Sbox_2_T22}), .c ({new_AGEMA_signal_5376, SubBytesIns_Inst_Sbox_2_T23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T24_U1 ( .a ({new_AGEMA_signal_4994, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_5372, SubBytesIns_Inst_Sbox_2_T10}), .c ({new_AGEMA_signal_5607, SubBytesIns_Inst_Sbox_2_T24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T25_U1 ( .a ({new_AGEMA_signal_5375, SubBytesIns_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_5374, SubBytesIns_Inst_Sbox_2_T17}), .c ({new_AGEMA_signal_5608, SubBytesIns_Inst_Sbox_2_T25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T26_U1 ( .a ({new_AGEMA_signal_4995, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_5185, SubBytesIns_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_5377, SubBytesIns_Inst_Sbox_2_T26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T27_U1 ( .a ({new_AGEMA_signal_4993, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5000, SubBytesIns_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_5188, SubBytesIns_Inst_Sbox_2_T27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T1_U1 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[28], ciphertext_s0[28]}), .c ({new_AGEMA_signal_5003, SubBytesIns_Inst_Sbox_3_T1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T2_U1 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_5004, SubBytesIns_Inst_Sbox_3_T2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T3_U1 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[25], ciphertext_s0[25]}), .c ({new_AGEMA_signal_5005, SubBytesIns_Inst_Sbox_3_T3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T4_U1 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_5006, SubBytesIns_Inst_Sbox_3_T4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T5_U1 ( .a ({ciphertext_s1[27], ciphertext_s0[27]}), .b ({ciphertext_s1[25], ciphertext_s0[25]}), .c ({new_AGEMA_signal_5007, SubBytesIns_Inst_Sbox_3_T5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T6_U1 ( .a ({new_AGEMA_signal_5003, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5007, SubBytesIns_Inst_Sbox_3_T5}), .c ({new_AGEMA_signal_5189, SubBytesIns_Inst_Sbox_3_T6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T7_U1 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({ciphertext_s1[29], ciphertext_s0[29]}), .c ({new_AGEMA_signal_5008, SubBytesIns_Inst_Sbox_3_T7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T8_U1 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({new_AGEMA_signal_5189, SubBytesIns_Inst_Sbox_3_T6}), .c ({new_AGEMA_signal_5384, SubBytesIns_Inst_Sbox_3_T8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T9_U1 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({new_AGEMA_signal_5008, SubBytesIns_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_5190, SubBytesIns_Inst_Sbox_3_T9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T10_U1 ( .a ({new_AGEMA_signal_5189, SubBytesIns_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_5008, SubBytesIns_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_5385, SubBytesIns_Inst_Sbox_3_T10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T11_U1 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_5009, SubBytesIns_Inst_Sbox_3_T11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T12_U1 ( .a ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_5010, SubBytesIns_Inst_Sbox_3_T12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T13_U1 ( .a ({new_AGEMA_signal_5005, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_5006, SubBytesIns_Inst_Sbox_3_T4}), .c ({new_AGEMA_signal_5191, SubBytesIns_Inst_Sbox_3_T13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T14_U1 ( .a ({new_AGEMA_signal_5189, SubBytesIns_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_5009, SubBytesIns_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_5386, SubBytesIns_Inst_Sbox_3_T14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T15_U1 ( .a ({new_AGEMA_signal_5007, SubBytesIns_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_5009, SubBytesIns_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_5192, SubBytesIns_Inst_Sbox_3_T15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T16_U1 ( .a ({new_AGEMA_signal_5007, SubBytesIns_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_5010, SubBytesIns_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_5193, SubBytesIns_Inst_Sbox_3_T16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T17_U1 ( .a ({new_AGEMA_signal_5190, SubBytesIns_Inst_Sbox_3_T9}), .b ({new_AGEMA_signal_5193, SubBytesIns_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_5387, SubBytesIns_Inst_Sbox_3_T17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T18_U1 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .c ({new_AGEMA_signal_5011, SubBytesIns_Inst_Sbox_3_T18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T19_U1 ( .a ({new_AGEMA_signal_5008, SubBytesIns_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_5011, SubBytesIns_Inst_Sbox_3_T18}), .c ({new_AGEMA_signal_5194, SubBytesIns_Inst_Sbox_3_T19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T20_U1 ( .a ({new_AGEMA_signal_5003, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5194, SubBytesIns_Inst_Sbox_3_T19}), .c ({new_AGEMA_signal_5388, SubBytesIns_Inst_Sbox_3_T20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T21_U1 ( .a ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .c ({new_AGEMA_signal_5012, SubBytesIns_Inst_Sbox_3_T21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T22_U1 ( .a ({new_AGEMA_signal_5008, SubBytesIns_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_5012, SubBytesIns_Inst_Sbox_3_T21}), .c ({new_AGEMA_signal_5195, SubBytesIns_Inst_Sbox_3_T22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T23_U1 ( .a ({new_AGEMA_signal_5004, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_5195, SubBytesIns_Inst_Sbox_3_T22}), .c ({new_AGEMA_signal_5389, SubBytesIns_Inst_Sbox_3_T23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T24_U1 ( .a ({new_AGEMA_signal_5004, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_5385, SubBytesIns_Inst_Sbox_3_T10}), .c ({new_AGEMA_signal_5616, SubBytesIns_Inst_Sbox_3_T24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T25_U1 ( .a ({new_AGEMA_signal_5388, SubBytesIns_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_5387, SubBytesIns_Inst_Sbox_3_T17}), .c ({new_AGEMA_signal_5617, SubBytesIns_Inst_Sbox_3_T25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T26_U1 ( .a ({new_AGEMA_signal_5005, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_5193, SubBytesIns_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_5390, SubBytesIns_Inst_Sbox_3_T26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T27_U1 ( .a ({new_AGEMA_signal_5003, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5010, SubBytesIns_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_5196, SubBytesIns_Inst_Sbox_3_T27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T1_U1 ( .a ({ciphertext_s1[39], ciphertext_s0[39]}), .b ({ciphertext_s1[36], ciphertext_s0[36]}), .c ({new_AGEMA_signal_5013, SubBytesIns_Inst_Sbox_4_T1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T2_U1 ( .a ({ciphertext_s1[39], ciphertext_s0[39]}), .b ({ciphertext_s1[34], ciphertext_s0[34]}), .c ({new_AGEMA_signal_5014, SubBytesIns_Inst_Sbox_4_T2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T3_U1 ( .a ({ciphertext_s1[39], ciphertext_s0[39]}), .b ({ciphertext_s1[33], ciphertext_s0[33]}), .c ({new_AGEMA_signal_5015, SubBytesIns_Inst_Sbox_4_T3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T4_U1 ( .a ({ciphertext_s1[36], ciphertext_s0[36]}), .b ({ciphertext_s1[34], ciphertext_s0[34]}), .c ({new_AGEMA_signal_5016, SubBytesIns_Inst_Sbox_4_T4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T5_U1 ( .a ({ciphertext_s1[35], ciphertext_s0[35]}), .b ({ciphertext_s1[33], ciphertext_s0[33]}), .c ({new_AGEMA_signal_5017, SubBytesIns_Inst_Sbox_4_T5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T6_U1 ( .a ({new_AGEMA_signal_5013, SubBytesIns_Inst_Sbox_4_T1}), .b ({new_AGEMA_signal_5017, SubBytesIns_Inst_Sbox_4_T5}), .c ({new_AGEMA_signal_5197, SubBytesIns_Inst_Sbox_4_T6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T7_U1 ( .a ({ciphertext_s1[38], ciphertext_s0[38]}), .b ({ciphertext_s1[37], ciphertext_s0[37]}), .c ({new_AGEMA_signal_5018, SubBytesIns_Inst_Sbox_4_T7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T8_U1 ( .a ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({new_AGEMA_signal_5197, SubBytesIns_Inst_Sbox_4_T6}), .c ({new_AGEMA_signal_5397, SubBytesIns_Inst_Sbox_4_T8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T9_U1 ( .a ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({new_AGEMA_signal_5018, SubBytesIns_Inst_Sbox_4_T7}), .c ({new_AGEMA_signal_5198, SubBytesIns_Inst_Sbox_4_T9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T10_U1 ( .a ({new_AGEMA_signal_5197, SubBytesIns_Inst_Sbox_4_T6}), .b ({new_AGEMA_signal_5018, SubBytesIns_Inst_Sbox_4_T7}), .c ({new_AGEMA_signal_5398, SubBytesIns_Inst_Sbox_4_T10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T11_U1 ( .a ({ciphertext_s1[38], ciphertext_s0[38]}), .b ({ciphertext_s1[34], ciphertext_s0[34]}), .c ({new_AGEMA_signal_5019, SubBytesIns_Inst_Sbox_4_T11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T12_U1 ( .a ({ciphertext_s1[37], ciphertext_s0[37]}), .b ({ciphertext_s1[34], ciphertext_s0[34]}), .c ({new_AGEMA_signal_5020, SubBytesIns_Inst_Sbox_4_T12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T13_U1 ( .a ({new_AGEMA_signal_5015, SubBytesIns_Inst_Sbox_4_T3}), .b ({new_AGEMA_signal_5016, SubBytesIns_Inst_Sbox_4_T4}), .c ({new_AGEMA_signal_5199, SubBytesIns_Inst_Sbox_4_T13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T14_U1 ( .a ({new_AGEMA_signal_5197, SubBytesIns_Inst_Sbox_4_T6}), .b ({new_AGEMA_signal_5019, SubBytesIns_Inst_Sbox_4_T11}), .c ({new_AGEMA_signal_5399, SubBytesIns_Inst_Sbox_4_T14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T15_U1 ( .a ({new_AGEMA_signal_5017, SubBytesIns_Inst_Sbox_4_T5}), .b ({new_AGEMA_signal_5019, SubBytesIns_Inst_Sbox_4_T11}), .c ({new_AGEMA_signal_5200, SubBytesIns_Inst_Sbox_4_T15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T16_U1 ( .a ({new_AGEMA_signal_5017, SubBytesIns_Inst_Sbox_4_T5}), .b ({new_AGEMA_signal_5020, SubBytesIns_Inst_Sbox_4_T12}), .c ({new_AGEMA_signal_5201, SubBytesIns_Inst_Sbox_4_T16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T17_U1 ( .a ({new_AGEMA_signal_5198, SubBytesIns_Inst_Sbox_4_T9}), .b ({new_AGEMA_signal_5201, SubBytesIns_Inst_Sbox_4_T16}), .c ({new_AGEMA_signal_5400, SubBytesIns_Inst_Sbox_4_T17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T18_U1 ( .a ({ciphertext_s1[36], ciphertext_s0[36]}), .b ({ciphertext_s1[32], ciphertext_s0[32]}), .c ({new_AGEMA_signal_5021, SubBytesIns_Inst_Sbox_4_T18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T19_U1 ( .a ({new_AGEMA_signal_5018, SubBytesIns_Inst_Sbox_4_T7}), .b ({new_AGEMA_signal_5021, SubBytesIns_Inst_Sbox_4_T18}), .c ({new_AGEMA_signal_5202, SubBytesIns_Inst_Sbox_4_T19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T20_U1 ( .a ({new_AGEMA_signal_5013, SubBytesIns_Inst_Sbox_4_T1}), .b ({new_AGEMA_signal_5202, SubBytesIns_Inst_Sbox_4_T19}), .c ({new_AGEMA_signal_5401, SubBytesIns_Inst_Sbox_4_T20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T21_U1 ( .a ({ciphertext_s1[33], ciphertext_s0[33]}), .b ({ciphertext_s1[32], ciphertext_s0[32]}), .c ({new_AGEMA_signal_5022, SubBytesIns_Inst_Sbox_4_T21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T22_U1 ( .a ({new_AGEMA_signal_5018, SubBytesIns_Inst_Sbox_4_T7}), .b ({new_AGEMA_signal_5022, SubBytesIns_Inst_Sbox_4_T21}), .c ({new_AGEMA_signal_5203, SubBytesIns_Inst_Sbox_4_T22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T23_U1 ( .a ({new_AGEMA_signal_5014, SubBytesIns_Inst_Sbox_4_T2}), .b ({new_AGEMA_signal_5203, SubBytesIns_Inst_Sbox_4_T22}), .c ({new_AGEMA_signal_5402, SubBytesIns_Inst_Sbox_4_T23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T24_U1 ( .a ({new_AGEMA_signal_5014, SubBytesIns_Inst_Sbox_4_T2}), .b ({new_AGEMA_signal_5398, SubBytesIns_Inst_Sbox_4_T10}), .c ({new_AGEMA_signal_5625, SubBytesIns_Inst_Sbox_4_T24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T25_U1 ( .a ({new_AGEMA_signal_5401, SubBytesIns_Inst_Sbox_4_T20}), .b ({new_AGEMA_signal_5400, SubBytesIns_Inst_Sbox_4_T17}), .c ({new_AGEMA_signal_5626, SubBytesIns_Inst_Sbox_4_T25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T26_U1 ( .a ({new_AGEMA_signal_5015, SubBytesIns_Inst_Sbox_4_T3}), .b ({new_AGEMA_signal_5201, SubBytesIns_Inst_Sbox_4_T16}), .c ({new_AGEMA_signal_5403, SubBytesIns_Inst_Sbox_4_T26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T27_U1 ( .a ({new_AGEMA_signal_5013, SubBytesIns_Inst_Sbox_4_T1}), .b ({new_AGEMA_signal_5020, SubBytesIns_Inst_Sbox_4_T12}), .c ({new_AGEMA_signal_5204, SubBytesIns_Inst_Sbox_4_T27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T1_U1 ( .a ({ciphertext_s1[47], ciphertext_s0[47]}), .b ({ciphertext_s1[44], ciphertext_s0[44]}), .c ({new_AGEMA_signal_5023, SubBytesIns_Inst_Sbox_5_T1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T2_U1 ( .a ({ciphertext_s1[47], ciphertext_s0[47]}), .b ({ciphertext_s1[42], ciphertext_s0[42]}), .c ({new_AGEMA_signal_5024, SubBytesIns_Inst_Sbox_5_T2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T3_U1 ( .a ({ciphertext_s1[47], ciphertext_s0[47]}), .b ({ciphertext_s1[41], ciphertext_s0[41]}), .c ({new_AGEMA_signal_5025, SubBytesIns_Inst_Sbox_5_T3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T4_U1 ( .a ({ciphertext_s1[44], ciphertext_s0[44]}), .b ({ciphertext_s1[42], ciphertext_s0[42]}), .c ({new_AGEMA_signal_5026, SubBytesIns_Inst_Sbox_5_T4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T5_U1 ( .a ({ciphertext_s1[43], ciphertext_s0[43]}), .b ({ciphertext_s1[41], ciphertext_s0[41]}), .c ({new_AGEMA_signal_5027, SubBytesIns_Inst_Sbox_5_T5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T6_U1 ( .a ({new_AGEMA_signal_5023, SubBytesIns_Inst_Sbox_5_T1}), .b ({new_AGEMA_signal_5027, SubBytesIns_Inst_Sbox_5_T5}), .c ({new_AGEMA_signal_5205, SubBytesIns_Inst_Sbox_5_T6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T7_U1 ( .a ({ciphertext_s1[46], ciphertext_s0[46]}), .b ({ciphertext_s1[45], ciphertext_s0[45]}), .c ({new_AGEMA_signal_5028, SubBytesIns_Inst_Sbox_5_T7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T8_U1 ( .a ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({new_AGEMA_signal_5205, SubBytesIns_Inst_Sbox_5_T6}), .c ({new_AGEMA_signal_5410, SubBytesIns_Inst_Sbox_5_T8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T9_U1 ( .a ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({new_AGEMA_signal_5028, SubBytesIns_Inst_Sbox_5_T7}), .c ({new_AGEMA_signal_5206, SubBytesIns_Inst_Sbox_5_T9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T10_U1 ( .a ({new_AGEMA_signal_5205, SubBytesIns_Inst_Sbox_5_T6}), .b ({new_AGEMA_signal_5028, SubBytesIns_Inst_Sbox_5_T7}), .c ({new_AGEMA_signal_5411, SubBytesIns_Inst_Sbox_5_T10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T11_U1 ( .a ({ciphertext_s1[46], ciphertext_s0[46]}), .b ({ciphertext_s1[42], ciphertext_s0[42]}), .c ({new_AGEMA_signal_5029, SubBytesIns_Inst_Sbox_5_T11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T12_U1 ( .a ({ciphertext_s1[45], ciphertext_s0[45]}), .b ({ciphertext_s1[42], ciphertext_s0[42]}), .c ({new_AGEMA_signal_5030, SubBytesIns_Inst_Sbox_5_T12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T13_U1 ( .a ({new_AGEMA_signal_5025, SubBytesIns_Inst_Sbox_5_T3}), .b ({new_AGEMA_signal_5026, SubBytesIns_Inst_Sbox_5_T4}), .c ({new_AGEMA_signal_5207, SubBytesIns_Inst_Sbox_5_T13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T14_U1 ( .a ({new_AGEMA_signal_5205, SubBytesIns_Inst_Sbox_5_T6}), .b ({new_AGEMA_signal_5029, SubBytesIns_Inst_Sbox_5_T11}), .c ({new_AGEMA_signal_5412, SubBytesIns_Inst_Sbox_5_T14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T15_U1 ( .a ({new_AGEMA_signal_5027, SubBytesIns_Inst_Sbox_5_T5}), .b ({new_AGEMA_signal_5029, SubBytesIns_Inst_Sbox_5_T11}), .c ({new_AGEMA_signal_5208, SubBytesIns_Inst_Sbox_5_T15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T16_U1 ( .a ({new_AGEMA_signal_5027, SubBytesIns_Inst_Sbox_5_T5}), .b ({new_AGEMA_signal_5030, SubBytesIns_Inst_Sbox_5_T12}), .c ({new_AGEMA_signal_5209, SubBytesIns_Inst_Sbox_5_T16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T17_U1 ( .a ({new_AGEMA_signal_5206, SubBytesIns_Inst_Sbox_5_T9}), .b ({new_AGEMA_signal_5209, SubBytesIns_Inst_Sbox_5_T16}), .c ({new_AGEMA_signal_5413, SubBytesIns_Inst_Sbox_5_T17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T18_U1 ( .a ({ciphertext_s1[44], ciphertext_s0[44]}), .b ({ciphertext_s1[40], ciphertext_s0[40]}), .c ({new_AGEMA_signal_5031, SubBytesIns_Inst_Sbox_5_T18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T19_U1 ( .a ({new_AGEMA_signal_5028, SubBytesIns_Inst_Sbox_5_T7}), .b ({new_AGEMA_signal_5031, SubBytesIns_Inst_Sbox_5_T18}), .c ({new_AGEMA_signal_5210, SubBytesIns_Inst_Sbox_5_T19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T20_U1 ( .a ({new_AGEMA_signal_5023, SubBytesIns_Inst_Sbox_5_T1}), .b ({new_AGEMA_signal_5210, SubBytesIns_Inst_Sbox_5_T19}), .c ({new_AGEMA_signal_5414, SubBytesIns_Inst_Sbox_5_T20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T21_U1 ( .a ({ciphertext_s1[41], ciphertext_s0[41]}), .b ({ciphertext_s1[40], ciphertext_s0[40]}), .c ({new_AGEMA_signal_5032, SubBytesIns_Inst_Sbox_5_T21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T22_U1 ( .a ({new_AGEMA_signal_5028, SubBytesIns_Inst_Sbox_5_T7}), .b ({new_AGEMA_signal_5032, SubBytesIns_Inst_Sbox_5_T21}), .c ({new_AGEMA_signal_5211, SubBytesIns_Inst_Sbox_5_T22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T23_U1 ( .a ({new_AGEMA_signal_5024, SubBytesIns_Inst_Sbox_5_T2}), .b ({new_AGEMA_signal_5211, SubBytesIns_Inst_Sbox_5_T22}), .c ({new_AGEMA_signal_5415, SubBytesIns_Inst_Sbox_5_T23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T24_U1 ( .a ({new_AGEMA_signal_5024, SubBytesIns_Inst_Sbox_5_T2}), .b ({new_AGEMA_signal_5411, SubBytesIns_Inst_Sbox_5_T10}), .c ({new_AGEMA_signal_5634, SubBytesIns_Inst_Sbox_5_T24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T25_U1 ( .a ({new_AGEMA_signal_5414, SubBytesIns_Inst_Sbox_5_T20}), .b ({new_AGEMA_signal_5413, SubBytesIns_Inst_Sbox_5_T17}), .c ({new_AGEMA_signal_5635, SubBytesIns_Inst_Sbox_5_T25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T26_U1 ( .a ({new_AGEMA_signal_5025, SubBytesIns_Inst_Sbox_5_T3}), .b ({new_AGEMA_signal_5209, SubBytesIns_Inst_Sbox_5_T16}), .c ({new_AGEMA_signal_5416, SubBytesIns_Inst_Sbox_5_T26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T27_U1 ( .a ({new_AGEMA_signal_5023, SubBytesIns_Inst_Sbox_5_T1}), .b ({new_AGEMA_signal_5030, SubBytesIns_Inst_Sbox_5_T12}), .c ({new_AGEMA_signal_5212, SubBytesIns_Inst_Sbox_5_T27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T1_U1 ( .a ({ciphertext_s1[55], ciphertext_s0[55]}), .b ({ciphertext_s1[52], ciphertext_s0[52]}), .c ({new_AGEMA_signal_5033, SubBytesIns_Inst_Sbox_6_T1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T2_U1 ( .a ({ciphertext_s1[55], ciphertext_s0[55]}), .b ({ciphertext_s1[50], ciphertext_s0[50]}), .c ({new_AGEMA_signal_5034, SubBytesIns_Inst_Sbox_6_T2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T3_U1 ( .a ({ciphertext_s1[55], ciphertext_s0[55]}), .b ({ciphertext_s1[49], ciphertext_s0[49]}), .c ({new_AGEMA_signal_5035, SubBytesIns_Inst_Sbox_6_T3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T4_U1 ( .a ({ciphertext_s1[52], ciphertext_s0[52]}), .b ({ciphertext_s1[50], ciphertext_s0[50]}), .c ({new_AGEMA_signal_5036, SubBytesIns_Inst_Sbox_6_T4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T5_U1 ( .a ({ciphertext_s1[51], ciphertext_s0[51]}), .b ({ciphertext_s1[49], ciphertext_s0[49]}), .c ({new_AGEMA_signal_5037, SubBytesIns_Inst_Sbox_6_T5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T6_U1 ( .a ({new_AGEMA_signal_5033, SubBytesIns_Inst_Sbox_6_T1}), .b ({new_AGEMA_signal_5037, SubBytesIns_Inst_Sbox_6_T5}), .c ({new_AGEMA_signal_5213, SubBytesIns_Inst_Sbox_6_T6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T7_U1 ( .a ({ciphertext_s1[54], ciphertext_s0[54]}), .b ({ciphertext_s1[53], ciphertext_s0[53]}), .c ({new_AGEMA_signal_5038, SubBytesIns_Inst_Sbox_6_T7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T8_U1 ( .a ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({new_AGEMA_signal_5213, SubBytesIns_Inst_Sbox_6_T6}), .c ({new_AGEMA_signal_5423, SubBytesIns_Inst_Sbox_6_T8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T9_U1 ( .a ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({new_AGEMA_signal_5038, SubBytesIns_Inst_Sbox_6_T7}), .c ({new_AGEMA_signal_5214, SubBytesIns_Inst_Sbox_6_T9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T10_U1 ( .a ({new_AGEMA_signal_5213, SubBytesIns_Inst_Sbox_6_T6}), .b ({new_AGEMA_signal_5038, SubBytesIns_Inst_Sbox_6_T7}), .c ({new_AGEMA_signal_5424, SubBytesIns_Inst_Sbox_6_T10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T11_U1 ( .a ({ciphertext_s1[54], ciphertext_s0[54]}), .b ({ciphertext_s1[50], ciphertext_s0[50]}), .c ({new_AGEMA_signal_5039, SubBytesIns_Inst_Sbox_6_T11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T12_U1 ( .a ({ciphertext_s1[53], ciphertext_s0[53]}), .b ({ciphertext_s1[50], ciphertext_s0[50]}), .c ({new_AGEMA_signal_5040, SubBytesIns_Inst_Sbox_6_T12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T13_U1 ( .a ({new_AGEMA_signal_5035, SubBytesIns_Inst_Sbox_6_T3}), .b ({new_AGEMA_signal_5036, SubBytesIns_Inst_Sbox_6_T4}), .c ({new_AGEMA_signal_5215, SubBytesIns_Inst_Sbox_6_T13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T14_U1 ( .a ({new_AGEMA_signal_5213, SubBytesIns_Inst_Sbox_6_T6}), .b ({new_AGEMA_signal_5039, SubBytesIns_Inst_Sbox_6_T11}), .c ({new_AGEMA_signal_5425, SubBytesIns_Inst_Sbox_6_T14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T15_U1 ( .a ({new_AGEMA_signal_5037, SubBytesIns_Inst_Sbox_6_T5}), .b ({new_AGEMA_signal_5039, SubBytesIns_Inst_Sbox_6_T11}), .c ({new_AGEMA_signal_5216, SubBytesIns_Inst_Sbox_6_T15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T16_U1 ( .a ({new_AGEMA_signal_5037, SubBytesIns_Inst_Sbox_6_T5}), .b ({new_AGEMA_signal_5040, SubBytesIns_Inst_Sbox_6_T12}), .c ({new_AGEMA_signal_5217, SubBytesIns_Inst_Sbox_6_T16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T17_U1 ( .a ({new_AGEMA_signal_5214, SubBytesIns_Inst_Sbox_6_T9}), .b ({new_AGEMA_signal_5217, SubBytesIns_Inst_Sbox_6_T16}), .c ({new_AGEMA_signal_5426, SubBytesIns_Inst_Sbox_6_T17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T18_U1 ( .a ({ciphertext_s1[52], ciphertext_s0[52]}), .b ({ciphertext_s1[48], ciphertext_s0[48]}), .c ({new_AGEMA_signal_5041, SubBytesIns_Inst_Sbox_6_T18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T19_U1 ( .a ({new_AGEMA_signal_5038, SubBytesIns_Inst_Sbox_6_T7}), .b ({new_AGEMA_signal_5041, SubBytesIns_Inst_Sbox_6_T18}), .c ({new_AGEMA_signal_5218, SubBytesIns_Inst_Sbox_6_T19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T20_U1 ( .a ({new_AGEMA_signal_5033, SubBytesIns_Inst_Sbox_6_T1}), .b ({new_AGEMA_signal_5218, SubBytesIns_Inst_Sbox_6_T19}), .c ({new_AGEMA_signal_5427, SubBytesIns_Inst_Sbox_6_T20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T21_U1 ( .a ({ciphertext_s1[49], ciphertext_s0[49]}), .b ({ciphertext_s1[48], ciphertext_s0[48]}), .c ({new_AGEMA_signal_5042, SubBytesIns_Inst_Sbox_6_T21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T22_U1 ( .a ({new_AGEMA_signal_5038, SubBytesIns_Inst_Sbox_6_T7}), .b ({new_AGEMA_signal_5042, SubBytesIns_Inst_Sbox_6_T21}), .c ({new_AGEMA_signal_5219, SubBytesIns_Inst_Sbox_6_T22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T23_U1 ( .a ({new_AGEMA_signal_5034, SubBytesIns_Inst_Sbox_6_T2}), .b ({new_AGEMA_signal_5219, SubBytesIns_Inst_Sbox_6_T22}), .c ({new_AGEMA_signal_5428, SubBytesIns_Inst_Sbox_6_T23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T24_U1 ( .a ({new_AGEMA_signal_5034, SubBytesIns_Inst_Sbox_6_T2}), .b ({new_AGEMA_signal_5424, SubBytesIns_Inst_Sbox_6_T10}), .c ({new_AGEMA_signal_5643, SubBytesIns_Inst_Sbox_6_T24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T25_U1 ( .a ({new_AGEMA_signal_5427, SubBytesIns_Inst_Sbox_6_T20}), .b ({new_AGEMA_signal_5426, SubBytesIns_Inst_Sbox_6_T17}), .c ({new_AGEMA_signal_5644, SubBytesIns_Inst_Sbox_6_T25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T26_U1 ( .a ({new_AGEMA_signal_5035, SubBytesIns_Inst_Sbox_6_T3}), .b ({new_AGEMA_signal_5217, SubBytesIns_Inst_Sbox_6_T16}), .c ({new_AGEMA_signal_5429, SubBytesIns_Inst_Sbox_6_T26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T27_U1 ( .a ({new_AGEMA_signal_5033, SubBytesIns_Inst_Sbox_6_T1}), .b ({new_AGEMA_signal_5040, SubBytesIns_Inst_Sbox_6_T12}), .c ({new_AGEMA_signal_5220, SubBytesIns_Inst_Sbox_6_T27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T1_U1 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[60], ciphertext_s0[60]}), .c ({new_AGEMA_signal_5043, SubBytesIns_Inst_Sbox_7_T1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T2_U1 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_5044, SubBytesIns_Inst_Sbox_7_T2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T3_U1 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[57], ciphertext_s0[57]}), .c ({new_AGEMA_signal_5045, SubBytesIns_Inst_Sbox_7_T3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T4_U1 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_5046, SubBytesIns_Inst_Sbox_7_T4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T5_U1 ( .a ({ciphertext_s1[59], ciphertext_s0[59]}), .b ({ciphertext_s1[57], ciphertext_s0[57]}), .c ({new_AGEMA_signal_5047, SubBytesIns_Inst_Sbox_7_T5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T6_U1 ( .a ({new_AGEMA_signal_5043, SubBytesIns_Inst_Sbox_7_T1}), .b ({new_AGEMA_signal_5047, SubBytesIns_Inst_Sbox_7_T5}), .c ({new_AGEMA_signal_5221, SubBytesIns_Inst_Sbox_7_T6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T7_U1 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({ciphertext_s1[61], ciphertext_s0[61]}), .c ({new_AGEMA_signal_5048, SubBytesIns_Inst_Sbox_7_T7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T8_U1 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({new_AGEMA_signal_5221, SubBytesIns_Inst_Sbox_7_T6}), .c ({new_AGEMA_signal_5436, SubBytesIns_Inst_Sbox_7_T8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T9_U1 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({new_AGEMA_signal_5048, SubBytesIns_Inst_Sbox_7_T7}), .c ({new_AGEMA_signal_5222, SubBytesIns_Inst_Sbox_7_T9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T10_U1 ( .a ({new_AGEMA_signal_5221, SubBytesIns_Inst_Sbox_7_T6}), .b ({new_AGEMA_signal_5048, SubBytesIns_Inst_Sbox_7_T7}), .c ({new_AGEMA_signal_5437, SubBytesIns_Inst_Sbox_7_T10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T11_U1 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_5049, SubBytesIns_Inst_Sbox_7_T11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T12_U1 ( .a ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_5050, SubBytesIns_Inst_Sbox_7_T12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T13_U1 ( .a ({new_AGEMA_signal_5045, SubBytesIns_Inst_Sbox_7_T3}), .b ({new_AGEMA_signal_5046, SubBytesIns_Inst_Sbox_7_T4}), .c ({new_AGEMA_signal_5223, SubBytesIns_Inst_Sbox_7_T13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T14_U1 ( .a ({new_AGEMA_signal_5221, SubBytesIns_Inst_Sbox_7_T6}), .b ({new_AGEMA_signal_5049, SubBytesIns_Inst_Sbox_7_T11}), .c ({new_AGEMA_signal_5438, SubBytesIns_Inst_Sbox_7_T14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T15_U1 ( .a ({new_AGEMA_signal_5047, SubBytesIns_Inst_Sbox_7_T5}), .b ({new_AGEMA_signal_5049, SubBytesIns_Inst_Sbox_7_T11}), .c ({new_AGEMA_signal_5224, SubBytesIns_Inst_Sbox_7_T15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T16_U1 ( .a ({new_AGEMA_signal_5047, SubBytesIns_Inst_Sbox_7_T5}), .b ({new_AGEMA_signal_5050, SubBytesIns_Inst_Sbox_7_T12}), .c ({new_AGEMA_signal_5225, SubBytesIns_Inst_Sbox_7_T16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T17_U1 ( .a ({new_AGEMA_signal_5222, SubBytesIns_Inst_Sbox_7_T9}), .b ({new_AGEMA_signal_5225, SubBytesIns_Inst_Sbox_7_T16}), .c ({new_AGEMA_signal_5439, SubBytesIns_Inst_Sbox_7_T17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T18_U1 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .c ({new_AGEMA_signal_5051, SubBytesIns_Inst_Sbox_7_T18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T19_U1 ( .a ({new_AGEMA_signal_5048, SubBytesIns_Inst_Sbox_7_T7}), .b ({new_AGEMA_signal_5051, SubBytesIns_Inst_Sbox_7_T18}), .c ({new_AGEMA_signal_5226, SubBytesIns_Inst_Sbox_7_T19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T20_U1 ( .a ({new_AGEMA_signal_5043, SubBytesIns_Inst_Sbox_7_T1}), .b ({new_AGEMA_signal_5226, SubBytesIns_Inst_Sbox_7_T19}), .c ({new_AGEMA_signal_5440, SubBytesIns_Inst_Sbox_7_T20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T21_U1 ( .a ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .c ({new_AGEMA_signal_5052, SubBytesIns_Inst_Sbox_7_T21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T22_U1 ( .a ({new_AGEMA_signal_5048, SubBytesIns_Inst_Sbox_7_T7}), .b ({new_AGEMA_signal_5052, SubBytesIns_Inst_Sbox_7_T21}), .c ({new_AGEMA_signal_5227, SubBytesIns_Inst_Sbox_7_T22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T23_U1 ( .a ({new_AGEMA_signal_5044, SubBytesIns_Inst_Sbox_7_T2}), .b ({new_AGEMA_signal_5227, SubBytesIns_Inst_Sbox_7_T22}), .c ({new_AGEMA_signal_5441, SubBytesIns_Inst_Sbox_7_T23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T24_U1 ( .a ({new_AGEMA_signal_5044, SubBytesIns_Inst_Sbox_7_T2}), .b ({new_AGEMA_signal_5437, SubBytesIns_Inst_Sbox_7_T10}), .c ({new_AGEMA_signal_5652, SubBytesIns_Inst_Sbox_7_T24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T25_U1 ( .a ({new_AGEMA_signal_5440, SubBytesIns_Inst_Sbox_7_T20}), .b ({new_AGEMA_signal_5439, SubBytesIns_Inst_Sbox_7_T17}), .c ({new_AGEMA_signal_5653, SubBytesIns_Inst_Sbox_7_T25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T26_U1 ( .a ({new_AGEMA_signal_5045, SubBytesIns_Inst_Sbox_7_T3}), .b ({new_AGEMA_signal_5225, SubBytesIns_Inst_Sbox_7_T16}), .c ({new_AGEMA_signal_5442, SubBytesIns_Inst_Sbox_7_T26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T27_U1 ( .a ({new_AGEMA_signal_5043, SubBytesIns_Inst_Sbox_7_T1}), .b ({new_AGEMA_signal_5050, SubBytesIns_Inst_Sbox_7_T12}), .c ({new_AGEMA_signal_5228, SubBytesIns_Inst_Sbox_7_T27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T1_U1 ( .a ({ciphertext_s1[71], ciphertext_s0[71]}), .b ({ciphertext_s1[68], ciphertext_s0[68]}), .c ({new_AGEMA_signal_5053, SubBytesIns_Inst_Sbox_8_T1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T2_U1 ( .a ({ciphertext_s1[71], ciphertext_s0[71]}), .b ({ciphertext_s1[66], ciphertext_s0[66]}), .c ({new_AGEMA_signal_5054, SubBytesIns_Inst_Sbox_8_T2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T3_U1 ( .a ({ciphertext_s1[71], ciphertext_s0[71]}), .b ({ciphertext_s1[65], ciphertext_s0[65]}), .c ({new_AGEMA_signal_5055, SubBytesIns_Inst_Sbox_8_T3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T4_U1 ( .a ({ciphertext_s1[68], ciphertext_s0[68]}), .b ({ciphertext_s1[66], ciphertext_s0[66]}), .c ({new_AGEMA_signal_5056, SubBytesIns_Inst_Sbox_8_T4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T5_U1 ( .a ({ciphertext_s1[67], ciphertext_s0[67]}), .b ({ciphertext_s1[65], ciphertext_s0[65]}), .c ({new_AGEMA_signal_5057, SubBytesIns_Inst_Sbox_8_T5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T6_U1 ( .a ({new_AGEMA_signal_5053, SubBytesIns_Inst_Sbox_8_T1}), .b ({new_AGEMA_signal_5057, SubBytesIns_Inst_Sbox_8_T5}), .c ({new_AGEMA_signal_5229, SubBytesIns_Inst_Sbox_8_T6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T7_U1 ( .a ({ciphertext_s1[70], ciphertext_s0[70]}), .b ({ciphertext_s1[69], ciphertext_s0[69]}), .c ({new_AGEMA_signal_5058, SubBytesIns_Inst_Sbox_8_T7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T8_U1 ( .a ({ciphertext_s1[64], ciphertext_s0[64]}), .b ({new_AGEMA_signal_5229, SubBytesIns_Inst_Sbox_8_T6}), .c ({new_AGEMA_signal_5449, SubBytesIns_Inst_Sbox_8_T8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T9_U1 ( .a ({ciphertext_s1[64], ciphertext_s0[64]}), .b ({new_AGEMA_signal_5058, SubBytesIns_Inst_Sbox_8_T7}), .c ({new_AGEMA_signal_5230, SubBytesIns_Inst_Sbox_8_T9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T10_U1 ( .a ({new_AGEMA_signal_5229, SubBytesIns_Inst_Sbox_8_T6}), .b ({new_AGEMA_signal_5058, SubBytesIns_Inst_Sbox_8_T7}), .c ({new_AGEMA_signal_5450, SubBytesIns_Inst_Sbox_8_T10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T11_U1 ( .a ({ciphertext_s1[70], ciphertext_s0[70]}), .b ({ciphertext_s1[66], ciphertext_s0[66]}), .c ({new_AGEMA_signal_5059, SubBytesIns_Inst_Sbox_8_T11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T12_U1 ( .a ({ciphertext_s1[69], ciphertext_s0[69]}), .b ({ciphertext_s1[66], ciphertext_s0[66]}), .c ({new_AGEMA_signal_5060, SubBytesIns_Inst_Sbox_8_T12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T13_U1 ( .a ({new_AGEMA_signal_5055, SubBytesIns_Inst_Sbox_8_T3}), .b ({new_AGEMA_signal_5056, SubBytesIns_Inst_Sbox_8_T4}), .c ({new_AGEMA_signal_5231, SubBytesIns_Inst_Sbox_8_T13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T14_U1 ( .a ({new_AGEMA_signal_5229, SubBytesIns_Inst_Sbox_8_T6}), .b ({new_AGEMA_signal_5059, SubBytesIns_Inst_Sbox_8_T11}), .c ({new_AGEMA_signal_5451, SubBytesIns_Inst_Sbox_8_T14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T15_U1 ( .a ({new_AGEMA_signal_5057, SubBytesIns_Inst_Sbox_8_T5}), .b ({new_AGEMA_signal_5059, SubBytesIns_Inst_Sbox_8_T11}), .c ({new_AGEMA_signal_5232, SubBytesIns_Inst_Sbox_8_T15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T16_U1 ( .a ({new_AGEMA_signal_5057, SubBytesIns_Inst_Sbox_8_T5}), .b ({new_AGEMA_signal_5060, SubBytesIns_Inst_Sbox_8_T12}), .c ({new_AGEMA_signal_5233, SubBytesIns_Inst_Sbox_8_T16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T17_U1 ( .a ({new_AGEMA_signal_5230, SubBytesIns_Inst_Sbox_8_T9}), .b ({new_AGEMA_signal_5233, SubBytesIns_Inst_Sbox_8_T16}), .c ({new_AGEMA_signal_5452, SubBytesIns_Inst_Sbox_8_T17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T18_U1 ( .a ({ciphertext_s1[68], ciphertext_s0[68]}), .b ({ciphertext_s1[64], ciphertext_s0[64]}), .c ({new_AGEMA_signal_5061, SubBytesIns_Inst_Sbox_8_T18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T19_U1 ( .a ({new_AGEMA_signal_5058, SubBytesIns_Inst_Sbox_8_T7}), .b ({new_AGEMA_signal_5061, SubBytesIns_Inst_Sbox_8_T18}), .c ({new_AGEMA_signal_5234, SubBytesIns_Inst_Sbox_8_T19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T20_U1 ( .a ({new_AGEMA_signal_5053, SubBytesIns_Inst_Sbox_8_T1}), .b ({new_AGEMA_signal_5234, SubBytesIns_Inst_Sbox_8_T19}), .c ({new_AGEMA_signal_5453, SubBytesIns_Inst_Sbox_8_T20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T21_U1 ( .a ({ciphertext_s1[65], ciphertext_s0[65]}), .b ({ciphertext_s1[64], ciphertext_s0[64]}), .c ({new_AGEMA_signal_5062, SubBytesIns_Inst_Sbox_8_T21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T22_U1 ( .a ({new_AGEMA_signal_5058, SubBytesIns_Inst_Sbox_8_T7}), .b ({new_AGEMA_signal_5062, SubBytesIns_Inst_Sbox_8_T21}), .c ({new_AGEMA_signal_5235, SubBytesIns_Inst_Sbox_8_T22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T23_U1 ( .a ({new_AGEMA_signal_5054, SubBytesIns_Inst_Sbox_8_T2}), .b ({new_AGEMA_signal_5235, SubBytesIns_Inst_Sbox_8_T22}), .c ({new_AGEMA_signal_5454, SubBytesIns_Inst_Sbox_8_T23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T24_U1 ( .a ({new_AGEMA_signal_5054, SubBytesIns_Inst_Sbox_8_T2}), .b ({new_AGEMA_signal_5450, SubBytesIns_Inst_Sbox_8_T10}), .c ({new_AGEMA_signal_5661, SubBytesIns_Inst_Sbox_8_T24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T25_U1 ( .a ({new_AGEMA_signal_5453, SubBytesIns_Inst_Sbox_8_T20}), .b ({new_AGEMA_signal_5452, SubBytesIns_Inst_Sbox_8_T17}), .c ({new_AGEMA_signal_5662, SubBytesIns_Inst_Sbox_8_T25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T26_U1 ( .a ({new_AGEMA_signal_5055, SubBytesIns_Inst_Sbox_8_T3}), .b ({new_AGEMA_signal_5233, SubBytesIns_Inst_Sbox_8_T16}), .c ({new_AGEMA_signal_5455, SubBytesIns_Inst_Sbox_8_T26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T27_U1 ( .a ({new_AGEMA_signal_5053, SubBytesIns_Inst_Sbox_8_T1}), .b ({new_AGEMA_signal_5060, SubBytesIns_Inst_Sbox_8_T12}), .c ({new_AGEMA_signal_5236, SubBytesIns_Inst_Sbox_8_T27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T1_U1 ( .a ({ciphertext_s1[79], ciphertext_s0[79]}), .b ({ciphertext_s1[76], ciphertext_s0[76]}), .c ({new_AGEMA_signal_5063, SubBytesIns_Inst_Sbox_9_T1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T2_U1 ( .a ({ciphertext_s1[79], ciphertext_s0[79]}), .b ({ciphertext_s1[74], ciphertext_s0[74]}), .c ({new_AGEMA_signal_5064, SubBytesIns_Inst_Sbox_9_T2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T3_U1 ( .a ({ciphertext_s1[79], ciphertext_s0[79]}), .b ({ciphertext_s1[73], ciphertext_s0[73]}), .c ({new_AGEMA_signal_5065, SubBytesIns_Inst_Sbox_9_T3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T4_U1 ( .a ({ciphertext_s1[76], ciphertext_s0[76]}), .b ({ciphertext_s1[74], ciphertext_s0[74]}), .c ({new_AGEMA_signal_5066, SubBytesIns_Inst_Sbox_9_T4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T5_U1 ( .a ({ciphertext_s1[75], ciphertext_s0[75]}), .b ({ciphertext_s1[73], ciphertext_s0[73]}), .c ({new_AGEMA_signal_5067, SubBytesIns_Inst_Sbox_9_T5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T6_U1 ( .a ({new_AGEMA_signal_5063, SubBytesIns_Inst_Sbox_9_T1}), .b ({new_AGEMA_signal_5067, SubBytesIns_Inst_Sbox_9_T5}), .c ({new_AGEMA_signal_5237, SubBytesIns_Inst_Sbox_9_T6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T7_U1 ( .a ({ciphertext_s1[78], ciphertext_s0[78]}), .b ({ciphertext_s1[77], ciphertext_s0[77]}), .c ({new_AGEMA_signal_5068, SubBytesIns_Inst_Sbox_9_T7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T8_U1 ( .a ({ciphertext_s1[72], ciphertext_s0[72]}), .b ({new_AGEMA_signal_5237, SubBytesIns_Inst_Sbox_9_T6}), .c ({new_AGEMA_signal_5462, SubBytesIns_Inst_Sbox_9_T8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T9_U1 ( .a ({ciphertext_s1[72], ciphertext_s0[72]}), .b ({new_AGEMA_signal_5068, SubBytesIns_Inst_Sbox_9_T7}), .c ({new_AGEMA_signal_5238, SubBytesIns_Inst_Sbox_9_T9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T10_U1 ( .a ({new_AGEMA_signal_5237, SubBytesIns_Inst_Sbox_9_T6}), .b ({new_AGEMA_signal_5068, SubBytesIns_Inst_Sbox_9_T7}), .c ({new_AGEMA_signal_5463, SubBytesIns_Inst_Sbox_9_T10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T11_U1 ( .a ({ciphertext_s1[78], ciphertext_s0[78]}), .b ({ciphertext_s1[74], ciphertext_s0[74]}), .c ({new_AGEMA_signal_5069, SubBytesIns_Inst_Sbox_9_T11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T12_U1 ( .a ({ciphertext_s1[77], ciphertext_s0[77]}), .b ({ciphertext_s1[74], ciphertext_s0[74]}), .c ({new_AGEMA_signal_5070, SubBytesIns_Inst_Sbox_9_T12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T13_U1 ( .a ({new_AGEMA_signal_5065, SubBytesIns_Inst_Sbox_9_T3}), .b ({new_AGEMA_signal_5066, SubBytesIns_Inst_Sbox_9_T4}), .c ({new_AGEMA_signal_5239, SubBytesIns_Inst_Sbox_9_T13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T14_U1 ( .a ({new_AGEMA_signal_5237, SubBytesIns_Inst_Sbox_9_T6}), .b ({new_AGEMA_signal_5069, SubBytesIns_Inst_Sbox_9_T11}), .c ({new_AGEMA_signal_5464, SubBytesIns_Inst_Sbox_9_T14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T15_U1 ( .a ({new_AGEMA_signal_5067, SubBytesIns_Inst_Sbox_9_T5}), .b ({new_AGEMA_signal_5069, SubBytesIns_Inst_Sbox_9_T11}), .c ({new_AGEMA_signal_5240, SubBytesIns_Inst_Sbox_9_T15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T16_U1 ( .a ({new_AGEMA_signal_5067, SubBytesIns_Inst_Sbox_9_T5}), .b ({new_AGEMA_signal_5070, SubBytesIns_Inst_Sbox_9_T12}), .c ({new_AGEMA_signal_5241, SubBytesIns_Inst_Sbox_9_T16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T17_U1 ( .a ({new_AGEMA_signal_5238, SubBytesIns_Inst_Sbox_9_T9}), .b ({new_AGEMA_signal_5241, SubBytesIns_Inst_Sbox_9_T16}), .c ({new_AGEMA_signal_5465, SubBytesIns_Inst_Sbox_9_T17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T18_U1 ( .a ({ciphertext_s1[76], ciphertext_s0[76]}), .b ({ciphertext_s1[72], ciphertext_s0[72]}), .c ({new_AGEMA_signal_5071, SubBytesIns_Inst_Sbox_9_T18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T19_U1 ( .a ({new_AGEMA_signal_5068, SubBytesIns_Inst_Sbox_9_T7}), .b ({new_AGEMA_signal_5071, SubBytesIns_Inst_Sbox_9_T18}), .c ({new_AGEMA_signal_5242, SubBytesIns_Inst_Sbox_9_T19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T20_U1 ( .a ({new_AGEMA_signal_5063, SubBytesIns_Inst_Sbox_9_T1}), .b ({new_AGEMA_signal_5242, SubBytesIns_Inst_Sbox_9_T19}), .c ({new_AGEMA_signal_5466, SubBytesIns_Inst_Sbox_9_T20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T21_U1 ( .a ({ciphertext_s1[73], ciphertext_s0[73]}), .b ({ciphertext_s1[72], ciphertext_s0[72]}), .c ({new_AGEMA_signal_5072, SubBytesIns_Inst_Sbox_9_T21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T22_U1 ( .a ({new_AGEMA_signal_5068, SubBytesIns_Inst_Sbox_9_T7}), .b ({new_AGEMA_signal_5072, SubBytesIns_Inst_Sbox_9_T21}), .c ({new_AGEMA_signal_5243, SubBytesIns_Inst_Sbox_9_T22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T23_U1 ( .a ({new_AGEMA_signal_5064, SubBytesIns_Inst_Sbox_9_T2}), .b ({new_AGEMA_signal_5243, SubBytesIns_Inst_Sbox_9_T22}), .c ({new_AGEMA_signal_5467, SubBytesIns_Inst_Sbox_9_T23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T24_U1 ( .a ({new_AGEMA_signal_5064, SubBytesIns_Inst_Sbox_9_T2}), .b ({new_AGEMA_signal_5463, SubBytesIns_Inst_Sbox_9_T10}), .c ({new_AGEMA_signal_5670, SubBytesIns_Inst_Sbox_9_T24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T25_U1 ( .a ({new_AGEMA_signal_5466, SubBytesIns_Inst_Sbox_9_T20}), .b ({new_AGEMA_signal_5465, SubBytesIns_Inst_Sbox_9_T17}), .c ({new_AGEMA_signal_5671, SubBytesIns_Inst_Sbox_9_T25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T26_U1 ( .a ({new_AGEMA_signal_5065, SubBytesIns_Inst_Sbox_9_T3}), .b ({new_AGEMA_signal_5241, SubBytesIns_Inst_Sbox_9_T16}), .c ({new_AGEMA_signal_5468, SubBytesIns_Inst_Sbox_9_T26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T27_U1 ( .a ({new_AGEMA_signal_5063, SubBytesIns_Inst_Sbox_9_T1}), .b ({new_AGEMA_signal_5070, SubBytesIns_Inst_Sbox_9_T12}), .c ({new_AGEMA_signal_5244, SubBytesIns_Inst_Sbox_9_T27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T1_U1 ( .a ({ciphertext_s1[87], ciphertext_s0[87]}), .b ({ciphertext_s1[84], ciphertext_s0[84]}), .c ({new_AGEMA_signal_5073, SubBytesIns_Inst_Sbox_10_T1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T2_U1 ( .a ({ciphertext_s1[87], ciphertext_s0[87]}), .b ({ciphertext_s1[82], ciphertext_s0[82]}), .c ({new_AGEMA_signal_5074, SubBytesIns_Inst_Sbox_10_T2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T3_U1 ( .a ({ciphertext_s1[87], ciphertext_s0[87]}), .b ({ciphertext_s1[81], ciphertext_s0[81]}), .c ({new_AGEMA_signal_5075, SubBytesIns_Inst_Sbox_10_T3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T4_U1 ( .a ({ciphertext_s1[84], ciphertext_s0[84]}), .b ({ciphertext_s1[82], ciphertext_s0[82]}), .c ({new_AGEMA_signal_5076, SubBytesIns_Inst_Sbox_10_T4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T5_U1 ( .a ({ciphertext_s1[83], ciphertext_s0[83]}), .b ({ciphertext_s1[81], ciphertext_s0[81]}), .c ({new_AGEMA_signal_5077, SubBytesIns_Inst_Sbox_10_T5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T6_U1 ( .a ({new_AGEMA_signal_5073, SubBytesIns_Inst_Sbox_10_T1}), .b ({new_AGEMA_signal_5077, SubBytesIns_Inst_Sbox_10_T5}), .c ({new_AGEMA_signal_5245, SubBytesIns_Inst_Sbox_10_T6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T7_U1 ( .a ({ciphertext_s1[86], ciphertext_s0[86]}), .b ({ciphertext_s1[85], ciphertext_s0[85]}), .c ({new_AGEMA_signal_5078, SubBytesIns_Inst_Sbox_10_T7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T8_U1 ( .a ({ciphertext_s1[80], ciphertext_s0[80]}), .b ({new_AGEMA_signal_5245, SubBytesIns_Inst_Sbox_10_T6}), .c ({new_AGEMA_signal_5475, SubBytesIns_Inst_Sbox_10_T8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T9_U1 ( .a ({ciphertext_s1[80], ciphertext_s0[80]}), .b ({new_AGEMA_signal_5078, SubBytesIns_Inst_Sbox_10_T7}), .c ({new_AGEMA_signal_5246, SubBytesIns_Inst_Sbox_10_T9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T10_U1 ( .a ({new_AGEMA_signal_5245, SubBytesIns_Inst_Sbox_10_T6}), .b ({new_AGEMA_signal_5078, SubBytesIns_Inst_Sbox_10_T7}), .c ({new_AGEMA_signal_5476, SubBytesIns_Inst_Sbox_10_T10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T11_U1 ( .a ({ciphertext_s1[86], ciphertext_s0[86]}), .b ({ciphertext_s1[82], ciphertext_s0[82]}), .c ({new_AGEMA_signal_5079, SubBytesIns_Inst_Sbox_10_T11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T12_U1 ( .a ({ciphertext_s1[85], ciphertext_s0[85]}), .b ({ciphertext_s1[82], ciphertext_s0[82]}), .c ({new_AGEMA_signal_5080, SubBytesIns_Inst_Sbox_10_T12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T13_U1 ( .a ({new_AGEMA_signal_5075, SubBytesIns_Inst_Sbox_10_T3}), .b ({new_AGEMA_signal_5076, SubBytesIns_Inst_Sbox_10_T4}), .c ({new_AGEMA_signal_5247, SubBytesIns_Inst_Sbox_10_T13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T14_U1 ( .a ({new_AGEMA_signal_5245, SubBytesIns_Inst_Sbox_10_T6}), .b ({new_AGEMA_signal_5079, SubBytesIns_Inst_Sbox_10_T11}), .c ({new_AGEMA_signal_5477, SubBytesIns_Inst_Sbox_10_T14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T15_U1 ( .a ({new_AGEMA_signal_5077, SubBytesIns_Inst_Sbox_10_T5}), .b ({new_AGEMA_signal_5079, SubBytesIns_Inst_Sbox_10_T11}), .c ({new_AGEMA_signal_5248, SubBytesIns_Inst_Sbox_10_T15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T16_U1 ( .a ({new_AGEMA_signal_5077, SubBytesIns_Inst_Sbox_10_T5}), .b ({new_AGEMA_signal_5080, SubBytesIns_Inst_Sbox_10_T12}), .c ({new_AGEMA_signal_5249, SubBytesIns_Inst_Sbox_10_T16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T17_U1 ( .a ({new_AGEMA_signal_5246, SubBytesIns_Inst_Sbox_10_T9}), .b ({new_AGEMA_signal_5249, SubBytesIns_Inst_Sbox_10_T16}), .c ({new_AGEMA_signal_5478, SubBytesIns_Inst_Sbox_10_T17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T18_U1 ( .a ({ciphertext_s1[84], ciphertext_s0[84]}), .b ({ciphertext_s1[80], ciphertext_s0[80]}), .c ({new_AGEMA_signal_5081, SubBytesIns_Inst_Sbox_10_T18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T19_U1 ( .a ({new_AGEMA_signal_5078, SubBytesIns_Inst_Sbox_10_T7}), .b ({new_AGEMA_signal_5081, SubBytesIns_Inst_Sbox_10_T18}), .c ({new_AGEMA_signal_5250, SubBytesIns_Inst_Sbox_10_T19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T20_U1 ( .a ({new_AGEMA_signal_5073, SubBytesIns_Inst_Sbox_10_T1}), .b ({new_AGEMA_signal_5250, SubBytesIns_Inst_Sbox_10_T19}), .c ({new_AGEMA_signal_5479, SubBytesIns_Inst_Sbox_10_T20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T21_U1 ( .a ({ciphertext_s1[81], ciphertext_s0[81]}), .b ({ciphertext_s1[80], ciphertext_s0[80]}), .c ({new_AGEMA_signal_5082, SubBytesIns_Inst_Sbox_10_T21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T22_U1 ( .a ({new_AGEMA_signal_5078, SubBytesIns_Inst_Sbox_10_T7}), .b ({new_AGEMA_signal_5082, SubBytesIns_Inst_Sbox_10_T21}), .c ({new_AGEMA_signal_5251, SubBytesIns_Inst_Sbox_10_T22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T23_U1 ( .a ({new_AGEMA_signal_5074, SubBytesIns_Inst_Sbox_10_T2}), .b ({new_AGEMA_signal_5251, SubBytesIns_Inst_Sbox_10_T22}), .c ({new_AGEMA_signal_5480, SubBytesIns_Inst_Sbox_10_T23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T24_U1 ( .a ({new_AGEMA_signal_5074, SubBytesIns_Inst_Sbox_10_T2}), .b ({new_AGEMA_signal_5476, SubBytesIns_Inst_Sbox_10_T10}), .c ({new_AGEMA_signal_5679, SubBytesIns_Inst_Sbox_10_T24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T25_U1 ( .a ({new_AGEMA_signal_5479, SubBytesIns_Inst_Sbox_10_T20}), .b ({new_AGEMA_signal_5478, SubBytesIns_Inst_Sbox_10_T17}), .c ({new_AGEMA_signal_5680, SubBytesIns_Inst_Sbox_10_T25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T26_U1 ( .a ({new_AGEMA_signal_5075, SubBytesIns_Inst_Sbox_10_T3}), .b ({new_AGEMA_signal_5249, SubBytesIns_Inst_Sbox_10_T16}), .c ({new_AGEMA_signal_5481, SubBytesIns_Inst_Sbox_10_T26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T27_U1 ( .a ({new_AGEMA_signal_5073, SubBytesIns_Inst_Sbox_10_T1}), .b ({new_AGEMA_signal_5080, SubBytesIns_Inst_Sbox_10_T12}), .c ({new_AGEMA_signal_5252, SubBytesIns_Inst_Sbox_10_T27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T1_U1 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[92], ciphertext_s0[92]}), .c ({new_AGEMA_signal_5083, SubBytesIns_Inst_Sbox_11_T1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T2_U1 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_5084, SubBytesIns_Inst_Sbox_11_T2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T3_U1 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[89], ciphertext_s0[89]}), .c ({new_AGEMA_signal_5085, SubBytesIns_Inst_Sbox_11_T3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T4_U1 ( .a ({ciphertext_s1[92], ciphertext_s0[92]}), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_5086, SubBytesIns_Inst_Sbox_11_T4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T5_U1 ( .a ({ciphertext_s1[91], ciphertext_s0[91]}), .b ({ciphertext_s1[89], ciphertext_s0[89]}), .c ({new_AGEMA_signal_5087, SubBytesIns_Inst_Sbox_11_T5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T6_U1 ( .a ({new_AGEMA_signal_5083, SubBytesIns_Inst_Sbox_11_T1}), .b ({new_AGEMA_signal_5087, SubBytesIns_Inst_Sbox_11_T5}), .c ({new_AGEMA_signal_5253, SubBytesIns_Inst_Sbox_11_T6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T7_U1 ( .a ({ciphertext_s1[94], ciphertext_s0[94]}), .b ({ciphertext_s1[93], ciphertext_s0[93]}), .c ({new_AGEMA_signal_5088, SubBytesIns_Inst_Sbox_11_T7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T8_U1 ( .a ({ciphertext_s1[88], ciphertext_s0[88]}), .b ({new_AGEMA_signal_5253, SubBytesIns_Inst_Sbox_11_T6}), .c ({new_AGEMA_signal_5488, SubBytesIns_Inst_Sbox_11_T8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T9_U1 ( .a ({ciphertext_s1[88], ciphertext_s0[88]}), .b ({new_AGEMA_signal_5088, SubBytesIns_Inst_Sbox_11_T7}), .c ({new_AGEMA_signal_5254, SubBytesIns_Inst_Sbox_11_T9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T10_U1 ( .a ({new_AGEMA_signal_5253, SubBytesIns_Inst_Sbox_11_T6}), .b ({new_AGEMA_signal_5088, SubBytesIns_Inst_Sbox_11_T7}), .c ({new_AGEMA_signal_5489, SubBytesIns_Inst_Sbox_11_T10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T11_U1 ( .a ({ciphertext_s1[94], ciphertext_s0[94]}), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_5089, SubBytesIns_Inst_Sbox_11_T11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T12_U1 ( .a ({ciphertext_s1[93], ciphertext_s0[93]}), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_5090, SubBytesIns_Inst_Sbox_11_T12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T13_U1 ( .a ({new_AGEMA_signal_5085, SubBytesIns_Inst_Sbox_11_T3}), .b ({new_AGEMA_signal_5086, SubBytesIns_Inst_Sbox_11_T4}), .c ({new_AGEMA_signal_5255, SubBytesIns_Inst_Sbox_11_T13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T14_U1 ( .a ({new_AGEMA_signal_5253, SubBytesIns_Inst_Sbox_11_T6}), .b ({new_AGEMA_signal_5089, SubBytesIns_Inst_Sbox_11_T11}), .c ({new_AGEMA_signal_5490, SubBytesIns_Inst_Sbox_11_T14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T15_U1 ( .a ({new_AGEMA_signal_5087, SubBytesIns_Inst_Sbox_11_T5}), .b ({new_AGEMA_signal_5089, SubBytesIns_Inst_Sbox_11_T11}), .c ({new_AGEMA_signal_5256, SubBytesIns_Inst_Sbox_11_T15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T16_U1 ( .a ({new_AGEMA_signal_5087, SubBytesIns_Inst_Sbox_11_T5}), .b ({new_AGEMA_signal_5090, SubBytesIns_Inst_Sbox_11_T12}), .c ({new_AGEMA_signal_5257, SubBytesIns_Inst_Sbox_11_T16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T17_U1 ( .a ({new_AGEMA_signal_5254, SubBytesIns_Inst_Sbox_11_T9}), .b ({new_AGEMA_signal_5257, SubBytesIns_Inst_Sbox_11_T16}), .c ({new_AGEMA_signal_5491, SubBytesIns_Inst_Sbox_11_T17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T18_U1 ( .a ({ciphertext_s1[92], ciphertext_s0[92]}), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .c ({new_AGEMA_signal_5091, SubBytesIns_Inst_Sbox_11_T18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T19_U1 ( .a ({new_AGEMA_signal_5088, SubBytesIns_Inst_Sbox_11_T7}), .b ({new_AGEMA_signal_5091, SubBytesIns_Inst_Sbox_11_T18}), .c ({new_AGEMA_signal_5258, SubBytesIns_Inst_Sbox_11_T19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T20_U1 ( .a ({new_AGEMA_signal_5083, SubBytesIns_Inst_Sbox_11_T1}), .b ({new_AGEMA_signal_5258, SubBytesIns_Inst_Sbox_11_T19}), .c ({new_AGEMA_signal_5492, SubBytesIns_Inst_Sbox_11_T20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T21_U1 ( .a ({ciphertext_s1[89], ciphertext_s0[89]}), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .c ({new_AGEMA_signal_5092, SubBytesIns_Inst_Sbox_11_T21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T22_U1 ( .a ({new_AGEMA_signal_5088, SubBytesIns_Inst_Sbox_11_T7}), .b ({new_AGEMA_signal_5092, SubBytesIns_Inst_Sbox_11_T21}), .c ({new_AGEMA_signal_5259, SubBytesIns_Inst_Sbox_11_T22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T23_U1 ( .a ({new_AGEMA_signal_5084, SubBytesIns_Inst_Sbox_11_T2}), .b ({new_AGEMA_signal_5259, SubBytesIns_Inst_Sbox_11_T22}), .c ({new_AGEMA_signal_5493, SubBytesIns_Inst_Sbox_11_T23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T24_U1 ( .a ({new_AGEMA_signal_5084, SubBytesIns_Inst_Sbox_11_T2}), .b ({new_AGEMA_signal_5489, SubBytesIns_Inst_Sbox_11_T10}), .c ({new_AGEMA_signal_5688, SubBytesIns_Inst_Sbox_11_T24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T25_U1 ( .a ({new_AGEMA_signal_5492, SubBytesIns_Inst_Sbox_11_T20}), .b ({new_AGEMA_signal_5491, SubBytesIns_Inst_Sbox_11_T17}), .c ({new_AGEMA_signal_5689, SubBytesIns_Inst_Sbox_11_T25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T26_U1 ( .a ({new_AGEMA_signal_5085, SubBytesIns_Inst_Sbox_11_T3}), .b ({new_AGEMA_signal_5257, SubBytesIns_Inst_Sbox_11_T16}), .c ({new_AGEMA_signal_5494, SubBytesIns_Inst_Sbox_11_T26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T27_U1 ( .a ({new_AGEMA_signal_5083, SubBytesIns_Inst_Sbox_11_T1}), .b ({new_AGEMA_signal_5090, SubBytesIns_Inst_Sbox_11_T12}), .c ({new_AGEMA_signal_5260, SubBytesIns_Inst_Sbox_11_T27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T1_U1 ( .a ({ciphertext_s1[103], ciphertext_s0[103]}), .b ({ciphertext_s1[100], ciphertext_s0[100]}), .c ({new_AGEMA_signal_5093, SubBytesIns_Inst_Sbox_12_T1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T2_U1 ( .a ({ciphertext_s1[103], ciphertext_s0[103]}), .b ({ciphertext_s1[98], ciphertext_s0[98]}), .c ({new_AGEMA_signal_5094, SubBytesIns_Inst_Sbox_12_T2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T3_U1 ( .a ({ciphertext_s1[103], ciphertext_s0[103]}), .b ({ciphertext_s1[97], ciphertext_s0[97]}), .c ({new_AGEMA_signal_5095, SubBytesIns_Inst_Sbox_12_T3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T4_U1 ( .a ({ciphertext_s1[100], ciphertext_s0[100]}), .b ({ciphertext_s1[98], ciphertext_s0[98]}), .c ({new_AGEMA_signal_5096, SubBytesIns_Inst_Sbox_12_T4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T5_U1 ( .a ({ciphertext_s1[99], ciphertext_s0[99]}), .b ({ciphertext_s1[97], ciphertext_s0[97]}), .c ({new_AGEMA_signal_5097, SubBytesIns_Inst_Sbox_12_T5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T6_U1 ( .a ({new_AGEMA_signal_5093, SubBytesIns_Inst_Sbox_12_T1}), .b ({new_AGEMA_signal_5097, SubBytesIns_Inst_Sbox_12_T5}), .c ({new_AGEMA_signal_5261, SubBytesIns_Inst_Sbox_12_T6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T7_U1 ( .a ({ciphertext_s1[102], ciphertext_s0[102]}), .b ({ciphertext_s1[101], ciphertext_s0[101]}), .c ({new_AGEMA_signal_5098, SubBytesIns_Inst_Sbox_12_T7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T8_U1 ( .a ({ciphertext_s1[96], ciphertext_s0[96]}), .b ({new_AGEMA_signal_5261, SubBytesIns_Inst_Sbox_12_T6}), .c ({new_AGEMA_signal_5501, SubBytesIns_Inst_Sbox_12_T8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T9_U1 ( .a ({ciphertext_s1[96], ciphertext_s0[96]}), .b ({new_AGEMA_signal_5098, SubBytesIns_Inst_Sbox_12_T7}), .c ({new_AGEMA_signal_5262, SubBytesIns_Inst_Sbox_12_T9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T10_U1 ( .a ({new_AGEMA_signal_5261, SubBytesIns_Inst_Sbox_12_T6}), .b ({new_AGEMA_signal_5098, SubBytesIns_Inst_Sbox_12_T7}), .c ({new_AGEMA_signal_5502, SubBytesIns_Inst_Sbox_12_T10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T11_U1 ( .a ({ciphertext_s1[102], ciphertext_s0[102]}), .b ({ciphertext_s1[98], ciphertext_s0[98]}), .c ({new_AGEMA_signal_5099, SubBytesIns_Inst_Sbox_12_T11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T12_U1 ( .a ({ciphertext_s1[101], ciphertext_s0[101]}), .b ({ciphertext_s1[98], ciphertext_s0[98]}), .c ({new_AGEMA_signal_5100, SubBytesIns_Inst_Sbox_12_T12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T13_U1 ( .a ({new_AGEMA_signal_5095, SubBytesIns_Inst_Sbox_12_T3}), .b ({new_AGEMA_signal_5096, SubBytesIns_Inst_Sbox_12_T4}), .c ({new_AGEMA_signal_5263, SubBytesIns_Inst_Sbox_12_T13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T14_U1 ( .a ({new_AGEMA_signal_5261, SubBytesIns_Inst_Sbox_12_T6}), .b ({new_AGEMA_signal_5099, SubBytesIns_Inst_Sbox_12_T11}), .c ({new_AGEMA_signal_5503, SubBytesIns_Inst_Sbox_12_T14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T15_U1 ( .a ({new_AGEMA_signal_5097, SubBytesIns_Inst_Sbox_12_T5}), .b ({new_AGEMA_signal_5099, SubBytesIns_Inst_Sbox_12_T11}), .c ({new_AGEMA_signal_5264, SubBytesIns_Inst_Sbox_12_T15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T16_U1 ( .a ({new_AGEMA_signal_5097, SubBytesIns_Inst_Sbox_12_T5}), .b ({new_AGEMA_signal_5100, SubBytesIns_Inst_Sbox_12_T12}), .c ({new_AGEMA_signal_5265, SubBytesIns_Inst_Sbox_12_T16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T17_U1 ( .a ({new_AGEMA_signal_5262, SubBytesIns_Inst_Sbox_12_T9}), .b ({new_AGEMA_signal_5265, SubBytesIns_Inst_Sbox_12_T16}), .c ({new_AGEMA_signal_5504, SubBytesIns_Inst_Sbox_12_T17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T18_U1 ( .a ({ciphertext_s1[100], ciphertext_s0[100]}), .b ({ciphertext_s1[96], ciphertext_s0[96]}), .c ({new_AGEMA_signal_5101, SubBytesIns_Inst_Sbox_12_T18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T19_U1 ( .a ({new_AGEMA_signal_5098, SubBytesIns_Inst_Sbox_12_T7}), .b ({new_AGEMA_signal_5101, SubBytesIns_Inst_Sbox_12_T18}), .c ({new_AGEMA_signal_5266, SubBytesIns_Inst_Sbox_12_T19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T20_U1 ( .a ({new_AGEMA_signal_5093, SubBytesIns_Inst_Sbox_12_T1}), .b ({new_AGEMA_signal_5266, SubBytesIns_Inst_Sbox_12_T19}), .c ({new_AGEMA_signal_5505, SubBytesIns_Inst_Sbox_12_T20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T21_U1 ( .a ({ciphertext_s1[97], ciphertext_s0[97]}), .b ({ciphertext_s1[96], ciphertext_s0[96]}), .c ({new_AGEMA_signal_5102, SubBytesIns_Inst_Sbox_12_T21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T22_U1 ( .a ({new_AGEMA_signal_5098, SubBytesIns_Inst_Sbox_12_T7}), .b ({new_AGEMA_signal_5102, SubBytesIns_Inst_Sbox_12_T21}), .c ({new_AGEMA_signal_5267, SubBytesIns_Inst_Sbox_12_T22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T23_U1 ( .a ({new_AGEMA_signal_5094, SubBytesIns_Inst_Sbox_12_T2}), .b ({new_AGEMA_signal_5267, SubBytesIns_Inst_Sbox_12_T22}), .c ({new_AGEMA_signal_5506, SubBytesIns_Inst_Sbox_12_T23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T24_U1 ( .a ({new_AGEMA_signal_5094, SubBytesIns_Inst_Sbox_12_T2}), .b ({new_AGEMA_signal_5502, SubBytesIns_Inst_Sbox_12_T10}), .c ({new_AGEMA_signal_5697, SubBytesIns_Inst_Sbox_12_T24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T25_U1 ( .a ({new_AGEMA_signal_5505, SubBytesIns_Inst_Sbox_12_T20}), .b ({new_AGEMA_signal_5504, SubBytesIns_Inst_Sbox_12_T17}), .c ({new_AGEMA_signal_5698, SubBytesIns_Inst_Sbox_12_T25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T26_U1 ( .a ({new_AGEMA_signal_5095, SubBytesIns_Inst_Sbox_12_T3}), .b ({new_AGEMA_signal_5265, SubBytesIns_Inst_Sbox_12_T16}), .c ({new_AGEMA_signal_5507, SubBytesIns_Inst_Sbox_12_T26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T27_U1 ( .a ({new_AGEMA_signal_5093, SubBytesIns_Inst_Sbox_12_T1}), .b ({new_AGEMA_signal_5100, SubBytesIns_Inst_Sbox_12_T12}), .c ({new_AGEMA_signal_5268, SubBytesIns_Inst_Sbox_12_T27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T1_U1 ( .a ({ciphertext_s1[111], ciphertext_s0[111]}), .b ({ciphertext_s1[108], ciphertext_s0[108]}), .c ({new_AGEMA_signal_5103, SubBytesIns_Inst_Sbox_13_T1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T2_U1 ( .a ({ciphertext_s1[111], ciphertext_s0[111]}), .b ({ciphertext_s1[106], ciphertext_s0[106]}), .c ({new_AGEMA_signal_5104, SubBytesIns_Inst_Sbox_13_T2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T3_U1 ( .a ({ciphertext_s1[111], ciphertext_s0[111]}), .b ({ciphertext_s1[105], ciphertext_s0[105]}), .c ({new_AGEMA_signal_5105, SubBytesIns_Inst_Sbox_13_T3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T4_U1 ( .a ({ciphertext_s1[108], ciphertext_s0[108]}), .b ({ciphertext_s1[106], ciphertext_s0[106]}), .c ({new_AGEMA_signal_5106, SubBytesIns_Inst_Sbox_13_T4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T5_U1 ( .a ({ciphertext_s1[107], ciphertext_s0[107]}), .b ({ciphertext_s1[105], ciphertext_s0[105]}), .c ({new_AGEMA_signal_5107, SubBytesIns_Inst_Sbox_13_T5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T6_U1 ( .a ({new_AGEMA_signal_5103, SubBytesIns_Inst_Sbox_13_T1}), .b ({new_AGEMA_signal_5107, SubBytesIns_Inst_Sbox_13_T5}), .c ({new_AGEMA_signal_5269, SubBytesIns_Inst_Sbox_13_T6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T7_U1 ( .a ({ciphertext_s1[110], ciphertext_s0[110]}), .b ({ciphertext_s1[109], ciphertext_s0[109]}), .c ({new_AGEMA_signal_5108, SubBytesIns_Inst_Sbox_13_T7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T8_U1 ( .a ({ciphertext_s1[104], ciphertext_s0[104]}), .b ({new_AGEMA_signal_5269, SubBytesIns_Inst_Sbox_13_T6}), .c ({new_AGEMA_signal_5514, SubBytesIns_Inst_Sbox_13_T8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T9_U1 ( .a ({ciphertext_s1[104], ciphertext_s0[104]}), .b ({new_AGEMA_signal_5108, SubBytesIns_Inst_Sbox_13_T7}), .c ({new_AGEMA_signal_5270, SubBytesIns_Inst_Sbox_13_T9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T10_U1 ( .a ({new_AGEMA_signal_5269, SubBytesIns_Inst_Sbox_13_T6}), .b ({new_AGEMA_signal_5108, SubBytesIns_Inst_Sbox_13_T7}), .c ({new_AGEMA_signal_5515, SubBytesIns_Inst_Sbox_13_T10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T11_U1 ( .a ({ciphertext_s1[110], ciphertext_s0[110]}), .b ({ciphertext_s1[106], ciphertext_s0[106]}), .c ({new_AGEMA_signal_5109, SubBytesIns_Inst_Sbox_13_T11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T12_U1 ( .a ({ciphertext_s1[109], ciphertext_s0[109]}), .b ({ciphertext_s1[106], ciphertext_s0[106]}), .c ({new_AGEMA_signal_5110, SubBytesIns_Inst_Sbox_13_T12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T13_U1 ( .a ({new_AGEMA_signal_5105, SubBytesIns_Inst_Sbox_13_T3}), .b ({new_AGEMA_signal_5106, SubBytesIns_Inst_Sbox_13_T4}), .c ({new_AGEMA_signal_5271, SubBytesIns_Inst_Sbox_13_T13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T14_U1 ( .a ({new_AGEMA_signal_5269, SubBytesIns_Inst_Sbox_13_T6}), .b ({new_AGEMA_signal_5109, SubBytesIns_Inst_Sbox_13_T11}), .c ({new_AGEMA_signal_5516, SubBytesIns_Inst_Sbox_13_T14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T15_U1 ( .a ({new_AGEMA_signal_5107, SubBytesIns_Inst_Sbox_13_T5}), .b ({new_AGEMA_signal_5109, SubBytesIns_Inst_Sbox_13_T11}), .c ({new_AGEMA_signal_5272, SubBytesIns_Inst_Sbox_13_T15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T16_U1 ( .a ({new_AGEMA_signal_5107, SubBytesIns_Inst_Sbox_13_T5}), .b ({new_AGEMA_signal_5110, SubBytesIns_Inst_Sbox_13_T12}), .c ({new_AGEMA_signal_5273, SubBytesIns_Inst_Sbox_13_T16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T17_U1 ( .a ({new_AGEMA_signal_5270, SubBytesIns_Inst_Sbox_13_T9}), .b ({new_AGEMA_signal_5273, SubBytesIns_Inst_Sbox_13_T16}), .c ({new_AGEMA_signal_5517, SubBytesIns_Inst_Sbox_13_T17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T18_U1 ( .a ({ciphertext_s1[108], ciphertext_s0[108]}), .b ({ciphertext_s1[104], ciphertext_s0[104]}), .c ({new_AGEMA_signal_5111, SubBytesIns_Inst_Sbox_13_T18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T19_U1 ( .a ({new_AGEMA_signal_5108, SubBytesIns_Inst_Sbox_13_T7}), .b ({new_AGEMA_signal_5111, SubBytesIns_Inst_Sbox_13_T18}), .c ({new_AGEMA_signal_5274, SubBytesIns_Inst_Sbox_13_T19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T20_U1 ( .a ({new_AGEMA_signal_5103, SubBytesIns_Inst_Sbox_13_T1}), .b ({new_AGEMA_signal_5274, SubBytesIns_Inst_Sbox_13_T19}), .c ({new_AGEMA_signal_5518, SubBytesIns_Inst_Sbox_13_T20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T21_U1 ( .a ({ciphertext_s1[105], ciphertext_s0[105]}), .b ({ciphertext_s1[104], ciphertext_s0[104]}), .c ({new_AGEMA_signal_5112, SubBytesIns_Inst_Sbox_13_T21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T22_U1 ( .a ({new_AGEMA_signal_5108, SubBytesIns_Inst_Sbox_13_T7}), .b ({new_AGEMA_signal_5112, SubBytesIns_Inst_Sbox_13_T21}), .c ({new_AGEMA_signal_5275, SubBytesIns_Inst_Sbox_13_T22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T23_U1 ( .a ({new_AGEMA_signal_5104, SubBytesIns_Inst_Sbox_13_T2}), .b ({new_AGEMA_signal_5275, SubBytesIns_Inst_Sbox_13_T22}), .c ({new_AGEMA_signal_5519, SubBytesIns_Inst_Sbox_13_T23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T24_U1 ( .a ({new_AGEMA_signal_5104, SubBytesIns_Inst_Sbox_13_T2}), .b ({new_AGEMA_signal_5515, SubBytesIns_Inst_Sbox_13_T10}), .c ({new_AGEMA_signal_5706, SubBytesIns_Inst_Sbox_13_T24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T25_U1 ( .a ({new_AGEMA_signal_5518, SubBytesIns_Inst_Sbox_13_T20}), .b ({new_AGEMA_signal_5517, SubBytesIns_Inst_Sbox_13_T17}), .c ({new_AGEMA_signal_5707, SubBytesIns_Inst_Sbox_13_T25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T26_U1 ( .a ({new_AGEMA_signal_5105, SubBytesIns_Inst_Sbox_13_T3}), .b ({new_AGEMA_signal_5273, SubBytesIns_Inst_Sbox_13_T16}), .c ({new_AGEMA_signal_5520, SubBytesIns_Inst_Sbox_13_T26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T27_U1 ( .a ({new_AGEMA_signal_5103, SubBytesIns_Inst_Sbox_13_T1}), .b ({new_AGEMA_signal_5110, SubBytesIns_Inst_Sbox_13_T12}), .c ({new_AGEMA_signal_5276, SubBytesIns_Inst_Sbox_13_T27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T1_U1 ( .a ({ciphertext_s1[119], ciphertext_s0[119]}), .b ({ciphertext_s1[116], ciphertext_s0[116]}), .c ({new_AGEMA_signal_5113, SubBytesIns_Inst_Sbox_14_T1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T2_U1 ( .a ({ciphertext_s1[119], ciphertext_s0[119]}), .b ({ciphertext_s1[114], ciphertext_s0[114]}), .c ({new_AGEMA_signal_5114, SubBytesIns_Inst_Sbox_14_T2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T3_U1 ( .a ({ciphertext_s1[119], ciphertext_s0[119]}), .b ({ciphertext_s1[113], ciphertext_s0[113]}), .c ({new_AGEMA_signal_5115, SubBytesIns_Inst_Sbox_14_T3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T4_U1 ( .a ({ciphertext_s1[116], ciphertext_s0[116]}), .b ({ciphertext_s1[114], ciphertext_s0[114]}), .c ({new_AGEMA_signal_5116, SubBytesIns_Inst_Sbox_14_T4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T5_U1 ( .a ({ciphertext_s1[115], ciphertext_s0[115]}), .b ({ciphertext_s1[113], ciphertext_s0[113]}), .c ({new_AGEMA_signal_5117, SubBytesIns_Inst_Sbox_14_T5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T6_U1 ( .a ({new_AGEMA_signal_5113, SubBytesIns_Inst_Sbox_14_T1}), .b ({new_AGEMA_signal_5117, SubBytesIns_Inst_Sbox_14_T5}), .c ({new_AGEMA_signal_5277, SubBytesIns_Inst_Sbox_14_T6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T7_U1 ( .a ({ciphertext_s1[118], ciphertext_s0[118]}), .b ({ciphertext_s1[117], ciphertext_s0[117]}), .c ({new_AGEMA_signal_5118, SubBytesIns_Inst_Sbox_14_T7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T8_U1 ( .a ({ciphertext_s1[112], ciphertext_s0[112]}), .b ({new_AGEMA_signal_5277, SubBytesIns_Inst_Sbox_14_T6}), .c ({new_AGEMA_signal_5527, SubBytesIns_Inst_Sbox_14_T8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T9_U1 ( .a ({ciphertext_s1[112], ciphertext_s0[112]}), .b ({new_AGEMA_signal_5118, SubBytesIns_Inst_Sbox_14_T7}), .c ({new_AGEMA_signal_5278, SubBytesIns_Inst_Sbox_14_T9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T10_U1 ( .a ({new_AGEMA_signal_5277, SubBytesIns_Inst_Sbox_14_T6}), .b ({new_AGEMA_signal_5118, SubBytesIns_Inst_Sbox_14_T7}), .c ({new_AGEMA_signal_5528, SubBytesIns_Inst_Sbox_14_T10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T11_U1 ( .a ({ciphertext_s1[118], ciphertext_s0[118]}), .b ({ciphertext_s1[114], ciphertext_s0[114]}), .c ({new_AGEMA_signal_5119, SubBytesIns_Inst_Sbox_14_T11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T12_U1 ( .a ({ciphertext_s1[117], ciphertext_s0[117]}), .b ({ciphertext_s1[114], ciphertext_s0[114]}), .c ({new_AGEMA_signal_5120, SubBytesIns_Inst_Sbox_14_T12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T13_U1 ( .a ({new_AGEMA_signal_5115, SubBytesIns_Inst_Sbox_14_T3}), .b ({new_AGEMA_signal_5116, SubBytesIns_Inst_Sbox_14_T4}), .c ({new_AGEMA_signal_5279, SubBytesIns_Inst_Sbox_14_T13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T14_U1 ( .a ({new_AGEMA_signal_5277, SubBytesIns_Inst_Sbox_14_T6}), .b ({new_AGEMA_signal_5119, SubBytesIns_Inst_Sbox_14_T11}), .c ({new_AGEMA_signal_5529, SubBytesIns_Inst_Sbox_14_T14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T15_U1 ( .a ({new_AGEMA_signal_5117, SubBytesIns_Inst_Sbox_14_T5}), .b ({new_AGEMA_signal_5119, SubBytesIns_Inst_Sbox_14_T11}), .c ({new_AGEMA_signal_5280, SubBytesIns_Inst_Sbox_14_T15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T16_U1 ( .a ({new_AGEMA_signal_5117, SubBytesIns_Inst_Sbox_14_T5}), .b ({new_AGEMA_signal_5120, SubBytesIns_Inst_Sbox_14_T12}), .c ({new_AGEMA_signal_5281, SubBytesIns_Inst_Sbox_14_T16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T17_U1 ( .a ({new_AGEMA_signal_5278, SubBytesIns_Inst_Sbox_14_T9}), .b ({new_AGEMA_signal_5281, SubBytesIns_Inst_Sbox_14_T16}), .c ({new_AGEMA_signal_5530, SubBytesIns_Inst_Sbox_14_T17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T18_U1 ( .a ({ciphertext_s1[116], ciphertext_s0[116]}), .b ({ciphertext_s1[112], ciphertext_s0[112]}), .c ({new_AGEMA_signal_5121, SubBytesIns_Inst_Sbox_14_T18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T19_U1 ( .a ({new_AGEMA_signal_5118, SubBytesIns_Inst_Sbox_14_T7}), .b ({new_AGEMA_signal_5121, SubBytesIns_Inst_Sbox_14_T18}), .c ({new_AGEMA_signal_5282, SubBytesIns_Inst_Sbox_14_T19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T20_U1 ( .a ({new_AGEMA_signal_5113, SubBytesIns_Inst_Sbox_14_T1}), .b ({new_AGEMA_signal_5282, SubBytesIns_Inst_Sbox_14_T19}), .c ({new_AGEMA_signal_5531, SubBytesIns_Inst_Sbox_14_T20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T21_U1 ( .a ({ciphertext_s1[113], ciphertext_s0[113]}), .b ({ciphertext_s1[112], ciphertext_s0[112]}), .c ({new_AGEMA_signal_5122, SubBytesIns_Inst_Sbox_14_T21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T22_U1 ( .a ({new_AGEMA_signal_5118, SubBytesIns_Inst_Sbox_14_T7}), .b ({new_AGEMA_signal_5122, SubBytesIns_Inst_Sbox_14_T21}), .c ({new_AGEMA_signal_5283, SubBytesIns_Inst_Sbox_14_T22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T23_U1 ( .a ({new_AGEMA_signal_5114, SubBytesIns_Inst_Sbox_14_T2}), .b ({new_AGEMA_signal_5283, SubBytesIns_Inst_Sbox_14_T22}), .c ({new_AGEMA_signal_5532, SubBytesIns_Inst_Sbox_14_T23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T24_U1 ( .a ({new_AGEMA_signal_5114, SubBytesIns_Inst_Sbox_14_T2}), .b ({new_AGEMA_signal_5528, SubBytesIns_Inst_Sbox_14_T10}), .c ({new_AGEMA_signal_5715, SubBytesIns_Inst_Sbox_14_T24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T25_U1 ( .a ({new_AGEMA_signal_5531, SubBytesIns_Inst_Sbox_14_T20}), .b ({new_AGEMA_signal_5530, SubBytesIns_Inst_Sbox_14_T17}), .c ({new_AGEMA_signal_5716, SubBytesIns_Inst_Sbox_14_T25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T26_U1 ( .a ({new_AGEMA_signal_5115, SubBytesIns_Inst_Sbox_14_T3}), .b ({new_AGEMA_signal_5281, SubBytesIns_Inst_Sbox_14_T16}), .c ({new_AGEMA_signal_5533, SubBytesIns_Inst_Sbox_14_T26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T27_U1 ( .a ({new_AGEMA_signal_5113, SubBytesIns_Inst_Sbox_14_T1}), .b ({new_AGEMA_signal_5120, SubBytesIns_Inst_Sbox_14_T12}), .c ({new_AGEMA_signal_5284, SubBytesIns_Inst_Sbox_14_T27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T1_U1 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[124], ciphertext_s0[124]}), .c ({new_AGEMA_signal_5123, SubBytesIns_Inst_Sbox_15_T1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T2_U1 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_5124, SubBytesIns_Inst_Sbox_15_T2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T3_U1 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[121], ciphertext_s0[121]}), .c ({new_AGEMA_signal_5125, SubBytesIns_Inst_Sbox_15_T3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T4_U1 ( .a ({ciphertext_s1[124], ciphertext_s0[124]}), .b ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_5126, SubBytesIns_Inst_Sbox_15_T4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T5_U1 ( .a ({ciphertext_s1[123], ciphertext_s0[123]}), .b ({ciphertext_s1[121], ciphertext_s0[121]}), .c ({new_AGEMA_signal_5127, SubBytesIns_Inst_Sbox_15_T5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T6_U1 ( .a ({new_AGEMA_signal_5123, SubBytesIns_Inst_Sbox_15_T1}), .b ({new_AGEMA_signal_5127, SubBytesIns_Inst_Sbox_15_T5}), .c ({new_AGEMA_signal_5285, SubBytesIns_Inst_Sbox_15_T6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T7_U1 ( .a ({ciphertext_s1[126], ciphertext_s0[126]}), .b ({ciphertext_s1[125], ciphertext_s0[125]}), .c ({new_AGEMA_signal_5128, SubBytesIns_Inst_Sbox_15_T7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T8_U1 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({new_AGEMA_signal_5285, SubBytesIns_Inst_Sbox_15_T6}), .c ({new_AGEMA_signal_5540, SubBytesIns_Inst_Sbox_15_T8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T9_U1 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({new_AGEMA_signal_5128, SubBytesIns_Inst_Sbox_15_T7}), .c ({new_AGEMA_signal_5286, SubBytesIns_Inst_Sbox_15_T9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T10_U1 ( .a ({new_AGEMA_signal_5285, SubBytesIns_Inst_Sbox_15_T6}), .b ({new_AGEMA_signal_5128, SubBytesIns_Inst_Sbox_15_T7}), .c ({new_AGEMA_signal_5541, SubBytesIns_Inst_Sbox_15_T10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T11_U1 ( .a ({ciphertext_s1[126], ciphertext_s0[126]}), .b ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_5129, SubBytesIns_Inst_Sbox_15_T11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T12_U1 ( .a ({ciphertext_s1[125], ciphertext_s0[125]}), .b ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_5130, SubBytesIns_Inst_Sbox_15_T12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T13_U1 ( .a ({new_AGEMA_signal_5125, SubBytesIns_Inst_Sbox_15_T3}), .b ({new_AGEMA_signal_5126, SubBytesIns_Inst_Sbox_15_T4}), .c ({new_AGEMA_signal_5287, SubBytesIns_Inst_Sbox_15_T13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T14_U1 ( .a ({new_AGEMA_signal_5285, SubBytesIns_Inst_Sbox_15_T6}), .b ({new_AGEMA_signal_5129, SubBytesIns_Inst_Sbox_15_T11}), .c ({new_AGEMA_signal_5542, SubBytesIns_Inst_Sbox_15_T14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T15_U1 ( .a ({new_AGEMA_signal_5127, SubBytesIns_Inst_Sbox_15_T5}), .b ({new_AGEMA_signal_5129, SubBytesIns_Inst_Sbox_15_T11}), .c ({new_AGEMA_signal_5288, SubBytesIns_Inst_Sbox_15_T15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T16_U1 ( .a ({new_AGEMA_signal_5127, SubBytesIns_Inst_Sbox_15_T5}), .b ({new_AGEMA_signal_5130, SubBytesIns_Inst_Sbox_15_T12}), .c ({new_AGEMA_signal_5289, SubBytesIns_Inst_Sbox_15_T16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T17_U1 ( .a ({new_AGEMA_signal_5286, SubBytesIns_Inst_Sbox_15_T9}), .b ({new_AGEMA_signal_5289, SubBytesIns_Inst_Sbox_15_T16}), .c ({new_AGEMA_signal_5543, SubBytesIns_Inst_Sbox_15_T17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T18_U1 ( .a ({ciphertext_s1[124], ciphertext_s0[124]}), .b ({ciphertext_s1[120], ciphertext_s0[120]}), .c ({new_AGEMA_signal_5131, SubBytesIns_Inst_Sbox_15_T18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T19_U1 ( .a ({new_AGEMA_signal_5128, SubBytesIns_Inst_Sbox_15_T7}), .b ({new_AGEMA_signal_5131, SubBytesIns_Inst_Sbox_15_T18}), .c ({new_AGEMA_signal_5290, SubBytesIns_Inst_Sbox_15_T19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T20_U1 ( .a ({new_AGEMA_signal_5123, SubBytesIns_Inst_Sbox_15_T1}), .b ({new_AGEMA_signal_5290, SubBytesIns_Inst_Sbox_15_T19}), .c ({new_AGEMA_signal_5544, SubBytesIns_Inst_Sbox_15_T20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T21_U1 ( .a ({ciphertext_s1[121], ciphertext_s0[121]}), .b ({ciphertext_s1[120], ciphertext_s0[120]}), .c ({new_AGEMA_signal_5132, SubBytesIns_Inst_Sbox_15_T21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T22_U1 ( .a ({new_AGEMA_signal_5128, SubBytesIns_Inst_Sbox_15_T7}), .b ({new_AGEMA_signal_5132, SubBytesIns_Inst_Sbox_15_T21}), .c ({new_AGEMA_signal_5291, SubBytesIns_Inst_Sbox_15_T22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T23_U1 ( .a ({new_AGEMA_signal_5124, SubBytesIns_Inst_Sbox_15_T2}), .b ({new_AGEMA_signal_5291, SubBytesIns_Inst_Sbox_15_T22}), .c ({new_AGEMA_signal_5545, SubBytesIns_Inst_Sbox_15_T23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T24_U1 ( .a ({new_AGEMA_signal_5124, SubBytesIns_Inst_Sbox_15_T2}), .b ({new_AGEMA_signal_5541, SubBytesIns_Inst_Sbox_15_T10}), .c ({new_AGEMA_signal_5724, SubBytesIns_Inst_Sbox_15_T24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T25_U1 ( .a ({new_AGEMA_signal_5544, SubBytesIns_Inst_Sbox_15_T20}), .b ({new_AGEMA_signal_5543, SubBytesIns_Inst_Sbox_15_T17}), .c ({new_AGEMA_signal_5725, SubBytesIns_Inst_Sbox_15_T25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T26_U1 ( .a ({new_AGEMA_signal_5125, SubBytesIns_Inst_Sbox_15_T3}), .b ({new_AGEMA_signal_5289, SubBytesIns_Inst_Sbox_15_T16}), .c ({new_AGEMA_signal_5546, SubBytesIns_Inst_Sbox_15_T26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T27_U1 ( .a ({new_AGEMA_signal_5123, SubBytesIns_Inst_Sbox_15_T1}), .b ({new_AGEMA_signal_5130, SubBytesIns_Inst_Sbox_15_T12}), .c ({new_AGEMA_signal_5292, SubBytesIns_Inst_Sbox_15_T27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T1_U1 ( .a ({new_AGEMA_signal_4679, RoundKey[23]}), .b ({new_AGEMA_signal_4670, RoundKey[20]}), .c ({new_AGEMA_signal_4933, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T2_U1 ( .a ({new_AGEMA_signal_4679, RoundKey[23]}), .b ({new_AGEMA_signal_4661, RoundKey[18]}), .c ({new_AGEMA_signal_4934, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T3_U1 ( .a ({new_AGEMA_signal_4679, RoundKey[23]}), .b ({new_AGEMA_signal_4658, RoundKey[17]}), .c ({new_AGEMA_signal_4935, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T4_U1 ( .a ({new_AGEMA_signal_4670, RoundKey[20]}), .b ({new_AGEMA_signal_4661, RoundKey[18]}), .c ({new_AGEMA_signal_4936, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T5_U1 ( .a ({new_AGEMA_signal_4664, RoundKey[19]}), .b ({new_AGEMA_signal_4658, RoundKey[17]}), .c ({new_AGEMA_signal_4937, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T6_U1 ( .a ({new_AGEMA_signal_4933, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_4937, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5}), .c ({new_AGEMA_signal_5133, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T7_U1 ( .a ({new_AGEMA_signal_4676, RoundKey[22]}), .b ({new_AGEMA_signal_4673, RoundKey[21]}), .c ({new_AGEMA_signal_4938, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T8_U1 ( .a ({new_AGEMA_signal_4655, RoundKey[16]}), .b ({new_AGEMA_signal_5133, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}), .c ({new_AGEMA_signal_5293, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T9_U1 ( .a ({new_AGEMA_signal_4655, RoundKey[16]}), .b ({new_AGEMA_signal_4938, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_5134, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T10_U1 ( .a ({new_AGEMA_signal_5133, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_4938, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_5294, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T11_U1 ( .a ({new_AGEMA_signal_4676, RoundKey[22]}), .b ({new_AGEMA_signal_4661, RoundKey[18]}), .c ({new_AGEMA_signal_4939, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T12_U1 ( .a ({new_AGEMA_signal_4673, RoundKey[21]}), .b ({new_AGEMA_signal_4661, RoundKey[18]}), .c ({new_AGEMA_signal_4940, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T13_U1 ( .a ({new_AGEMA_signal_4935, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_4936, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4}), .c ({new_AGEMA_signal_5135, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T14_U1 ( .a ({new_AGEMA_signal_5133, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_4939, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_5295, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T15_U1 ( .a ({new_AGEMA_signal_4937, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_4939, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_5136, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T16_U1 ( .a ({new_AGEMA_signal_4937, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_4940, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_5137, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T17_U1 ( .a ({new_AGEMA_signal_5134, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9}), .b ({new_AGEMA_signal_5137, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_5296, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T18_U1 ( .a ({new_AGEMA_signal_4670, RoundKey[20]}), .b ({new_AGEMA_signal_4655, RoundKey[16]}), .c ({new_AGEMA_signal_4941, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T19_U1 ( .a ({new_AGEMA_signal_4938, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_4941, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T18}), .c ({new_AGEMA_signal_5138, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T20_U1 ( .a ({new_AGEMA_signal_4933, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_5138, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19}), .c ({new_AGEMA_signal_5297, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T21_U1 ( .a ({new_AGEMA_signal_4658, RoundKey[17]}), .b ({new_AGEMA_signal_4655, RoundKey[16]}), .c ({new_AGEMA_signal_4942, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T22_U1 ( .a ({new_AGEMA_signal_4938, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_4942, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T21}), .c ({new_AGEMA_signal_5139, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T23_U1 ( .a ({new_AGEMA_signal_4934, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_5139, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22}), .c ({new_AGEMA_signal_5298, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T24_U1 ( .a ({new_AGEMA_signal_4934, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_5294, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10}), .c ({new_AGEMA_signal_5553, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T25_U1 ( .a ({new_AGEMA_signal_5297, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_5296, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17}), .c ({new_AGEMA_signal_5554, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T26_U1 ( .a ({new_AGEMA_signal_4935, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_5137, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_5299, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T27_U1 ( .a ({new_AGEMA_signal_4933, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_4940, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_5140, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T1_U1 ( .a ({new_AGEMA_signal_4652, RoundKey[15]}), .b ({new_AGEMA_signal_4643, RoundKey[12]}), .c ({new_AGEMA_signal_4943, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T2_U1 ( .a ({new_AGEMA_signal_4652, RoundKey[15]}), .b ({new_AGEMA_signal_4583, RoundKey[10]}), .c ({new_AGEMA_signal_4944, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T3_U1 ( .a ({new_AGEMA_signal_4652, RoundKey[15]}), .b ({new_AGEMA_signal_4931, RoundKey[9]}), .c ({new_AGEMA_signal_4945, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T4_U1 ( .a ({new_AGEMA_signal_4643, RoundKey[12]}), .b ({new_AGEMA_signal_4583, RoundKey[10]}), .c ({new_AGEMA_signal_4946, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T5_U1 ( .a ({new_AGEMA_signal_4616, RoundKey[11]}), .b ({new_AGEMA_signal_4931, RoundKey[9]}), .c ({new_AGEMA_signal_4947, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T6_U1 ( .a ({new_AGEMA_signal_4943, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_4947, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5}), .c ({new_AGEMA_signal_5141, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T7_U1 ( .a ({new_AGEMA_signal_4649, RoundKey[14]}), .b ({new_AGEMA_signal_4646, RoundKey[13]}), .c ({new_AGEMA_signal_4948, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T8_U1 ( .a ({new_AGEMA_signal_4898, RoundKey[8]}), .b ({new_AGEMA_signal_5141, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}), .c ({new_AGEMA_signal_5306, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T9_U1 ( .a ({new_AGEMA_signal_4898, RoundKey[8]}), .b ({new_AGEMA_signal_4948, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_5142, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T10_U1 ( .a ({new_AGEMA_signal_5141, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_4948, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_5307, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T11_U1 ( .a ({new_AGEMA_signal_4649, RoundKey[14]}), .b ({new_AGEMA_signal_4583, RoundKey[10]}), .c ({new_AGEMA_signal_4949, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T12_U1 ( .a ({new_AGEMA_signal_4646, RoundKey[13]}), .b ({new_AGEMA_signal_4583, RoundKey[10]}), .c ({new_AGEMA_signal_4950, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T13_U1 ( .a ({new_AGEMA_signal_4945, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_4946, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4}), .c ({new_AGEMA_signal_5143, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T14_U1 ( .a ({new_AGEMA_signal_5141, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_4949, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_5308, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T15_U1 ( .a ({new_AGEMA_signal_4947, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_4949, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_5144, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T16_U1 ( .a ({new_AGEMA_signal_4947, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_4950, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_5145, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T17_U1 ( .a ({new_AGEMA_signal_5142, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9}), .b ({new_AGEMA_signal_5145, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_5309, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T18_U1 ( .a ({new_AGEMA_signal_4643, RoundKey[12]}), .b ({new_AGEMA_signal_4898, RoundKey[8]}), .c ({new_AGEMA_signal_4951, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T19_U1 ( .a ({new_AGEMA_signal_4948, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_4951, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T18}), .c ({new_AGEMA_signal_5146, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T20_U1 ( .a ({new_AGEMA_signal_4943, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_5146, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19}), .c ({new_AGEMA_signal_5310, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T21_U1 ( .a ({new_AGEMA_signal_4931, RoundKey[9]}), .b ({new_AGEMA_signal_4898, RoundKey[8]}), .c ({new_AGEMA_signal_4952, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T22_U1 ( .a ({new_AGEMA_signal_4948, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_4952, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T21}), .c ({new_AGEMA_signal_5147, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T23_U1 ( .a ({new_AGEMA_signal_4944, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_5147, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22}), .c ({new_AGEMA_signal_5311, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T24_U1 ( .a ({new_AGEMA_signal_4944, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_5307, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10}), .c ({new_AGEMA_signal_5562, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T25_U1 ( .a ({new_AGEMA_signal_5310, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_5309, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17}), .c ({new_AGEMA_signal_5563, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T26_U1 ( .a ({new_AGEMA_signal_4945, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_5145, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_5312, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T27_U1 ( .a ({new_AGEMA_signal_4943, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_4950, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_5148, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T1_U1 ( .a ({new_AGEMA_signal_4865, RoundKey[7]}), .b ({new_AGEMA_signal_4766, RoundKey[4]}), .c ({new_AGEMA_signal_4953, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T2_U1 ( .a ({new_AGEMA_signal_4865, RoundKey[7]}), .b ({new_AGEMA_signal_4700, RoundKey[2]}), .c ({new_AGEMA_signal_4954, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T3_U1 ( .a ({new_AGEMA_signal_4865, RoundKey[7]}), .b ({new_AGEMA_signal_4667, RoundKey[1]}), .c ({new_AGEMA_signal_4955, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T4_U1 ( .a ({new_AGEMA_signal_4766, RoundKey[4]}), .b ({new_AGEMA_signal_4700, RoundKey[2]}), .c ({new_AGEMA_signal_4956, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T5_U1 ( .a ({new_AGEMA_signal_4733, RoundKey[3]}), .b ({new_AGEMA_signal_4667, RoundKey[1]}), .c ({new_AGEMA_signal_4957, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T6_U1 ( .a ({new_AGEMA_signal_4953, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_4957, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5}), .c ({new_AGEMA_signal_5149, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T7_U1 ( .a ({new_AGEMA_signal_4832, RoundKey[6]}), .b ({new_AGEMA_signal_4799, RoundKey[5]}), .c ({new_AGEMA_signal_4958, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T8_U1 ( .a ({new_AGEMA_signal_4550, RoundKey[0]}), .b ({new_AGEMA_signal_5149, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}), .c ({new_AGEMA_signal_5319, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T9_U1 ( .a ({new_AGEMA_signal_4550, RoundKey[0]}), .b ({new_AGEMA_signal_4958, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_5150, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T10_U1 ( .a ({new_AGEMA_signal_5149, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_4958, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_5320, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T11_U1 ( .a ({new_AGEMA_signal_4832, RoundKey[6]}), .b ({new_AGEMA_signal_4700, RoundKey[2]}), .c ({new_AGEMA_signal_4959, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T12_U1 ( .a ({new_AGEMA_signal_4799, RoundKey[5]}), .b ({new_AGEMA_signal_4700, RoundKey[2]}), .c ({new_AGEMA_signal_4960, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T13_U1 ( .a ({new_AGEMA_signal_4955, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_4956, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4}), .c ({new_AGEMA_signal_5151, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T14_U1 ( .a ({new_AGEMA_signal_5149, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_4959, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_5321, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T15_U1 ( .a ({new_AGEMA_signal_4957, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_4959, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_5152, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T16_U1 ( .a ({new_AGEMA_signal_4957, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_4960, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_5153, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T17_U1 ( .a ({new_AGEMA_signal_5150, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9}), .b ({new_AGEMA_signal_5153, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_5322, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T18_U1 ( .a ({new_AGEMA_signal_4766, RoundKey[4]}), .b ({new_AGEMA_signal_4550, RoundKey[0]}), .c ({new_AGEMA_signal_4961, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T19_U1 ( .a ({new_AGEMA_signal_4958, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_4961, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T18}), .c ({new_AGEMA_signal_5154, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T20_U1 ( .a ({new_AGEMA_signal_4953, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5154, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19}), .c ({new_AGEMA_signal_5323, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T21_U1 ( .a ({new_AGEMA_signal_4667, RoundKey[1]}), .b ({new_AGEMA_signal_4550, RoundKey[0]}), .c ({new_AGEMA_signal_4962, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T22_U1 ( .a ({new_AGEMA_signal_4958, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_4962, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T21}), .c ({new_AGEMA_signal_5155, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T23_U1 ( .a ({new_AGEMA_signal_4954, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_5155, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22}), .c ({new_AGEMA_signal_5324, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T24_U1 ( .a ({new_AGEMA_signal_4954, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_5320, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10}), .c ({new_AGEMA_signal_5571, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T25_U1 ( .a ({new_AGEMA_signal_5323, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_5322, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17}), .c ({new_AGEMA_signal_5572, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T26_U1 ( .a ({new_AGEMA_signal_4955, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_5153, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_5325, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T27_U1 ( .a ({new_AGEMA_signal_4953, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_4960, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_5156, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T1_U1 ( .a ({new_AGEMA_signal_4706, RoundKey[31]}), .b ({new_AGEMA_signal_4694, RoundKey[28]}), .c ({new_AGEMA_signal_4963, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T2_U1 ( .a ({new_AGEMA_signal_4706, RoundKey[31]}), .b ({new_AGEMA_signal_4688, RoundKey[26]}), .c ({new_AGEMA_signal_4964, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T3_U1 ( .a ({new_AGEMA_signal_4706, RoundKey[31]}), .b ({new_AGEMA_signal_4685, RoundKey[25]}), .c ({new_AGEMA_signal_4965, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T4_U1 ( .a ({new_AGEMA_signal_4694, RoundKey[28]}), .b ({new_AGEMA_signal_4688, RoundKey[26]}), .c ({new_AGEMA_signal_4966, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T5_U1 ( .a ({new_AGEMA_signal_4691, RoundKey[27]}), .b ({new_AGEMA_signal_4685, RoundKey[25]}), .c ({new_AGEMA_signal_4967, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T6_U1 ( .a ({new_AGEMA_signal_4963, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_4967, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5}), .c ({new_AGEMA_signal_5157, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T7_U1 ( .a ({new_AGEMA_signal_4703, RoundKey[30]}), .b ({new_AGEMA_signal_4697, RoundKey[29]}), .c ({new_AGEMA_signal_4968, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T8_U1 ( .a ({new_AGEMA_signal_4682, RoundKey[24]}), .b ({new_AGEMA_signal_5157, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}), .c ({new_AGEMA_signal_5332, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T9_U1 ( .a ({new_AGEMA_signal_4682, RoundKey[24]}), .b ({new_AGEMA_signal_4968, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_5158, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T10_U1 ( .a ({new_AGEMA_signal_5157, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_4968, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_5333, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T11_U1 ( .a ({new_AGEMA_signal_4703, RoundKey[30]}), .b ({new_AGEMA_signal_4688, RoundKey[26]}), .c ({new_AGEMA_signal_4969, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T12_U1 ( .a ({new_AGEMA_signal_4697, RoundKey[29]}), .b ({new_AGEMA_signal_4688, RoundKey[26]}), .c ({new_AGEMA_signal_4970, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T13_U1 ( .a ({new_AGEMA_signal_4965, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_4966, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4}), .c ({new_AGEMA_signal_5159, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T14_U1 ( .a ({new_AGEMA_signal_5157, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_4969, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_5334, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T15_U1 ( .a ({new_AGEMA_signal_4967, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_4969, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_5160, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T16_U1 ( .a ({new_AGEMA_signal_4967, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_4970, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_5161, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T17_U1 ( .a ({new_AGEMA_signal_5158, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9}), .b ({new_AGEMA_signal_5161, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_5335, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T18_U1 ( .a ({new_AGEMA_signal_4694, RoundKey[28]}), .b ({new_AGEMA_signal_4682, RoundKey[24]}), .c ({new_AGEMA_signal_4971, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T19_U1 ( .a ({new_AGEMA_signal_4968, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_4971, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T18}), .c ({new_AGEMA_signal_5162, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T20_U1 ( .a ({new_AGEMA_signal_4963, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5162, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19}), .c ({new_AGEMA_signal_5336, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T21_U1 ( .a ({new_AGEMA_signal_4685, RoundKey[25]}), .b ({new_AGEMA_signal_4682, RoundKey[24]}), .c ({new_AGEMA_signal_4972, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T22_U1 ( .a ({new_AGEMA_signal_4968, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_4972, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T21}), .c ({new_AGEMA_signal_5163, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T23_U1 ( .a ({new_AGEMA_signal_4964, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_5163, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22}), .c ({new_AGEMA_signal_5337, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T24_U1 ( .a ({new_AGEMA_signal_4964, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_5333, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10}), .c ({new_AGEMA_signal_5580, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T25_U1 ( .a ({new_AGEMA_signal_5336, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_5335, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17}), .c ({new_AGEMA_signal_5581, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T26_U1 ( .a ({new_AGEMA_signal_4965, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_5161, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_5338, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T27_U1 ( .a ({new_AGEMA_signal_4963, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_4970, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_5164, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27}) ) ;
    INV_X1 RoundCounterIns_U14 ( .A (RoundCounterIns_n13), .ZN (RoundCounterIns_n1) ) ;
    MUX2_X1 RoundCounterIns_U13 ( .S (RoundCounterIns_n5), .A (RoundCounterIns_n12), .B (RoundCounterIns_n11), .Z (RoundCounterIns_n13) ) ;
    NOR2_X1 RoundCounterIns_U12 ( .A1 (reset), .A2 (RoundCounterIns_n10), .ZN (RoundCounterIns_N8) ) ;
    XNOR2_X1 RoundCounterIns_U11 ( .A (RoundCounter[0]), .B (RoundCounter[1]), .ZN (RoundCounterIns_n10) ) ;
    MUX2_X1 RoundCounterIns_U10 ( .S (RoundCounter[3]), .A (RoundCounterIns_n9), .B (RoundCounterIns_n8), .Z (RoundCounterIns_N10) ) ;
    NAND2_X1 RoundCounterIns_U9 ( .A1 (RoundCounterIns_n12), .A2 (RoundCounterIns_n7), .ZN (RoundCounterIns_n8) ) ;
    NAND2_X1 RoundCounterIns_U8 ( .A1 (RoundCounterIns_n5), .A2 (RoundCounterIns_n2), .ZN (RoundCounterIns_n7) ) ;
    NOR2_X1 RoundCounterIns_U7 ( .A1 (RoundCounterIns_n4), .A2 (RoundCounterIns_N7), .ZN (RoundCounterIns_n12) ) ;
    NOR2_X1 RoundCounterIns_U6 ( .A1 (RoundCounter[1]), .A2 (reset), .ZN (RoundCounterIns_n4) ) ;
    NOR2_X1 RoundCounterIns_U5 ( .A1 (RoundCounterIns_n5), .A2 (RoundCounterIns_n11), .ZN (RoundCounterIns_n9) ) ;
    NAND2_X1 RoundCounterIns_U4 ( .A1 (RoundCounter[1]), .A2 (RoundCounterIns_n3), .ZN (RoundCounterIns_n11) ) ;
    NOR2_X1 RoundCounterIns_U3 ( .A1 (reset), .A2 (RoundCounterIns_n6), .ZN (RoundCounterIns_n3) ) ;
    NOR2_X1 RoundCounterIns_U2 ( .A1 (reset), .A2 (RoundCounter[0]), .ZN (RoundCounterIns_N7) ) ;
    INV_X1 RoundCounterIns_U1 ( .A (reset), .ZN (RoundCounterIns_n2) ) ;
    INV_X1 RoundCounterIns_count_reg_0__U1 ( .A (RoundCounter[0]), .ZN (RoundCounterIns_n6) ) ;
    INV_X1 RoundCounterIns_count_reg_2__U1 ( .A (RoundCounter[2]), .ZN (RoundCounterIns_n5) ) ;

    /* cells in depth 1 */
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M1_U1 ( .a ({new_AGEMA_signal_5167, SubBytesIns_Inst_Sbox_0_T13}), .b ({new_AGEMA_signal_5165, SubBytesIns_Inst_Sbox_0_T6}), .clk (clk), .r ({Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_5352, SubBytesIns_Inst_Sbox_0_M1}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M2_U1 ( .a ({new_AGEMA_signal_5350, SubBytesIns_Inst_Sbox_0_T23}), .b ({new_AGEMA_signal_5345, SubBytesIns_Inst_Sbox_0_T8}), .clk (clk), .r ({Fresh[3], Fresh[2]}), .c ({new_AGEMA_signal_5591, SubBytesIns_Inst_Sbox_0_M2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M3_U1 ( .a ({new_AGEMA_signal_10062, new_AGEMA_signal_10061}), .b ({new_AGEMA_signal_5352, SubBytesIns_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_5592, SubBytesIns_Inst_Sbox_0_M3}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M4_U1 ( .a ({new_AGEMA_signal_5170, SubBytesIns_Inst_Sbox_0_T19}), .b ({ciphertext_s1[0], ciphertext_s0[0]}), .clk (clk), .r ({Fresh[5], Fresh[4]}), .c ({new_AGEMA_signal_5353, SubBytesIns_Inst_Sbox_0_M4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M5_U1 ( .a ({new_AGEMA_signal_5353, SubBytesIns_Inst_Sbox_0_M4}), .b ({new_AGEMA_signal_5352, SubBytesIns_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_5593, SubBytesIns_Inst_Sbox_0_M5}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M6_U1 ( .a ({new_AGEMA_signal_4975, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_5169, SubBytesIns_Inst_Sbox_0_T16}), .clk (clk), .r ({Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_5354, SubBytesIns_Inst_Sbox_0_M6}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M7_U1 ( .a ({new_AGEMA_signal_5171, SubBytesIns_Inst_Sbox_0_T22}), .b ({new_AGEMA_signal_5166, SubBytesIns_Inst_Sbox_0_T9}), .clk (clk), .r ({Fresh[9], Fresh[8]}), .c ({new_AGEMA_signal_5355, SubBytesIns_Inst_Sbox_0_M7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M8_U1 ( .a ({new_AGEMA_signal_10064, new_AGEMA_signal_10063}), .b ({new_AGEMA_signal_5354, SubBytesIns_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_5594, SubBytesIns_Inst_Sbox_0_M8}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M9_U1 ( .a ({new_AGEMA_signal_5349, SubBytesIns_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_5348, SubBytesIns_Inst_Sbox_0_T17}), .clk (clk), .r ({Fresh[11], Fresh[10]}), .c ({new_AGEMA_signal_5595, SubBytesIns_Inst_Sbox_0_M9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M10_U1 ( .a ({new_AGEMA_signal_5595, SubBytesIns_Inst_Sbox_0_M9}), .b ({new_AGEMA_signal_5354, SubBytesIns_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_5753, SubBytesIns_Inst_Sbox_0_M10}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M11_U1 ( .a ({new_AGEMA_signal_4973, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_5168, SubBytesIns_Inst_Sbox_0_T15}), .clk (clk), .r ({Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_5356, SubBytesIns_Inst_Sbox_0_M11}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M12_U1 ( .a ({new_AGEMA_signal_4976, SubBytesIns_Inst_Sbox_0_T4}), .b ({new_AGEMA_signal_5172, SubBytesIns_Inst_Sbox_0_T27}), .clk (clk), .r ({Fresh[15], Fresh[14]}), .c ({new_AGEMA_signal_5357, SubBytesIns_Inst_Sbox_0_M12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M13_U1 ( .a ({new_AGEMA_signal_5357, SubBytesIns_Inst_Sbox_0_M12}), .b ({new_AGEMA_signal_5356, SubBytesIns_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_5596, SubBytesIns_Inst_Sbox_0_M13}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M14_U1 ( .a ({new_AGEMA_signal_4974, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_5346, SubBytesIns_Inst_Sbox_0_T10}), .clk (clk), .r ({Fresh[17], Fresh[16]}), .c ({new_AGEMA_signal_5597, SubBytesIns_Inst_Sbox_0_M14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M15_U1 ( .a ({new_AGEMA_signal_5597, SubBytesIns_Inst_Sbox_0_M14}), .b ({new_AGEMA_signal_5356, SubBytesIns_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_5754, SubBytesIns_Inst_Sbox_0_M15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M16_U1 ( .a ({new_AGEMA_signal_5592, SubBytesIns_Inst_Sbox_0_M3}), .b ({new_AGEMA_signal_5591, SubBytesIns_Inst_Sbox_0_M2}), .c ({new_AGEMA_signal_5755, SubBytesIns_Inst_Sbox_0_M16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M17_U1 ( .a ({new_AGEMA_signal_5593, SubBytesIns_Inst_Sbox_0_M5}), .b ({new_AGEMA_signal_10066, new_AGEMA_signal_10065}), .c ({new_AGEMA_signal_5756, SubBytesIns_Inst_Sbox_0_M17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M18_U1 ( .a ({new_AGEMA_signal_5594, SubBytesIns_Inst_Sbox_0_M8}), .b ({new_AGEMA_signal_5355, SubBytesIns_Inst_Sbox_0_M7}), .c ({new_AGEMA_signal_5757, SubBytesIns_Inst_Sbox_0_M18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M19_U1 ( .a ({new_AGEMA_signal_5753, SubBytesIns_Inst_Sbox_0_M10}), .b ({new_AGEMA_signal_5754, SubBytesIns_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_5849, SubBytesIns_Inst_Sbox_0_M19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M20_U1 ( .a ({new_AGEMA_signal_5755, SubBytesIns_Inst_Sbox_0_M16}), .b ({new_AGEMA_signal_5596, SubBytesIns_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_5850, SubBytesIns_Inst_Sbox_0_M20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M21_U1 ( .a ({new_AGEMA_signal_5756, SubBytesIns_Inst_Sbox_0_M17}), .b ({new_AGEMA_signal_5754, SubBytesIns_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_5851, SubBytesIns_Inst_Sbox_0_M21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M22_U1 ( .a ({new_AGEMA_signal_5757, SubBytesIns_Inst_Sbox_0_M18}), .b ({new_AGEMA_signal_5596, SubBytesIns_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_5852, SubBytesIns_Inst_Sbox_0_M22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M23_U1 ( .a ({new_AGEMA_signal_5849, SubBytesIns_Inst_Sbox_0_M19}), .b ({new_AGEMA_signal_10068, new_AGEMA_signal_10067}), .c ({new_AGEMA_signal_5929, SubBytesIns_Inst_Sbox_0_M23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M24_U1 ( .a ({new_AGEMA_signal_5852, SubBytesIns_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_5929, SubBytesIns_Inst_Sbox_0_M23}), .c ({new_AGEMA_signal_6013, SubBytesIns_Inst_Sbox_0_M24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M27_U1 ( .a ({new_AGEMA_signal_5850, SubBytesIns_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_5851, SubBytesIns_Inst_Sbox_0_M21}), .c ({new_AGEMA_signal_5931, SubBytesIns_Inst_Sbox_0_M27}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M1_U1 ( .a ({new_AGEMA_signal_5175, SubBytesIns_Inst_Sbox_1_T13}), .b ({new_AGEMA_signal_5173, SubBytesIns_Inst_Sbox_1_T6}), .clk (clk), .r ({Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_5365, SubBytesIns_Inst_Sbox_1_M1}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M2_U1 ( .a ({new_AGEMA_signal_5363, SubBytesIns_Inst_Sbox_1_T23}), .b ({new_AGEMA_signal_5358, SubBytesIns_Inst_Sbox_1_T8}), .clk (clk), .r ({Fresh[21], Fresh[20]}), .c ({new_AGEMA_signal_5600, SubBytesIns_Inst_Sbox_1_M2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M3_U1 ( .a ({new_AGEMA_signal_10070, new_AGEMA_signal_10069}), .b ({new_AGEMA_signal_5365, SubBytesIns_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_5601, SubBytesIns_Inst_Sbox_1_M3}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M4_U1 ( .a ({new_AGEMA_signal_5178, SubBytesIns_Inst_Sbox_1_T19}), .b ({ciphertext_s1[8], ciphertext_s0[8]}), .clk (clk), .r ({Fresh[23], Fresh[22]}), .c ({new_AGEMA_signal_5366, SubBytesIns_Inst_Sbox_1_M4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M5_U1 ( .a ({new_AGEMA_signal_5366, SubBytesIns_Inst_Sbox_1_M4}), .b ({new_AGEMA_signal_5365, SubBytesIns_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_5602, SubBytesIns_Inst_Sbox_1_M5}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M6_U1 ( .a ({new_AGEMA_signal_4985, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_5177, SubBytesIns_Inst_Sbox_1_T16}), .clk (clk), .r ({Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_5367, SubBytesIns_Inst_Sbox_1_M6}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M7_U1 ( .a ({new_AGEMA_signal_5179, SubBytesIns_Inst_Sbox_1_T22}), .b ({new_AGEMA_signal_5174, SubBytesIns_Inst_Sbox_1_T9}), .clk (clk), .r ({Fresh[27], Fresh[26]}), .c ({new_AGEMA_signal_5368, SubBytesIns_Inst_Sbox_1_M7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M8_U1 ( .a ({new_AGEMA_signal_10072, new_AGEMA_signal_10071}), .b ({new_AGEMA_signal_5367, SubBytesIns_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_5603, SubBytesIns_Inst_Sbox_1_M8}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M9_U1 ( .a ({new_AGEMA_signal_5362, SubBytesIns_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_5361, SubBytesIns_Inst_Sbox_1_T17}), .clk (clk), .r ({Fresh[29], Fresh[28]}), .c ({new_AGEMA_signal_5604, SubBytesIns_Inst_Sbox_1_M9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M10_U1 ( .a ({new_AGEMA_signal_5604, SubBytesIns_Inst_Sbox_1_M9}), .b ({new_AGEMA_signal_5367, SubBytesIns_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_5758, SubBytesIns_Inst_Sbox_1_M10}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M11_U1 ( .a ({new_AGEMA_signal_4983, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_5176, SubBytesIns_Inst_Sbox_1_T15}), .clk (clk), .r ({Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_5369, SubBytesIns_Inst_Sbox_1_M11}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M12_U1 ( .a ({new_AGEMA_signal_4986, SubBytesIns_Inst_Sbox_1_T4}), .b ({new_AGEMA_signal_5180, SubBytesIns_Inst_Sbox_1_T27}), .clk (clk), .r ({Fresh[33], Fresh[32]}), .c ({new_AGEMA_signal_5370, SubBytesIns_Inst_Sbox_1_M12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M13_U1 ( .a ({new_AGEMA_signal_5370, SubBytesIns_Inst_Sbox_1_M12}), .b ({new_AGEMA_signal_5369, SubBytesIns_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_5605, SubBytesIns_Inst_Sbox_1_M13}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M14_U1 ( .a ({new_AGEMA_signal_4984, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_5359, SubBytesIns_Inst_Sbox_1_T10}), .clk (clk), .r ({Fresh[35], Fresh[34]}), .c ({new_AGEMA_signal_5606, SubBytesIns_Inst_Sbox_1_M14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M15_U1 ( .a ({new_AGEMA_signal_5606, SubBytesIns_Inst_Sbox_1_M14}), .b ({new_AGEMA_signal_5369, SubBytesIns_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_5759, SubBytesIns_Inst_Sbox_1_M15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M16_U1 ( .a ({new_AGEMA_signal_5601, SubBytesIns_Inst_Sbox_1_M3}), .b ({new_AGEMA_signal_5600, SubBytesIns_Inst_Sbox_1_M2}), .c ({new_AGEMA_signal_5760, SubBytesIns_Inst_Sbox_1_M16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M17_U1 ( .a ({new_AGEMA_signal_5602, SubBytesIns_Inst_Sbox_1_M5}), .b ({new_AGEMA_signal_10074, new_AGEMA_signal_10073}), .c ({new_AGEMA_signal_5761, SubBytesIns_Inst_Sbox_1_M17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M18_U1 ( .a ({new_AGEMA_signal_5603, SubBytesIns_Inst_Sbox_1_M8}), .b ({new_AGEMA_signal_5368, SubBytesIns_Inst_Sbox_1_M7}), .c ({new_AGEMA_signal_5762, SubBytesIns_Inst_Sbox_1_M18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M19_U1 ( .a ({new_AGEMA_signal_5758, SubBytesIns_Inst_Sbox_1_M10}), .b ({new_AGEMA_signal_5759, SubBytesIns_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_5853, SubBytesIns_Inst_Sbox_1_M19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M20_U1 ( .a ({new_AGEMA_signal_5760, SubBytesIns_Inst_Sbox_1_M16}), .b ({new_AGEMA_signal_5605, SubBytesIns_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_5854, SubBytesIns_Inst_Sbox_1_M20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M21_U1 ( .a ({new_AGEMA_signal_5761, SubBytesIns_Inst_Sbox_1_M17}), .b ({new_AGEMA_signal_5759, SubBytesIns_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_5855, SubBytesIns_Inst_Sbox_1_M21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M22_U1 ( .a ({new_AGEMA_signal_5762, SubBytesIns_Inst_Sbox_1_M18}), .b ({new_AGEMA_signal_5605, SubBytesIns_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_5856, SubBytesIns_Inst_Sbox_1_M22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M23_U1 ( .a ({new_AGEMA_signal_5853, SubBytesIns_Inst_Sbox_1_M19}), .b ({new_AGEMA_signal_10076, new_AGEMA_signal_10075}), .c ({new_AGEMA_signal_5933, SubBytesIns_Inst_Sbox_1_M23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M24_U1 ( .a ({new_AGEMA_signal_5856, SubBytesIns_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_5933, SubBytesIns_Inst_Sbox_1_M23}), .c ({new_AGEMA_signal_6018, SubBytesIns_Inst_Sbox_1_M24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M27_U1 ( .a ({new_AGEMA_signal_5854, SubBytesIns_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_5855, SubBytesIns_Inst_Sbox_1_M21}), .c ({new_AGEMA_signal_5935, SubBytesIns_Inst_Sbox_1_M27}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M1_U1 ( .a ({new_AGEMA_signal_5183, SubBytesIns_Inst_Sbox_2_T13}), .b ({new_AGEMA_signal_5181, SubBytesIns_Inst_Sbox_2_T6}), .clk (clk), .r ({Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_5378, SubBytesIns_Inst_Sbox_2_M1}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M2_U1 ( .a ({new_AGEMA_signal_5376, SubBytesIns_Inst_Sbox_2_T23}), .b ({new_AGEMA_signal_5371, SubBytesIns_Inst_Sbox_2_T8}), .clk (clk), .r ({Fresh[39], Fresh[38]}), .c ({new_AGEMA_signal_5609, SubBytesIns_Inst_Sbox_2_M2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M3_U1 ( .a ({new_AGEMA_signal_10078, new_AGEMA_signal_10077}), .b ({new_AGEMA_signal_5378, SubBytesIns_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_5610, SubBytesIns_Inst_Sbox_2_M3}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M4_U1 ( .a ({new_AGEMA_signal_5186, SubBytesIns_Inst_Sbox_2_T19}), .b ({ciphertext_s1[16], ciphertext_s0[16]}), .clk (clk), .r ({Fresh[41], Fresh[40]}), .c ({new_AGEMA_signal_5379, SubBytesIns_Inst_Sbox_2_M4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M5_U1 ( .a ({new_AGEMA_signal_5379, SubBytesIns_Inst_Sbox_2_M4}), .b ({new_AGEMA_signal_5378, SubBytesIns_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_5611, SubBytesIns_Inst_Sbox_2_M5}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M6_U1 ( .a ({new_AGEMA_signal_4995, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_5185, SubBytesIns_Inst_Sbox_2_T16}), .clk (clk), .r ({Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_5380, SubBytesIns_Inst_Sbox_2_M6}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M7_U1 ( .a ({new_AGEMA_signal_5187, SubBytesIns_Inst_Sbox_2_T22}), .b ({new_AGEMA_signal_5182, SubBytesIns_Inst_Sbox_2_T9}), .clk (clk), .r ({Fresh[45], Fresh[44]}), .c ({new_AGEMA_signal_5381, SubBytesIns_Inst_Sbox_2_M7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M8_U1 ( .a ({new_AGEMA_signal_10080, new_AGEMA_signal_10079}), .b ({new_AGEMA_signal_5380, SubBytesIns_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_5612, SubBytesIns_Inst_Sbox_2_M8}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M9_U1 ( .a ({new_AGEMA_signal_5375, SubBytesIns_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_5374, SubBytesIns_Inst_Sbox_2_T17}), .clk (clk), .r ({Fresh[47], Fresh[46]}), .c ({new_AGEMA_signal_5613, SubBytesIns_Inst_Sbox_2_M9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M10_U1 ( .a ({new_AGEMA_signal_5613, SubBytesIns_Inst_Sbox_2_M9}), .b ({new_AGEMA_signal_5380, SubBytesIns_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_5763, SubBytesIns_Inst_Sbox_2_M10}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M11_U1 ( .a ({new_AGEMA_signal_4993, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5184, SubBytesIns_Inst_Sbox_2_T15}), .clk (clk), .r ({Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_5382, SubBytesIns_Inst_Sbox_2_M11}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M12_U1 ( .a ({new_AGEMA_signal_4996, SubBytesIns_Inst_Sbox_2_T4}), .b ({new_AGEMA_signal_5188, SubBytesIns_Inst_Sbox_2_T27}), .clk (clk), .r ({Fresh[51], Fresh[50]}), .c ({new_AGEMA_signal_5383, SubBytesIns_Inst_Sbox_2_M12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M13_U1 ( .a ({new_AGEMA_signal_5383, SubBytesIns_Inst_Sbox_2_M12}), .b ({new_AGEMA_signal_5382, SubBytesIns_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_5614, SubBytesIns_Inst_Sbox_2_M13}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M14_U1 ( .a ({new_AGEMA_signal_4994, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_5372, SubBytesIns_Inst_Sbox_2_T10}), .clk (clk), .r ({Fresh[53], Fresh[52]}), .c ({new_AGEMA_signal_5615, SubBytesIns_Inst_Sbox_2_M14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M15_U1 ( .a ({new_AGEMA_signal_5615, SubBytesIns_Inst_Sbox_2_M14}), .b ({new_AGEMA_signal_5382, SubBytesIns_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_5764, SubBytesIns_Inst_Sbox_2_M15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M16_U1 ( .a ({new_AGEMA_signal_5610, SubBytesIns_Inst_Sbox_2_M3}), .b ({new_AGEMA_signal_5609, SubBytesIns_Inst_Sbox_2_M2}), .c ({new_AGEMA_signal_5765, SubBytesIns_Inst_Sbox_2_M16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M17_U1 ( .a ({new_AGEMA_signal_5611, SubBytesIns_Inst_Sbox_2_M5}), .b ({new_AGEMA_signal_10082, new_AGEMA_signal_10081}), .c ({new_AGEMA_signal_5766, SubBytesIns_Inst_Sbox_2_M17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M18_U1 ( .a ({new_AGEMA_signal_5612, SubBytesIns_Inst_Sbox_2_M8}), .b ({new_AGEMA_signal_5381, SubBytesIns_Inst_Sbox_2_M7}), .c ({new_AGEMA_signal_5767, SubBytesIns_Inst_Sbox_2_M18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M19_U1 ( .a ({new_AGEMA_signal_5763, SubBytesIns_Inst_Sbox_2_M10}), .b ({new_AGEMA_signal_5764, SubBytesIns_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_5857, SubBytesIns_Inst_Sbox_2_M19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M20_U1 ( .a ({new_AGEMA_signal_5765, SubBytesIns_Inst_Sbox_2_M16}), .b ({new_AGEMA_signal_5614, SubBytesIns_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_5858, SubBytesIns_Inst_Sbox_2_M20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M21_U1 ( .a ({new_AGEMA_signal_5766, SubBytesIns_Inst_Sbox_2_M17}), .b ({new_AGEMA_signal_5764, SubBytesIns_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_5859, SubBytesIns_Inst_Sbox_2_M21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M22_U1 ( .a ({new_AGEMA_signal_5767, SubBytesIns_Inst_Sbox_2_M18}), .b ({new_AGEMA_signal_5614, SubBytesIns_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_5860, SubBytesIns_Inst_Sbox_2_M22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M23_U1 ( .a ({new_AGEMA_signal_5857, SubBytesIns_Inst_Sbox_2_M19}), .b ({new_AGEMA_signal_10084, new_AGEMA_signal_10083}), .c ({new_AGEMA_signal_5937, SubBytesIns_Inst_Sbox_2_M23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M24_U1 ( .a ({new_AGEMA_signal_5860, SubBytesIns_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_5937, SubBytesIns_Inst_Sbox_2_M23}), .c ({new_AGEMA_signal_6023, SubBytesIns_Inst_Sbox_2_M24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M27_U1 ( .a ({new_AGEMA_signal_5858, SubBytesIns_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_5859, SubBytesIns_Inst_Sbox_2_M21}), .c ({new_AGEMA_signal_5939, SubBytesIns_Inst_Sbox_2_M27}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M1_U1 ( .a ({new_AGEMA_signal_5191, SubBytesIns_Inst_Sbox_3_T13}), .b ({new_AGEMA_signal_5189, SubBytesIns_Inst_Sbox_3_T6}), .clk (clk), .r ({Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_5391, SubBytesIns_Inst_Sbox_3_M1}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M2_U1 ( .a ({new_AGEMA_signal_5389, SubBytesIns_Inst_Sbox_3_T23}), .b ({new_AGEMA_signal_5384, SubBytesIns_Inst_Sbox_3_T8}), .clk (clk), .r ({Fresh[57], Fresh[56]}), .c ({new_AGEMA_signal_5618, SubBytesIns_Inst_Sbox_3_M2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M3_U1 ( .a ({new_AGEMA_signal_10086, new_AGEMA_signal_10085}), .b ({new_AGEMA_signal_5391, SubBytesIns_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_5619, SubBytesIns_Inst_Sbox_3_M3}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M4_U1 ( .a ({new_AGEMA_signal_5194, SubBytesIns_Inst_Sbox_3_T19}), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .clk (clk), .r ({Fresh[59], Fresh[58]}), .c ({new_AGEMA_signal_5392, SubBytesIns_Inst_Sbox_3_M4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M5_U1 ( .a ({new_AGEMA_signal_5392, SubBytesIns_Inst_Sbox_3_M4}), .b ({new_AGEMA_signal_5391, SubBytesIns_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_5620, SubBytesIns_Inst_Sbox_3_M5}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M6_U1 ( .a ({new_AGEMA_signal_5005, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_5193, SubBytesIns_Inst_Sbox_3_T16}), .clk (clk), .r ({Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_5393, SubBytesIns_Inst_Sbox_3_M6}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M7_U1 ( .a ({new_AGEMA_signal_5195, SubBytesIns_Inst_Sbox_3_T22}), .b ({new_AGEMA_signal_5190, SubBytesIns_Inst_Sbox_3_T9}), .clk (clk), .r ({Fresh[63], Fresh[62]}), .c ({new_AGEMA_signal_5394, SubBytesIns_Inst_Sbox_3_M7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M8_U1 ( .a ({new_AGEMA_signal_10088, new_AGEMA_signal_10087}), .b ({new_AGEMA_signal_5393, SubBytesIns_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_5621, SubBytesIns_Inst_Sbox_3_M8}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M9_U1 ( .a ({new_AGEMA_signal_5388, SubBytesIns_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_5387, SubBytesIns_Inst_Sbox_3_T17}), .clk (clk), .r ({Fresh[65], Fresh[64]}), .c ({new_AGEMA_signal_5622, SubBytesIns_Inst_Sbox_3_M9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M10_U1 ( .a ({new_AGEMA_signal_5622, SubBytesIns_Inst_Sbox_3_M9}), .b ({new_AGEMA_signal_5393, SubBytesIns_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_5768, SubBytesIns_Inst_Sbox_3_M10}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M11_U1 ( .a ({new_AGEMA_signal_5003, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5192, SubBytesIns_Inst_Sbox_3_T15}), .clk (clk), .r ({Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_5395, SubBytesIns_Inst_Sbox_3_M11}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M12_U1 ( .a ({new_AGEMA_signal_5006, SubBytesIns_Inst_Sbox_3_T4}), .b ({new_AGEMA_signal_5196, SubBytesIns_Inst_Sbox_3_T27}), .clk (clk), .r ({Fresh[69], Fresh[68]}), .c ({new_AGEMA_signal_5396, SubBytesIns_Inst_Sbox_3_M12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M13_U1 ( .a ({new_AGEMA_signal_5396, SubBytesIns_Inst_Sbox_3_M12}), .b ({new_AGEMA_signal_5395, SubBytesIns_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_5623, SubBytesIns_Inst_Sbox_3_M13}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M14_U1 ( .a ({new_AGEMA_signal_5004, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_5385, SubBytesIns_Inst_Sbox_3_T10}), .clk (clk), .r ({Fresh[71], Fresh[70]}), .c ({new_AGEMA_signal_5624, SubBytesIns_Inst_Sbox_3_M14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M15_U1 ( .a ({new_AGEMA_signal_5624, SubBytesIns_Inst_Sbox_3_M14}), .b ({new_AGEMA_signal_5395, SubBytesIns_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_5769, SubBytesIns_Inst_Sbox_3_M15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M16_U1 ( .a ({new_AGEMA_signal_5619, SubBytesIns_Inst_Sbox_3_M3}), .b ({new_AGEMA_signal_5618, SubBytesIns_Inst_Sbox_3_M2}), .c ({new_AGEMA_signal_5770, SubBytesIns_Inst_Sbox_3_M16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M17_U1 ( .a ({new_AGEMA_signal_5620, SubBytesIns_Inst_Sbox_3_M5}), .b ({new_AGEMA_signal_10090, new_AGEMA_signal_10089}), .c ({new_AGEMA_signal_5771, SubBytesIns_Inst_Sbox_3_M17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M18_U1 ( .a ({new_AGEMA_signal_5621, SubBytesIns_Inst_Sbox_3_M8}), .b ({new_AGEMA_signal_5394, SubBytesIns_Inst_Sbox_3_M7}), .c ({new_AGEMA_signal_5772, SubBytesIns_Inst_Sbox_3_M18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M19_U1 ( .a ({new_AGEMA_signal_5768, SubBytesIns_Inst_Sbox_3_M10}), .b ({new_AGEMA_signal_5769, SubBytesIns_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_5861, SubBytesIns_Inst_Sbox_3_M19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M20_U1 ( .a ({new_AGEMA_signal_5770, SubBytesIns_Inst_Sbox_3_M16}), .b ({new_AGEMA_signal_5623, SubBytesIns_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_5862, SubBytesIns_Inst_Sbox_3_M20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M21_U1 ( .a ({new_AGEMA_signal_5771, SubBytesIns_Inst_Sbox_3_M17}), .b ({new_AGEMA_signal_5769, SubBytesIns_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_5863, SubBytesIns_Inst_Sbox_3_M21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M22_U1 ( .a ({new_AGEMA_signal_5772, SubBytesIns_Inst_Sbox_3_M18}), .b ({new_AGEMA_signal_5623, SubBytesIns_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_5864, SubBytesIns_Inst_Sbox_3_M22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M23_U1 ( .a ({new_AGEMA_signal_5861, SubBytesIns_Inst_Sbox_3_M19}), .b ({new_AGEMA_signal_10092, new_AGEMA_signal_10091}), .c ({new_AGEMA_signal_5941, SubBytesIns_Inst_Sbox_3_M23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M24_U1 ( .a ({new_AGEMA_signal_5864, SubBytesIns_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_5941, SubBytesIns_Inst_Sbox_3_M23}), .c ({new_AGEMA_signal_6028, SubBytesIns_Inst_Sbox_3_M24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M27_U1 ( .a ({new_AGEMA_signal_5862, SubBytesIns_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_5863, SubBytesIns_Inst_Sbox_3_M21}), .c ({new_AGEMA_signal_5943, SubBytesIns_Inst_Sbox_3_M27}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M1_U1 ( .a ({new_AGEMA_signal_5199, SubBytesIns_Inst_Sbox_4_T13}), .b ({new_AGEMA_signal_5197, SubBytesIns_Inst_Sbox_4_T6}), .clk (clk), .r ({Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_5404, SubBytesIns_Inst_Sbox_4_M1}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M2_U1 ( .a ({new_AGEMA_signal_5402, SubBytesIns_Inst_Sbox_4_T23}), .b ({new_AGEMA_signal_5397, SubBytesIns_Inst_Sbox_4_T8}), .clk (clk), .r ({Fresh[75], Fresh[74]}), .c ({new_AGEMA_signal_5627, SubBytesIns_Inst_Sbox_4_M2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M3_U1 ( .a ({new_AGEMA_signal_10094, new_AGEMA_signal_10093}), .b ({new_AGEMA_signal_5404, SubBytesIns_Inst_Sbox_4_M1}), .c ({new_AGEMA_signal_5628, SubBytesIns_Inst_Sbox_4_M3}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M4_U1 ( .a ({new_AGEMA_signal_5202, SubBytesIns_Inst_Sbox_4_T19}), .b ({ciphertext_s1[32], ciphertext_s0[32]}), .clk (clk), .r ({Fresh[77], Fresh[76]}), .c ({new_AGEMA_signal_5405, SubBytesIns_Inst_Sbox_4_M4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M5_U1 ( .a ({new_AGEMA_signal_5405, SubBytesIns_Inst_Sbox_4_M4}), .b ({new_AGEMA_signal_5404, SubBytesIns_Inst_Sbox_4_M1}), .c ({new_AGEMA_signal_5629, SubBytesIns_Inst_Sbox_4_M5}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M6_U1 ( .a ({new_AGEMA_signal_5015, SubBytesIns_Inst_Sbox_4_T3}), .b ({new_AGEMA_signal_5201, SubBytesIns_Inst_Sbox_4_T16}), .clk (clk), .r ({Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_5406, SubBytesIns_Inst_Sbox_4_M6}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M7_U1 ( .a ({new_AGEMA_signal_5203, SubBytesIns_Inst_Sbox_4_T22}), .b ({new_AGEMA_signal_5198, SubBytesIns_Inst_Sbox_4_T9}), .clk (clk), .r ({Fresh[81], Fresh[80]}), .c ({new_AGEMA_signal_5407, SubBytesIns_Inst_Sbox_4_M7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M8_U1 ( .a ({new_AGEMA_signal_10096, new_AGEMA_signal_10095}), .b ({new_AGEMA_signal_5406, SubBytesIns_Inst_Sbox_4_M6}), .c ({new_AGEMA_signal_5630, SubBytesIns_Inst_Sbox_4_M8}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M9_U1 ( .a ({new_AGEMA_signal_5401, SubBytesIns_Inst_Sbox_4_T20}), .b ({new_AGEMA_signal_5400, SubBytesIns_Inst_Sbox_4_T17}), .clk (clk), .r ({Fresh[83], Fresh[82]}), .c ({new_AGEMA_signal_5631, SubBytesIns_Inst_Sbox_4_M9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M10_U1 ( .a ({new_AGEMA_signal_5631, SubBytesIns_Inst_Sbox_4_M9}), .b ({new_AGEMA_signal_5406, SubBytesIns_Inst_Sbox_4_M6}), .c ({new_AGEMA_signal_5773, SubBytesIns_Inst_Sbox_4_M10}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M11_U1 ( .a ({new_AGEMA_signal_5013, SubBytesIns_Inst_Sbox_4_T1}), .b ({new_AGEMA_signal_5200, SubBytesIns_Inst_Sbox_4_T15}), .clk (clk), .r ({Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_5408, SubBytesIns_Inst_Sbox_4_M11}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M12_U1 ( .a ({new_AGEMA_signal_5016, SubBytesIns_Inst_Sbox_4_T4}), .b ({new_AGEMA_signal_5204, SubBytesIns_Inst_Sbox_4_T27}), .clk (clk), .r ({Fresh[87], Fresh[86]}), .c ({new_AGEMA_signal_5409, SubBytesIns_Inst_Sbox_4_M12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M13_U1 ( .a ({new_AGEMA_signal_5409, SubBytesIns_Inst_Sbox_4_M12}), .b ({new_AGEMA_signal_5408, SubBytesIns_Inst_Sbox_4_M11}), .c ({new_AGEMA_signal_5632, SubBytesIns_Inst_Sbox_4_M13}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M14_U1 ( .a ({new_AGEMA_signal_5014, SubBytesIns_Inst_Sbox_4_T2}), .b ({new_AGEMA_signal_5398, SubBytesIns_Inst_Sbox_4_T10}), .clk (clk), .r ({Fresh[89], Fresh[88]}), .c ({new_AGEMA_signal_5633, SubBytesIns_Inst_Sbox_4_M14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M15_U1 ( .a ({new_AGEMA_signal_5633, SubBytesIns_Inst_Sbox_4_M14}), .b ({new_AGEMA_signal_5408, SubBytesIns_Inst_Sbox_4_M11}), .c ({new_AGEMA_signal_5774, SubBytesIns_Inst_Sbox_4_M15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M16_U1 ( .a ({new_AGEMA_signal_5628, SubBytesIns_Inst_Sbox_4_M3}), .b ({new_AGEMA_signal_5627, SubBytesIns_Inst_Sbox_4_M2}), .c ({new_AGEMA_signal_5775, SubBytesIns_Inst_Sbox_4_M16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M17_U1 ( .a ({new_AGEMA_signal_5629, SubBytesIns_Inst_Sbox_4_M5}), .b ({new_AGEMA_signal_10098, new_AGEMA_signal_10097}), .c ({new_AGEMA_signal_5776, SubBytesIns_Inst_Sbox_4_M17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M18_U1 ( .a ({new_AGEMA_signal_5630, SubBytesIns_Inst_Sbox_4_M8}), .b ({new_AGEMA_signal_5407, SubBytesIns_Inst_Sbox_4_M7}), .c ({new_AGEMA_signal_5777, SubBytesIns_Inst_Sbox_4_M18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M19_U1 ( .a ({new_AGEMA_signal_5773, SubBytesIns_Inst_Sbox_4_M10}), .b ({new_AGEMA_signal_5774, SubBytesIns_Inst_Sbox_4_M15}), .c ({new_AGEMA_signal_5865, SubBytesIns_Inst_Sbox_4_M19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M20_U1 ( .a ({new_AGEMA_signal_5775, SubBytesIns_Inst_Sbox_4_M16}), .b ({new_AGEMA_signal_5632, SubBytesIns_Inst_Sbox_4_M13}), .c ({new_AGEMA_signal_5866, SubBytesIns_Inst_Sbox_4_M20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M21_U1 ( .a ({new_AGEMA_signal_5776, SubBytesIns_Inst_Sbox_4_M17}), .b ({new_AGEMA_signal_5774, SubBytesIns_Inst_Sbox_4_M15}), .c ({new_AGEMA_signal_5867, SubBytesIns_Inst_Sbox_4_M21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M22_U1 ( .a ({new_AGEMA_signal_5777, SubBytesIns_Inst_Sbox_4_M18}), .b ({new_AGEMA_signal_5632, SubBytesIns_Inst_Sbox_4_M13}), .c ({new_AGEMA_signal_5868, SubBytesIns_Inst_Sbox_4_M22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M23_U1 ( .a ({new_AGEMA_signal_5865, SubBytesIns_Inst_Sbox_4_M19}), .b ({new_AGEMA_signal_10100, new_AGEMA_signal_10099}), .c ({new_AGEMA_signal_5945, SubBytesIns_Inst_Sbox_4_M23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M24_U1 ( .a ({new_AGEMA_signal_5868, SubBytesIns_Inst_Sbox_4_M22}), .b ({new_AGEMA_signal_5945, SubBytesIns_Inst_Sbox_4_M23}), .c ({new_AGEMA_signal_6033, SubBytesIns_Inst_Sbox_4_M24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M27_U1 ( .a ({new_AGEMA_signal_5866, SubBytesIns_Inst_Sbox_4_M20}), .b ({new_AGEMA_signal_5867, SubBytesIns_Inst_Sbox_4_M21}), .c ({new_AGEMA_signal_5947, SubBytesIns_Inst_Sbox_4_M27}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M1_U1 ( .a ({new_AGEMA_signal_5207, SubBytesIns_Inst_Sbox_5_T13}), .b ({new_AGEMA_signal_5205, SubBytesIns_Inst_Sbox_5_T6}), .clk (clk), .r ({Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_5417, SubBytesIns_Inst_Sbox_5_M1}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M2_U1 ( .a ({new_AGEMA_signal_5415, SubBytesIns_Inst_Sbox_5_T23}), .b ({new_AGEMA_signal_5410, SubBytesIns_Inst_Sbox_5_T8}), .clk (clk), .r ({Fresh[93], Fresh[92]}), .c ({new_AGEMA_signal_5636, SubBytesIns_Inst_Sbox_5_M2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M3_U1 ( .a ({new_AGEMA_signal_10102, new_AGEMA_signal_10101}), .b ({new_AGEMA_signal_5417, SubBytesIns_Inst_Sbox_5_M1}), .c ({new_AGEMA_signal_5637, SubBytesIns_Inst_Sbox_5_M3}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M4_U1 ( .a ({new_AGEMA_signal_5210, SubBytesIns_Inst_Sbox_5_T19}), .b ({ciphertext_s1[40], ciphertext_s0[40]}), .clk (clk), .r ({Fresh[95], Fresh[94]}), .c ({new_AGEMA_signal_5418, SubBytesIns_Inst_Sbox_5_M4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M5_U1 ( .a ({new_AGEMA_signal_5418, SubBytesIns_Inst_Sbox_5_M4}), .b ({new_AGEMA_signal_5417, SubBytesIns_Inst_Sbox_5_M1}), .c ({new_AGEMA_signal_5638, SubBytesIns_Inst_Sbox_5_M5}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M6_U1 ( .a ({new_AGEMA_signal_5025, SubBytesIns_Inst_Sbox_5_T3}), .b ({new_AGEMA_signal_5209, SubBytesIns_Inst_Sbox_5_T16}), .clk (clk), .r ({Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_5419, SubBytesIns_Inst_Sbox_5_M6}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M7_U1 ( .a ({new_AGEMA_signal_5211, SubBytesIns_Inst_Sbox_5_T22}), .b ({new_AGEMA_signal_5206, SubBytesIns_Inst_Sbox_5_T9}), .clk (clk), .r ({Fresh[99], Fresh[98]}), .c ({new_AGEMA_signal_5420, SubBytesIns_Inst_Sbox_5_M7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M8_U1 ( .a ({new_AGEMA_signal_10104, new_AGEMA_signal_10103}), .b ({new_AGEMA_signal_5419, SubBytesIns_Inst_Sbox_5_M6}), .c ({new_AGEMA_signal_5639, SubBytesIns_Inst_Sbox_5_M8}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M9_U1 ( .a ({new_AGEMA_signal_5414, SubBytesIns_Inst_Sbox_5_T20}), .b ({new_AGEMA_signal_5413, SubBytesIns_Inst_Sbox_5_T17}), .clk (clk), .r ({Fresh[101], Fresh[100]}), .c ({new_AGEMA_signal_5640, SubBytesIns_Inst_Sbox_5_M9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M10_U1 ( .a ({new_AGEMA_signal_5640, SubBytesIns_Inst_Sbox_5_M9}), .b ({new_AGEMA_signal_5419, SubBytesIns_Inst_Sbox_5_M6}), .c ({new_AGEMA_signal_5778, SubBytesIns_Inst_Sbox_5_M10}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M11_U1 ( .a ({new_AGEMA_signal_5023, SubBytesIns_Inst_Sbox_5_T1}), .b ({new_AGEMA_signal_5208, SubBytesIns_Inst_Sbox_5_T15}), .clk (clk), .r ({Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_5421, SubBytesIns_Inst_Sbox_5_M11}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M12_U1 ( .a ({new_AGEMA_signal_5026, SubBytesIns_Inst_Sbox_5_T4}), .b ({new_AGEMA_signal_5212, SubBytesIns_Inst_Sbox_5_T27}), .clk (clk), .r ({Fresh[105], Fresh[104]}), .c ({new_AGEMA_signal_5422, SubBytesIns_Inst_Sbox_5_M12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M13_U1 ( .a ({new_AGEMA_signal_5422, SubBytesIns_Inst_Sbox_5_M12}), .b ({new_AGEMA_signal_5421, SubBytesIns_Inst_Sbox_5_M11}), .c ({new_AGEMA_signal_5641, SubBytesIns_Inst_Sbox_5_M13}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M14_U1 ( .a ({new_AGEMA_signal_5024, SubBytesIns_Inst_Sbox_5_T2}), .b ({new_AGEMA_signal_5411, SubBytesIns_Inst_Sbox_5_T10}), .clk (clk), .r ({Fresh[107], Fresh[106]}), .c ({new_AGEMA_signal_5642, SubBytesIns_Inst_Sbox_5_M14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M15_U1 ( .a ({new_AGEMA_signal_5642, SubBytesIns_Inst_Sbox_5_M14}), .b ({new_AGEMA_signal_5421, SubBytesIns_Inst_Sbox_5_M11}), .c ({new_AGEMA_signal_5779, SubBytesIns_Inst_Sbox_5_M15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M16_U1 ( .a ({new_AGEMA_signal_5637, SubBytesIns_Inst_Sbox_5_M3}), .b ({new_AGEMA_signal_5636, SubBytesIns_Inst_Sbox_5_M2}), .c ({new_AGEMA_signal_5780, SubBytesIns_Inst_Sbox_5_M16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M17_U1 ( .a ({new_AGEMA_signal_5638, SubBytesIns_Inst_Sbox_5_M5}), .b ({new_AGEMA_signal_10106, new_AGEMA_signal_10105}), .c ({new_AGEMA_signal_5781, SubBytesIns_Inst_Sbox_5_M17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M18_U1 ( .a ({new_AGEMA_signal_5639, SubBytesIns_Inst_Sbox_5_M8}), .b ({new_AGEMA_signal_5420, SubBytesIns_Inst_Sbox_5_M7}), .c ({new_AGEMA_signal_5782, SubBytesIns_Inst_Sbox_5_M18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M19_U1 ( .a ({new_AGEMA_signal_5778, SubBytesIns_Inst_Sbox_5_M10}), .b ({new_AGEMA_signal_5779, SubBytesIns_Inst_Sbox_5_M15}), .c ({new_AGEMA_signal_5869, SubBytesIns_Inst_Sbox_5_M19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M20_U1 ( .a ({new_AGEMA_signal_5780, SubBytesIns_Inst_Sbox_5_M16}), .b ({new_AGEMA_signal_5641, SubBytesIns_Inst_Sbox_5_M13}), .c ({new_AGEMA_signal_5870, SubBytesIns_Inst_Sbox_5_M20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M21_U1 ( .a ({new_AGEMA_signal_5781, SubBytesIns_Inst_Sbox_5_M17}), .b ({new_AGEMA_signal_5779, SubBytesIns_Inst_Sbox_5_M15}), .c ({new_AGEMA_signal_5871, SubBytesIns_Inst_Sbox_5_M21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M22_U1 ( .a ({new_AGEMA_signal_5782, SubBytesIns_Inst_Sbox_5_M18}), .b ({new_AGEMA_signal_5641, SubBytesIns_Inst_Sbox_5_M13}), .c ({new_AGEMA_signal_5872, SubBytesIns_Inst_Sbox_5_M22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M23_U1 ( .a ({new_AGEMA_signal_5869, SubBytesIns_Inst_Sbox_5_M19}), .b ({new_AGEMA_signal_10108, new_AGEMA_signal_10107}), .c ({new_AGEMA_signal_5949, SubBytesIns_Inst_Sbox_5_M23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M24_U1 ( .a ({new_AGEMA_signal_5872, SubBytesIns_Inst_Sbox_5_M22}), .b ({new_AGEMA_signal_5949, SubBytesIns_Inst_Sbox_5_M23}), .c ({new_AGEMA_signal_6038, SubBytesIns_Inst_Sbox_5_M24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M27_U1 ( .a ({new_AGEMA_signal_5870, SubBytesIns_Inst_Sbox_5_M20}), .b ({new_AGEMA_signal_5871, SubBytesIns_Inst_Sbox_5_M21}), .c ({new_AGEMA_signal_5951, SubBytesIns_Inst_Sbox_5_M27}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M1_U1 ( .a ({new_AGEMA_signal_5215, SubBytesIns_Inst_Sbox_6_T13}), .b ({new_AGEMA_signal_5213, SubBytesIns_Inst_Sbox_6_T6}), .clk (clk), .r ({Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_5430, SubBytesIns_Inst_Sbox_6_M1}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M2_U1 ( .a ({new_AGEMA_signal_5428, SubBytesIns_Inst_Sbox_6_T23}), .b ({new_AGEMA_signal_5423, SubBytesIns_Inst_Sbox_6_T8}), .clk (clk), .r ({Fresh[111], Fresh[110]}), .c ({new_AGEMA_signal_5645, SubBytesIns_Inst_Sbox_6_M2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M3_U1 ( .a ({new_AGEMA_signal_10110, new_AGEMA_signal_10109}), .b ({new_AGEMA_signal_5430, SubBytesIns_Inst_Sbox_6_M1}), .c ({new_AGEMA_signal_5646, SubBytesIns_Inst_Sbox_6_M3}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M4_U1 ( .a ({new_AGEMA_signal_5218, SubBytesIns_Inst_Sbox_6_T19}), .b ({ciphertext_s1[48], ciphertext_s0[48]}), .clk (clk), .r ({Fresh[113], Fresh[112]}), .c ({new_AGEMA_signal_5431, SubBytesIns_Inst_Sbox_6_M4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M5_U1 ( .a ({new_AGEMA_signal_5431, SubBytesIns_Inst_Sbox_6_M4}), .b ({new_AGEMA_signal_5430, SubBytesIns_Inst_Sbox_6_M1}), .c ({new_AGEMA_signal_5647, SubBytesIns_Inst_Sbox_6_M5}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M6_U1 ( .a ({new_AGEMA_signal_5035, SubBytesIns_Inst_Sbox_6_T3}), .b ({new_AGEMA_signal_5217, SubBytesIns_Inst_Sbox_6_T16}), .clk (clk), .r ({Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_5432, SubBytesIns_Inst_Sbox_6_M6}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M7_U1 ( .a ({new_AGEMA_signal_5219, SubBytesIns_Inst_Sbox_6_T22}), .b ({new_AGEMA_signal_5214, SubBytesIns_Inst_Sbox_6_T9}), .clk (clk), .r ({Fresh[117], Fresh[116]}), .c ({new_AGEMA_signal_5433, SubBytesIns_Inst_Sbox_6_M7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M8_U1 ( .a ({new_AGEMA_signal_10112, new_AGEMA_signal_10111}), .b ({new_AGEMA_signal_5432, SubBytesIns_Inst_Sbox_6_M6}), .c ({new_AGEMA_signal_5648, SubBytesIns_Inst_Sbox_6_M8}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M9_U1 ( .a ({new_AGEMA_signal_5427, SubBytesIns_Inst_Sbox_6_T20}), .b ({new_AGEMA_signal_5426, SubBytesIns_Inst_Sbox_6_T17}), .clk (clk), .r ({Fresh[119], Fresh[118]}), .c ({new_AGEMA_signal_5649, SubBytesIns_Inst_Sbox_6_M9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M10_U1 ( .a ({new_AGEMA_signal_5649, SubBytesIns_Inst_Sbox_6_M9}), .b ({new_AGEMA_signal_5432, SubBytesIns_Inst_Sbox_6_M6}), .c ({new_AGEMA_signal_5783, SubBytesIns_Inst_Sbox_6_M10}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M11_U1 ( .a ({new_AGEMA_signal_5033, SubBytesIns_Inst_Sbox_6_T1}), .b ({new_AGEMA_signal_5216, SubBytesIns_Inst_Sbox_6_T15}), .clk (clk), .r ({Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_5434, SubBytesIns_Inst_Sbox_6_M11}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M12_U1 ( .a ({new_AGEMA_signal_5036, SubBytesIns_Inst_Sbox_6_T4}), .b ({new_AGEMA_signal_5220, SubBytesIns_Inst_Sbox_6_T27}), .clk (clk), .r ({Fresh[123], Fresh[122]}), .c ({new_AGEMA_signal_5435, SubBytesIns_Inst_Sbox_6_M12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M13_U1 ( .a ({new_AGEMA_signal_5435, SubBytesIns_Inst_Sbox_6_M12}), .b ({new_AGEMA_signal_5434, SubBytesIns_Inst_Sbox_6_M11}), .c ({new_AGEMA_signal_5650, SubBytesIns_Inst_Sbox_6_M13}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M14_U1 ( .a ({new_AGEMA_signal_5034, SubBytesIns_Inst_Sbox_6_T2}), .b ({new_AGEMA_signal_5424, SubBytesIns_Inst_Sbox_6_T10}), .clk (clk), .r ({Fresh[125], Fresh[124]}), .c ({new_AGEMA_signal_5651, SubBytesIns_Inst_Sbox_6_M14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M15_U1 ( .a ({new_AGEMA_signal_5651, SubBytesIns_Inst_Sbox_6_M14}), .b ({new_AGEMA_signal_5434, SubBytesIns_Inst_Sbox_6_M11}), .c ({new_AGEMA_signal_5784, SubBytesIns_Inst_Sbox_6_M15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M16_U1 ( .a ({new_AGEMA_signal_5646, SubBytesIns_Inst_Sbox_6_M3}), .b ({new_AGEMA_signal_5645, SubBytesIns_Inst_Sbox_6_M2}), .c ({new_AGEMA_signal_5785, SubBytesIns_Inst_Sbox_6_M16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M17_U1 ( .a ({new_AGEMA_signal_5647, SubBytesIns_Inst_Sbox_6_M5}), .b ({new_AGEMA_signal_10114, new_AGEMA_signal_10113}), .c ({new_AGEMA_signal_5786, SubBytesIns_Inst_Sbox_6_M17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M18_U1 ( .a ({new_AGEMA_signal_5648, SubBytesIns_Inst_Sbox_6_M8}), .b ({new_AGEMA_signal_5433, SubBytesIns_Inst_Sbox_6_M7}), .c ({new_AGEMA_signal_5787, SubBytesIns_Inst_Sbox_6_M18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M19_U1 ( .a ({new_AGEMA_signal_5783, SubBytesIns_Inst_Sbox_6_M10}), .b ({new_AGEMA_signal_5784, SubBytesIns_Inst_Sbox_6_M15}), .c ({new_AGEMA_signal_5873, SubBytesIns_Inst_Sbox_6_M19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M20_U1 ( .a ({new_AGEMA_signal_5785, SubBytesIns_Inst_Sbox_6_M16}), .b ({new_AGEMA_signal_5650, SubBytesIns_Inst_Sbox_6_M13}), .c ({new_AGEMA_signal_5874, SubBytesIns_Inst_Sbox_6_M20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M21_U1 ( .a ({new_AGEMA_signal_5786, SubBytesIns_Inst_Sbox_6_M17}), .b ({new_AGEMA_signal_5784, SubBytesIns_Inst_Sbox_6_M15}), .c ({new_AGEMA_signal_5875, SubBytesIns_Inst_Sbox_6_M21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M22_U1 ( .a ({new_AGEMA_signal_5787, SubBytesIns_Inst_Sbox_6_M18}), .b ({new_AGEMA_signal_5650, SubBytesIns_Inst_Sbox_6_M13}), .c ({new_AGEMA_signal_5876, SubBytesIns_Inst_Sbox_6_M22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M23_U1 ( .a ({new_AGEMA_signal_5873, SubBytesIns_Inst_Sbox_6_M19}), .b ({new_AGEMA_signal_10116, new_AGEMA_signal_10115}), .c ({new_AGEMA_signal_5953, SubBytesIns_Inst_Sbox_6_M23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M24_U1 ( .a ({new_AGEMA_signal_5876, SubBytesIns_Inst_Sbox_6_M22}), .b ({new_AGEMA_signal_5953, SubBytesIns_Inst_Sbox_6_M23}), .c ({new_AGEMA_signal_6043, SubBytesIns_Inst_Sbox_6_M24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M27_U1 ( .a ({new_AGEMA_signal_5874, SubBytesIns_Inst_Sbox_6_M20}), .b ({new_AGEMA_signal_5875, SubBytesIns_Inst_Sbox_6_M21}), .c ({new_AGEMA_signal_5955, SubBytesIns_Inst_Sbox_6_M27}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M1_U1 ( .a ({new_AGEMA_signal_5223, SubBytesIns_Inst_Sbox_7_T13}), .b ({new_AGEMA_signal_5221, SubBytesIns_Inst_Sbox_7_T6}), .clk (clk), .r ({Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_5443, SubBytesIns_Inst_Sbox_7_M1}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M2_U1 ( .a ({new_AGEMA_signal_5441, SubBytesIns_Inst_Sbox_7_T23}), .b ({new_AGEMA_signal_5436, SubBytesIns_Inst_Sbox_7_T8}), .clk (clk), .r ({Fresh[129], Fresh[128]}), .c ({new_AGEMA_signal_5654, SubBytesIns_Inst_Sbox_7_M2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M3_U1 ( .a ({new_AGEMA_signal_10118, new_AGEMA_signal_10117}), .b ({new_AGEMA_signal_5443, SubBytesIns_Inst_Sbox_7_M1}), .c ({new_AGEMA_signal_5655, SubBytesIns_Inst_Sbox_7_M3}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M4_U1 ( .a ({new_AGEMA_signal_5226, SubBytesIns_Inst_Sbox_7_T19}), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .clk (clk), .r ({Fresh[131], Fresh[130]}), .c ({new_AGEMA_signal_5444, SubBytesIns_Inst_Sbox_7_M4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M5_U1 ( .a ({new_AGEMA_signal_5444, SubBytesIns_Inst_Sbox_7_M4}), .b ({new_AGEMA_signal_5443, SubBytesIns_Inst_Sbox_7_M1}), .c ({new_AGEMA_signal_5656, SubBytesIns_Inst_Sbox_7_M5}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M6_U1 ( .a ({new_AGEMA_signal_5045, SubBytesIns_Inst_Sbox_7_T3}), .b ({new_AGEMA_signal_5225, SubBytesIns_Inst_Sbox_7_T16}), .clk (clk), .r ({Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_5445, SubBytesIns_Inst_Sbox_7_M6}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M7_U1 ( .a ({new_AGEMA_signal_5227, SubBytesIns_Inst_Sbox_7_T22}), .b ({new_AGEMA_signal_5222, SubBytesIns_Inst_Sbox_7_T9}), .clk (clk), .r ({Fresh[135], Fresh[134]}), .c ({new_AGEMA_signal_5446, SubBytesIns_Inst_Sbox_7_M7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M8_U1 ( .a ({new_AGEMA_signal_10120, new_AGEMA_signal_10119}), .b ({new_AGEMA_signal_5445, SubBytesIns_Inst_Sbox_7_M6}), .c ({new_AGEMA_signal_5657, SubBytesIns_Inst_Sbox_7_M8}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M9_U1 ( .a ({new_AGEMA_signal_5440, SubBytesIns_Inst_Sbox_7_T20}), .b ({new_AGEMA_signal_5439, SubBytesIns_Inst_Sbox_7_T17}), .clk (clk), .r ({Fresh[137], Fresh[136]}), .c ({new_AGEMA_signal_5658, SubBytesIns_Inst_Sbox_7_M9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M10_U1 ( .a ({new_AGEMA_signal_5658, SubBytesIns_Inst_Sbox_7_M9}), .b ({new_AGEMA_signal_5445, SubBytesIns_Inst_Sbox_7_M6}), .c ({new_AGEMA_signal_5788, SubBytesIns_Inst_Sbox_7_M10}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M11_U1 ( .a ({new_AGEMA_signal_5043, SubBytesIns_Inst_Sbox_7_T1}), .b ({new_AGEMA_signal_5224, SubBytesIns_Inst_Sbox_7_T15}), .clk (clk), .r ({Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_5447, SubBytesIns_Inst_Sbox_7_M11}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M12_U1 ( .a ({new_AGEMA_signal_5046, SubBytesIns_Inst_Sbox_7_T4}), .b ({new_AGEMA_signal_5228, SubBytesIns_Inst_Sbox_7_T27}), .clk (clk), .r ({Fresh[141], Fresh[140]}), .c ({new_AGEMA_signal_5448, SubBytesIns_Inst_Sbox_7_M12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M13_U1 ( .a ({new_AGEMA_signal_5448, SubBytesIns_Inst_Sbox_7_M12}), .b ({new_AGEMA_signal_5447, SubBytesIns_Inst_Sbox_7_M11}), .c ({new_AGEMA_signal_5659, SubBytesIns_Inst_Sbox_7_M13}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M14_U1 ( .a ({new_AGEMA_signal_5044, SubBytesIns_Inst_Sbox_7_T2}), .b ({new_AGEMA_signal_5437, SubBytesIns_Inst_Sbox_7_T10}), .clk (clk), .r ({Fresh[143], Fresh[142]}), .c ({new_AGEMA_signal_5660, SubBytesIns_Inst_Sbox_7_M14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M15_U1 ( .a ({new_AGEMA_signal_5660, SubBytesIns_Inst_Sbox_7_M14}), .b ({new_AGEMA_signal_5447, SubBytesIns_Inst_Sbox_7_M11}), .c ({new_AGEMA_signal_5789, SubBytesIns_Inst_Sbox_7_M15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M16_U1 ( .a ({new_AGEMA_signal_5655, SubBytesIns_Inst_Sbox_7_M3}), .b ({new_AGEMA_signal_5654, SubBytesIns_Inst_Sbox_7_M2}), .c ({new_AGEMA_signal_5790, SubBytesIns_Inst_Sbox_7_M16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M17_U1 ( .a ({new_AGEMA_signal_5656, SubBytesIns_Inst_Sbox_7_M5}), .b ({new_AGEMA_signal_10122, new_AGEMA_signal_10121}), .c ({new_AGEMA_signal_5791, SubBytesIns_Inst_Sbox_7_M17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M18_U1 ( .a ({new_AGEMA_signal_5657, SubBytesIns_Inst_Sbox_7_M8}), .b ({new_AGEMA_signal_5446, SubBytesIns_Inst_Sbox_7_M7}), .c ({new_AGEMA_signal_5792, SubBytesIns_Inst_Sbox_7_M18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M19_U1 ( .a ({new_AGEMA_signal_5788, SubBytesIns_Inst_Sbox_7_M10}), .b ({new_AGEMA_signal_5789, SubBytesIns_Inst_Sbox_7_M15}), .c ({new_AGEMA_signal_5877, SubBytesIns_Inst_Sbox_7_M19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M20_U1 ( .a ({new_AGEMA_signal_5790, SubBytesIns_Inst_Sbox_7_M16}), .b ({new_AGEMA_signal_5659, SubBytesIns_Inst_Sbox_7_M13}), .c ({new_AGEMA_signal_5878, SubBytesIns_Inst_Sbox_7_M20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M21_U1 ( .a ({new_AGEMA_signal_5791, SubBytesIns_Inst_Sbox_7_M17}), .b ({new_AGEMA_signal_5789, SubBytesIns_Inst_Sbox_7_M15}), .c ({new_AGEMA_signal_5879, SubBytesIns_Inst_Sbox_7_M21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M22_U1 ( .a ({new_AGEMA_signal_5792, SubBytesIns_Inst_Sbox_7_M18}), .b ({new_AGEMA_signal_5659, SubBytesIns_Inst_Sbox_7_M13}), .c ({new_AGEMA_signal_5880, SubBytesIns_Inst_Sbox_7_M22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M23_U1 ( .a ({new_AGEMA_signal_5877, SubBytesIns_Inst_Sbox_7_M19}), .b ({new_AGEMA_signal_10124, new_AGEMA_signal_10123}), .c ({new_AGEMA_signal_5957, SubBytesIns_Inst_Sbox_7_M23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M24_U1 ( .a ({new_AGEMA_signal_5880, SubBytesIns_Inst_Sbox_7_M22}), .b ({new_AGEMA_signal_5957, SubBytesIns_Inst_Sbox_7_M23}), .c ({new_AGEMA_signal_6048, SubBytesIns_Inst_Sbox_7_M24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M27_U1 ( .a ({new_AGEMA_signal_5878, SubBytesIns_Inst_Sbox_7_M20}), .b ({new_AGEMA_signal_5879, SubBytesIns_Inst_Sbox_7_M21}), .c ({new_AGEMA_signal_5959, SubBytesIns_Inst_Sbox_7_M27}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M1_U1 ( .a ({new_AGEMA_signal_5231, SubBytesIns_Inst_Sbox_8_T13}), .b ({new_AGEMA_signal_5229, SubBytesIns_Inst_Sbox_8_T6}), .clk (clk), .r ({Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_5456, SubBytesIns_Inst_Sbox_8_M1}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M2_U1 ( .a ({new_AGEMA_signal_5454, SubBytesIns_Inst_Sbox_8_T23}), .b ({new_AGEMA_signal_5449, SubBytesIns_Inst_Sbox_8_T8}), .clk (clk), .r ({Fresh[147], Fresh[146]}), .c ({new_AGEMA_signal_5663, SubBytesIns_Inst_Sbox_8_M2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M3_U1 ( .a ({new_AGEMA_signal_10126, new_AGEMA_signal_10125}), .b ({new_AGEMA_signal_5456, SubBytesIns_Inst_Sbox_8_M1}), .c ({new_AGEMA_signal_5664, SubBytesIns_Inst_Sbox_8_M3}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M4_U1 ( .a ({new_AGEMA_signal_5234, SubBytesIns_Inst_Sbox_8_T19}), .b ({ciphertext_s1[64], ciphertext_s0[64]}), .clk (clk), .r ({Fresh[149], Fresh[148]}), .c ({new_AGEMA_signal_5457, SubBytesIns_Inst_Sbox_8_M4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M5_U1 ( .a ({new_AGEMA_signal_5457, SubBytesIns_Inst_Sbox_8_M4}), .b ({new_AGEMA_signal_5456, SubBytesIns_Inst_Sbox_8_M1}), .c ({new_AGEMA_signal_5665, SubBytesIns_Inst_Sbox_8_M5}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M6_U1 ( .a ({new_AGEMA_signal_5055, SubBytesIns_Inst_Sbox_8_T3}), .b ({new_AGEMA_signal_5233, SubBytesIns_Inst_Sbox_8_T16}), .clk (clk), .r ({Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_5458, SubBytesIns_Inst_Sbox_8_M6}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M7_U1 ( .a ({new_AGEMA_signal_5235, SubBytesIns_Inst_Sbox_8_T22}), .b ({new_AGEMA_signal_5230, SubBytesIns_Inst_Sbox_8_T9}), .clk (clk), .r ({Fresh[153], Fresh[152]}), .c ({new_AGEMA_signal_5459, SubBytesIns_Inst_Sbox_8_M7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M8_U1 ( .a ({new_AGEMA_signal_10128, new_AGEMA_signal_10127}), .b ({new_AGEMA_signal_5458, SubBytesIns_Inst_Sbox_8_M6}), .c ({new_AGEMA_signal_5666, SubBytesIns_Inst_Sbox_8_M8}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M9_U1 ( .a ({new_AGEMA_signal_5453, SubBytesIns_Inst_Sbox_8_T20}), .b ({new_AGEMA_signal_5452, SubBytesIns_Inst_Sbox_8_T17}), .clk (clk), .r ({Fresh[155], Fresh[154]}), .c ({new_AGEMA_signal_5667, SubBytesIns_Inst_Sbox_8_M9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M10_U1 ( .a ({new_AGEMA_signal_5667, SubBytesIns_Inst_Sbox_8_M9}), .b ({new_AGEMA_signal_5458, SubBytesIns_Inst_Sbox_8_M6}), .c ({new_AGEMA_signal_5793, SubBytesIns_Inst_Sbox_8_M10}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M11_U1 ( .a ({new_AGEMA_signal_5053, SubBytesIns_Inst_Sbox_8_T1}), .b ({new_AGEMA_signal_5232, SubBytesIns_Inst_Sbox_8_T15}), .clk (clk), .r ({Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_5460, SubBytesIns_Inst_Sbox_8_M11}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M12_U1 ( .a ({new_AGEMA_signal_5056, SubBytesIns_Inst_Sbox_8_T4}), .b ({new_AGEMA_signal_5236, SubBytesIns_Inst_Sbox_8_T27}), .clk (clk), .r ({Fresh[159], Fresh[158]}), .c ({new_AGEMA_signal_5461, SubBytesIns_Inst_Sbox_8_M12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M13_U1 ( .a ({new_AGEMA_signal_5461, SubBytesIns_Inst_Sbox_8_M12}), .b ({new_AGEMA_signal_5460, SubBytesIns_Inst_Sbox_8_M11}), .c ({new_AGEMA_signal_5668, SubBytesIns_Inst_Sbox_8_M13}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M14_U1 ( .a ({new_AGEMA_signal_5054, SubBytesIns_Inst_Sbox_8_T2}), .b ({new_AGEMA_signal_5450, SubBytesIns_Inst_Sbox_8_T10}), .clk (clk), .r ({Fresh[161], Fresh[160]}), .c ({new_AGEMA_signal_5669, SubBytesIns_Inst_Sbox_8_M14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M15_U1 ( .a ({new_AGEMA_signal_5669, SubBytesIns_Inst_Sbox_8_M14}), .b ({new_AGEMA_signal_5460, SubBytesIns_Inst_Sbox_8_M11}), .c ({new_AGEMA_signal_5794, SubBytesIns_Inst_Sbox_8_M15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M16_U1 ( .a ({new_AGEMA_signal_5664, SubBytesIns_Inst_Sbox_8_M3}), .b ({new_AGEMA_signal_5663, SubBytesIns_Inst_Sbox_8_M2}), .c ({new_AGEMA_signal_5795, SubBytesIns_Inst_Sbox_8_M16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M17_U1 ( .a ({new_AGEMA_signal_5665, SubBytesIns_Inst_Sbox_8_M5}), .b ({new_AGEMA_signal_10130, new_AGEMA_signal_10129}), .c ({new_AGEMA_signal_5796, SubBytesIns_Inst_Sbox_8_M17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M18_U1 ( .a ({new_AGEMA_signal_5666, SubBytesIns_Inst_Sbox_8_M8}), .b ({new_AGEMA_signal_5459, SubBytesIns_Inst_Sbox_8_M7}), .c ({new_AGEMA_signal_5797, SubBytesIns_Inst_Sbox_8_M18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M19_U1 ( .a ({new_AGEMA_signal_5793, SubBytesIns_Inst_Sbox_8_M10}), .b ({new_AGEMA_signal_5794, SubBytesIns_Inst_Sbox_8_M15}), .c ({new_AGEMA_signal_5881, SubBytesIns_Inst_Sbox_8_M19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M20_U1 ( .a ({new_AGEMA_signal_5795, SubBytesIns_Inst_Sbox_8_M16}), .b ({new_AGEMA_signal_5668, SubBytesIns_Inst_Sbox_8_M13}), .c ({new_AGEMA_signal_5882, SubBytesIns_Inst_Sbox_8_M20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M21_U1 ( .a ({new_AGEMA_signal_5796, SubBytesIns_Inst_Sbox_8_M17}), .b ({new_AGEMA_signal_5794, SubBytesIns_Inst_Sbox_8_M15}), .c ({new_AGEMA_signal_5883, SubBytesIns_Inst_Sbox_8_M21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M22_U1 ( .a ({new_AGEMA_signal_5797, SubBytesIns_Inst_Sbox_8_M18}), .b ({new_AGEMA_signal_5668, SubBytesIns_Inst_Sbox_8_M13}), .c ({new_AGEMA_signal_5884, SubBytesIns_Inst_Sbox_8_M22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M23_U1 ( .a ({new_AGEMA_signal_5881, SubBytesIns_Inst_Sbox_8_M19}), .b ({new_AGEMA_signal_10132, new_AGEMA_signal_10131}), .c ({new_AGEMA_signal_5961, SubBytesIns_Inst_Sbox_8_M23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M24_U1 ( .a ({new_AGEMA_signal_5884, SubBytesIns_Inst_Sbox_8_M22}), .b ({new_AGEMA_signal_5961, SubBytesIns_Inst_Sbox_8_M23}), .c ({new_AGEMA_signal_6053, SubBytesIns_Inst_Sbox_8_M24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M27_U1 ( .a ({new_AGEMA_signal_5882, SubBytesIns_Inst_Sbox_8_M20}), .b ({new_AGEMA_signal_5883, SubBytesIns_Inst_Sbox_8_M21}), .c ({new_AGEMA_signal_5963, SubBytesIns_Inst_Sbox_8_M27}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M1_U1 ( .a ({new_AGEMA_signal_5239, SubBytesIns_Inst_Sbox_9_T13}), .b ({new_AGEMA_signal_5237, SubBytesIns_Inst_Sbox_9_T6}), .clk (clk), .r ({Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_5469, SubBytesIns_Inst_Sbox_9_M1}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M2_U1 ( .a ({new_AGEMA_signal_5467, SubBytesIns_Inst_Sbox_9_T23}), .b ({new_AGEMA_signal_5462, SubBytesIns_Inst_Sbox_9_T8}), .clk (clk), .r ({Fresh[165], Fresh[164]}), .c ({new_AGEMA_signal_5672, SubBytesIns_Inst_Sbox_9_M2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M3_U1 ( .a ({new_AGEMA_signal_10134, new_AGEMA_signal_10133}), .b ({new_AGEMA_signal_5469, SubBytesIns_Inst_Sbox_9_M1}), .c ({new_AGEMA_signal_5673, SubBytesIns_Inst_Sbox_9_M3}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M4_U1 ( .a ({new_AGEMA_signal_5242, SubBytesIns_Inst_Sbox_9_T19}), .b ({ciphertext_s1[72], ciphertext_s0[72]}), .clk (clk), .r ({Fresh[167], Fresh[166]}), .c ({new_AGEMA_signal_5470, SubBytesIns_Inst_Sbox_9_M4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M5_U1 ( .a ({new_AGEMA_signal_5470, SubBytesIns_Inst_Sbox_9_M4}), .b ({new_AGEMA_signal_5469, SubBytesIns_Inst_Sbox_9_M1}), .c ({new_AGEMA_signal_5674, SubBytesIns_Inst_Sbox_9_M5}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M6_U1 ( .a ({new_AGEMA_signal_5065, SubBytesIns_Inst_Sbox_9_T3}), .b ({new_AGEMA_signal_5241, SubBytesIns_Inst_Sbox_9_T16}), .clk (clk), .r ({Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_5471, SubBytesIns_Inst_Sbox_9_M6}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M7_U1 ( .a ({new_AGEMA_signal_5243, SubBytesIns_Inst_Sbox_9_T22}), .b ({new_AGEMA_signal_5238, SubBytesIns_Inst_Sbox_9_T9}), .clk (clk), .r ({Fresh[171], Fresh[170]}), .c ({new_AGEMA_signal_5472, SubBytesIns_Inst_Sbox_9_M7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M8_U1 ( .a ({new_AGEMA_signal_10136, new_AGEMA_signal_10135}), .b ({new_AGEMA_signal_5471, SubBytesIns_Inst_Sbox_9_M6}), .c ({new_AGEMA_signal_5675, SubBytesIns_Inst_Sbox_9_M8}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M9_U1 ( .a ({new_AGEMA_signal_5466, SubBytesIns_Inst_Sbox_9_T20}), .b ({new_AGEMA_signal_5465, SubBytesIns_Inst_Sbox_9_T17}), .clk (clk), .r ({Fresh[173], Fresh[172]}), .c ({new_AGEMA_signal_5676, SubBytesIns_Inst_Sbox_9_M9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M10_U1 ( .a ({new_AGEMA_signal_5676, SubBytesIns_Inst_Sbox_9_M9}), .b ({new_AGEMA_signal_5471, SubBytesIns_Inst_Sbox_9_M6}), .c ({new_AGEMA_signal_5798, SubBytesIns_Inst_Sbox_9_M10}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M11_U1 ( .a ({new_AGEMA_signal_5063, SubBytesIns_Inst_Sbox_9_T1}), .b ({new_AGEMA_signal_5240, SubBytesIns_Inst_Sbox_9_T15}), .clk (clk), .r ({Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_5473, SubBytesIns_Inst_Sbox_9_M11}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M12_U1 ( .a ({new_AGEMA_signal_5066, SubBytesIns_Inst_Sbox_9_T4}), .b ({new_AGEMA_signal_5244, SubBytesIns_Inst_Sbox_9_T27}), .clk (clk), .r ({Fresh[177], Fresh[176]}), .c ({new_AGEMA_signal_5474, SubBytesIns_Inst_Sbox_9_M12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M13_U1 ( .a ({new_AGEMA_signal_5474, SubBytesIns_Inst_Sbox_9_M12}), .b ({new_AGEMA_signal_5473, SubBytesIns_Inst_Sbox_9_M11}), .c ({new_AGEMA_signal_5677, SubBytesIns_Inst_Sbox_9_M13}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M14_U1 ( .a ({new_AGEMA_signal_5064, SubBytesIns_Inst_Sbox_9_T2}), .b ({new_AGEMA_signal_5463, SubBytesIns_Inst_Sbox_9_T10}), .clk (clk), .r ({Fresh[179], Fresh[178]}), .c ({new_AGEMA_signal_5678, SubBytesIns_Inst_Sbox_9_M14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M15_U1 ( .a ({new_AGEMA_signal_5678, SubBytesIns_Inst_Sbox_9_M14}), .b ({new_AGEMA_signal_5473, SubBytesIns_Inst_Sbox_9_M11}), .c ({new_AGEMA_signal_5799, SubBytesIns_Inst_Sbox_9_M15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M16_U1 ( .a ({new_AGEMA_signal_5673, SubBytesIns_Inst_Sbox_9_M3}), .b ({new_AGEMA_signal_5672, SubBytesIns_Inst_Sbox_9_M2}), .c ({new_AGEMA_signal_5800, SubBytesIns_Inst_Sbox_9_M16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M17_U1 ( .a ({new_AGEMA_signal_5674, SubBytesIns_Inst_Sbox_9_M5}), .b ({new_AGEMA_signal_10138, new_AGEMA_signal_10137}), .c ({new_AGEMA_signal_5801, SubBytesIns_Inst_Sbox_9_M17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M18_U1 ( .a ({new_AGEMA_signal_5675, SubBytesIns_Inst_Sbox_9_M8}), .b ({new_AGEMA_signal_5472, SubBytesIns_Inst_Sbox_9_M7}), .c ({new_AGEMA_signal_5802, SubBytesIns_Inst_Sbox_9_M18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M19_U1 ( .a ({new_AGEMA_signal_5798, SubBytesIns_Inst_Sbox_9_M10}), .b ({new_AGEMA_signal_5799, SubBytesIns_Inst_Sbox_9_M15}), .c ({new_AGEMA_signal_5885, SubBytesIns_Inst_Sbox_9_M19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M20_U1 ( .a ({new_AGEMA_signal_5800, SubBytesIns_Inst_Sbox_9_M16}), .b ({new_AGEMA_signal_5677, SubBytesIns_Inst_Sbox_9_M13}), .c ({new_AGEMA_signal_5886, SubBytesIns_Inst_Sbox_9_M20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M21_U1 ( .a ({new_AGEMA_signal_5801, SubBytesIns_Inst_Sbox_9_M17}), .b ({new_AGEMA_signal_5799, SubBytesIns_Inst_Sbox_9_M15}), .c ({new_AGEMA_signal_5887, SubBytesIns_Inst_Sbox_9_M21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M22_U1 ( .a ({new_AGEMA_signal_5802, SubBytesIns_Inst_Sbox_9_M18}), .b ({new_AGEMA_signal_5677, SubBytesIns_Inst_Sbox_9_M13}), .c ({new_AGEMA_signal_5888, SubBytesIns_Inst_Sbox_9_M22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M23_U1 ( .a ({new_AGEMA_signal_5885, SubBytesIns_Inst_Sbox_9_M19}), .b ({new_AGEMA_signal_10140, new_AGEMA_signal_10139}), .c ({new_AGEMA_signal_5965, SubBytesIns_Inst_Sbox_9_M23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M24_U1 ( .a ({new_AGEMA_signal_5888, SubBytesIns_Inst_Sbox_9_M22}), .b ({new_AGEMA_signal_5965, SubBytesIns_Inst_Sbox_9_M23}), .c ({new_AGEMA_signal_6058, SubBytesIns_Inst_Sbox_9_M24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M27_U1 ( .a ({new_AGEMA_signal_5886, SubBytesIns_Inst_Sbox_9_M20}), .b ({new_AGEMA_signal_5887, SubBytesIns_Inst_Sbox_9_M21}), .c ({new_AGEMA_signal_5967, SubBytesIns_Inst_Sbox_9_M27}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M1_U1 ( .a ({new_AGEMA_signal_5247, SubBytesIns_Inst_Sbox_10_T13}), .b ({new_AGEMA_signal_5245, SubBytesIns_Inst_Sbox_10_T6}), .clk (clk), .r ({Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_5482, SubBytesIns_Inst_Sbox_10_M1}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M2_U1 ( .a ({new_AGEMA_signal_5480, SubBytesIns_Inst_Sbox_10_T23}), .b ({new_AGEMA_signal_5475, SubBytesIns_Inst_Sbox_10_T8}), .clk (clk), .r ({Fresh[183], Fresh[182]}), .c ({new_AGEMA_signal_5681, SubBytesIns_Inst_Sbox_10_M2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M3_U1 ( .a ({new_AGEMA_signal_10142, new_AGEMA_signal_10141}), .b ({new_AGEMA_signal_5482, SubBytesIns_Inst_Sbox_10_M1}), .c ({new_AGEMA_signal_5682, SubBytesIns_Inst_Sbox_10_M3}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M4_U1 ( .a ({new_AGEMA_signal_5250, SubBytesIns_Inst_Sbox_10_T19}), .b ({ciphertext_s1[80], ciphertext_s0[80]}), .clk (clk), .r ({Fresh[185], Fresh[184]}), .c ({new_AGEMA_signal_5483, SubBytesIns_Inst_Sbox_10_M4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M5_U1 ( .a ({new_AGEMA_signal_5483, SubBytesIns_Inst_Sbox_10_M4}), .b ({new_AGEMA_signal_5482, SubBytesIns_Inst_Sbox_10_M1}), .c ({new_AGEMA_signal_5683, SubBytesIns_Inst_Sbox_10_M5}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M6_U1 ( .a ({new_AGEMA_signal_5075, SubBytesIns_Inst_Sbox_10_T3}), .b ({new_AGEMA_signal_5249, SubBytesIns_Inst_Sbox_10_T16}), .clk (clk), .r ({Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_5484, SubBytesIns_Inst_Sbox_10_M6}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M7_U1 ( .a ({new_AGEMA_signal_5251, SubBytesIns_Inst_Sbox_10_T22}), .b ({new_AGEMA_signal_5246, SubBytesIns_Inst_Sbox_10_T9}), .clk (clk), .r ({Fresh[189], Fresh[188]}), .c ({new_AGEMA_signal_5485, SubBytesIns_Inst_Sbox_10_M7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M8_U1 ( .a ({new_AGEMA_signal_10144, new_AGEMA_signal_10143}), .b ({new_AGEMA_signal_5484, SubBytesIns_Inst_Sbox_10_M6}), .c ({new_AGEMA_signal_5684, SubBytesIns_Inst_Sbox_10_M8}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M9_U1 ( .a ({new_AGEMA_signal_5479, SubBytesIns_Inst_Sbox_10_T20}), .b ({new_AGEMA_signal_5478, SubBytesIns_Inst_Sbox_10_T17}), .clk (clk), .r ({Fresh[191], Fresh[190]}), .c ({new_AGEMA_signal_5685, SubBytesIns_Inst_Sbox_10_M9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M10_U1 ( .a ({new_AGEMA_signal_5685, SubBytesIns_Inst_Sbox_10_M9}), .b ({new_AGEMA_signal_5484, SubBytesIns_Inst_Sbox_10_M6}), .c ({new_AGEMA_signal_5803, SubBytesIns_Inst_Sbox_10_M10}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M11_U1 ( .a ({new_AGEMA_signal_5073, SubBytesIns_Inst_Sbox_10_T1}), .b ({new_AGEMA_signal_5248, SubBytesIns_Inst_Sbox_10_T15}), .clk (clk), .r ({Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_5486, SubBytesIns_Inst_Sbox_10_M11}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M12_U1 ( .a ({new_AGEMA_signal_5076, SubBytesIns_Inst_Sbox_10_T4}), .b ({new_AGEMA_signal_5252, SubBytesIns_Inst_Sbox_10_T27}), .clk (clk), .r ({Fresh[195], Fresh[194]}), .c ({new_AGEMA_signal_5487, SubBytesIns_Inst_Sbox_10_M12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M13_U1 ( .a ({new_AGEMA_signal_5487, SubBytesIns_Inst_Sbox_10_M12}), .b ({new_AGEMA_signal_5486, SubBytesIns_Inst_Sbox_10_M11}), .c ({new_AGEMA_signal_5686, SubBytesIns_Inst_Sbox_10_M13}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M14_U1 ( .a ({new_AGEMA_signal_5074, SubBytesIns_Inst_Sbox_10_T2}), .b ({new_AGEMA_signal_5476, SubBytesIns_Inst_Sbox_10_T10}), .clk (clk), .r ({Fresh[197], Fresh[196]}), .c ({new_AGEMA_signal_5687, SubBytesIns_Inst_Sbox_10_M14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M15_U1 ( .a ({new_AGEMA_signal_5687, SubBytesIns_Inst_Sbox_10_M14}), .b ({new_AGEMA_signal_5486, SubBytesIns_Inst_Sbox_10_M11}), .c ({new_AGEMA_signal_5804, SubBytesIns_Inst_Sbox_10_M15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M16_U1 ( .a ({new_AGEMA_signal_5682, SubBytesIns_Inst_Sbox_10_M3}), .b ({new_AGEMA_signal_5681, SubBytesIns_Inst_Sbox_10_M2}), .c ({new_AGEMA_signal_5805, SubBytesIns_Inst_Sbox_10_M16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M17_U1 ( .a ({new_AGEMA_signal_5683, SubBytesIns_Inst_Sbox_10_M5}), .b ({new_AGEMA_signal_10146, new_AGEMA_signal_10145}), .c ({new_AGEMA_signal_5806, SubBytesIns_Inst_Sbox_10_M17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M18_U1 ( .a ({new_AGEMA_signal_5684, SubBytesIns_Inst_Sbox_10_M8}), .b ({new_AGEMA_signal_5485, SubBytesIns_Inst_Sbox_10_M7}), .c ({new_AGEMA_signal_5807, SubBytesIns_Inst_Sbox_10_M18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M19_U1 ( .a ({new_AGEMA_signal_5803, SubBytesIns_Inst_Sbox_10_M10}), .b ({new_AGEMA_signal_5804, SubBytesIns_Inst_Sbox_10_M15}), .c ({new_AGEMA_signal_5889, SubBytesIns_Inst_Sbox_10_M19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M20_U1 ( .a ({new_AGEMA_signal_5805, SubBytesIns_Inst_Sbox_10_M16}), .b ({new_AGEMA_signal_5686, SubBytesIns_Inst_Sbox_10_M13}), .c ({new_AGEMA_signal_5890, SubBytesIns_Inst_Sbox_10_M20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M21_U1 ( .a ({new_AGEMA_signal_5806, SubBytesIns_Inst_Sbox_10_M17}), .b ({new_AGEMA_signal_5804, SubBytesIns_Inst_Sbox_10_M15}), .c ({new_AGEMA_signal_5891, SubBytesIns_Inst_Sbox_10_M21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M22_U1 ( .a ({new_AGEMA_signal_5807, SubBytesIns_Inst_Sbox_10_M18}), .b ({new_AGEMA_signal_5686, SubBytesIns_Inst_Sbox_10_M13}), .c ({new_AGEMA_signal_5892, SubBytesIns_Inst_Sbox_10_M22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M23_U1 ( .a ({new_AGEMA_signal_5889, SubBytesIns_Inst_Sbox_10_M19}), .b ({new_AGEMA_signal_10148, new_AGEMA_signal_10147}), .c ({new_AGEMA_signal_5969, SubBytesIns_Inst_Sbox_10_M23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M24_U1 ( .a ({new_AGEMA_signal_5892, SubBytesIns_Inst_Sbox_10_M22}), .b ({new_AGEMA_signal_5969, SubBytesIns_Inst_Sbox_10_M23}), .c ({new_AGEMA_signal_6063, SubBytesIns_Inst_Sbox_10_M24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M27_U1 ( .a ({new_AGEMA_signal_5890, SubBytesIns_Inst_Sbox_10_M20}), .b ({new_AGEMA_signal_5891, SubBytesIns_Inst_Sbox_10_M21}), .c ({new_AGEMA_signal_5971, SubBytesIns_Inst_Sbox_10_M27}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M1_U1 ( .a ({new_AGEMA_signal_5255, SubBytesIns_Inst_Sbox_11_T13}), .b ({new_AGEMA_signal_5253, SubBytesIns_Inst_Sbox_11_T6}), .clk (clk), .r ({Fresh[199], Fresh[198]}), .c ({new_AGEMA_signal_5495, SubBytesIns_Inst_Sbox_11_M1}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M2_U1 ( .a ({new_AGEMA_signal_5493, SubBytesIns_Inst_Sbox_11_T23}), .b ({new_AGEMA_signal_5488, SubBytesIns_Inst_Sbox_11_T8}), .clk (clk), .r ({Fresh[201], Fresh[200]}), .c ({new_AGEMA_signal_5690, SubBytesIns_Inst_Sbox_11_M2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M3_U1 ( .a ({new_AGEMA_signal_10150, new_AGEMA_signal_10149}), .b ({new_AGEMA_signal_5495, SubBytesIns_Inst_Sbox_11_M1}), .c ({new_AGEMA_signal_5691, SubBytesIns_Inst_Sbox_11_M3}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M4_U1 ( .a ({new_AGEMA_signal_5258, SubBytesIns_Inst_Sbox_11_T19}), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .clk (clk), .r ({Fresh[203], Fresh[202]}), .c ({new_AGEMA_signal_5496, SubBytesIns_Inst_Sbox_11_M4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M5_U1 ( .a ({new_AGEMA_signal_5496, SubBytesIns_Inst_Sbox_11_M4}), .b ({new_AGEMA_signal_5495, SubBytesIns_Inst_Sbox_11_M1}), .c ({new_AGEMA_signal_5692, SubBytesIns_Inst_Sbox_11_M5}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M6_U1 ( .a ({new_AGEMA_signal_5085, SubBytesIns_Inst_Sbox_11_T3}), .b ({new_AGEMA_signal_5257, SubBytesIns_Inst_Sbox_11_T16}), .clk (clk), .r ({Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_5497, SubBytesIns_Inst_Sbox_11_M6}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M7_U1 ( .a ({new_AGEMA_signal_5259, SubBytesIns_Inst_Sbox_11_T22}), .b ({new_AGEMA_signal_5254, SubBytesIns_Inst_Sbox_11_T9}), .clk (clk), .r ({Fresh[207], Fresh[206]}), .c ({new_AGEMA_signal_5498, SubBytesIns_Inst_Sbox_11_M7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M8_U1 ( .a ({new_AGEMA_signal_10152, new_AGEMA_signal_10151}), .b ({new_AGEMA_signal_5497, SubBytesIns_Inst_Sbox_11_M6}), .c ({new_AGEMA_signal_5693, SubBytesIns_Inst_Sbox_11_M8}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M9_U1 ( .a ({new_AGEMA_signal_5492, SubBytesIns_Inst_Sbox_11_T20}), .b ({new_AGEMA_signal_5491, SubBytesIns_Inst_Sbox_11_T17}), .clk (clk), .r ({Fresh[209], Fresh[208]}), .c ({new_AGEMA_signal_5694, SubBytesIns_Inst_Sbox_11_M9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M10_U1 ( .a ({new_AGEMA_signal_5694, SubBytesIns_Inst_Sbox_11_M9}), .b ({new_AGEMA_signal_5497, SubBytesIns_Inst_Sbox_11_M6}), .c ({new_AGEMA_signal_5808, SubBytesIns_Inst_Sbox_11_M10}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M11_U1 ( .a ({new_AGEMA_signal_5083, SubBytesIns_Inst_Sbox_11_T1}), .b ({new_AGEMA_signal_5256, SubBytesIns_Inst_Sbox_11_T15}), .clk (clk), .r ({Fresh[211], Fresh[210]}), .c ({new_AGEMA_signal_5499, SubBytesIns_Inst_Sbox_11_M11}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M12_U1 ( .a ({new_AGEMA_signal_5086, SubBytesIns_Inst_Sbox_11_T4}), .b ({new_AGEMA_signal_5260, SubBytesIns_Inst_Sbox_11_T27}), .clk (clk), .r ({Fresh[213], Fresh[212]}), .c ({new_AGEMA_signal_5500, SubBytesIns_Inst_Sbox_11_M12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M13_U1 ( .a ({new_AGEMA_signal_5500, SubBytesIns_Inst_Sbox_11_M12}), .b ({new_AGEMA_signal_5499, SubBytesIns_Inst_Sbox_11_M11}), .c ({new_AGEMA_signal_5695, SubBytesIns_Inst_Sbox_11_M13}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M14_U1 ( .a ({new_AGEMA_signal_5084, SubBytesIns_Inst_Sbox_11_T2}), .b ({new_AGEMA_signal_5489, SubBytesIns_Inst_Sbox_11_T10}), .clk (clk), .r ({Fresh[215], Fresh[214]}), .c ({new_AGEMA_signal_5696, SubBytesIns_Inst_Sbox_11_M14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M15_U1 ( .a ({new_AGEMA_signal_5696, SubBytesIns_Inst_Sbox_11_M14}), .b ({new_AGEMA_signal_5499, SubBytesIns_Inst_Sbox_11_M11}), .c ({new_AGEMA_signal_5809, SubBytesIns_Inst_Sbox_11_M15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M16_U1 ( .a ({new_AGEMA_signal_5691, SubBytesIns_Inst_Sbox_11_M3}), .b ({new_AGEMA_signal_5690, SubBytesIns_Inst_Sbox_11_M2}), .c ({new_AGEMA_signal_5810, SubBytesIns_Inst_Sbox_11_M16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M17_U1 ( .a ({new_AGEMA_signal_5692, SubBytesIns_Inst_Sbox_11_M5}), .b ({new_AGEMA_signal_10154, new_AGEMA_signal_10153}), .c ({new_AGEMA_signal_5811, SubBytesIns_Inst_Sbox_11_M17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M18_U1 ( .a ({new_AGEMA_signal_5693, SubBytesIns_Inst_Sbox_11_M8}), .b ({new_AGEMA_signal_5498, SubBytesIns_Inst_Sbox_11_M7}), .c ({new_AGEMA_signal_5812, SubBytesIns_Inst_Sbox_11_M18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M19_U1 ( .a ({new_AGEMA_signal_5808, SubBytesIns_Inst_Sbox_11_M10}), .b ({new_AGEMA_signal_5809, SubBytesIns_Inst_Sbox_11_M15}), .c ({new_AGEMA_signal_5893, SubBytesIns_Inst_Sbox_11_M19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M20_U1 ( .a ({new_AGEMA_signal_5810, SubBytesIns_Inst_Sbox_11_M16}), .b ({new_AGEMA_signal_5695, SubBytesIns_Inst_Sbox_11_M13}), .c ({new_AGEMA_signal_5894, SubBytesIns_Inst_Sbox_11_M20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M21_U1 ( .a ({new_AGEMA_signal_5811, SubBytesIns_Inst_Sbox_11_M17}), .b ({new_AGEMA_signal_5809, SubBytesIns_Inst_Sbox_11_M15}), .c ({new_AGEMA_signal_5895, SubBytesIns_Inst_Sbox_11_M21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M22_U1 ( .a ({new_AGEMA_signal_5812, SubBytesIns_Inst_Sbox_11_M18}), .b ({new_AGEMA_signal_5695, SubBytesIns_Inst_Sbox_11_M13}), .c ({new_AGEMA_signal_5896, SubBytesIns_Inst_Sbox_11_M22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M23_U1 ( .a ({new_AGEMA_signal_5893, SubBytesIns_Inst_Sbox_11_M19}), .b ({new_AGEMA_signal_10156, new_AGEMA_signal_10155}), .c ({new_AGEMA_signal_5973, SubBytesIns_Inst_Sbox_11_M23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M24_U1 ( .a ({new_AGEMA_signal_5896, SubBytesIns_Inst_Sbox_11_M22}), .b ({new_AGEMA_signal_5973, SubBytesIns_Inst_Sbox_11_M23}), .c ({new_AGEMA_signal_6068, SubBytesIns_Inst_Sbox_11_M24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M27_U1 ( .a ({new_AGEMA_signal_5894, SubBytesIns_Inst_Sbox_11_M20}), .b ({new_AGEMA_signal_5895, SubBytesIns_Inst_Sbox_11_M21}), .c ({new_AGEMA_signal_5975, SubBytesIns_Inst_Sbox_11_M27}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M1_U1 ( .a ({new_AGEMA_signal_5263, SubBytesIns_Inst_Sbox_12_T13}), .b ({new_AGEMA_signal_5261, SubBytesIns_Inst_Sbox_12_T6}), .clk (clk), .r ({Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_5508, SubBytesIns_Inst_Sbox_12_M1}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M2_U1 ( .a ({new_AGEMA_signal_5506, SubBytesIns_Inst_Sbox_12_T23}), .b ({new_AGEMA_signal_5501, SubBytesIns_Inst_Sbox_12_T8}), .clk (clk), .r ({Fresh[219], Fresh[218]}), .c ({new_AGEMA_signal_5699, SubBytesIns_Inst_Sbox_12_M2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M3_U1 ( .a ({new_AGEMA_signal_10158, new_AGEMA_signal_10157}), .b ({new_AGEMA_signal_5508, SubBytesIns_Inst_Sbox_12_M1}), .c ({new_AGEMA_signal_5700, SubBytesIns_Inst_Sbox_12_M3}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M4_U1 ( .a ({new_AGEMA_signal_5266, SubBytesIns_Inst_Sbox_12_T19}), .b ({ciphertext_s1[96], ciphertext_s0[96]}), .clk (clk), .r ({Fresh[221], Fresh[220]}), .c ({new_AGEMA_signal_5509, SubBytesIns_Inst_Sbox_12_M4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M5_U1 ( .a ({new_AGEMA_signal_5509, SubBytesIns_Inst_Sbox_12_M4}), .b ({new_AGEMA_signal_5508, SubBytesIns_Inst_Sbox_12_M1}), .c ({new_AGEMA_signal_5701, SubBytesIns_Inst_Sbox_12_M5}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M6_U1 ( .a ({new_AGEMA_signal_5095, SubBytesIns_Inst_Sbox_12_T3}), .b ({new_AGEMA_signal_5265, SubBytesIns_Inst_Sbox_12_T16}), .clk (clk), .r ({Fresh[223], Fresh[222]}), .c ({new_AGEMA_signal_5510, SubBytesIns_Inst_Sbox_12_M6}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M7_U1 ( .a ({new_AGEMA_signal_5267, SubBytesIns_Inst_Sbox_12_T22}), .b ({new_AGEMA_signal_5262, SubBytesIns_Inst_Sbox_12_T9}), .clk (clk), .r ({Fresh[225], Fresh[224]}), .c ({new_AGEMA_signal_5511, SubBytesIns_Inst_Sbox_12_M7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M8_U1 ( .a ({new_AGEMA_signal_10160, new_AGEMA_signal_10159}), .b ({new_AGEMA_signal_5510, SubBytesIns_Inst_Sbox_12_M6}), .c ({new_AGEMA_signal_5702, SubBytesIns_Inst_Sbox_12_M8}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M9_U1 ( .a ({new_AGEMA_signal_5505, SubBytesIns_Inst_Sbox_12_T20}), .b ({new_AGEMA_signal_5504, SubBytesIns_Inst_Sbox_12_T17}), .clk (clk), .r ({Fresh[227], Fresh[226]}), .c ({new_AGEMA_signal_5703, SubBytesIns_Inst_Sbox_12_M9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M10_U1 ( .a ({new_AGEMA_signal_5703, SubBytesIns_Inst_Sbox_12_M9}), .b ({new_AGEMA_signal_5510, SubBytesIns_Inst_Sbox_12_M6}), .c ({new_AGEMA_signal_5813, SubBytesIns_Inst_Sbox_12_M10}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M11_U1 ( .a ({new_AGEMA_signal_5093, SubBytesIns_Inst_Sbox_12_T1}), .b ({new_AGEMA_signal_5264, SubBytesIns_Inst_Sbox_12_T15}), .clk (clk), .r ({Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_5512, SubBytesIns_Inst_Sbox_12_M11}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M12_U1 ( .a ({new_AGEMA_signal_5096, SubBytesIns_Inst_Sbox_12_T4}), .b ({new_AGEMA_signal_5268, SubBytesIns_Inst_Sbox_12_T27}), .clk (clk), .r ({Fresh[231], Fresh[230]}), .c ({new_AGEMA_signal_5513, SubBytesIns_Inst_Sbox_12_M12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M13_U1 ( .a ({new_AGEMA_signal_5513, SubBytesIns_Inst_Sbox_12_M12}), .b ({new_AGEMA_signal_5512, SubBytesIns_Inst_Sbox_12_M11}), .c ({new_AGEMA_signal_5704, SubBytesIns_Inst_Sbox_12_M13}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M14_U1 ( .a ({new_AGEMA_signal_5094, SubBytesIns_Inst_Sbox_12_T2}), .b ({new_AGEMA_signal_5502, SubBytesIns_Inst_Sbox_12_T10}), .clk (clk), .r ({Fresh[233], Fresh[232]}), .c ({new_AGEMA_signal_5705, SubBytesIns_Inst_Sbox_12_M14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M15_U1 ( .a ({new_AGEMA_signal_5705, SubBytesIns_Inst_Sbox_12_M14}), .b ({new_AGEMA_signal_5512, SubBytesIns_Inst_Sbox_12_M11}), .c ({new_AGEMA_signal_5814, SubBytesIns_Inst_Sbox_12_M15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M16_U1 ( .a ({new_AGEMA_signal_5700, SubBytesIns_Inst_Sbox_12_M3}), .b ({new_AGEMA_signal_5699, SubBytesIns_Inst_Sbox_12_M2}), .c ({new_AGEMA_signal_5815, SubBytesIns_Inst_Sbox_12_M16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M17_U1 ( .a ({new_AGEMA_signal_5701, SubBytesIns_Inst_Sbox_12_M5}), .b ({new_AGEMA_signal_10162, new_AGEMA_signal_10161}), .c ({new_AGEMA_signal_5816, SubBytesIns_Inst_Sbox_12_M17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M18_U1 ( .a ({new_AGEMA_signal_5702, SubBytesIns_Inst_Sbox_12_M8}), .b ({new_AGEMA_signal_5511, SubBytesIns_Inst_Sbox_12_M7}), .c ({new_AGEMA_signal_5817, SubBytesIns_Inst_Sbox_12_M18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M19_U1 ( .a ({new_AGEMA_signal_5813, SubBytesIns_Inst_Sbox_12_M10}), .b ({new_AGEMA_signal_5814, SubBytesIns_Inst_Sbox_12_M15}), .c ({new_AGEMA_signal_5897, SubBytesIns_Inst_Sbox_12_M19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M20_U1 ( .a ({new_AGEMA_signal_5815, SubBytesIns_Inst_Sbox_12_M16}), .b ({new_AGEMA_signal_5704, SubBytesIns_Inst_Sbox_12_M13}), .c ({new_AGEMA_signal_5898, SubBytesIns_Inst_Sbox_12_M20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M21_U1 ( .a ({new_AGEMA_signal_5816, SubBytesIns_Inst_Sbox_12_M17}), .b ({new_AGEMA_signal_5814, SubBytesIns_Inst_Sbox_12_M15}), .c ({new_AGEMA_signal_5899, SubBytesIns_Inst_Sbox_12_M21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M22_U1 ( .a ({new_AGEMA_signal_5817, SubBytesIns_Inst_Sbox_12_M18}), .b ({new_AGEMA_signal_5704, SubBytesIns_Inst_Sbox_12_M13}), .c ({new_AGEMA_signal_5900, SubBytesIns_Inst_Sbox_12_M22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M23_U1 ( .a ({new_AGEMA_signal_5897, SubBytesIns_Inst_Sbox_12_M19}), .b ({new_AGEMA_signal_10164, new_AGEMA_signal_10163}), .c ({new_AGEMA_signal_5977, SubBytesIns_Inst_Sbox_12_M23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M24_U1 ( .a ({new_AGEMA_signal_5900, SubBytesIns_Inst_Sbox_12_M22}), .b ({new_AGEMA_signal_5977, SubBytesIns_Inst_Sbox_12_M23}), .c ({new_AGEMA_signal_6073, SubBytesIns_Inst_Sbox_12_M24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M27_U1 ( .a ({new_AGEMA_signal_5898, SubBytesIns_Inst_Sbox_12_M20}), .b ({new_AGEMA_signal_5899, SubBytesIns_Inst_Sbox_12_M21}), .c ({new_AGEMA_signal_5979, SubBytesIns_Inst_Sbox_12_M27}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M1_U1 ( .a ({new_AGEMA_signal_5271, SubBytesIns_Inst_Sbox_13_T13}), .b ({new_AGEMA_signal_5269, SubBytesIns_Inst_Sbox_13_T6}), .clk (clk), .r ({Fresh[235], Fresh[234]}), .c ({new_AGEMA_signal_5521, SubBytesIns_Inst_Sbox_13_M1}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M2_U1 ( .a ({new_AGEMA_signal_5519, SubBytesIns_Inst_Sbox_13_T23}), .b ({new_AGEMA_signal_5514, SubBytesIns_Inst_Sbox_13_T8}), .clk (clk), .r ({Fresh[237], Fresh[236]}), .c ({new_AGEMA_signal_5708, SubBytesIns_Inst_Sbox_13_M2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M3_U1 ( .a ({new_AGEMA_signal_10166, new_AGEMA_signal_10165}), .b ({new_AGEMA_signal_5521, SubBytesIns_Inst_Sbox_13_M1}), .c ({new_AGEMA_signal_5709, SubBytesIns_Inst_Sbox_13_M3}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M4_U1 ( .a ({new_AGEMA_signal_5274, SubBytesIns_Inst_Sbox_13_T19}), .b ({ciphertext_s1[104], ciphertext_s0[104]}), .clk (clk), .r ({Fresh[239], Fresh[238]}), .c ({new_AGEMA_signal_5522, SubBytesIns_Inst_Sbox_13_M4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M5_U1 ( .a ({new_AGEMA_signal_5522, SubBytesIns_Inst_Sbox_13_M4}), .b ({new_AGEMA_signal_5521, SubBytesIns_Inst_Sbox_13_M1}), .c ({new_AGEMA_signal_5710, SubBytesIns_Inst_Sbox_13_M5}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M6_U1 ( .a ({new_AGEMA_signal_5105, SubBytesIns_Inst_Sbox_13_T3}), .b ({new_AGEMA_signal_5273, SubBytesIns_Inst_Sbox_13_T16}), .clk (clk), .r ({Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_5523, SubBytesIns_Inst_Sbox_13_M6}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M7_U1 ( .a ({new_AGEMA_signal_5275, SubBytesIns_Inst_Sbox_13_T22}), .b ({new_AGEMA_signal_5270, SubBytesIns_Inst_Sbox_13_T9}), .clk (clk), .r ({Fresh[243], Fresh[242]}), .c ({new_AGEMA_signal_5524, SubBytesIns_Inst_Sbox_13_M7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M8_U1 ( .a ({new_AGEMA_signal_10168, new_AGEMA_signal_10167}), .b ({new_AGEMA_signal_5523, SubBytesIns_Inst_Sbox_13_M6}), .c ({new_AGEMA_signal_5711, SubBytesIns_Inst_Sbox_13_M8}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M9_U1 ( .a ({new_AGEMA_signal_5518, SubBytesIns_Inst_Sbox_13_T20}), .b ({new_AGEMA_signal_5517, SubBytesIns_Inst_Sbox_13_T17}), .clk (clk), .r ({Fresh[245], Fresh[244]}), .c ({new_AGEMA_signal_5712, SubBytesIns_Inst_Sbox_13_M9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M10_U1 ( .a ({new_AGEMA_signal_5712, SubBytesIns_Inst_Sbox_13_M9}), .b ({new_AGEMA_signal_5523, SubBytesIns_Inst_Sbox_13_M6}), .c ({new_AGEMA_signal_5818, SubBytesIns_Inst_Sbox_13_M10}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M11_U1 ( .a ({new_AGEMA_signal_5103, SubBytesIns_Inst_Sbox_13_T1}), .b ({new_AGEMA_signal_5272, SubBytesIns_Inst_Sbox_13_T15}), .clk (clk), .r ({Fresh[247], Fresh[246]}), .c ({new_AGEMA_signal_5525, SubBytesIns_Inst_Sbox_13_M11}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M12_U1 ( .a ({new_AGEMA_signal_5106, SubBytesIns_Inst_Sbox_13_T4}), .b ({new_AGEMA_signal_5276, SubBytesIns_Inst_Sbox_13_T27}), .clk (clk), .r ({Fresh[249], Fresh[248]}), .c ({new_AGEMA_signal_5526, SubBytesIns_Inst_Sbox_13_M12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M13_U1 ( .a ({new_AGEMA_signal_5526, SubBytesIns_Inst_Sbox_13_M12}), .b ({new_AGEMA_signal_5525, SubBytesIns_Inst_Sbox_13_M11}), .c ({new_AGEMA_signal_5713, SubBytesIns_Inst_Sbox_13_M13}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M14_U1 ( .a ({new_AGEMA_signal_5104, SubBytesIns_Inst_Sbox_13_T2}), .b ({new_AGEMA_signal_5515, SubBytesIns_Inst_Sbox_13_T10}), .clk (clk), .r ({Fresh[251], Fresh[250]}), .c ({new_AGEMA_signal_5714, SubBytesIns_Inst_Sbox_13_M14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M15_U1 ( .a ({new_AGEMA_signal_5714, SubBytesIns_Inst_Sbox_13_M14}), .b ({new_AGEMA_signal_5525, SubBytesIns_Inst_Sbox_13_M11}), .c ({new_AGEMA_signal_5819, SubBytesIns_Inst_Sbox_13_M15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M16_U1 ( .a ({new_AGEMA_signal_5709, SubBytesIns_Inst_Sbox_13_M3}), .b ({new_AGEMA_signal_5708, SubBytesIns_Inst_Sbox_13_M2}), .c ({new_AGEMA_signal_5820, SubBytesIns_Inst_Sbox_13_M16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M17_U1 ( .a ({new_AGEMA_signal_5710, SubBytesIns_Inst_Sbox_13_M5}), .b ({new_AGEMA_signal_10170, new_AGEMA_signal_10169}), .c ({new_AGEMA_signal_5821, SubBytesIns_Inst_Sbox_13_M17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M18_U1 ( .a ({new_AGEMA_signal_5711, SubBytesIns_Inst_Sbox_13_M8}), .b ({new_AGEMA_signal_5524, SubBytesIns_Inst_Sbox_13_M7}), .c ({new_AGEMA_signal_5822, SubBytesIns_Inst_Sbox_13_M18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M19_U1 ( .a ({new_AGEMA_signal_5818, SubBytesIns_Inst_Sbox_13_M10}), .b ({new_AGEMA_signal_5819, SubBytesIns_Inst_Sbox_13_M15}), .c ({new_AGEMA_signal_5901, SubBytesIns_Inst_Sbox_13_M19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M20_U1 ( .a ({new_AGEMA_signal_5820, SubBytesIns_Inst_Sbox_13_M16}), .b ({new_AGEMA_signal_5713, SubBytesIns_Inst_Sbox_13_M13}), .c ({new_AGEMA_signal_5902, SubBytesIns_Inst_Sbox_13_M20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M21_U1 ( .a ({new_AGEMA_signal_5821, SubBytesIns_Inst_Sbox_13_M17}), .b ({new_AGEMA_signal_5819, SubBytesIns_Inst_Sbox_13_M15}), .c ({new_AGEMA_signal_5903, SubBytesIns_Inst_Sbox_13_M21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M22_U1 ( .a ({new_AGEMA_signal_5822, SubBytesIns_Inst_Sbox_13_M18}), .b ({new_AGEMA_signal_5713, SubBytesIns_Inst_Sbox_13_M13}), .c ({new_AGEMA_signal_5904, SubBytesIns_Inst_Sbox_13_M22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M23_U1 ( .a ({new_AGEMA_signal_5901, SubBytesIns_Inst_Sbox_13_M19}), .b ({new_AGEMA_signal_10172, new_AGEMA_signal_10171}), .c ({new_AGEMA_signal_5981, SubBytesIns_Inst_Sbox_13_M23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M24_U1 ( .a ({new_AGEMA_signal_5904, SubBytesIns_Inst_Sbox_13_M22}), .b ({new_AGEMA_signal_5981, SubBytesIns_Inst_Sbox_13_M23}), .c ({new_AGEMA_signal_6078, SubBytesIns_Inst_Sbox_13_M24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M27_U1 ( .a ({new_AGEMA_signal_5902, SubBytesIns_Inst_Sbox_13_M20}), .b ({new_AGEMA_signal_5903, SubBytesIns_Inst_Sbox_13_M21}), .c ({new_AGEMA_signal_5983, SubBytesIns_Inst_Sbox_13_M27}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M1_U1 ( .a ({new_AGEMA_signal_5279, SubBytesIns_Inst_Sbox_14_T13}), .b ({new_AGEMA_signal_5277, SubBytesIns_Inst_Sbox_14_T6}), .clk (clk), .r ({Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_5534, SubBytesIns_Inst_Sbox_14_M1}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M2_U1 ( .a ({new_AGEMA_signal_5532, SubBytesIns_Inst_Sbox_14_T23}), .b ({new_AGEMA_signal_5527, SubBytesIns_Inst_Sbox_14_T8}), .clk (clk), .r ({Fresh[255], Fresh[254]}), .c ({new_AGEMA_signal_5717, SubBytesIns_Inst_Sbox_14_M2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M3_U1 ( .a ({new_AGEMA_signal_10174, new_AGEMA_signal_10173}), .b ({new_AGEMA_signal_5534, SubBytesIns_Inst_Sbox_14_M1}), .c ({new_AGEMA_signal_5718, SubBytesIns_Inst_Sbox_14_M3}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M4_U1 ( .a ({new_AGEMA_signal_5282, SubBytesIns_Inst_Sbox_14_T19}), .b ({ciphertext_s1[112], ciphertext_s0[112]}), .clk (clk), .r ({Fresh[257], Fresh[256]}), .c ({new_AGEMA_signal_5535, SubBytesIns_Inst_Sbox_14_M4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M5_U1 ( .a ({new_AGEMA_signal_5535, SubBytesIns_Inst_Sbox_14_M4}), .b ({new_AGEMA_signal_5534, SubBytesIns_Inst_Sbox_14_M1}), .c ({new_AGEMA_signal_5719, SubBytesIns_Inst_Sbox_14_M5}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M6_U1 ( .a ({new_AGEMA_signal_5115, SubBytesIns_Inst_Sbox_14_T3}), .b ({new_AGEMA_signal_5281, SubBytesIns_Inst_Sbox_14_T16}), .clk (clk), .r ({Fresh[259], Fresh[258]}), .c ({new_AGEMA_signal_5536, SubBytesIns_Inst_Sbox_14_M6}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M7_U1 ( .a ({new_AGEMA_signal_5283, SubBytesIns_Inst_Sbox_14_T22}), .b ({new_AGEMA_signal_5278, SubBytesIns_Inst_Sbox_14_T9}), .clk (clk), .r ({Fresh[261], Fresh[260]}), .c ({new_AGEMA_signal_5537, SubBytesIns_Inst_Sbox_14_M7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M8_U1 ( .a ({new_AGEMA_signal_10176, new_AGEMA_signal_10175}), .b ({new_AGEMA_signal_5536, SubBytesIns_Inst_Sbox_14_M6}), .c ({new_AGEMA_signal_5720, SubBytesIns_Inst_Sbox_14_M8}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M9_U1 ( .a ({new_AGEMA_signal_5531, SubBytesIns_Inst_Sbox_14_T20}), .b ({new_AGEMA_signal_5530, SubBytesIns_Inst_Sbox_14_T17}), .clk (clk), .r ({Fresh[263], Fresh[262]}), .c ({new_AGEMA_signal_5721, SubBytesIns_Inst_Sbox_14_M9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M10_U1 ( .a ({new_AGEMA_signal_5721, SubBytesIns_Inst_Sbox_14_M9}), .b ({new_AGEMA_signal_5536, SubBytesIns_Inst_Sbox_14_M6}), .c ({new_AGEMA_signal_5823, SubBytesIns_Inst_Sbox_14_M10}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M11_U1 ( .a ({new_AGEMA_signal_5113, SubBytesIns_Inst_Sbox_14_T1}), .b ({new_AGEMA_signal_5280, SubBytesIns_Inst_Sbox_14_T15}), .clk (clk), .r ({Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_5538, SubBytesIns_Inst_Sbox_14_M11}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M12_U1 ( .a ({new_AGEMA_signal_5116, SubBytesIns_Inst_Sbox_14_T4}), .b ({new_AGEMA_signal_5284, SubBytesIns_Inst_Sbox_14_T27}), .clk (clk), .r ({Fresh[267], Fresh[266]}), .c ({new_AGEMA_signal_5539, SubBytesIns_Inst_Sbox_14_M12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M13_U1 ( .a ({new_AGEMA_signal_5539, SubBytesIns_Inst_Sbox_14_M12}), .b ({new_AGEMA_signal_5538, SubBytesIns_Inst_Sbox_14_M11}), .c ({new_AGEMA_signal_5722, SubBytesIns_Inst_Sbox_14_M13}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M14_U1 ( .a ({new_AGEMA_signal_5114, SubBytesIns_Inst_Sbox_14_T2}), .b ({new_AGEMA_signal_5528, SubBytesIns_Inst_Sbox_14_T10}), .clk (clk), .r ({Fresh[269], Fresh[268]}), .c ({new_AGEMA_signal_5723, SubBytesIns_Inst_Sbox_14_M14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M15_U1 ( .a ({new_AGEMA_signal_5723, SubBytesIns_Inst_Sbox_14_M14}), .b ({new_AGEMA_signal_5538, SubBytesIns_Inst_Sbox_14_M11}), .c ({new_AGEMA_signal_5824, SubBytesIns_Inst_Sbox_14_M15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M16_U1 ( .a ({new_AGEMA_signal_5718, SubBytesIns_Inst_Sbox_14_M3}), .b ({new_AGEMA_signal_5717, SubBytesIns_Inst_Sbox_14_M2}), .c ({new_AGEMA_signal_5825, SubBytesIns_Inst_Sbox_14_M16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M17_U1 ( .a ({new_AGEMA_signal_5719, SubBytesIns_Inst_Sbox_14_M5}), .b ({new_AGEMA_signal_10178, new_AGEMA_signal_10177}), .c ({new_AGEMA_signal_5826, SubBytesIns_Inst_Sbox_14_M17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M18_U1 ( .a ({new_AGEMA_signal_5720, SubBytesIns_Inst_Sbox_14_M8}), .b ({new_AGEMA_signal_5537, SubBytesIns_Inst_Sbox_14_M7}), .c ({new_AGEMA_signal_5827, SubBytesIns_Inst_Sbox_14_M18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M19_U1 ( .a ({new_AGEMA_signal_5823, SubBytesIns_Inst_Sbox_14_M10}), .b ({new_AGEMA_signal_5824, SubBytesIns_Inst_Sbox_14_M15}), .c ({new_AGEMA_signal_5905, SubBytesIns_Inst_Sbox_14_M19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M20_U1 ( .a ({new_AGEMA_signal_5825, SubBytesIns_Inst_Sbox_14_M16}), .b ({new_AGEMA_signal_5722, SubBytesIns_Inst_Sbox_14_M13}), .c ({new_AGEMA_signal_5906, SubBytesIns_Inst_Sbox_14_M20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M21_U1 ( .a ({new_AGEMA_signal_5826, SubBytesIns_Inst_Sbox_14_M17}), .b ({new_AGEMA_signal_5824, SubBytesIns_Inst_Sbox_14_M15}), .c ({new_AGEMA_signal_5907, SubBytesIns_Inst_Sbox_14_M21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M22_U1 ( .a ({new_AGEMA_signal_5827, SubBytesIns_Inst_Sbox_14_M18}), .b ({new_AGEMA_signal_5722, SubBytesIns_Inst_Sbox_14_M13}), .c ({new_AGEMA_signal_5908, SubBytesIns_Inst_Sbox_14_M22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M23_U1 ( .a ({new_AGEMA_signal_5905, SubBytesIns_Inst_Sbox_14_M19}), .b ({new_AGEMA_signal_10180, new_AGEMA_signal_10179}), .c ({new_AGEMA_signal_5985, SubBytesIns_Inst_Sbox_14_M23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M24_U1 ( .a ({new_AGEMA_signal_5908, SubBytesIns_Inst_Sbox_14_M22}), .b ({new_AGEMA_signal_5985, SubBytesIns_Inst_Sbox_14_M23}), .c ({new_AGEMA_signal_6083, SubBytesIns_Inst_Sbox_14_M24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M27_U1 ( .a ({new_AGEMA_signal_5906, SubBytesIns_Inst_Sbox_14_M20}), .b ({new_AGEMA_signal_5907, SubBytesIns_Inst_Sbox_14_M21}), .c ({new_AGEMA_signal_5987, SubBytesIns_Inst_Sbox_14_M27}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M1_U1 ( .a ({new_AGEMA_signal_5287, SubBytesIns_Inst_Sbox_15_T13}), .b ({new_AGEMA_signal_5285, SubBytesIns_Inst_Sbox_15_T6}), .clk (clk), .r ({Fresh[271], Fresh[270]}), .c ({new_AGEMA_signal_5547, SubBytesIns_Inst_Sbox_15_M1}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M2_U1 ( .a ({new_AGEMA_signal_5545, SubBytesIns_Inst_Sbox_15_T23}), .b ({new_AGEMA_signal_5540, SubBytesIns_Inst_Sbox_15_T8}), .clk (clk), .r ({Fresh[273], Fresh[272]}), .c ({new_AGEMA_signal_5726, SubBytesIns_Inst_Sbox_15_M2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M3_U1 ( .a ({new_AGEMA_signal_10182, new_AGEMA_signal_10181}), .b ({new_AGEMA_signal_5547, SubBytesIns_Inst_Sbox_15_M1}), .c ({new_AGEMA_signal_5727, SubBytesIns_Inst_Sbox_15_M3}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M4_U1 ( .a ({new_AGEMA_signal_5290, SubBytesIns_Inst_Sbox_15_T19}), .b ({ciphertext_s1[120], ciphertext_s0[120]}), .clk (clk), .r ({Fresh[275], Fresh[274]}), .c ({new_AGEMA_signal_5548, SubBytesIns_Inst_Sbox_15_M4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M5_U1 ( .a ({new_AGEMA_signal_5548, SubBytesIns_Inst_Sbox_15_M4}), .b ({new_AGEMA_signal_5547, SubBytesIns_Inst_Sbox_15_M1}), .c ({new_AGEMA_signal_5728, SubBytesIns_Inst_Sbox_15_M5}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M6_U1 ( .a ({new_AGEMA_signal_5125, SubBytesIns_Inst_Sbox_15_T3}), .b ({new_AGEMA_signal_5289, SubBytesIns_Inst_Sbox_15_T16}), .clk (clk), .r ({Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_5549, SubBytesIns_Inst_Sbox_15_M6}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M7_U1 ( .a ({new_AGEMA_signal_5291, SubBytesIns_Inst_Sbox_15_T22}), .b ({new_AGEMA_signal_5286, SubBytesIns_Inst_Sbox_15_T9}), .clk (clk), .r ({Fresh[279], Fresh[278]}), .c ({new_AGEMA_signal_5550, SubBytesIns_Inst_Sbox_15_M7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M8_U1 ( .a ({new_AGEMA_signal_10184, new_AGEMA_signal_10183}), .b ({new_AGEMA_signal_5549, SubBytesIns_Inst_Sbox_15_M6}), .c ({new_AGEMA_signal_5729, SubBytesIns_Inst_Sbox_15_M8}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M9_U1 ( .a ({new_AGEMA_signal_5544, SubBytesIns_Inst_Sbox_15_T20}), .b ({new_AGEMA_signal_5543, SubBytesIns_Inst_Sbox_15_T17}), .clk (clk), .r ({Fresh[281], Fresh[280]}), .c ({new_AGEMA_signal_5730, SubBytesIns_Inst_Sbox_15_M9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M10_U1 ( .a ({new_AGEMA_signal_5730, SubBytesIns_Inst_Sbox_15_M9}), .b ({new_AGEMA_signal_5549, SubBytesIns_Inst_Sbox_15_M6}), .c ({new_AGEMA_signal_5828, SubBytesIns_Inst_Sbox_15_M10}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M11_U1 ( .a ({new_AGEMA_signal_5123, SubBytesIns_Inst_Sbox_15_T1}), .b ({new_AGEMA_signal_5288, SubBytesIns_Inst_Sbox_15_T15}), .clk (clk), .r ({Fresh[283], Fresh[282]}), .c ({new_AGEMA_signal_5551, SubBytesIns_Inst_Sbox_15_M11}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M12_U1 ( .a ({new_AGEMA_signal_5126, SubBytesIns_Inst_Sbox_15_T4}), .b ({new_AGEMA_signal_5292, SubBytesIns_Inst_Sbox_15_T27}), .clk (clk), .r ({Fresh[285], Fresh[284]}), .c ({new_AGEMA_signal_5552, SubBytesIns_Inst_Sbox_15_M12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M13_U1 ( .a ({new_AGEMA_signal_5552, SubBytesIns_Inst_Sbox_15_M12}), .b ({new_AGEMA_signal_5551, SubBytesIns_Inst_Sbox_15_M11}), .c ({new_AGEMA_signal_5731, SubBytesIns_Inst_Sbox_15_M13}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M14_U1 ( .a ({new_AGEMA_signal_5124, SubBytesIns_Inst_Sbox_15_T2}), .b ({new_AGEMA_signal_5541, SubBytesIns_Inst_Sbox_15_T10}), .clk (clk), .r ({Fresh[287], Fresh[286]}), .c ({new_AGEMA_signal_5732, SubBytesIns_Inst_Sbox_15_M14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M15_U1 ( .a ({new_AGEMA_signal_5732, SubBytesIns_Inst_Sbox_15_M14}), .b ({new_AGEMA_signal_5551, SubBytesIns_Inst_Sbox_15_M11}), .c ({new_AGEMA_signal_5829, SubBytesIns_Inst_Sbox_15_M15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M16_U1 ( .a ({new_AGEMA_signal_5727, SubBytesIns_Inst_Sbox_15_M3}), .b ({new_AGEMA_signal_5726, SubBytesIns_Inst_Sbox_15_M2}), .c ({new_AGEMA_signal_5830, SubBytesIns_Inst_Sbox_15_M16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M17_U1 ( .a ({new_AGEMA_signal_5728, SubBytesIns_Inst_Sbox_15_M5}), .b ({new_AGEMA_signal_10186, new_AGEMA_signal_10185}), .c ({new_AGEMA_signal_5831, SubBytesIns_Inst_Sbox_15_M17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M18_U1 ( .a ({new_AGEMA_signal_5729, SubBytesIns_Inst_Sbox_15_M8}), .b ({new_AGEMA_signal_5550, SubBytesIns_Inst_Sbox_15_M7}), .c ({new_AGEMA_signal_5832, SubBytesIns_Inst_Sbox_15_M18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M19_U1 ( .a ({new_AGEMA_signal_5828, SubBytesIns_Inst_Sbox_15_M10}), .b ({new_AGEMA_signal_5829, SubBytesIns_Inst_Sbox_15_M15}), .c ({new_AGEMA_signal_5909, SubBytesIns_Inst_Sbox_15_M19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M20_U1 ( .a ({new_AGEMA_signal_5830, SubBytesIns_Inst_Sbox_15_M16}), .b ({new_AGEMA_signal_5731, SubBytesIns_Inst_Sbox_15_M13}), .c ({new_AGEMA_signal_5910, SubBytesIns_Inst_Sbox_15_M20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M21_U1 ( .a ({new_AGEMA_signal_5831, SubBytesIns_Inst_Sbox_15_M17}), .b ({new_AGEMA_signal_5829, SubBytesIns_Inst_Sbox_15_M15}), .c ({new_AGEMA_signal_5911, SubBytesIns_Inst_Sbox_15_M21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M22_U1 ( .a ({new_AGEMA_signal_5832, SubBytesIns_Inst_Sbox_15_M18}), .b ({new_AGEMA_signal_5731, SubBytesIns_Inst_Sbox_15_M13}), .c ({new_AGEMA_signal_5912, SubBytesIns_Inst_Sbox_15_M22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M23_U1 ( .a ({new_AGEMA_signal_5909, SubBytesIns_Inst_Sbox_15_M19}), .b ({new_AGEMA_signal_10188, new_AGEMA_signal_10187}), .c ({new_AGEMA_signal_5989, SubBytesIns_Inst_Sbox_15_M23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M24_U1 ( .a ({new_AGEMA_signal_5912, SubBytesIns_Inst_Sbox_15_M22}), .b ({new_AGEMA_signal_5989, SubBytesIns_Inst_Sbox_15_M23}), .c ({new_AGEMA_signal_6088, SubBytesIns_Inst_Sbox_15_M24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M27_U1 ( .a ({new_AGEMA_signal_5910, SubBytesIns_Inst_Sbox_15_M20}), .b ({new_AGEMA_signal_5911, SubBytesIns_Inst_Sbox_15_M21}), .c ({new_AGEMA_signal_5991, SubBytesIns_Inst_Sbox_15_M27}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M1_U1 ( .a ({new_AGEMA_signal_5135, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13}), .b ({new_AGEMA_signal_5133, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}), .clk (clk), .r ({Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_5300, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M2_U1 ( .a ({new_AGEMA_signal_5298, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23}), .b ({new_AGEMA_signal_5293, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8}), .clk (clk), .r ({Fresh[291], Fresh[290]}), .c ({new_AGEMA_signal_5555, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M3_U1 ( .a ({new_AGEMA_signal_10190, new_AGEMA_signal_10189}), .b ({new_AGEMA_signal_5300, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_5556, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M3}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M4_U1 ( .a ({new_AGEMA_signal_5138, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19}), .b ({new_AGEMA_signal_4655, RoundKey[16]}), .clk (clk), .r ({Fresh[293], Fresh[292]}), .c ({new_AGEMA_signal_5301, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M5_U1 ( .a ({new_AGEMA_signal_5301, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M4}), .b ({new_AGEMA_signal_5300, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_5557, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M5}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M6_U1 ( .a ({new_AGEMA_signal_4935, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_5137, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16}), .clk (clk), .r ({Fresh[295], Fresh[294]}), .c ({new_AGEMA_signal_5302, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M7_U1 ( .a ({new_AGEMA_signal_5139, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22}), .b ({new_AGEMA_signal_5134, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9}), .clk (clk), .r ({Fresh[297], Fresh[296]}), .c ({new_AGEMA_signal_5303, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M8_U1 ( .a ({new_AGEMA_signal_10192, new_AGEMA_signal_10191}), .b ({new_AGEMA_signal_5302, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_5558, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M8}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M9_U1 ( .a ({new_AGEMA_signal_5297, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_5296, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17}), .clk (clk), .r ({Fresh[299], Fresh[298]}), .c ({new_AGEMA_signal_5559, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M10_U1 ( .a ({new_AGEMA_signal_5559, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M9}), .b ({new_AGEMA_signal_5302, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_5733, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M10}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M11_U1 ( .a ({new_AGEMA_signal_4933, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_5136, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15}), .clk (clk), .r ({Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_5304, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M12_U1 ( .a ({new_AGEMA_signal_4936, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4}), .b ({new_AGEMA_signal_5140, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27}), .clk (clk), .r ({Fresh[303], Fresh[302]}), .c ({new_AGEMA_signal_5305, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M13_U1 ( .a ({new_AGEMA_signal_5305, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M12}), .b ({new_AGEMA_signal_5304, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_5560, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M14_U1 ( .a ({new_AGEMA_signal_4934, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_5294, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10}), .clk (clk), .r ({Fresh[305], Fresh[304]}), .c ({new_AGEMA_signal_5561, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M15_U1 ( .a ({new_AGEMA_signal_5561, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M14}), .b ({new_AGEMA_signal_5304, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_5734, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M16_U1 ( .a ({new_AGEMA_signal_5556, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M3}), .b ({new_AGEMA_signal_5555, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M2}), .c ({new_AGEMA_signal_5735, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M17_U1 ( .a ({new_AGEMA_signal_5557, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M5}), .b ({new_AGEMA_signal_10194, new_AGEMA_signal_10193}), .c ({new_AGEMA_signal_5736, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M18_U1 ( .a ({new_AGEMA_signal_5558, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M8}), .b ({new_AGEMA_signal_5303, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M7}), .c ({new_AGEMA_signal_5737, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M19_U1 ( .a ({new_AGEMA_signal_5733, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M10}), .b ({new_AGEMA_signal_5734, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_5833, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M20_U1 ( .a ({new_AGEMA_signal_5735, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M16}), .b ({new_AGEMA_signal_5560, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_5834, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M21_U1 ( .a ({new_AGEMA_signal_5736, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M17}), .b ({new_AGEMA_signal_5734, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_5835, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M22_U1 ( .a ({new_AGEMA_signal_5737, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M18}), .b ({new_AGEMA_signal_5560, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_5836, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M23_U1 ( .a ({new_AGEMA_signal_5833, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M19}), .b ({new_AGEMA_signal_10196, new_AGEMA_signal_10195}), .c ({new_AGEMA_signal_5913, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M24_U1 ( .a ({new_AGEMA_signal_5836, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_5913, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23}), .c ({new_AGEMA_signal_5993, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M27_U1 ( .a ({new_AGEMA_signal_5834, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_5835, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21}), .c ({new_AGEMA_signal_5915, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M1_U1 ( .a ({new_AGEMA_signal_5143, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13}), .b ({new_AGEMA_signal_5141, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}), .clk (clk), .r ({Fresh[307], Fresh[306]}), .c ({new_AGEMA_signal_5313, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M2_U1 ( .a ({new_AGEMA_signal_5311, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23}), .b ({new_AGEMA_signal_5306, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8}), .clk (clk), .r ({Fresh[309], Fresh[308]}), .c ({new_AGEMA_signal_5564, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M3_U1 ( .a ({new_AGEMA_signal_10198, new_AGEMA_signal_10197}), .b ({new_AGEMA_signal_5313, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_5565, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M3}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M4_U1 ( .a ({new_AGEMA_signal_5146, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19}), .b ({new_AGEMA_signal_4898, RoundKey[8]}), .clk (clk), .r ({Fresh[311], Fresh[310]}), .c ({new_AGEMA_signal_5314, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M5_U1 ( .a ({new_AGEMA_signal_5314, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M4}), .b ({new_AGEMA_signal_5313, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_5566, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M5}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M6_U1 ( .a ({new_AGEMA_signal_4945, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_5145, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16}), .clk (clk), .r ({Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_5315, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M7_U1 ( .a ({new_AGEMA_signal_5147, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22}), .b ({new_AGEMA_signal_5142, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9}), .clk (clk), .r ({Fresh[315], Fresh[314]}), .c ({new_AGEMA_signal_5316, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M8_U1 ( .a ({new_AGEMA_signal_10200, new_AGEMA_signal_10199}), .b ({new_AGEMA_signal_5315, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_5567, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M8}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M9_U1 ( .a ({new_AGEMA_signal_5310, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_5309, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17}), .clk (clk), .r ({Fresh[317], Fresh[316]}), .c ({new_AGEMA_signal_5568, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M10_U1 ( .a ({new_AGEMA_signal_5568, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M9}), .b ({new_AGEMA_signal_5315, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_5738, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M10}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M11_U1 ( .a ({new_AGEMA_signal_4943, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_5144, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15}), .clk (clk), .r ({Fresh[319], Fresh[318]}), .c ({new_AGEMA_signal_5317, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M12_U1 ( .a ({new_AGEMA_signal_4946, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4}), .b ({new_AGEMA_signal_5148, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27}), .clk (clk), .r ({Fresh[321], Fresh[320]}), .c ({new_AGEMA_signal_5318, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M13_U1 ( .a ({new_AGEMA_signal_5318, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M12}), .b ({new_AGEMA_signal_5317, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_5569, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M14_U1 ( .a ({new_AGEMA_signal_4944, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_5307, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10}), .clk (clk), .r ({Fresh[323], Fresh[322]}), .c ({new_AGEMA_signal_5570, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M15_U1 ( .a ({new_AGEMA_signal_5570, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M14}), .b ({new_AGEMA_signal_5317, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_5739, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M16_U1 ( .a ({new_AGEMA_signal_5565, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M3}), .b ({new_AGEMA_signal_5564, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M2}), .c ({new_AGEMA_signal_5740, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M17_U1 ( .a ({new_AGEMA_signal_5566, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M5}), .b ({new_AGEMA_signal_10202, new_AGEMA_signal_10201}), .c ({new_AGEMA_signal_5741, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M18_U1 ( .a ({new_AGEMA_signal_5567, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M8}), .b ({new_AGEMA_signal_5316, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M7}), .c ({new_AGEMA_signal_5742, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M19_U1 ( .a ({new_AGEMA_signal_5738, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M10}), .b ({new_AGEMA_signal_5739, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_5837, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M20_U1 ( .a ({new_AGEMA_signal_5740, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M16}), .b ({new_AGEMA_signal_5569, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_5838, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M21_U1 ( .a ({new_AGEMA_signal_5741, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M17}), .b ({new_AGEMA_signal_5739, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_5839, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M22_U1 ( .a ({new_AGEMA_signal_5742, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M18}), .b ({new_AGEMA_signal_5569, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_5840, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M23_U1 ( .a ({new_AGEMA_signal_5837, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M19}), .b ({new_AGEMA_signal_10204, new_AGEMA_signal_10203}), .c ({new_AGEMA_signal_5917, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M24_U1 ( .a ({new_AGEMA_signal_5840, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_5917, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23}), .c ({new_AGEMA_signal_5998, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M27_U1 ( .a ({new_AGEMA_signal_5838, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_5839, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21}), .c ({new_AGEMA_signal_5919, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M1_U1 ( .a ({new_AGEMA_signal_5151, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13}), .b ({new_AGEMA_signal_5149, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}), .clk (clk), .r ({Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_5326, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M2_U1 ( .a ({new_AGEMA_signal_5324, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23}), .b ({new_AGEMA_signal_5319, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8}), .clk (clk), .r ({Fresh[327], Fresh[326]}), .c ({new_AGEMA_signal_5573, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M3_U1 ( .a ({new_AGEMA_signal_10206, new_AGEMA_signal_10205}), .b ({new_AGEMA_signal_5326, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_5574, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M3}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M4_U1 ( .a ({new_AGEMA_signal_5154, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19}), .b ({new_AGEMA_signal_4550, RoundKey[0]}), .clk (clk), .r ({Fresh[329], Fresh[328]}), .c ({new_AGEMA_signal_5327, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M5_U1 ( .a ({new_AGEMA_signal_5327, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M4}), .b ({new_AGEMA_signal_5326, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_5575, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M5}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M6_U1 ( .a ({new_AGEMA_signal_4955, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_5153, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16}), .clk (clk), .r ({Fresh[331], Fresh[330]}), .c ({new_AGEMA_signal_5328, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M7_U1 ( .a ({new_AGEMA_signal_5155, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22}), .b ({new_AGEMA_signal_5150, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9}), .clk (clk), .r ({Fresh[333], Fresh[332]}), .c ({new_AGEMA_signal_5329, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M8_U1 ( .a ({new_AGEMA_signal_10208, new_AGEMA_signal_10207}), .b ({new_AGEMA_signal_5328, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_5576, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M8}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M9_U1 ( .a ({new_AGEMA_signal_5323, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_5322, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17}), .clk (clk), .r ({Fresh[335], Fresh[334]}), .c ({new_AGEMA_signal_5577, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M10_U1 ( .a ({new_AGEMA_signal_5577, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M9}), .b ({new_AGEMA_signal_5328, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_5743, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M10}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M11_U1 ( .a ({new_AGEMA_signal_4953, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5152, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15}), .clk (clk), .r ({Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_5330, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M12_U1 ( .a ({new_AGEMA_signal_4956, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4}), .b ({new_AGEMA_signal_5156, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27}), .clk (clk), .r ({Fresh[339], Fresh[338]}), .c ({new_AGEMA_signal_5331, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M13_U1 ( .a ({new_AGEMA_signal_5331, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M12}), .b ({new_AGEMA_signal_5330, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_5578, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M14_U1 ( .a ({new_AGEMA_signal_4954, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_5320, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10}), .clk (clk), .r ({Fresh[341], Fresh[340]}), .c ({new_AGEMA_signal_5579, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M15_U1 ( .a ({new_AGEMA_signal_5579, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M14}), .b ({new_AGEMA_signal_5330, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_5744, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M16_U1 ( .a ({new_AGEMA_signal_5574, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M3}), .b ({new_AGEMA_signal_5573, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M2}), .c ({new_AGEMA_signal_5745, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M17_U1 ( .a ({new_AGEMA_signal_5575, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M5}), .b ({new_AGEMA_signal_10210, new_AGEMA_signal_10209}), .c ({new_AGEMA_signal_5746, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M18_U1 ( .a ({new_AGEMA_signal_5576, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M8}), .b ({new_AGEMA_signal_5329, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M7}), .c ({new_AGEMA_signal_5747, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M19_U1 ( .a ({new_AGEMA_signal_5743, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M10}), .b ({new_AGEMA_signal_5744, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_5841, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M20_U1 ( .a ({new_AGEMA_signal_5745, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M16}), .b ({new_AGEMA_signal_5578, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_5842, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M21_U1 ( .a ({new_AGEMA_signal_5746, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M17}), .b ({new_AGEMA_signal_5744, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_5843, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M22_U1 ( .a ({new_AGEMA_signal_5747, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M18}), .b ({new_AGEMA_signal_5578, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_5844, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M23_U1 ( .a ({new_AGEMA_signal_5841, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M19}), .b ({new_AGEMA_signal_10212, new_AGEMA_signal_10211}), .c ({new_AGEMA_signal_5921, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M24_U1 ( .a ({new_AGEMA_signal_5844, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_5921, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23}), .c ({new_AGEMA_signal_6003, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M27_U1 ( .a ({new_AGEMA_signal_5842, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_5843, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21}), .c ({new_AGEMA_signal_5923, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M1_U1 ( .a ({new_AGEMA_signal_5159, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13}), .b ({new_AGEMA_signal_5157, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}), .clk (clk), .r ({Fresh[343], Fresh[342]}), .c ({new_AGEMA_signal_5339, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M2_U1 ( .a ({new_AGEMA_signal_5337, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23}), .b ({new_AGEMA_signal_5332, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8}), .clk (clk), .r ({Fresh[345], Fresh[344]}), .c ({new_AGEMA_signal_5582, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M3_U1 ( .a ({new_AGEMA_signal_10214, new_AGEMA_signal_10213}), .b ({new_AGEMA_signal_5339, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_5583, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M3}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M4_U1 ( .a ({new_AGEMA_signal_5162, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19}), .b ({new_AGEMA_signal_4682, RoundKey[24]}), .clk (clk), .r ({Fresh[347], Fresh[346]}), .c ({new_AGEMA_signal_5340, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M5_U1 ( .a ({new_AGEMA_signal_5340, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M4}), .b ({new_AGEMA_signal_5339, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_5584, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M5}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M6_U1 ( .a ({new_AGEMA_signal_4965, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_5161, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16}), .clk (clk), .r ({Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_5341, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M7_U1 ( .a ({new_AGEMA_signal_5163, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22}), .b ({new_AGEMA_signal_5158, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9}), .clk (clk), .r ({Fresh[351], Fresh[350]}), .c ({new_AGEMA_signal_5342, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M8_U1 ( .a ({new_AGEMA_signal_10216, new_AGEMA_signal_10215}), .b ({new_AGEMA_signal_5341, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_5585, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M8}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M9_U1 ( .a ({new_AGEMA_signal_5336, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_5335, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17}), .clk (clk), .r ({Fresh[353], Fresh[352]}), .c ({new_AGEMA_signal_5586, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M10_U1 ( .a ({new_AGEMA_signal_5586, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M9}), .b ({new_AGEMA_signal_5341, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_5748, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M10}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M11_U1 ( .a ({new_AGEMA_signal_4963, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5160, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15}), .clk (clk), .r ({Fresh[355], Fresh[354]}), .c ({new_AGEMA_signal_5343, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M12_U1 ( .a ({new_AGEMA_signal_4966, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4}), .b ({new_AGEMA_signal_5164, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27}), .clk (clk), .r ({Fresh[357], Fresh[356]}), .c ({new_AGEMA_signal_5344, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M13_U1 ( .a ({new_AGEMA_signal_5344, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M12}), .b ({new_AGEMA_signal_5343, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_5587, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M14_U1 ( .a ({new_AGEMA_signal_4964, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_5333, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10}), .clk (clk), .r ({Fresh[359], Fresh[358]}), .c ({new_AGEMA_signal_5588, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M15_U1 ( .a ({new_AGEMA_signal_5588, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M14}), .b ({new_AGEMA_signal_5343, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_5749, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M16_U1 ( .a ({new_AGEMA_signal_5583, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M3}), .b ({new_AGEMA_signal_5582, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M2}), .c ({new_AGEMA_signal_5750, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M17_U1 ( .a ({new_AGEMA_signal_5584, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M5}), .b ({new_AGEMA_signal_10218, new_AGEMA_signal_10217}), .c ({new_AGEMA_signal_5751, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M18_U1 ( .a ({new_AGEMA_signal_5585, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M8}), .b ({new_AGEMA_signal_5342, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M7}), .c ({new_AGEMA_signal_5752, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M19_U1 ( .a ({new_AGEMA_signal_5748, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M10}), .b ({new_AGEMA_signal_5749, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_5845, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M20_U1 ( .a ({new_AGEMA_signal_5750, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M16}), .b ({new_AGEMA_signal_5587, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_5846, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M21_U1 ( .a ({new_AGEMA_signal_5751, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M17}), .b ({new_AGEMA_signal_5749, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_5847, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M22_U1 ( .a ({new_AGEMA_signal_5752, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M18}), .b ({new_AGEMA_signal_5587, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_5848, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M23_U1 ( .a ({new_AGEMA_signal_5845, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M19}), .b ({new_AGEMA_signal_10220, new_AGEMA_signal_10219}), .c ({new_AGEMA_signal_5925, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M24_U1 ( .a ({new_AGEMA_signal_5848, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_5925, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23}), .c ({new_AGEMA_signal_6008, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M27_U1 ( .a ({new_AGEMA_signal_5846, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_5847, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21}), .c ({new_AGEMA_signal_5927, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27}) ) ;
    buf_clk new_AGEMA_reg_buffer_4209 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T14), .Q (new_AGEMA_signal_10061) ) ;
    buf_clk new_AGEMA_reg_buffer_4210 ( .C (clk), .D (new_AGEMA_signal_5347), .Q (new_AGEMA_signal_10062) ) ;
    buf_clk new_AGEMA_reg_buffer_4211 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T26), .Q (new_AGEMA_signal_10063) ) ;
    buf_clk new_AGEMA_reg_buffer_4212 ( .C (clk), .D (new_AGEMA_signal_5351), .Q (new_AGEMA_signal_10064) ) ;
    buf_clk new_AGEMA_reg_buffer_4213 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T24), .Q (new_AGEMA_signal_10065) ) ;
    buf_clk new_AGEMA_reg_buffer_4214 ( .C (clk), .D (new_AGEMA_signal_5589), .Q (new_AGEMA_signal_10066) ) ;
    buf_clk new_AGEMA_reg_buffer_4215 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T25), .Q (new_AGEMA_signal_10067) ) ;
    buf_clk new_AGEMA_reg_buffer_4216 ( .C (clk), .D (new_AGEMA_signal_5590), .Q (new_AGEMA_signal_10068) ) ;
    buf_clk new_AGEMA_reg_buffer_4217 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T14), .Q (new_AGEMA_signal_10069) ) ;
    buf_clk new_AGEMA_reg_buffer_4218 ( .C (clk), .D (new_AGEMA_signal_5360), .Q (new_AGEMA_signal_10070) ) ;
    buf_clk new_AGEMA_reg_buffer_4219 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T26), .Q (new_AGEMA_signal_10071) ) ;
    buf_clk new_AGEMA_reg_buffer_4220 ( .C (clk), .D (new_AGEMA_signal_5364), .Q (new_AGEMA_signal_10072) ) ;
    buf_clk new_AGEMA_reg_buffer_4221 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T24), .Q (new_AGEMA_signal_10073) ) ;
    buf_clk new_AGEMA_reg_buffer_4222 ( .C (clk), .D (new_AGEMA_signal_5598), .Q (new_AGEMA_signal_10074) ) ;
    buf_clk new_AGEMA_reg_buffer_4223 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T25), .Q (new_AGEMA_signal_10075) ) ;
    buf_clk new_AGEMA_reg_buffer_4224 ( .C (clk), .D (new_AGEMA_signal_5599), .Q (new_AGEMA_signal_10076) ) ;
    buf_clk new_AGEMA_reg_buffer_4225 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T14), .Q (new_AGEMA_signal_10077) ) ;
    buf_clk new_AGEMA_reg_buffer_4226 ( .C (clk), .D (new_AGEMA_signal_5373), .Q (new_AGEMA_signal_10078) ) ;
    buf_clk new_AGEMA_reg_buffer_4227 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T26), .Q (new_AGEMA_signal_10079) ) ;
    buf_clk new_AGEMA_reg_buffer_4228 ( .C (clk), .D (new_AGEMA_signal_5377), .Q (new_AGEMA_signal_10080) ) ;
    buf_clk new_AGEMA_reg_buffer_4229 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T24), .Q (new_AGEMA_signal_10081) ) ;
    buf_clk new_AGEMA_reg_buffer_4230 ( .C (clk), .D (new_AGEMA_signal_5607), .Q (new_AGEMA_signal_10082) ) ;
    buf_clk new_AGEMA_reg_buffer_4231 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T25), .Q (new_AGEMA_signal_10083) ) ;
    buf_clk new_AGEMA_reg_buffer_4232 ( .C (clk), .D (new_AGEMA_signal_5608), .Q (new_AGEMA_signal_10084) ) ;
    buf_clk new_AGEMA_reg_buffer_4233 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T14), .Q (new_AGEMA_signal_10085) ) ;
    buf_clk new_AGEMA_reg_buffer_4234 ( .C (clk), .D (new_AGEMA_signal_5386), .Q (new_AGEMA_signal_10086) ) ;
    buf_clk new_AGEMA_reg_buffer_4235 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T26), .Q (new_AGEMA_signal_10087) ) ;
    buf_clk new_AGEMA_reg_buffer_4236 ( .C (clk), .D (new_AGEMA_signal_5390), .Q (new_AGEMA_signal_10088) ) ;
    buf_clk new_AGEMA_reg_buffer_4237 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T24), .Q (new_AGEMA_signal_10089) ) ;
    buf_clk new_AGEMA_reg_buffer_4238 ( .C (clk), .D (new_AGEMA_signal_5616), .Q (new_AGEMA_signal_10090) ) ;
    buf_clk new_AGEMA_reg_buffer_4239 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T25), .Q (new_AGEMA_signal_10091) ) ;
    buf_clk new_AGEMA_reg_buffer_4240 ( .C (clk), .D (new_AGEMA_signal_5617), .Q (new_AGEMA_signal_10092) ) ;
    buf_clk new_AGEMA_reg_buffer_4241 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T14), .Q (new_AGEMA_signal_10093) ) ;
    buf_clk new_AGEMA_reg_buffer_4242 ( .C (clk), .D (new_AGEMA_signal_5399), .Q (new_AGEMA_signal_10094) ) ;
    buf_clk new_AGEMA_reg_buffer_4243 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T26), .Q (new_AGEMA_signal_10095) ) ;
    buf_clk new_AGEMA_reg_buffer_4244 ( .C (clk), .D (new_AGEMA_signal_5403), .Q (new_AGEMA_signal_10096) ) ;
    buf_clk new_AGEMA_reg_buffer_4245 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T24), .Q (new_AGEMA_signal_10097) ) ;
    buf_clk new_AGEMA_reg_buffer_4246 ( .C (clk), .D (new_AGEMA_signal_5625), .Q (new_AGEMA_signal_10098) ) ;
    buf_clk new_AGEMA_reg_buffer_4247 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T25), .Q (new_AGEMA_signal_10099) ) ;
    buf_clk new_AGEMA_reg_buffer_4248 ( .C (clk), .D (new_AGEMA_signal_5626), .Q (new_AGEMA_signal_10100) ) ;
    buf_clk new_AGEMA_reg_buffer_4249 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T14), .Q (new_AGEMA_signal_10101) ) ;
    buf_clk new_AGEMA_reg_buffer_4250 ( .C (clk), .D (new_AGEMA_signal_5412), .Q (new_AGEMA_signal_10102) ) ;
    buf_clk new_AGEMA_reg_buffer_4251 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T26), .Q (new_AGEMA_signal_10103) ) ;
    buf_clk new_AGEMA_reg_buffer_4252 ( .C (clk), .D (new_AGEMA_signal_5416), .Q (new_AGEMA_signal_10104) ) ;
    buf_clk new_AGEMA_reg_buffer_4253 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T24), .Q (new_AGEMA_signal_10105) ) ;
    buf_clk new_AGEMA_reg_buffer_4254 ( .C (clk), .D (new_AGEMA_signal_5634), .Q (new_AGEMA_signal_10106) ) ;
    buf_clk new_AGEMA_reg_buffer_4255 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T25), .Q (new_AGEMA_signal_10107) ) ;
    buf_clk new_AGEMA_reg_buffer_4256 ( .C (clk), .D (new_AGEMA_signal_5635), .Q (new_AGEMA_signal_10108) ) ;
    buf_clk new_AGEMA_reg_buffer_4257 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T14), .Q (new_AGEMA_signal_10109) ) ;
    buf_clk new_AGEMA_reg_buffer_4258 ( .C (clk), .D (new_AGEMA_signal_5425), .Q (new_AGEMA_signal_10110) ) ;
    buf_clk new_AGEMA_reg_buffer_4259 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T26), .Q (new_AGEMA_signal_10111) ) ;
    buf_clk new_AGEMA_reg_buffer_4260 ( .C (clk), .D (new_AGEMA_signal_5429), .Q (new_AGEMA_signal_10112) ) ;
    buf_clk new_AGEMA_reg_buffer_4261 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T24), .Q (new_AGEMA_signal_10113) ) ;
    buf_clk new_AGEMA_reg_buffer_4262 ( .C (clk), .D (new_AGEMA_signal_5643), .Q (new_AGEMA_signal_10114) ) ;
    buf_clk new_AGEMA_reg_buffer_4263 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T25), .Q (new_AGEMA_signal_10115) ) ;
    buf_clk new_AGEMA_reg_buffer_4264 ( .C (clk), .D (new_AGEMA_signal_5644), .Q (new_AGEMA_signal_10116) ) ;
    buf_clk new_AGEMA_reg_buffer_4265 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T14), .Q (new_AGEMA_signal_10117) ) ;
    buf_clk new_AGEMA_reg_buffer_4266 ( .C (clk), .D (new_AGEMA_signal_5438), .Q (new_AGEMA_signal_10118) ) ;
    buf_clk new_AGEMA_reg_buffer_4267 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T26), .Q (new_AGEMA_signal_10119) ) ;
    buf_clk new_AGEMA_reg_buffer_4268 ( .C (clk), .D (new_AGEMA_signal_5442), .Q (new_AGEMA_signal_10120) ) ;
    buf_clk new_AGEMA_reg_buffer_4269 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T24), .Q (new_AGEMA_signal_10121) ) ;
    buf_clk new_AGEMA_reg_buffer_4270 ( .C (clk), .D (new_AGEMA_signal_5652), .Q (new_AGEMA_signal_10122) ) ;
    buf_clk new_AGEMA_reg_buffer_4271 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T25), .Q (new_AGEMA_signal_10123) ) ;
    buf_clk new_AGEMA_reg_buffer_4272 ( .C (clk), .D (new_AGEMA_signal_5653), .Q (new_AGEMA_signal_10124) ) ;
    buf_clk new_AGEMA_reg_buffer_4273 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T14), .Q (new_AGEMA_signal_10125) ) ;
    buf_clk new_AGEMA_reg_buffer_4274 ( .C (clk), .D (new_AGEMA_signal_5451), .Q (new_AGEMA_signal_10126) ) ;
    buf_clk new_AGEMA_reg_buffer_4275 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T26), .Q (new_AGEMA_signal_10127) ) ;
    buf_clk new_AGEMA_reg_buffer_4276 ( .C (clk), .D (new_AGEMA_signal_5455), .Q (new_AGEMA_signal_10128) ) ;
    buf_clk new_AGEMA_reg_buffer_4277 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T24), .Q (new_AGEMA_signal_10129) ) ;
    buf_clk new_AGEMA_reg_buffer_4278 ( .C (clk), .D (new_AGEMA_signal_5661), .Q (new_AGEMA_signal_10130) ) ;
    buf_clk new_AGEMA_reg_buffer_4279 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T25), .Q (new_AGEMA_signal_10131) ) ;
    buf_clk new_AGEMA_reg_buffer_4280 ( .C (clk), .D (new_AGEMA_signal_5662), .Q (new_AGEMA_signal_10132) ) ;
    buf_clk new_AGEMA_reg_buffer_4281 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T14), .Q (new_AGEMA_signal_10133) ) ;
    buf_clk new_AGEMA_reg_buffer_4282 ( .C (clk), .D (new_AGEMA_signal_5464), .Q (new_AGEMA_signal_10134) ) ;
    buf_clk new_AGEMA_reg_buffer_4283 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T26), .Q (new_AGEMA_signal_10135) ) ;
    buf_clk new_AGEMA_reg_buffer_4284 ( .C (clk), .D (new_AGEMA_signal_5468), .Q (new_AGEMA_signal_10136) ) ;
    buf_clk new_AGEMA_reg_buffer_4285 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T24), .Q (new_AGEMA_signal_10137) ) ;
    buf_clk new_AGEMA_reg_buffer_4286 ( .C (clk), .D (new_AGEMA_signal_5670), .Q (new_AGEMA_signal_10138) ) ;
    buf_clk new_AGEMA_reg_buffer_4287 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T25), .Q (new_AGEMA_signal_10139) ) ;
    buf_clk new_AGEMA_reg_buffer_4288 ( .C (clk), .D (new_AGEMA_signal_5671), .Q (new_AGEMA_signal_10140) ) ;
    buf_clk new_AGEMA_reg_buffer_4289 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T14), .Q (new_AGEMA_signal_10141) ) ;
    buf_clk new_AGEMA_reg_buffer_4290 ( .C (clk), .D (new_AGEMA_signal_5477), .Q (new_AGEMA_signal_10142) ) ;
    buf_clk new_AGEMA_reg_buffer_4291 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T26), .Q (new_AGEMA_signal_10143) ) ;
    buf_clk new_AGEMA_reg_buffer_4292 ( .C (clk), .D (new_AGEMA_signal_5481), .Q (new_AGEMA_signal_10144) ) ;
    buf_clk new_AGEMA_reg_buffer_4293 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T24), .Q (new_AGEMA_signal_10145) ) ;
    buf_clk new_AGEMA_reg_buffer_4294 ( .C (clk), .D (new_AGEMA_signal_5679), .Q (new_AGEMA_signal_10146) ) ;
    buf_clk new_AGEMA_reg_buffer_4295 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T25), .Q (new_AGEMA_signal_10147) ) ;
    buf_clk new_AGEMA_reg_buffer_4296 ( .C (clk), .D (new_AGEMA_signal_5680), .Q (new_AGEMA_signal_10148) ) ;
    buf_clk new_AGEMA_reg_buffer_4297 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T14), .Q (new_AGEMA_signal_10149) ) ;
    buf_clk new_AGEMA_reg_buffer_4298 ( .C (clk), .D (new_AGEMA_signal_5490), .Q (new_AGEMA_signal_10150) ) ;
    buf_clk new_AGEMA_reg_buffer_4299 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T26), .Q (new_AGEMA_signal_10151) ) ;
    buf_clk new_AGEMA_reg_buffer_4300 ( .C (clk), .D (new_AGEMA_signal_5494), .Q (new_AGEMA_signal_10152) ) ;
    buf_clk new_AGEMA_reg_buffer_4301 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T24), .Q (new_AGEMA_signal_10153) ) ;
    buf_clk new_AGEMA_reg_buffer_4302 ( .C (clk), .D (new_AGEMA_signal_5688), .Q (new_AGEMA_signal_10154) ) ;
    buf_clk new_AGEMA_reg_buffer_4303 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T25), .Q (new_AGEMA_signal_10155) ) ;
    buf_clk new_AGEMA_reg_buffer_4304 ( .C (clk), .D (new_AGEMA_signal_5689), .Q (new_AGEMA_signal_10156) ) ;
    buf_clk new_AGEMA_reg_buffer_4305 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T14), .Q (new_AGEMA_signal_10157) ) ;
    buf_clk new_AGEMA_reg_buffer_4306 ( .C (clk), .D (new_AGEMA_signal_5503), .Q (new_AGEMA_signal_10158) ) ;
    buf_clk new_AGEMA_reg_buffer_4307 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T26), .Q (new_AGEMA_signal_10159) ) ;
    buf_clk new_AGEMA_reg_buffer_4308 ( .C (clk), .D (new_AGEMA_signal_5507), .Q (new_AGEMA_signal_10160) ) ;
    buf_clk new_AGEMA_reg_buffer_4309 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T24), .Q (new_AGEMA_signal_10161) ) ;
    buf_clk new_AGEMA_reg_buffer_4310 ( .C (clk), .D (new_AGEMA_signal_5697), .Q (new_AGEMA_signal_10162) ) ;
    buf_clk new_AGEMA_reg_buffer_4311 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T25), .Q (new_AGEMA_signal_10163) ) ;
    buf_clk new_AGEMA_reg_buffer_4312 ( .C (clk), .D (new_AGEMA_signal_5698), .Q (new_AGEMA_signal_10164) ) ;
    buf_clk new_AGEMA_reg_buffer_4313 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T14), .Q (new_AGEMA_signal_10165) ) ;
    buf_clk new_AGEMA_reg_buffer_4314 ( .C (clk), .D (new_AGEMA_signal_5516), .Q (new_AGEMA_signal_10166) ) ;
    buf_clk new_AGEMA_reg_buffer_4315 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T26), .Q (new_AGEMA_signal_10167) ) ;
    buf_clk new_AGEMA_reg_buffer_4316 ( .C (clk), .D (new_AGEMA_signal_5520), .Q (new_AGEMA_signal_10168) ) ;
    buf_clk new_AGEMA_reg_buffer_4317 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T24), .Q (new_AGEMA_signal_10169) ) ;
    buf_clk new_AGEMA_reg_buffer_4318 ( .C (clk), .D (new_AGEMA_signal_5706), .Q (new_AGEMA_signal_10170) ) ;
    buf_clk new_AGEMA_reg_buffer_4319 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T25), .Q (new_AGEMA_signal_10171) ) ;
    buf_clk new_AGEMA_reg_buffer_4320 ( .C (clk), .D (new_AGEMA_signal_5707), .Q (new_AGEMA_signal_10172) ) ;
    buf_clk new_AGEMA_reg_buffer_4321 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T14), .Q (new_AGEMA_signal_10173) ) ;
    buf_clk new_AGEMA_reg_buffer_4322 ( .C (clk), .D (new_AGEMA_signal_5529), .Q (new_AGEMA_signal_10174) ) ;
    buf_clk new_AGEMA_reg_buffer_4323 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T26), .Q (new_AGEMA_signal_10175) ) ;
    buf_clk new_AGEMA_reg_buffer_4324 ( .C (clk), .D (new_AGEMA_signal_5533), .Q (new_AGEMA_signal_10176) ) ;
    buf_clk new_AGEMA_reg_buffer_4325 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T24), .Q (new_AGEMA_signal_10177) ) ;
    buf_clk new_AGEMA_reg_buffer_4326 ( .C (clk), .D (new_AGEMA_signal_5715), .Q (new_AGEMA_signal_10178) ) ;
    buf_clk new_AGEMA_reg_buffer_4327 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T25), .Q (new_AGEMA_signal_10179) ) ;
    buf_clk new_AGEMA_reg_buffer_4328 ( .C (clk), .D (new_AGEMA_signal_5716), .Q (new_AGEMA_signal_10180) ) ;
    buf_clk new_AGEMA_reg_buffer_4329 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T14), .Q (new_AGEMA_signal_10181) ) ;
    buf_clk new_AGEMA_reg_buffer_4330 ( .C (clk), .D (new_AGEMA_signal_5542), .Q (new_AGEMA_signal_10182) ) ;
    buf_clk new_AGEMA_reg_buffer_4331 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T26), .Q (new_AGEMA_signal_10183) ) ;
    buf_clk new_AGEMA_reg_buffer_4332 ( .C (clk), .D (new_AGEMA_signal_5546), .Q (new_AGEMA_signal_10184) ) ;
    buf_clk new_AGEMA_reg_buffer_4333 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T24), .Q (new_AGEMA_signal_10185) ) ;
    buf_clk new_AGEMA_reg_buffer_4334 ( .C (clk), .D (new_AGEMA_signal_5724), .Q (new_AGEMA_signal_10186) ) ;
    buf_clk new_AGEMA_reg_buffer_4335 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T25), .Q (new_AGEMA_signal_10187) ) ;
    buf_clk new_AGEMA_reg_buffer_4336 ( .C (clk), .D (new_AGEMA_signal_5725), .Q (new_AGEMA_signal_10188) ) ;
    buf_clk new_AGEMA_reg_buffer_4337 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T14), .Q (new_AGEMA_signal_10189) ) ;
    buf_clk new_AGEMA_reg_buffer_4338 ( .C (clk), .D (new_AGEMA_signal_5295), .Q (new_AGEMA_signal_10190) ) ;
    buf_clk new_AGEMA_reg_buffer_4339 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T26), .Q (new_AGEMA_signal_10191) ) ;
    buf_clk new_AGEMA_reg_buffer_4340 ( .C (clk), .D (new_AGEMA_signal_5299), .Q (new_AGEMA_signal_10192) ) ;
    buf_clk new_AGEMA_reg_buffer_4341 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T24), .Q (new_AGEMA_signal_10193) ) ;
    buf_clk new_AGEMA_reg_buffer_4342 ( .C (clk), .D (new_AGEMA_signal_5553), .Q (new_AGEMA_signal_10194) ) ;
    buf_clk new_AGEMA_reg_buffer_4343 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T25), .Q (new_AGEMA_signal_10195) ) ;
    buf_clk new_AGEMA_reg_buffer_4344 ( .C (clk), .D (new_AGEMA_signal_5554), .Q (new_AGEMA_signal_10196) ) ;
    buf_clk new_AGEMA_reg_buffer_4345 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T14), .Q (new_AGEMA_signal_10197) ) ;
    buf_clk new_AGEMA_reg_buffer_4346 ( .C (clk), .D (new_AGEMA_signal_5308), .Q (new_AGEMA_signal_10198) ) ;
    buf_clk new_AGEMA_reg_buffer_4347 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T26), .Q (new_AGEMA_signal_10199) ) ;
    buf_clk new_AGEMA_reg_buffer_4348 ( .C (clk), .D (new_AGEMA_signal_5312), .Q (new_AGEMA_signal_10200) ) ;
    buf_clk new_AGEMA_reg_buffer_4349 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T24), .Q (new_AGEMA_signal_10201) ) ;
    buf_clk new_AGEMA_reg_buffer_4350 ( .C (clk), .D (new_AGEMA_signal_5562), .Q (new_AGEMA_signal_10202) ) ;
    buf_clk new_AGEMA_reg_buffer_4351 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T25), .Q (new_AGEMA_signal_10203) ) ;
    buf_clk new_AGEMA_reg_buffer_4352 ( .C (clk), .D (new_AGEMA_signal_5563), .Q (new_AGEMA_signal_10204) ) ;
    buf_clk new_AGEMA_reg_buffer_4353 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T14), .Q (new_AGEMA_signal_10205) ) ;
    buf_clk new_AGEMA_reg_buffer_4354 ( .C (clk), .D (new_AGEMA_signal_5321), .Q (new_AGEMA_signal_10206) ) ;
    buf_clk new_AGEMA_reg_buffer_4355 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T26), .Q (new_AGEMA_signal_10207) ) ;
    buf_clk new_AGEMA_reg_buffer_4356 ( .C (clk), .D (new_AGEMA_signal_5325), .Q (new_AGEMA_signal_10208) ) ;
    buf_clk new_AGEMA_reg_buffer_4357 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T24), .Q (new_AGEMA_signal_10209) ) ;
    buf_clk new_AGEMA_reg_buffer_4358 ( .C (clk), .D (new_AGEMA_signal_5571), .Q (new_AGEMA_signal_10210) ) ;
    buf_clk new_AGEMA_reg_buffer_4359 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T25), .Q (new_AGEMA_signal_10211) ) ;
    buf_clk new_AGEMA_reg_buffer_4360 ( .C (clk), .D (new_AGEMA_signal_5572), .Q (new_AGEMA_signal_10212) ) ;
    buf_clk new_AGEMA_reg_buffer_4361 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T14), .Q (new_AGEMA_signal_10213) ) ;
    buf_clk new_AGEMA_reg_buffer_4362 ( .C (clk), .D (new_AGEMA_signal_5334), .Q (new_AGEMA_signal_10214) ) ;
    buf_clk new_AGEMA_reg_buffer_4363 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T26), .Q (new_AGEMA_signal_10215) ) ;
    buf_clk new_AGEMA_reg_buffer_4364 ( .C (clk), .D (new_AGEMA_signal_5338), .Q (new_AGEMA_signal_10216) ) ;
    buf_clk new_AGEMA_reg_buffer_4365 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T24), .Q (new_AGEMA_signal_10217) ) ;
    buf_clk new_AGEMA_reg_buffer_4366 ( .C (clk), .D (new_AGEMA_signal_5580), .Q (new_AGEMA_signal_10218) ) ;
    buf_clk new_AGEMA_reg_buffer_4367 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T25), .Q (new_AGEMA_signal_10219) ) ;
    buf_clk new_AGEMA_reg_buffer_4368 ( .C (clk), .D (new_AGEMA_signal_5581), .Q (new_AGEMA_signal_10220) ) ;
    buf_clk new_AGEMA_reg_buffer_4689 ( .C (clk), .D (n321), .Q (new_AGEMA_signal_10541) ) ;
    buf_clk new_AGEMA_reg_buffer_4693 ( .C (clk), .D (n315), .Q (new_AGEMA_signal_10545) ) ;
    buf_clk new_AGEMA_reg_buffer_4697 ( .C (clk), .D (n316), .Q (new_AGEMA_signal_10549) ) ;
    buf_clk new_AGEMA_reg_buffer_4701 ( .C (clk), .D (n317), .Q (new_AGEMA_signal_10553) ) ;
    buf_clk new_AGEMA_reg_buffer_4705 ( .C (clk), .D (n318), .Q (new_AGEMA_signal_10557) ) ;
    buf_clk new_AGEMA_reg_buffer_4709 ( .C (clk), .D (n319), .Q (new_AGEMA_signal_10561) ) ;
    buf_clk new_AGEMA_reg_buffer_4713 ( .C (clk), .D (n320), .Q (new_AGEMA_signal_10565) ) ;
    buf_clk new_AGEMA_reg_buffer_4717 ( .C (clk), .D (reset), .Q (new_AGEMA_signal_10569) ) ;
    buf_clk new_AGEMA_reg_buffer_4721 ( .C (clk), .D (plaintext_s0[0]), .Q (new_AGEMA_signal_10573) ) ;
    buf_clk new_AGEMA_reg_buffer_4725 ( .C (clk), .D (plaintext_s1[0]), .Q (new_AGEMA_signal_10577) ) ;
    buf_clk new_AGEMA_reg_buffer_4729 ( .C (clk), .D (plaintext_s0[1]), .Q (new_AGEMA_signal_10581) ) ;
    buf_clk new_AGEMA_reg_buffer_4733 ( .C (clk), .D (plaintext_s1[1]), .Q (new_AGEMA_signal_10585) ) ;
    buf_clk new_AGEMA_reg_buffer_4737 ( .C (clk), .D (plaintext_s0[2]), .Q (new_AGEMA_signal_10589) ) ;
    buf_clk new_AGEMA_reg_buffer_4741 ( .C (clk), .D (plaintext_s1[2]), .Q (new_AGEMA_signal_10593) ) ;
    buf_clk new_AGEMA_reg_buffer_4745 ( .C (clk), .D (plaintext_s0[3]), .Q (new_AGEMA_signal_10597) ) ;
    buf_clk new_AGEMA_reg_buffer_4749 ( .C (clk), .D (plaintext_s1[3]), .Q (new_AGEMA_signal_10601) ) ;
    buf_clk new_AGEMA_reg_buffer_4753 ( .C (clk), .D (plaintext_s0[4]), .Q (new_AGEMA_signal_10605) ) ;
    buf_clk new_AGEMA_reg_buffer_4757 ( .C (clk), .D (plaintext_s1[4]), .Q (new_AGEMA_signal_10609) ) ;
    buf_clk new_AGEMA_reg_buffer_4761 ( .C (clk), .D (plaintext_s0[5]), .Q (new_AGEMA_signal_10613) ) ;
    buf_clk new_AGEMA_reg_buffer_4765 ( .C (clk), .D (plaintext_s1[5]), .Q (new_AGEMA_signal_10617) ) ;
    buf_clk new_AGEMA_reg_buffer_4769 ( .C (clk), .D (plaintext_s0[6]), .Q (new_AGEMA_signal_10621) ) ;
    buf_clk new_AGEMA_reg_buffer_4773 ( .C (clk), .D (plaintext_s1[6]), .Q (new_AGEMA_signal_10625) ) ;
    buf_clk new_AGEMA_reg_buffer_4777 ( .C (clk), .D (plaintext_s0[7]), .Q (new_AGEMA_signal_10629) ) ;
    buf_clk new_AGEMA_reg_buffer_4781 ( .C (clk), .D (plaintext_s1[7]), .Q (new_AGEMA_signal_10633) ) ;
    buf_clk new_AGEMA_reg_buffer_4785 ( .C (clk), .D (plaintext_s0[8]), .Q (new_AGEMA_signal_10637) ) ;
    buf_clk new_AGEMA_reg_buffer_4789 ( .C (clk), .D (plaintext_s1[8]), .Q (new_AGEMA_signal_10641) ) ;
    buf_clk new_AGEMA_reg_buffer_4793 ( .C (clk), .D (plaintext_s0[9]), .Q (new_AGEMA_signal_10645) ) ;
    buf_clk new_AGEMA_reg_buffer_4797 ( .C (clk), .D (plaintext_s1[9]), .Q (new_AGEMA_signal_10649) ) ;
    buf_clk new_AGEMA_reg_buffer_4801 ( .C (clk), .D (plaintext_s0[10]), .Q (new_AGEMA_signal_10653) ) ;
    buf_clk new_AGEMA_reg_buffer_4805 ( .C (clk), .D (plaintext_s1[10]), .Q (new_AGEMA_signal_10657) ) ;
    buf_clk new_AGEMA_reg_buffer_4809 ( .C (clk), .D (plaintext_s0[11]), .Q (new_AGEMA_signal_10661) ) ;
    buf_clk new_AGEMA_reg_buffer_4813 ( .C (clk), .D (plaintext_s1[11]), .Q (new_AGEMA_signal_10665) ) ;
    buf_clk new_AGEMA_reg_buffer_4817 ( .C (clk), .D (plaintext_s0[12]), .Q (new_AGEMA_signal_10669) ) ;
    buf_clk new_AGEMA_reg_buffer_4821 ( .C (clk), .D (plaintext_s1[12]), .Q (new_AGEMA_signal_10673) ) ;
    buf_clk new_AGEMA_reg_buffer_4825 ( .C (clk), .D (plaintext_s0[13]), .Q (new_AGEMA_signal_10677) ) ;
    buf_clk new_AGEMA_reg_buffer_4829 ( .C (clk), .D (plaintext_s1[13]), .Q (new_AGEMA_signal_10681) ) ;
    buf_clk new_AGEMA_reg_buffer_4833 ( .C (clk), .D (plaintext_s0[14]), .Q (new_AGEMA_signal_10685) ) ;
    buf_clk new_AGEMA_reg_buffer_4837 ( .C (clk), .D (plaintext_s1[14]), .Q (new_AGEMA_signal_10689) ) ;
    buf_clk new_AGEMA_reg_buffer_4841 ( .C (clk), .D (plaintext_s0[15]), .Q (new_AGEMA_signal_10693) ) ;
    buf_clk new_AGEMA_reg_buffer_4845 ( .C (clk), .D (plaintext_s1[15]), .Q (new_AGEMA_signal_10697) ) ;
    buf_clk new_AGEMA_reg_buffer_4849 ( .C (clk), .D (plaintext_s0[16]), .Q (new_AGEMA_signal_10701) ) ;
    buf_clk new_AGEMA_reg_buffer_4853 ( .C (clk), .D (plaintext_s1[16]), .Q (new_AGEMA_signal_10705) ) ;
    buf_clk new_AGEMA_reg_buffer_4857 ( .C (clk), .D (plaintext_s0[17]), .Q (new_AGEMA_signal_10709) ) ;
    buf_clk new_AGEMA_reg_buffer_4861 ( .C (clk), .D (plaintext_s1[17]), .Q (new_AGEMA_signal_10713) ) ;
    buf_clk new_AGEMA_reg_buffer_4865 ( .C (clk), .D (plaintext_s0[18]), .Q (new_AGEMA_signal_10717) ) ;
    buf_clk new_AGEMA_reg_buffer_4869 ( .C (clk), .D (plaintext_s1[18]), .Q (new_AGEMA_signal_10721) ) ;
    buf_clk new_AGEMA_reg_buffer_4873 ( .C (clk), .D (plaintext_s0[19]), .Q (new_AGEMA_signal_10725) ) ;
    buf_clk new_AGEMA_reg_buffer_4877 ( .C (clk), .D (plaintext_s1[19]), .Q (new_AGEMA_signal_10729) ) ;
    buf_clk new_AGEMA_reg_buffer_4881 ( .C (clk), .D (plaintext_s0[20]), .Q (new_AGEMA_signal_10733) ) ;
    buf_clk new_AGEMA_reg_buffer_4885 ( .C (clk), .D (plaintext_s1[20]), .Q (new_AGEMA_signal_10737) ) ;
    buf_clk new_AGEMA_reg_buffer_4889 ( .C (clk), .D (plaintext_s0[21]), .Q (new_AGEMA_signal_10741) ) ;
    buf_clk new_AGEMA_reg_buffer_4893 ( .C (clk), .D (plaintext_s1[21]), .Q (new_AGEMA_signal_10745) ) ;
    buf_clk new_AGEMA_reg_buffer_4897 ( .C (clk), .D (plaintext_s0[22]), .Q (new_AGEMA_signal_10749) ) ;
    buf_clk new_AGEMA_reg_buffer_4901 ( .C (clk), .D (plaintext_s1[22]), .Q (new_AGEMA_signal_10753) ) ;
    buf_clk new_AGEMA_reg_buffer_4905 ( .C (clk), .D (plaintext_s0[23]), .Q (new_AGEMA_signal_10757) ) ;
    buf_clk new_AGEMA_reg_buffer_4909 ( .C (clk), .D (plaintext_s1[23]), .Q (new_AGEMA_signal_10761) ) ;
    buf_clk new_AGEMA_reg_buffer_4913 ( .C (clk), .D (plaintext_s0[24]), .Q (new_AGEMA_signal_10765) ) ;
    buf_clk new_AGEMA_reg_buffer_4917 ( .C (clk), .D (plaintext_s1[24]), .Q (new_AGEMA_signal_10769) ) ;
    buf_clk new_AGEMA_reg_buffer_4921 ( .C (clk), .D (plaintext_s0[25]), .Q (new_AGEMA_signal_10773) ) ;
    buf_clk new_AGEMA_reg_buffer_4925 ( .C (clk), .D (plaintext_s1[25]), .Q (new_AGEMA_signal_10777) ) ;
    buf_clk new_AGEMA_reg_buffer_4929 ( .C (clk), .D (plaintext_s0[26]), .Q (new_AGEMA_signal_10781) ) ;
    buf_clk new_AGEMA_reg_buffer_4933 ( .C (clk), .D (plaintext_s1[26]), .Q (new_AGEMA_signal_10785) ) ;
    buf_clk new_AGEMA_reg_buffer_4937 ( .C (clk), .D (plaintext_s0[27]), .Q (new_AGEMA_signal_10789) ) ;
    buf_clk new_AGEMA_reg_buffer_4941 ( .C (clk), .D (plaintext_s1[27]), .Q (new_AGEMA_signal_10793) ) ;
    buf_clk new_AGEMA_reg_buffer_4945 ( .C (clk), .D (plaintext_s0[28]), .Q (new_AGEMA_signal_10797) ) ;
    buf_clk new_AGEMA_reg_buffer_4949 ( .C (clk), .D (plaintext_s1[28]), .Q (new_AGEMA_signal_10801) ) ;
    buf_clk new_AGEMA_reg_buffer_4953 ( .C (clk), .D (plaintext_s0[29]), .Q (new_AGEMA_signal_10805) ) ;
    buf_clk new_AGEMA_reg_buffer_4957 ( .C (clk), .D (plaintext_s1[29]), .Q (new_AGEMA_signal_10809) ) ;
    buf_clk new_AGEMA_reg_buffer_4961 ( .C (clk), .D (plaintext_s0[30]), .Q (new_AGEMA_signal_10813) ) ;
    buf_clk new_AGEMA_reg_buffer_4965 ( .C (clk), .D (plaintext_s1[30]), .Q (new_AGEMA_signal_10817) ) ;
    buf_clk new_AGEMA_reg_buffer_4969 ( .C (clk), .D (plaintext_s0[31]), .Q (new_AGEMA_signal_10821) ) ;
    buf_clk new_AGEMA_reg_buffer_4973 ( .C (clk), .D (plaintext_s1[31]), .Q (new_AGEMA_signal_10825) ) ;
    buf_clk new_AGEMA_reg_buffer_4977 ( .C (clk), .D (plaintext_s0[32]), .Q (new_AGEMA_signal_10829) ) ;
    buf_clk new_AGEMA_reg_buffer_4981 ( .C (clk), .D (plaintext_s1[32]), .Q (new_AGEMA_signal_10833) ) ;
    buf_clk new_AGEMA_reg_buffer_4985 ( .C (clk), .D (plaintext_s0[33]), .Q (new_AGEMA_signal_10837) ) ;
    buf_clk new_AGEMA_reg_buffer_4989 ( .C (clk), .D (plaintext_s1[33]), .Q (new_AGEMA_signal_10841) ) ;
    buf_clk new_AGEMA_reg_buffer_4993 ( .C (clk), .D (plaintext_s0[34]), .Q (new_AGEMA_signal_10845) ) ;
    buf_clk new_AGEMA_reg_buffer_4997 ( .C (clk), .D (plaintext_s1[34]), .Q (new_AGEMA_signal_10849) ) ;
    buf_clk new_AGEMA_reg_buffer_5001 ( .C (clk), .D (plaintext_s0[35]), .Q (new_AGEMA_signal_10853) ) ;
    buf_clk new_AGEMA_reg_buffer_5005 ( .C (clk), .D (plaintext_s1[35]), .Q (new_AGEMA_signal_10857) ) ;
    buf_clk new_AGEMA_reg_buffer_5009 ( .C (clk), .D (plaintext_s0[36]), .Q (new_AGEMA_signal_10861) ) ;
    buf_clk new_AGEMA_reg_buffer_5013 ( .C (clk), .D (plaintext_s1[36]), .Q (new_AGEMA_signal_10865) ) ;
    buf_clk new_AGEMA_reg_buffer_5017 ( .C (clk), .D (plaintext_s0[37]), .Q (new_AGEMA_signal_10869) ) ;
    buf_clk new_AGEMA_reg_buffer_5021 ( .C (clk), .D (plaintext_s1[37]), .Q (new_AGEMA_signal_10873) ) ;
    buf_clk new_AGEMA_reg_buffer_5025 ( .C (clk), .D (plaintext_s0[38]), .Q (new_AGEMA_signal_10877) ) ;
    buf_clk new_AGEMA_reg_buffer_5029 ( .C (clk), .D (plaintext_s1[38]), .Q (new_AGEMA_signal_10881) ) ;
    buf_clk new_AGEMA_reg_buffer_5033 ( .C (clk), .D (plaintext_s0[39]), .Q (new_AGEMA_signal_10885) ) ;
    buf_clk new_AGEMA_reg_buffer_5037 ( .C (clk), .D (plaintext_s1[39]), .Q (new_AGEMA_signal_10889) ) ;
    buf_clk new_AGEMA_reg_buffer_5041 ( .C (clk), .D (plaintext_s0[40]), .Q (new_AGEMA_signal_10893) ) ;
    buf_clk new_AGEMA_reg_buffer_5045 ( .C (clk), .D (plaintext_s1[40]), .Q (new_AGEMA_signal_10897) ) ;
    buf_clk new_AGEMA_reg_buffer_5049 ( .C (clk), .D (plaintext_s0[41]), .Q (new_AGEMA_signal_10901) ) ;
    buf_clk new_AGEMA_reg_buffer_5053 ( .C (clk), .D (plaintext_s1[41]), .Q (new_AGEMA_signal_10905) ) ;
    buf_clk new_AGEMA_reg_buffer_5057 ( .C (clk), .D (plaintext_s0[42]), .Q (new_AGEMA_signal_10909) ) ;
    buf_clk new_AGEMA_reg_buffer_5061 ( .C (clk), .D (plaintext_s1[42]), .Q (new_AGEMA_signal_10913) ) ;
    buf_clk new_AGEMA_reg_buffer_5065 ( .C (clk), .D (plaintext_s0[43]), .Q (new_AGEMA_signal_10917) ) ;
    buf_clk new_AGEMA_reg_buffer_5069 ( .C (clk), .D (plaintext_s1[43]), .Q (new_AGEMA_signal_10921) ) ;
    buf_clk new_AGEMA_reg_buffer_5073 ( .C (clk), .D (plaintext_s0[44]), .Q (new_AGEMA_signal_10925) ) ;
    buf_clk new_AGEMA_reg_buffer_5077 ( .C (clk), .D (plaintext_s1[44]), .Q (new_AGEMA_signal_10929) ) ;
    buf_clk new_AGEMA_reg_buffer_5081 ( .C (clk), .D (plaintext_s0[45]), .Q (new_AGEMA_signal_10933) ) ;
    buf_clk new_AGEMA_reg_buffer_5085 ( .C (clk), .D (plaintext_s1[45]), .Q (new_AGEMA_signal_10937) ) ;
    buf_clk new_AGEMA_reg_buffer_5089 ( .C (clk), .D (plaintext_s0[46]), .Q (new_AGEMA_signal_10941) ) ;
    buf_clk new_AGEMA_reg_buffer_5093 ( .C (clk), .D (plaintext_s1[46]), .Q (new_AGEMA_signal_10945) ) ;
    buf_clk new_AGEMA_reg_buffer_5097 ( .C (clk), .D (plaintext_s0[47]), .Q (new_AGEMA_signal_10949) ) ;
    buf_clk new_AGEMA_reg_buffer_5101 ( .C (clk), .D (plaintext_s1[47]), .Q (new_AGEMA_signal_10953) ) ;
    buf_clk new_AGEMA_reg_buffer_5105 ( .C (clk), .D (plaintext_s0[48]), .Q (new_AGEMA_signal_10957) ) ;
    buf_clk new_AGEMA_reg_buffer_5109 ( .C (clk), .D (plaintext_s1[48]), .Q (new_AGEMA_signal_10961) ) ;
    buf_clk new_AGEMA_reg_buffer_5113 ( .C (clk), .D (plaintext_s0[49]), .Q (new_AGEMA_signal_10965) ) ;
    buf_clk new_AGEMA_reg_buffer_5117 ( .C (clk), .D (plaintext_s1[49]), .Q (new_AGEMA_signal_10969) ) ;
    buf_clk new_AGEMA_reg_buffer_5121 ( .C (clk), .D (plaintext_s0[50]), .Q (new_AGEMA_signal_10973) ) ;
    buf_clk new_AGEMA_reg_buffer_5125 ( .C (clk), .D (plaintext_s1[50]), .Q (new_AGEMA_signal_10977) ) ;
    buf_clk new_AGEMA_reg_buffer_5129 ( .C (clk), .D (plaintext_s0[51]), .Q (new_AGEMA_signal_10981) ) ;
    buf_clk new_AGEMA_reg_buffer_5133 ( .C (clk), .D (plaintext_s1[51]), .Q (new_AGEMA_signal_10985) ) ;
    buf_clk new_AGEMA_reg_buffer_5137 ( .C (clk), .D (plaintext_s0[52]), .Q (new_AGEMA_signal_10989) ) ;
    buf_clk new_AGEMA_reg_buffer_5141 ( .C (clk), .D (plaintext_s1[52]), .Q (new_AGEMA_signal_10993) ) ;
    buf_clk new_AGEMA_reg_buffer_5145 ( .C (clk), .D (plaintext_s0[53]), .Q (new_AGEMA_signal_10997) ) ;
    buf_clk new_AGEMA_reg_buffer_5149 ( .C (clk), .D (plaintext_s1[53]), .Q (new_AGEMA_signal_11001) ) ;
    buf_clk new_AGEMA_reg_buffer_5153 ( .C (clk), .D (plaintext_s0[54]), .Q (new_AGEMA_signal_11005) ) ;
    buf_clk new_AGEMA_reg_buffer_5157 ( .C (clk), .D (plaintext_s1[54]), .Q (new_AGEMA_signal_11009) ) ;
    buf_clk new_AGEMA_reg_buffer_5161 ( .C (clk), .D (plaintext_s0[55]), .Q (new_AGEMA_signal_11013) ) ;
    buf_clk new_AGEMA_reg_buffer_5165 ( .C (clk), .D (plaintext_s1[55]), .Q (new_AGEMA_signal_11017) ) ;
    buf_clk new_AGEMA_reg_buffer_5169 ( .C (clk), .D (plaintext_s0[56]), .Q (new_AGEMA_signal_11021) ) ;
    buf_clk new_AGEMA_reg_buffer_5173 ( .C (clk), .D (plaintext_s1[56]), .Q (new_AGEMA_signal_11025) ) ;
    buf_clk new_AGEMA_reg_buffer_5177 ( .C (clk), .D (plaintext_s0[57]), .Q (new_AGEMA_signal_11029) ) ;
    buf_clk new_AGEMA_reg_buffer_5181 ( .C (clk), .D (plaintext_s1[57]), .Q (new_AGEMA_signal_11033) ) ;
    buf_clk new_AGEMA_reg_buffer_5185 ( .C (clk), .D (plaintext_s0[58]), .Q (new_AGEMA_signal_11037) ) ;
    buf_clk new_AGEMA_reg_buffer_5189 ( .C (clk), .D (plaintext_s1[58]), .Q (new_AGEMA_signal_11041) ) ;
    buf_clk new_AGEMA_reg_buffer_5193 ( .C (clk), .D (plaintext_s0[59]), .Q (new_AGEMA_signal_11045) ) ;
    buf_clk new_AGEMA_reg_buffer_5197 ( .C (clk), .D (plaintext_s1[59]), .Q (new_AGEMA_signal_11049) ) ;
    buf_clk new_AGEMA_reg_buffer_5201 ( .C (clk), .D (plaintext_s0[60]), .Q (new_AGEMA_signal_11053) ) ;
    buf_clk new_AGEMA_reg_buffer_5205 ( .C (clk), .D (plaintext_s1[60]), .Q (new_AGEMA_signal_11057) ) ;
    buf_clk new_AGEMA_reg_buffer_5209 ( .C (clk), .D (plaintext_s0[61]), .Q (new_AGEMA_signal_11061) ) ;
    buf_clk new_AGEMA_reg_buffer_5213 ( .C (clk), .D (plaintext_s1[61]), .Q (new_AGEMA_signal_11065) ) ;
    buf_clk new_AGEMA_reg_buffer_5217 ( .C (clk), .D (plaintext_s0[62]), .Q (new_AGEMA_signal_11069) ) ;
    buf_clk new_AGEMA_reg_buffer_5221 ( .C (clk), .D (plaintext_s1[62]), .Q (new_AGEMA_signal_11073) ) ;
    buf_clk new_AGEMA_reg_buffer_5225 ( .C (clk), .D (plaintext_s0[63]), .Q (new_AGEMA_signal_11077) ) ;
    buf_clk new_AGEMA_reg_buffer_5229 ( .C (clk), .D (plaintext_s1[63]), .Q (new_AGEMA_signal_11081) ) ;
    buf_clk new_AGEMA_reg_buffer_5233 ( .C (clk), .D (plaintext_s0[64]), .Q (new_AGEMA_signal_11085) ) ;
    buf_clk new_AGEMA_reg_buffer_5237 ( .C (clk), .D (plaintext_s1[64]), .Q (new_AGEMA_signal_11089) ) ;
    buf_clk new_AGEMA_reg_buffer_5241 ( .C (clk), .D (plaintext_s0[65]), .Q (new_AGEMA_signal_11093) ) ;
    buf_clk new_AGEMA_reg_buffer_5245 ( .C (clk), .D (plaintext_s1[65]), .Q (new_AGEMA_signal_11097) ) ;
    buf_clk new_AGEMA_reg_buffer_5249 ( .C (clk), .D (plaintext_s0[66]), .Q (new_AGEMA_signal_11101) ) ;
    buf_clk new_AGEMA_reg_buffer_5253 ( .C (clk), .D (plaintext_s1[66]), .Q (new_AGEMA_signal_11105) ) ;
    buf_clk new_AGEMA_reg_buffer_5257 ( .C (clk), .D (plaintext_s0[67]), .Q (new_AGEMA_signal_11109) ) ;
    buf_clk new_AGEMA_reg_buffer_5261 ( .C (clk), .D (plaintext_s1[67]), .Q (new_AGEMA_signal_11113) ) ;
    buf_clk new_AGEMA_reg_buffer_5265 ( .C (clk), .D (plaintext_s0[68]), .Q (new_AGEMA_signal_11117) ) ;
    buf_clk new_AGEMA_reg_buffer_5269 ( .C (clk), .D (plaintext_s1[68]), .Q (new_AGEMA_signal_11121) ) ;
    buf_clk new_AGEMA_reg_buffer_5273 ( .C (clk), .D (plaintext_s0[69]), .Q (new_AGEMA_signal_11125) ) ;
    buf_clk new_AGEMA_reg_buffer_5277 ( .C (clk), .D (plaintext_s1[69]), .Q (new_AGEMA_signal_11129) ) ;
    buf_clk new_AGEMA_reg_buffer_5281 ( .C (clk), .D (plaintext_s0[70]), .Q (new_AGEMA_signal_11133) ) ;
    buf_clk new_AGEMA_reg_buffer_5285 ( .C (clk), .D (plaintext_s1[70]), .Q (new_AGEMA_signal_11137) ) ;
    buf_clk new_AGEMA_reg_buffer_5289 ( .C (clk), .D (plaintext_s0[71]), .Q (new_AGEMA_signal_11141) ) ;
    buf_clk new_AGEMA_reg_buffer_5293 ( .C (clk), .D (plaintext_s1[71]), .Q (new_AGEMA_signal_11145) ) ;
    buf_clk new_AGEMA_reg_buffer_5297 ( .C (clk), .D (plaintext_s0[72]), .Q (new_AGEMA_signal_11149) ) ;
    buf_clk new_AGEMA_reg_buffer_5301 ( .C (clk), .D (plaintext_s1[72]), .Q (new_AGEMA_signal_11153) ) ;
    buf_clk new_AGEMA_reg_buffer_5305 ( .C (clk), .D (plaintext_s0[73]), .Q (new_AGEMA_signal_11157) ) ;
    buf_clk new_AGEMA_reg_buffer_5309 ( .C (clk), .D (plaintext_s1[73]), .Q (new_AGEMA_signal_11161) ) ;
    buf_clk new_AGEMA_reg_buffer_5313 ( .C (clk), .D (plaintext_s0[74]), .Q (new_AGEMA_signal_11165) ) ;
    buf_clk new_AGEMA_reg_buffer_5317 ( .C (clk), .D (plaintext_s1[74]), .Q (new_AGEMA_signal_11169) ) ;
    buf_clk new_AGEMA_reg_buffer_5321 ( .C (clk), .D (plaintext_s0[75]), .Q (new_AGEMA_signal_11173) ) ;
    buf_clk new_AGEMA_reg_buffer_5325 ( .C (clk), .D (plaintext_s1[75]), .Q (new_AGEMA_signal_11177) ) ;
    buf_clk new_AGEMA_reg_buffer_5329 ( .C (clk), .D (plaintext_s0[76]), .Q (new_AGEMA_signal_11181) ) ;
    buf_clk new_AGEMA_reg_buffer_5333 ( .C (clk), .D (plaintext_s1[76]), .Q (new_AGEMA_signal_11185) ) ;
    buf_clk new_AGEMA_reg_buffer_5337 ( .C (clk), .D (plaintext_s0[77]), .Q (new_AGEMA_signal_11189) ) ;
    buf_clk new_AGEMA_reg_buffer_5341 ( .C (clk), .D (plaintext_s1[77]), .Q (new_AGEMA_signal_11193) ) ;
    buf_clk new_AGEMA_reg_buffer_5345 ( .C (clk), .D (plaintext_s0[78]), .Q (new_AGEMA_signal_11197) ) ;
    buf_clk new_AGEMA_reg_buffer_5349 ( .C (clk), .D (plaintext_s1[78]), .Q (new_AGEMA_signal_11201) ) ;
    buf_clk new_AGEMA_reg_buffer_5353 ( .C (clk), .D (plaintext_s0[79]), .Q (new_AGEMA_signal_11205) ) ;
    buf_clk new_AGEMA_reg_buffer_5357 ( .C (clk), .D (plaintext_s1[79]), .Q (new_AGEMA_signal_11209) ) ;
    buf_clk new_AGEMA_reg_buffer_5361 ( .C (clk), .D (plaintext_s0[80]), .Q (new_AGEMA_signal_11213) ) ;
    buf_clk new_AGEMA_reg_buffer_5365 ( .C (clk), .D (plaintext_s1[80]), .Q (new_AGEMA_signal_11217) ) ;
    buf_clk new_AGEMA_reg_buffer_5369 ( .C (clk), .D (plaintext_s0[81]), .Q (new_AGEMA_signal_11221) ) ;
    buf_clk new_AGEMA_reg_buffer_5373 ( .C (clk), .D (plaintext_s1[81]), .Q (new_AGEMA_signal_11225) ) ;
    buf_clk new_AGEMA_reg_buffer_5377 ( .C (clk), .D (plaintext_s0[82]), .Q (new_AGEMA_signal_11229) ) ;
    buf_clk new_AGEMA_reg_buffer_5381 ( .C (clk), .D (plaintext_s1[82]), .Q (new_AGEMA_signal_11233) ) ;
    buf_clk new_AGEMA_reg_buffer_5385 ( .C (clk), .D (plaintext_s0[83]), .Q (new_AGEMA_signal_11237) ) ;
    buf_clk new_AGEMA_reg_buffer_5389 ( .C (clk), .D (plaintext_s1[83]), .Q (new_AGEMA_signal_11241) ) ;
    buf_clk new_AGEMA_reg_buffer_5393 ( .C (clk), .D (plaintext_s0[84]), .Q (new_AGEMA_signal_11245) ) ;
    buf_clk new_AGEMA_reg_buffer_5397 ( .C (clk), .D (plaintext_s1[84]), .Q (new_AGEMA_signal_11249) ) ;
    buf_clk new_AGEMA_reg_buffer_5401 ( .C (clk), .D (plaintext_s0[85]), .Q (new_AGEMA_signal_11253) ) ;
    buf_clk new_AGEMA_reg_buffer_5405 ( .C (clk), .D (plaintext_s1[85]), .Q (new_AGEMA_signal_11257) ) ;
    buf_clk new_AGEMA_reg_buffer_5409 ( .C (clk), .D (plaintext_s0[86]), .Q (new_AGEMA_signal_11261) ) ;
    buf_clk new_AGEMA_reg_buffer_5413 ( .C (clk), .D (plaintext_s1[86]), .Q (new_AGEMA_signal_11265) ) ;
    buf_clk new_AGEMA_reg_buffer_5417 ( .C (clk), .D (plaintext_s0[87]), .Q (new_AGEMA_signal_11269) ) ;
    buf_clk new_AGEMA_reg_buffer_5421 ( .C (clk), .D (plaintext_s1[87]), .Q (new_AGEMA_signal_11273) ) ;
    buf_clk new_AGEMA_reg_buffer_5425 ( .C (clk), .D (plaintext_s0[88]), .Q (new_AGEMA_signal_11277) ) ;
    buf_clk new_AGEMA_reg_buffer_5429 ( .C (clk), .D (plaintext_s1[88]), .Q (new_AGEMA_signal_11281) ) ;
    buf_clk new_AGEMA_reg_buffer_5433 ( .C (clk), .D (plaintext_s0[89]), .Q (new_AGEMA_signal_11285) ) ;
    buf_clk new_AGEMA_reg_buffer_5437 ( .C (clk), .D (plaintext_s1[89]), .Q (new_AGEMA_signal_11289) ) ;
    buf_clk new_AGEMA_reg_buffer_5441 ( .C (clk), .D (plaintext_s0[90]), .Q (new_AGEMA_signal_11293) ) ;
    buf_clk new_AGEMA_reg_buffer_5445 ( .C (clk), .D (plaintext_s1[90]), .Q (new_AGEMA_signal_11297) ) ;
    buf_clk new_AGEMA_reg_buffer_5449 ( .C (clk), .D (plaintext_s0[91]), .Q (new_AGEMA_signal_11301) ) ;
    buf_clk new_AGEMA_reg_buffer_5453 ( .C (clk), .D (plaintext_s1[91]), .Q (new_AGEMA_signal_11305) ) ;
    buf_clk new_AGEMA_reg_buffer_5457 ( .C (clk), .D (plaintext_s0[92]), .Q (new_AGEMA_signal_11309) ) ;
    buf_clk new_AGEMA_reg_buffer_5461 ( .C (clk), .D (plaintext_s1[92]), .Q (new_AGEMA_signal_11313) ) ;
    buf_clk new_AGEMA_reg_buffer_5465 ( .C (clk), .D (plaintext_s0[93]), .Q (new_AGEMA_signal_11317) ) ;
    buf_clk new_AGEMA_reg_buffer_5469 ( .C (clk), .D (plaintext_s1[93]), .Q (new_AGEMA_signal_11321) ) ;
    buf_clk new_AGEMA_reg_buffer_5473 ( .C (clk), .D (plaintext_s0[94]), .Q (new_AGEMA_signal_11325) ) ;
    buf_clk new_AGEMA_reg_buffer_5477 ( .C (clk), .D (plaintext_s1[94]), .Q (new_AGEMA_signal_11329) ) ;
    buf_clk new_AGEMA_reg_buffer_5481 ( .C (clk), .D (plaintext_s0[95]), .Q (new_AGEMA_signal_11333) ) ;
    buf_clk new_AGEMA_reg_buffer_5485 ( .C (clk), .D (plaintext_s1[95]), .Q (new_AGEMA_signal_11337) ) ;
    buf_clk new_AGEMA_reg_buffer_5489 ( .C (clk), .D (plaintext_s0[96]), .Q (new_AGEMA_signal_11341) ) ;
    buf_clk new_AGEMA_reg_buffer_5493 ( .C (clk), .D (plaintext_s1[96]), .Q (new_AGEMA_signal_11345) ) ;
    buf_clk new_AGEMA_reg_buffer_5497 ( .C (clk), .D (plaintext_s0[97]), .Q (new_AGEMA_signal_11349) ) ;
    buf_clk new_AGEMA_reg_buffer_5501 ( .C (clk), .D (plaintext_s1[97]), .Q (new_AGEMA_signal_11353) ) ;
    buf_clk new_AGEMA_reg_buffer_5505 ( .C (clk), .D (plaintext_s0[98]), .Q (new_AGEMA_signal_11357) ) ;
    buf_clk new_AGEMA_reg_buffer_5509 ( .C (clk), .D (plaintext_s1[98]), .Q (new_AGEMA_signal_11361) ) ;
    buf_clk new_AGEMA_reg_buffer_5513 ( .C (clk), .D (plaintext_s0[99]), .Q (new_AGEMA_signal_11365) ) ;
    buf_clk new_AGEMA_reg_buffer_5517 ( .C (clk), .D (plaintext_s1[99]), .Q (new_AGEMA_signal_11369) ) ;
    buf_clk new_AGEMA_reg_buffer_5521 ( .C (clk), .D (plaintext_s0[100]), .Q (new_AGEMA_signal_11373) ) ;
    buf_clk new_AGEMA_reg_buffer_5525 ( .C (clk), .D (plaintext_s1[100]), .Q (new_AGEMA_signal_11377) ) ;
    buf_clk new_AGEMA_reg_buffer_5529 ( .C (clk), .D (plaintext_s0[101]), .Q (new_AGEMA_signal_11381) ) ;
    buf_clk new_AGEMA_reg_buffer_5533 ( .C (clk), .D (plaintext_s1[101]), .Q (new_AGEMA_signal_11385) ) ;
    buf_clk new_AGEMA_reg_buffer_5537 ( .C (clk), .D (plaintext_s0[102]), .Q (new_AGEMA_signal_11389) ) ;
    buf_clk new_AGEMA_reg_buffer_5541 ( .C (clk), .D (plaintext_s1[102]), .Q (new_AGEMA_signal_11393) ) ;
    buf_clk new_AGEMA_reg_buffer_5545 ( .C (clk), .D (plaintext_s0[103]), .Q (new_AGEMA_signal_11397) ) ;
    buf_clk new_AGEMA_reg_buffer_5549 ( .C (clk), .D (plaintext_s1[103]), .Q (new_AGEMA_signal_11401) ) ;
    buf_clk new_AGEMA_reg_buffer_5553 ( .C (clk), .D (plaintext_s0[104]), .Q (new_AGEMA_signal_11405) ) ;
    buf_clk new_AGEMA_reg_buffer_5557 ( .C (clk), .D (plaintext_s1[104]), .Q (new_AGEMA_signal_11409) ) ;
    buf_clk new_AGEMA_reg_buffer_5561 ( .C (clk), .D (plaintext_s0[105]), .Q (new_AGEMA_signal_11413) ) ;
    buf_clk new_AGEMA_reg_buffer_5565 ( .C (clk), .D (plaintext_s1[105]), .Q (new_AGEMA_signal_11417) ) ;
    buf_clk new_AGEMA_reg_buffer_5569 ( .C (clk), .D (plaintext_s0[106]), .Q (new_AGEMA_signal_11421) ) ;
    buf_clk new_AGEMA_reg_buffer_5573 ( .C (clk), .D (plaintext_s1[106]), .Q (new_AGEMA_signal_11425) ) ;
    buf_clk new_AGEMA_reg_buffer_5577 ( .C (clk), .D (plaintext_s0[107]), .Q (new_AGEMA_signal_11429) ) ;
    buf_clk new_AGEMA_reg_buffer_5581 ( .C (clk), .D (plaintext_s1[107]), .Q (new_AGEMA_signal_11433) ) ;
    buf_clk new_AGEMA_reg_buffer_5585 ( .C (clk), .D (plaintext_s0[108]), .Q (new_AGEMA_signal_11437) ) ;
    buf_clk new_AGEMA_reg_buffer_5589 ( .C (clk), .D (plaintext_s1[108]), .Q (new_AGEMA_signal_11441) ) ;
    buf_clk new_AGEMA_reg_buffer_5593 ( .C (clk), .D (plaintext_s0[109]), .Q (new_AGEMA_signal_11445) ) ;
    buf_clk new_AGEMA_reg_buffer_5597 ( .C (clk), .D (plaintext_s1[109]), .Q (new_AGEMA_signal_11449) ) ;
    buf_clk new_AGEMA_reg_buffer_5601 ( .C (clk), .D (plaintext_s0[110]), .Q (new_AGEMA_signal_11453) ) ;
    buf_clk new_AGEMA_reg_buffer_5605 ( .C (clk), .D (plaintext_s1[110]), .Q (new_AGEMA_signal_11457) ) ;
    buf_clk new_AGEMA_reg_buffer_5609 ( .C (clk), .D (plaintext_s0[111]), .Q (new_AGEMA_signal_11461) ) ;
    buf_clk new_AGEMA_reg_buffer_5613 ( .C (clk), .D (plaintext_s1[111]), .Q (new_AGEMA_signal_11465) ) ;
    buf_clk new_AGEMA_reg_buffer_5617 ( .C (clk), .D (plaintext_s0[112]), .Q (new_AGEMA_signal_11469) ) ;
    buf_clk new_AGEMA_reg_buffer_5621 ( .C (clk), .D (plaintext_s1[112]), .Q (new_AGEMA_signal_11473) ) ;
    buf_clk new_AGEMA_reg_buffer_5625 ( .C (clk), .D (plaintext_s0[113]), .Q (new_AGEMA_signal_11477) ) ;
    buf_clk new_AGEMA_reg_buffer_5629 ( .C (clk), .D (plaintext_s1[113]), .Q (new_AGEMA_signal_11481) ) ;
    buf_clk new_AGEMA_reg_buffer_5633 ( .C (clk), .D (plaintext_s0[114]), .Q (new_AGEMA_signal_11485) ) ;
    buf_clk new_AGEMA_reg_buffer_5637 ( .C (clk), .D (plaintext_s1[114]), .Q (new_AGEMA_signal_11489) ) ;
    buf_clk new_AGEMA_reg_buffer_5641 ( .C (clk), .D (plaintext_s0[115]), .Q (new_AGEMA_signal_11493) ) ;
    buf_clk new_AGEMA_reg_buffer_5645 ( .C (clk), .D (plaintext_s1[115]), .Q (new_AGEMA_signal_11497) ) ;
    buf_clk new_AGEMA_reg_buffer_5649 ( .C (clk), .D (plaintext_s0[116]), .Q (new_AGEMA_signal_11501) ) ;
    buf_clk new_AGEMA_reg_buffer_5653 ( .C (clk), .D (plaintext_s1[116]), .Q (new_AGEMA_signal_11505) ) ;
    buf_clk new_AGEMA_reg_buffer_5657 ( .C (clk), .D (plaintext_s0[117]), .Q (new_AGEMA_signal_11509) ) ;
    buf_clk new_AGEMA_reg_buffer_5661 ( .C (clk), .D (plaintext_s1[117]), .Q (new_AGEMA_signal_11513) ) ;
    buf_clk new_AGEMA_reg_buffer_5665 ( .C (clk), .D (plaintext_s0[118]), .Q (new_AGEMA_signal_11517) ) ;
    buf_clk new_AGEMA_reg_buffer_5669 ( .C (clk), .D (plaintext_s1[118]), .Q (new_AGEMA_signal_11521) ) ;
    buf_clk new_AGEMA_reg_buffer_5673 ( .C (clk), .D (plaintext_s0[119]), .Q (new_AGEMA_signal_11525) ) ;
    buf_clk new_AGEMA_reg_buffer_5677 ( .C (clk), .D (plaintext_s1[119]), .Q (new_AGEMA_signal_11529) ) ;
    buf_clk new_AGEMA_reg_buffer_5681 ( .C (clk), .D (plaintext_s0[120]), .Q (new_AGEMA_signal_11533) ) ;
    buf_clk new_AGEMA_reg_buffer_5685 ( .C (clk), .D (plaintext_s1[120]), .Q (new_AGEMA_signal_11537) ) ;
    buf_clk new_AGEMA_reg_buffer_5689 ( .C (clk), .D (plaintext_s0[121]), .Q (new_AGEMA_signal_11541) ) ;
    buf_clk new_AGEMA_reg_buffer_5693 ( .C (clk), .D (plaintext_s1[121]), .Q (new_AGEMA_signal_11545) ) ;
    buf_clk new_AGEMA_reg_buffer_5697 ( .C (clk), .D (plaintext_s0[122]), .Q (new_AGEMA_signal_11549) ) ;
    buf_clk new_AGEMA_reg_buffer_5701 ( .C (clk), .D (plaintext_s1[122]), .Q (new_AGEMA_signal_11553) ) ;
    buf_clk new_AGEMA_reg_buffer_5705 ( .C (clk), .D (plaintext_s0[123]), .Q (new_AGEMA_signal_11557) ) ;
    buf_clk new_AGEMA_reg_buffer_5709 ( .C (clk), .D (plaintext_s1[123]), .Q (new_AGEMA_signal_11561) ) ;
    buf_clk new_AGEMA_reg_buffer_5713 ( .C (clk), .D (plaintext_s0[124]), .Q (new_AGEMA_signal_11565) ) ;
    buf_clk new_AGEMA_reg_buffer_5717 ( .C (clk), .D (plaintext_s1[124]), .Q (new_AGEMA_signal_11569) ) ;
    buf_clk new_AGEMA_reg_buffer_5721 ( .C (clk), .D (plaintext_s0[125]), .Q (new_AGEMA_signal_11573) ) ;
    buf_clk new_AGEMA_reg_buffer_5725 ( .C (clk), .D (plaintext_s1[125]), .Q (new_AGEMA_signal_11577) ) ;
    buf_clk new_AGEMA_reg_buffer_5729 ( .C (clk), .D (plaintext_s0[126]), .Q (new_AGEMA_signal_11581) ) ;
    buf_clk new_AGEMA_reg_buffer_5733 ( .C (clk), .D (plaintext_s1[126]), .Q (new_AGEMA_signal_11585) ) ;
    buf_clk new_AGEMA_reg_buffer_5737 ( .C (clk), .D (plaintext_s0[127]), .Q (new_AGEMA_signal_11589) ) ;
    buf_clk new_AGEMA_reg_buffer_5741 ( .C (clk), .D (plaintext_s1[127]), .Q (new_AGEMA_signal_11593) ) ;
    buf_clk new_AGEMA_reg_buffer_5745 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T6), .Q (new_AGEMA_signal_11597) ) ;
    buf_clk new_AGEMA_reg_buffer_5748 ( .C (clk), .D (new_AGEMA_signal_5165), .Q (new_AGEMA_signal_11600) ) ;
    buf_clk new_AGEMA_reg_buffer_5751 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T8), .Q (new_AGEMA_signal_11603) ) ;
    buf_clk new_AGEMA_reg_buffer_5754 ( .C (clk), .D (new_AGEMA_signal_5345), .Q (new_AGEMA_signal_11606) ) ;
    buf_clk new_AGEMA_reg_buffer_5757 ( .C (clk), .D (ciphertext_s0[0]), .Q (new_AGEMA_signal_11609) ) ;
    buf_clk new_AGEMA_reg_buffer_5760 ( .C (clk), .D (ciphertext_s1[0]), .Q (new_AGEMA_signal_11612) ) ;
    buf_clk new_AGEMA_reg_buffer_5763 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T16), .Q (new_AGEMA_signal_11615) ) ;
    buf_clk new_AGEMA_reg_buffer_5766 ( .C (clk), .D (new_AGEMA_signal_5169), .Q (new_AGEMA_signal_11618) ) ;
    buf_clk new_AGEMA_reg_buffer_5769 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T9), .Q (new_AGEMA_signal_11621) ) ;
    buf_clk new_AGEMA_reg_buffer_5772 ( .C (clk), .D (new_AGEMA_signal_5166), .Q (new_AGEMA_signal_11624) ) ;
    buf_clk new_AGEMA_reg_buffer_5775 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T17), .Q (new_AGEMA_signal_11627) ) ;
    buf_clk new_AGEMA_reg_buffer_5778 ( .C (clk), .D (new_AGEMA_signal_5348), .Q (new_AGEMA_signal_11630) ) ;
    buf_clk new_AGEMA_reg_buffer_5781 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T15), .Q (new_AGEMA_signal_11633) ) ;
    buf_clk new_AGEMA_reg_buffer_5784 ( .C (clk), .D (new_AGEMA_signal_5168), .Q (new_AGEMA_signal_11636) ) ;
    buf_clk new_AGEMA_reg_buffer_5787 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T27), .Q (new_AGEMA_signal_11639) ) ;
    buf_clk new_AGEMA_reg_buffer_5790 ( .C (clk), .D (new_AGEMA_signal_5172), .Q (new_AGEMA_signal_11642) ) ;
    buf_clk new_AGEMA_reg_buffer_5793 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T10), .Q (new_AGEMA_signal_11645) ) ;
    buf_clk new_AGEMA_reg_buffer_5796 ( .C (clk), .D (new_AGEMA_signal_5346), .Q (new_AGEMA_signal_11648) ) ;
    buf_clk new_AGEMA_reg_buffer_5799 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T13), .Q (new_AGEMA_signal_11651) ) ;
    buf_clk new_AGEMA_reg_buffer_5802 ( .C (clk), .D (new_AGEMA_signal_5167), .Q (new_AGEMA_signal_11654) ) ;
    buf_clk new_AGEMA_reg_buffer_5805 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T23), .Q (new_AGEMA_signal_11657) ) ;
    buf_clk new_AGEMA_reg_buffer_5808 ( .C (clk), .D (new_AGEMA_signal_5350), .Q (new_AGEMA_signal_11660) ) ;
    buf_clk new_AGEMA_reg_buffer_5811 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T19), .Q (new_AGEMA_signal_11663) ) ;
    buf_clk new_AGEMA_reg_buffer_5814 ( .C (clk), .D (new_AGEMA_signal_5170), .Q (new_AGEMA_signal_11666) ) ;
    buf_clk new_AGEMA_reg_buffer_5817 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T3), .Q (new_AGEMA_signal_11669) ) ;
    buf_clk new_AGEMA_reg_buffer_5820 ( .C (clk), .D (new_AGEMA_signal_4975), .Q (new_AGEMA_signal_11672) ) ;
    buf_clk new_AGEMA_reg_buffer_5823 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T22), .Q (new_AGEMA_signal_11675) ) ;
    buf_clk new_AGEMA_reg_buffer_5826 ( .C (clk), .D (new_AGEMA_signal_5171), .Q (new_AGEMA_signal_11678) ) ;
    buf_clk new_AGEMA_reg_buffer_5829 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T20), .Q (new_AGEMA_signal_11681) ) ;
    buf_clk new_AGEMA_reg_buffer_5832 ( .C (clk), .D (new_AGEMA_signal_5349), .Q (new_AGEMA_signal_11684) ) ;
    buf_clk new_AGEMA_reg_buffer_5835 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T1), .Q (new_AGEMA_signal_11687) ) ;
    buf_clk new_AGEMA_reg_buffer_5838 ( .C (clk), .D (new_AGEMA_signal_4973), .Q (new_AGEMA_signal_11690) ) ;
    buf_clk new_AGEMA_reg_buffer_5841 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T4), .Q (new_AGEMA_signal_11693) ) ;
    buf_clk new_AGEMA_reg_buffer_5844 ( .C (clk), .D (new_AGEMA_signal_4976), .Q (new_AGEMA_signal_11696) ) ;
    buf_clk new_AGEMA_reg_buffer_5847 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T2), .Q (new_AGEMA_signal_11699) ) ;
    buf_clk new_AGEMA_reg_buffer_5850 ( .C (clk), .D (new_AGEMA_signal_4974), .Q (new_AGEMA_signal_11702) ) ;
    buf_clk new_AGEMA_reg_buffer_5853 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T6), .Q (new_AGEMA_signal_11705) ) ;
    buf_clk new_AGEMA_reg_buffer_5856 ( .C (clk), .D (new_AGEMA_signal_5173), .Q (new_AGEMA_signal_11708) ) ;
    buf_clk new_AGEMA_reg_buffer_5859 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T8), .Q (new_AGEMA_signal_11711) ) ;
    buf_clk new_AGEMA_reg_buffer_5862 ( .C (clk), .D (new_AGEMA_signal_5358), .Q (new_AGEMA_signal_11714) ) ;
    buf_clk new_AGEMA_reg_buffer_5865 ( .C (clk), .D (ciphertext_s0[8]), .Q (new_AGEMA_signal_11717) ) ;
    buf_clk new_AGEMA_reg_buffer_5868 ( .C (clk), .D (ciphertext_s1[8]), .Q (new_AGEMA_signal_11720) ) ;
    buf_clk new_AGEMA_reg_buffer_5871 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T16), .Q (new_AGEMA_signal_11723) ) ;
    buf_clk new_AGEMA_reg_buffer_5874 ( .C (clk), .D (new_AGEMA_signal_5177), .Q (new_AGEMA_signal_11726) ) ;
    buf_clk new_AGEMA_reg_buffer_5877 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T9), .Q (new_AGEMA_signal_11729) ) ;
    buf_clk new_AGEMA_reg_buffer_5880 ( .C (clk), .D (new_AGEMA_signal_5174), .Q (new_AGEMA_signal_11732) ) ;
    buf_clk new_AGEMA_reg_buffer_5883 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T17), .Q (new_AGEMA_signal_11735) ) ;
    buf_clk new_AGEMA_reg_buffer_5886 ( .C (clk), .D (new_AGEMA_signal_5361), .Q (new_AGEMA_signal_11738) ) ;
    buf_clk new_AGEMA_reg_buffer_5889 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T15), .Q (new_AGEMA_signal_11741) ) ;
    buf_clk new_AGEMA_reg_buffer_5892 ( .C (clk), .D (new_AGEMA_signal_5176), .Q (new_AGEMA_signal_11744) ) ;
    buf_clk new_AGEMA_reg_buffer_5895 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T27), .Q (new_AGEMA_signal_11747) ) ;
    buf_clk new_AGEMA_reg_buffer_5898 ( .C (clk), .D (new_AGEMA_signal_5180), .Q (new_AGEMA_signal_11750) ) ;
    buf_clk new_AGEMA_reg_buffer_5901 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T10), .Q (new_AGEMA_signal_11753) ) ;
    buf_clk new_AGEMA_reg_buffer_5904 ( .C (clk), .D (new_AGEMA_signal_5359), .Q (new_AGEMA_signal_11756) ) ;
    buf_clk new_AGEMA_reg_buffer_5907 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T13), .Q (new_AGEMA_signal_11759) ) ;
    buf_clk new_AGEMA_reg_buffer_5910 ( .C (clk), .D (new_AGEMA_signal_5175), .Q (new_AGEMA_signal_11762) ) ;
    buf_clk new_AGEMA_reg_buffer_5913 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T23), .Q (new_AGEMA_signal_11765) ) ;
    buf_clk new_AGEMA_reg_buffer_5916 ( .C (clk), .D (new_AGEMA_signal_5363), .Q (new_AGEMA_signal_11768) ) ;
    buf_clk new_AGEMA_reg_buffer_5919 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T19), .Q (new_AGEMA_signal_11771) ) ;
    buf_clk new_AGEMA_reg_buffer_5922 ( .C (clk), .D (new_AGEMA_signal_5178), .Q (new_AGEMA_signal_11774) ) ;
    buf_clk new_AGEMA_reg_buffer_5925 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T3), .Q (new_AGEMA_signal_11777) ) ;
    buf_clk new_AGEMA_reg_buffer_5928 ( .C (clk), .D (new_AGEMA_signal_4985), .Q (new_AGEMA_signal_11780) ) ;
    buf_clk new_AGEMA_reg_buffer_5931 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T22), .Q (new_AGEMA_signal_11783) ) ;
    buf_clk new_AGEMA_reg_buffer_5934 ( .C (clk), .D (new_AGEMA_signal_5179), .Q (new_AGEMA_signal_11786) ) ;
    buf_clk new_AGEMA_reg_buffer_5937 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T20), .Q (new_AGEMA_signal_11789) ) ;
    buf_clk new_AGEMA_reg_buffer_5940 ( .C (clk), .D (new_AGEMA_signal_5362), .Q (new_AGEMA_signal_11792) ) ;
    buf_clk new_AGEMA_reg_buffer_5943 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T1), .Q (new_AGEMA_signal_11795) ) ;
    buf_clk new_AGEMA_reg_buffer_5946 ( .C (clk), .D (new_AGEMA_signal_4983), .Q (new_AGEMA_signal_11798) ) ;
    buf_clk new_AGEMA_reg_buffer_5949 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T4), .Q (new_AGEMA_signal_11801) ) ;
    buf_clk new_AGEMA_reg_buffer_5952 ( .C (clk), .D (new_AGEMA_signal_4986), .Q (new_AGEMA_signal_11804) ) ;
    buf_clk new_AGEMA_reg_buffer_5955 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T2), .Q (new_AGEMA_signal_11807) ) ;
    buf_clk new_AGEMA_reg_buffer_5958 ( .C (clk), .D (new_AGEMA_signal_4984), .Q (new_AGEMA_signal_11810) ) ;
    buf_clk new_AGEMA_reg_buffer_5961 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T6), .Q (new_AGEMA_signal_11813) ) ;
    buf_clk new_AGEMA_reg_buffer_5964 ( .C (clk), .D (new_AGEMA_signal_5181), .Q (new_AGEMA_signal_11816) ) ;
    buf_clk new_AGEMA_reg_buffer_5967 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T8), .Q (new_AGEMA_signal_11819) ) ;
    buf_clk new_AGEMA_reg_buffer_5970 ( .C (clk), .D (new_AGEMA_signal_5371), .Q (new_AGEMA_signal_11822) ) ;
    buf_clk new_AGEMA_reg_buffer_5973 ( .C (clk), .D (ciphertext_s0[16]), .Q (new_AGEMA_signal_11825) ) ;
    buf_clk new_AGEMA_reg_buffer_5976 ( .C (clk), .D (ciphertext_s1[16]), .Q (new_AGEMA_signal_11828) ) ;
    buf_clk new_AGEMA_reg_buffer_5979 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T16), .Q (new_AGEMA_signal_11831) ) ;
    buf_clk new_AGEMA_reg_buffer_5982 ( .C (clk), .D (new_AGEMA_signal_5185), .Q (new_AGEMA_signal_11834) ) ;
    buf_clk new_AGEMA_reg_buffer_5985 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T9), .Q (new_AGEMA_signal_11837) ) ;
    buf_clk new_AGEMA_reg_buffer_5988 ( .C (clk), .D (new_AGEMA_signal_5182), .Q (new_AGEMA_signal_11840) ) ;
    buf_clk new_AGEMA_reg_buffer_5991 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T17), .Q (new_AGEMA_signal_11843) ) ;
    buf_clk new_AGEMA_reg_buffer_5994 ( .C (clk), .D (new_AGEMA_signal_5374), .Q (new_AGEMA_signal_11846) ) ;
    buf_clk new_AGEMA_reg_buffer_5997 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T15), .Q (new_AGEMA_signal_11849) ) ;
    buf_clk new_AGEMA_reg_buffer_6000 ( .C (clk), .D (new_AGEMA_signal_5184), .Q (new_AGEMA_signal_11852) ) ;
    buf_clk new_AGEMA_reg_buffer_6003 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T27), .Q (new_AGEMA_signal_11855) ) ;
    buf_clk new_AGEMA_reg_buffer_6006 ( .C (clk), .D (new_AGEMA_signal_5188), .Q (new_AGEMA_signal_11858) ) ;
    buf_clk new_AGEMA_reg_buffer_6009 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T10), .Q (new_AGEMA_signal_11861) ) ;
    buf_clk new_AGEMA_reg_buffer_6012 ( .C (clk), .D (new_AGEMA_signal_5372), .Q (new_AGEMA_signal_11864) ) ;
    buf_clk new_AGEMA_reg_buffer_6015 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T13), .Q (new_AGEMA_signal_11867) ) ;
    buf_clk new_AGEMA_reg_buffer_6018 ( .C (clk), .D (new_AGEMA_signal_5183), .Q (new_AGEMA_signal_11870) ) ;
    buf_clk new_AGEMA_reg_buffer_6021 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T23), .Q (new_AGEMA_signal_11873) ) ;
    buf_clk new_AGEMA_reg_buffer_6024 ( .C (clk), .D (new_AGEMA_signal_5376), .Q (new_AGEMA_signal_11876) ) ;
    buf_clk new_AGEMA_reg_buffer_6027 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T19), .Q (new_AGEMA_signal_11879) ) ;
    buf_clk new_AGEMA_reg_buffer_6030 ( .C (clk), .D (new_AGEMA_signal_5186), .Q (new_AGEMA_signal_11882) ) ;
    buf_clk new_AGEMA_reg_buffer_6033 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T3), .Q (new_AGEMA_signal_11885) ) ;
    buf_clk new_AGEMA_reg_buffer_6036 ( .C (clk), .D (new_AGEMA_signal_4995), .Q (new_AGEMA_signal_11888) ) ;
    buf_clk new_AGEMA_reg_buffer_6039 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T22), .Q (new_AGEMA_signal_11891) ) ;
    buf_clk new_AGEMA_reg_buffer_6042 ( .C (clk), .D (new_AGEMA_signal_5187), .Q (new_AGEMA_signal_11894) ) ;
    buf_clk new_AGEMA_reg_buffer_6045 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T20), .Q (new_AGEMA_signal_11897) ) ;
    buf_clk new_AGEMA_reg_buffer_6048 ( .C (clk), .D (new_AGEMA_signal_5375), .Q (new_AGEMA_signal_11900) ) ;
    buf_clk new_AGEMA_reg_buffer_6051 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T1), .Q (new_AGEMA_signal_11903) ) ;
    buf_clk new_AGEMA_reg_buffer_6054 ( .C (clk), .D (new_AGEMA_signal_4993), .Q (new_AGEMA_signal_11906) ) ;
    buf_clk new_AGEMA_reg_buffer_6057 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T4), .Q (new_AGEMA_signal_11909) ) ;
    buf_clk new_AGEMA_reg_buffer_6060 ( .C (clk), .D (new_AGEMA_signal_4996), .Q (new_AGEMA_signal_11912) ) ;
    buf_clk new_AGEMA_reg_buffer_6063 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T2), .Q (new_AGEMA_signal_11915) ) ;
    buf_clk new_AGEMA_reg_buffer_6066 ( .C (clk), .D (new_AGEMA_signal_4994), .Q (new_AGEMA_signal_11918) ) ;
    buf_clk new_AGEMA_reg_buffer_6069 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T6), .Q (new_AGEMA_signal_11921) ) ;
    buf_clk new_AGEMA_reg_buffer_6072 ( .C (clk), .D (new_AGEMA_signal_5189), .Q (new_AGEMA_signal_11924) ) ;
    buf_clk new_AGEMA_reg_buffer_6075 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T8), .Q (new_AGEMA_signal_11927) ) ;
    buf_clk new_AGEMA_reg_buffer_6078 ( .C (clk), .D (new_AGEMA_signal_5384), .Q (new_AGEMA_signal_11930) ) ;
    buf_clk new_AGEMA_reg_buffer_6081 ( .C (clk), .D (ciphertext_s0[24]), .Q (new_AGEMA_signal_11933) ) ;
    buf_clk new_AGEMA_reg_buffer_6084 ( .C (clk), .D (ciphertext_s1[24]), .Q (new_AGEMA_signal_11936) ) ;
    buf_clk new_AGEMA_reg_buffer_6087 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T16), .Q (new_AGEMA_signal_11939) ) ;
    buf_clk new_AGEMA_reg_buffer_6090 ( .C (clk), .D (new_AGEMA_signal_5193), .Q (new_AGEMA_signal_11942) ) ;
    buf_clk new_AGEMA_reg_buffer_6093 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T9), .Q (new_AGEMA_signal_11945) ) ;
    buf_clk new_AGEMA_reg_buffer_6096 ( .C (clk), .D (new_AGEMA_signal_5190), .Q (new_AGEMA_signal_11948) ) ;
    buf_clk new_AGEMA_reg_buffer_6099 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T17), .Q (new_AGEMA_signal_11951) ) ;
    buf_clk new_AGEMA_reg_buffer_6102 ( .C (clk), .D (new_AGEMA_signal_5387), .Q (new_AGEMA_signal_11954) ) ;
    buf_clk new_AGEMA_reg_buffer_6105 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T15), .Q (new_AGEMA_signal_11957) ) ;
    buf_clk new_AGEMA_reg_buffer_6108 ( .C (clk), .D (new_AGEMA_signal_5192), .Q (new_AGEMA_signal_11960) ) ;
    buf_clk new_AGEMA_reg_buffer_6111 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T27), .Q (new_AGEMA_signal_11963) ) ;
    buf_clk new_AGEMA_reg_buffer_6114 ( .C (clk), .D (new_AGEMA_signal_5196), .Q (new_AGEMA_signal_11966) ) ;
    buf_clk new_AGEMA_reg_buffer_6117 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T10), .Q (new_AGEMA_signal_11969) ) ;
    buf_clk new_AGEMA_reg_buffer_6120 ( .C (clk), .D (new_AGEMA_signal_5385), .Q (new_AGEMA_signal_11972) ) ;
    buf_clk new_AGEMA_reg_buffer_6123 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T13), .Q (new_AGEMA_signal_11975) ) ;
    buf_clk new_AGEMA_reg_buffer_6126 ( .C (clk), .D (new_AGEMA_signal_5191), .Q (new_AGEMA_signal_11978) ) ;
    buf_clk new_AGEMA_reg_buffer_6129 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T23), .Q (new_AGEMA_signal_11981) ) ;
    buf_clk new_AGEMA_reg_buffer_6132 ( .C (clk), .D (new_AGEMA_signal_5389), .Q (new_AGEMA_signal_11984) ) ;
    buf_clk new_AGEMA_reg_buffer_6135 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T19), .Q (new_AGEMA_signal_11987) ) ;
    buf_clk new_AGEMA_reg_buffer_6138 ( .C (clk), .D (new_AGEMA_signal_5194), .Q (new_AGEMA_signal_11990) ) ;
    buf_clk new_AGEMA_reg_buffer_6141 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T3), .Q (new_AGEMA_signal_11993) ) ;
    buf_clk new_AGEMA_reg_buffer_6144 ( .C (clk), .D (new_AGEMA_signal_5005), .Q (new_AGEMA_signal_11996) ) ;
    buf_clk new_AGEMA_reg_buffer_6147 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T22), .Q (new_AGEMA_signal_11999) ) ;
    buf_clk new_AGEMA_reg_buffer_6150 ( .C (clk), .D (new_AGEMA_signal_5195), .Q (new_AGEMA_signal_12002) ) ;
    buf_clk new_AGEMA_reg_buffer_6153 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T20), .Q (new_AGEMA_signal_12005) ) ;
    buf_clk new_AGEMA_reg_buffer_6156 ( .C (clk), .D (new_AGEMA_signal_5388), .Q (new_AGEMA_signal_12008) ) ;
    buf_clk new_AGEMA_reg_buffer_6159 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T1), .Q (new_AGEMA_signal_12011) ) ;
    buf_clk new_AGEMA_reg_buffer_6162 ( .C (clk), .D (new_AGEMA_signal_5003), .Q (new_AGEMA_signal_12014) ) ;
    buf_clk new_AGEMA_reg_buffer_6165 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T4), .Q (new_AGEMA_signal_12017) ) ;
    buf_clk new_AGEMA_reg_buffer_6168 ( .C (clk), .D (new_AGEMA_signal_5006), .Q (new_AGEMA_signal_12020) ) ;
    buf_clk new_AGEMA_reg_buffer_6171 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T2), .Q (new_AGEMA_signal_12023) ) ;
    buf_clk new_AGEMA_reg_buffer_6174 ( .C (clk), .D (new_AGEMA_signal_5004), .Q (new_AGEMA_signal_12026) ) ;
    buf_clk new_AGEMA_reg_buffer_6177 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T6), .Q (new_AGEMA_signal_12029) ) ;
    buf_clk new_AGEMA_reg_buffer_6180 ( .C (clk), .D (new_AGEMA_signal_5197), .Q (new_AGEMA_signal_12032) ) ;
    buf_clk new_AGEMA_reg_buffer_6183 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T8), .Q (new_AGEMA_signal_12035) ) ;
    buf_clk new_AGEMA_reg_buffer_6186 ( .C (clk), .D (new_AGEMA_signal_5397), .Q (new_AGEMA_signal_12038) ) ;
    buf_clk new_AGEMA_reg_buffer_6189 ( .C (clk), .D (ciphertext_s0[32]), .Q (new_AGEMA_signal_12041) ) ;
    buf_clk new_AGEMA_reg_buffer_6192 ( .C (clk), .D (ciphertext_s1[32]), .Q (new_AGEMA_signal_12044) ) ;
    buf_clk new_AGEMA_reg_buffer_6195 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T16), .Q (new_AGEMA_signal_12047) ) ;
    buf_clk new_AGEMA_reg_buffer_6198 ( .C (clk), .D (new_AGEMA_signal_5201), .Q (new_AGEMA_signal_12050) ) ;
    buf_clk new_AGEMA_reg_buffer_6201 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T9), .Q (new_AGEMA_signal_12053) ) ;
    buf_clk new_AGEMA_reg_buffer_6204 ( .C (clk), .D (new_AGEMA_signal_5198), .Q (new_AGEMA_signal_12056) ) ;
    buf_clk new_AGEMA_reg_buffer_6207 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T17), .Q (new_AGEMA_signal_12059) ) ;
    buf_clk new_AGEMA_reg_buffer_6210 ( .C (clk), .D (new_AGEMA_signal_5400), .Q (new_AGEMA_signal_12062) ) ;
    buf_clk new_AGEMA_reg_buffer_6213 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T15), .Q (new_AGEMA_signal_12065) ) ;
    buf_clk new_AGEMA_reg_buffer_6216 ( .C (clk), .D (new_AGEMA_signal_5200), .Q (new_AGEMA_signal_12068) ) ;
    buf_clk new_AGEMA_reg_buffer_6219 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T27), .Q (new_AGEMA_signal_12071) ) ;
    buf_clk new_AGEMA_reg_buffer_6222 ( .C (clk), .D (new_AGEMA_signal_5204), .Q (new_AGEMA_signal_12074) ) ;
    buf_clk new_AGEMA_reg_buffer_6225 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T10), .Q (new_AGEMA_signal_12077) ) ;
    buf_clk new_AGEMA_reg_buffer_6228 ( .C (clk), .D (new_AGEMA_signal_5398), .Q (new_AGEMA_signal_12080) ) ;
    buf_clk new_AGEMA_reg_buffer_6231 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T13), .Q (new_AGEMA_signal_12083) ) ;
    buf_clk new_AGEMA_reg_buffer_6234 ( .C (clk), .D (new_AGEMA_signal_5199), .Q (new_AGEMA_signal_12086) ) ;
    buf_clk new_AGEMA_reg_buffer_6237 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T23), .Q (new_AGEMA_signal_12089) ) ;
    buf_clk new_AGEMA_reg_buffer_6240 ( .C (clk), .D (new_AGEMA_signal_5402), .Q (new_AGEMA_signal_12092) ) ;
    buf_clk new_AGEMA_reg_buffer_6243 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T19), .Q (new_AGEMA_signal_12095) ) ;
    buf_clk new_AGEMA_reg_buffer_6246 ( .C (clk), .D (new_AGEMA_signal_5202), .Q (new_AGEMA_signal_12098) ) ;
    buf_clk new_AGEMA_reg_buffer_6249 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T3), .Q (new_AGEMA_signal_12101) ) ;
    buf_clk new_AGEMA_reg_buffer_6252 ( .C (clk), .D (new_AGEMA_signal_5015), .Q (new_AGEMA_signal_12104) ) ;
    buf_clk new_AGEMA_reg_buffer_6255 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T22), .Q (new_AGEMA_signal_12107) ) ;
    buf_clk new_AGEMA_reg_buffer_6258 ( .C (clk), .D (new_AGEMA_signal_5203), .Q (new_AGEMA_signal_12110) ) ;
    buf_clk new_AGEMA_reg_buffer_6261 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T20), .Q (new_AGEMA_signal_12113) ) ;
    buf_clk new_AGEMA_reg_buffer_6264 ( .C (clk), .D (new_AGEMA_signal_5401), .Q (new_AGEMA_signal_12116) ) ;
    buf_clk new_AGEMA_reg_buffer_6267 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T1), .Q (new_AGEMA_signal_12119) ) ;
    buf_clk new_AGEMA_reg_buffer_6270 ( .C (clk), .D (new_AGEMA_signal_5013), .Q (new_AGEMA_signal_12122) ) ;
    buf_clk new_AGEMA_reg_buffer_6273 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T4), .Q (new_AGEMA_signal_12125) ) ;
    buf_clk new_AGEMA_reg_buffer_6276 ( .C (clk), .D (new_AGEMA_signal_5016), .Q (new_AGEMA_signal_12128) ) ;
    buf_clk new_AGEMA_reg_buffer_6279 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T2), .Q (new_AGEMA_signal_12131) ) ;
    buf_clk new_AGEMA_reg_buffer_6282 ( .C (clk), .D (new_AGEMA_signal_5014), .Q (new_AGEMA_signal_12134) ) ;
    buf_clk new_AGEMA_reg_buffer_6285 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T6), .Q (new_AGEMA_signal_12137) ) ;
    buf_clk new_AGEMA_reg_buffer_6288 ( .C (clk), .D (new_AGEMA_signal_5205), .Q (new_AGEMA_signal_12140) ) ;
    buf_clk new_AGEMA_reg_buffer_6291 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T8), .Q (new_AGEMA_signal_12143) ) ;
    buf_clk new_AGEMA_reg_buffer_6294 ( .C (clk), .D (new_AGEMA_signal_5410), .Q (new_AGEMA_signal_12146) ) ;
    buf_clk new_AGEMA_reg_buffer_6297 ( .C (clk), .D (ciphertext_s0[40]), .Q (new_AGEMA_signal_12149) ) ;
    buf_clk new_AGEMA_reg_buffer_6300 ( .C (clk), .D (ciphertext_s1[40]), .Q (new_AGEMA_signal_12152) ) ;
    buf_clk new_AGEMA_reg_buffer_6303 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T16), .Q (new_AGEMA_signal_12155) ) ;
    buf_clk new_AGEMA_reg_buffer_6306 ( .C (clk), .D (new_AGEMA_signal_5209), .Q (new_AGEMA_signal_12158) ) ;
    buf_clk new_AGEMA_reg_buffer_6309 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T9), .Q (new_AGEMA_signal_12161) ) ;
    buf_clk new_AGEMA_reg_buffer_6312 ( .C (clk), .D (new_AGEMA_signal_5206), .Q (new_AGEMA_signal_12164) ) ;
    buf_clk new_AGEMA_reg_buffer_6315 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T17), .Q (new_AGEMA_signal_12167) ) ;
    buf_clk new_AGEMA_reg_buffer_6318 ( .C (clk), .D (new_AGEMA_signal_5413), .Q (new_AGEMA_signal_12170) ) ;
    buf_clk new_AGEMA_reg_buffer_6321 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T15), .Q (new_AGEMA_signal_12173) ) ;
    buf_clk new_AGEMA_reg_buffer_6324 ( .C (clk), .D (new_AGEMA_signal_5208), .Q (new_AGEMA_signal_12176) ) ;
    buf_clk new_AGEMA_reg_buffer_6327 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T27), .Q (new_AGEMA_signal_12179) ) ;
    buf_clk new_AGEMA_reg_buffer_6330 ( .C (clk), .D (new_AGEMA_signal_5212), .Q (new_AGEMA_signal_12182) ) ;
    buf_clk new_AGEMA_reg_buffer_6333 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T10), .Q (new_AGEMA_signal_12185) ) ;
    buf_clk new_AGEMA_reg_buffer_6336 ( .C (clk), .D (new_AGEMA_signal_5411), .Q (new_AGEMA_signal_12188) ) ;
    buf_clk new_AGEMA_reg_buffer_6339 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T13), .Q (new_AGEMA_signal_12191) ) ;
    buf_clk new_AGEMA_reg_buffer_6342 ( .C (clk), .D (new_AGEMA_signal_5207), .Q (new_AGEMA_signal_12194) ) ;
    buf_clk new_AGEMA_reg_buffer_6345 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T23), .Q (new_AGEMA_signal_12197) ) ;
    buf_clk new_AGEMA_reg_buffer_6348 ( .C (clk), .D (new_AGEMA_signal_5415), .Q (new_AGEMA_signal_12200) ) ;
    buf_clk new_AGEMA_reg_buffer_6351 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T19), .Q (new_AGEMA_signal_12203) ) ;
    buf_clk new_AGEMA_reg_buffer_6354 ( .C (clk), .D (new_AGEMA_signal_5210), .Q (new_AGEMA_signal_12206) ) ;
    buf_clk new_AGEMA_reg_buffer_6357 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T3), .Q (new_AGEMA_signal_12209) ) ;
    buf_clk new_AGEMA_reg_buffer_6360 ( .C (clk), .D (new_AGEMA_signal_5025), .Q (new_AGEMA_signal_12212) ) ;
    buf_clk new_AGEMA_reg_buffer_6363 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T22), .Q (new_AGEMA_signal_12215) ) ;
    buf_clk new_AGEMA_reg_buffer_6366 ( .C (clk), .D (new_AGEMA_signal_5211), .Q (new_AGEMA_signal_12218) ) ;
    buf_clk new_AGEMA_reg_buffer_6369 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T20), .Q (new_AGEMA_signal_12221) ) ;
    buf_clk new_AGEMA_reg_buffer_6372 ( .C (clk), .D (new_AGEMA_signal_5414), .Q (new_AGEMA_signal_12224) ) ;
    buf_clk new_AGEMA_reg_buffer_6375 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T1), .Q (new_AGEMA_signal_12227) ) ;
    buf_clk new_AGEMA_reg_buffer_6378 ( .C (clk), .D (new_AGEMA_signal_5023), .Q (new_AGEMA_signal_12230) ) ;
    buf_clk new_AGEMA_reg_buffer_6381 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T4), .Q (new_AGEMA_signal_12233) ) ;
    buf_clk new_AGEMA_reg_buffer_6384 ( .C (clk), .D (new_AGEMA_signal_5026), .Q (new_AGEMA_signal_12236) ) ;
    buf_clk new_AGEMA_reg_buffer_6387 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T2), .Q (new_AGEMA_signal_12239) ) ;
    buf_clk new_AGEMA_reg_buffer_6390 ( .C (clk), .D (new_AGEMA_signal_5024), .Q (new_AGEMA_signal_12242) ) ;
    buf_clk new_AGEMA_reg_buffer_6393 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T6), .Q (new_AGEMA_signal_12245) ) ;
    buf_clk new_AGEMA_reg_buffer_6396 ( .C (clk), .D (new_AGEMA_signal_5213), .Q (new_AGEMA_signal_12248) ) ;
    buf_clk new_AGEMA_reg_buffer_6399 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T8), .Q (new_AGEMA_signal_12251) ) ;
    buf_clk new_AGEMA_reg_buffer_6402 ( .C (clk), .D (new_AGEMA_signal_5423), .Q (new_AGEMA_signal_12254) ) ;
    buf_clk new_AGEMA_reg_buffer_6405 ( .C (clk), .D (ciphertext_s0[48]), .Q (new_AGEMA_signal_12257) ) ;
    buf_clk new_AGEMA_reg_buffer_6408 ( .C (clk), .D (ciphertext_s1[48]), .Q (new_AGEMA_signal_12260) ) ;
    buf_clk new_AGEMA_reg_buffer_6411 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T16), .Q (new_AGEMA_signal_12263) ) ;
    buf_clk new_AGEMA_reg_buffer_6414 ( .C (clk), .D (new_AGEMA_signal_5217), .Q (new_AGEMA_signal_12266) ) ;
    buf_clk new_AGEMA_reg_buffer_6417 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T9), .Q (new_AGEMA_signal_12269) ) ;
    buf_clk new_AGEMA_reg_buffer_6420 ( .C (clk), .D (new_AGEMA_signal_5214), .Q (new_AGEMA_signal_12272) ) ;
    buf_clk new_AGEMA_reg_buffer_6423 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T17), .Q (new_AGEMA_signal_12275) ) ;
    buf_clk new_AGEMA_reg_buffer_6426 ( .C (clk), .D (new_AGEMA_signal_5426), .Q (new_AGEMA_signal_12278) ) ;
    buf_clk new_AGEMA_reg_buffer_6429 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T15), .Q (new_AGEMA_signal_12281) ) ;
    buf_clk new_AGEMA_reg_buffer_6432 ( .C (clk), .D (new_AGEMA_signal_5216), .Q (new_AGEMA_signal_12284) ) ;
    buf_clk new_AGEMA_reg_buffer_6435 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T27), .Q (new_AGEMA_signal_12287) ) ;
    buf_clk new_AGEMA_reg_buffer_6438 ( .C (clk), .D (new_AGEMA_signal_5220), .Q (new_AGEMA_signal_12290) ) ;
    buf_clk new_AGEMA_reg_buffer_6441 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T10), .Q (new_AGEMA_signal_12293) ) ;
    buf_clk new_AGEMA_reg_buffer_6444 ( .C (clk), .D (new_AGEMA_signal_5424), .Q (new_AGEMA_signal_12296) ) ;
    buf_clk new_AGEMA_reg_buffer_6447 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T13), .Q (new_AGEMA_signal_12299) ) ;
    buf_clk new_AGEMA_reg_buffer_6450 ( .C (clk), .D (new_AGEMA_signal_5215), .Q (new_AGEMA_signal_12302) ) ;
    buf_clk new_AGEMA_reg_buffer_6453 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T23), .Q (new_AGEMA_signal_12305) ) ;
    buf_clk new_AGEMA_reg_buffer_6456 ( .C (clk), .D (new_AGEMA_signal_5428), .Q (new_AGEMA_signal_12308) ) ;
    buf_clk new_AGEMA_reg_buffer_6459 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T19), .Q (new_AGEMA_signal_12311) ) ;
    buf_clk new_AGEMA_reg_buffer_6462 ( .C (clk), .D (new_AGEMA_signal_5218), .Q (new_AGEMA_signal_12314) ) ;
    buf_clk new_AGEMA_reg_buffer_6465 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T3), .Q (new_AGEMA_signal_12317) ) ;
    buf_clk new_AGEMA_reg_buffer_6468 ( .C (clk), .D (new_AGEMA_signal_5035), .Q (new_AGEMA_signal_12320) ) ;
    buf_clk new_AGEMA_reg_buffer_6471 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T22), .Q (new_AGEMA_signal_12323) ) ;
    buf_clk new_AGEMA_reg_buffer_6474 ( .C (clk), .D (new_AGEMA_signal_5219), .Q (new_AGEMA_signal_12326) ) ;
    buf_clk new_AGEMA_reg_buffer_6477 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T20), .Q (new_AGEMA_signal_12329) ) ;
    buf_clk new_AGEMA_reg_buffer_6480 ( .C (clk), .D (new_AGEMA_signal_5427), .Q (new_AGEMA_signal_12332) ) ;
    buf_clk new_AGEMA_reg_buffer_6483 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T1), .Q (new_AGEMA_signal_12335) ) ;
    buf_clk new_AGEMA_reg_buffer_6486 ( .C (clk), .D (new_AGEMA_signal_5033), .Q (new_AGEMA_signal_12338) ) ;
    buf_clk new_AGEMA_reg_buffer_6489 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T4), .Q (new_AGEMA_signal_12341) ) ;
    buf_clk new_AGEMA_reg_buffer_6492 ( .C (clk), .D (new_AGEMA_signal_5036), .Q (new_AGEMA_signal_12344) ) ;
    buf_clk new_AGEMA_reg_buffer_6495 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T2), .Q (new_AGEMA_signal_12347) ) ;
    buf_clk new_AGEMA_reg_buffer_6498 ( .C (clk), .D (new_AGEMA_signal_5034), .Q (new_AGEMA_signal_12350) ) ;
    buf_clk new_AGEMA_reg_buffer_6501 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T6), .Q (new_AGEMA_signal_12353) ) ;
    buf_clk new_AGEMA_reg_buffer_6504 ( .C (clk), .D (new_AGEMA_signal_5221), .Q (new_AGEMA_signal_12356) ) ;
    buf_clk new_AGEMA_reg_buffer_6507 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T8), .Q (new_AGEMA_signal_12359) ) ;
    buf_clk new_AGEMA_reg_buffer_6510 ( .C (clk), .D (new_AGEMA_signal_5436), .Q (new_AGEMA_signal_12362) ) ;
    buf_clk new_AGEMA_reg_buffer_6513 ( .C (clk), .D (ciphertext_s0[56]), .Q (new_AGEMA_signal_12365) ) ;
    buf_clk new_AGEMA_reg_buffer_6516 ( .C (clk), .D (ciphertext_s1[56]), .Q (new_AGEMA_signal_12368) ) ;
    buf_clk new_AGEMA_reg_buffer_6519 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T16), .Q (new_AGEMA_signal_12371) ) ;
    buf_clk new_AGEMA_reg_buffer_6522 ( .C (clk), .D (new_AGEMA_signal_5225), .Q (new_AGEMA_signal_12374) ) ;
    buf_clk new_AGEMA_reg_buffer_6525 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T9), .Q (new_AGEMA_signal_12377) ) ;
    buf_clk new_AGEMA_reg_buffer_6528 ( .C (clk), .D (new_AGEMA_signal_5222), .Q (new_AGEMA_signal_12380) ) ;
    buf_clk new_AGEMA_reg_buffer_6531 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T17), .Q (new_AGEMA_signal_12383) ) ;
    buf_clk new_AGEMA_reg_buffer_6534 ( .C (clk), .D (new_AGEMA_signal_5439), .Q (new_AGEMA_signal_12386) ) ;
    buf_clk new_AGEMA_reg_buffer_6537 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T15), .Q (new_AGEMA_signal_12389) ) ;
    buf_clk new_AGEMA_reg_buffer_6540 ( .C (clk), .D (new_AGEMA_signal_5224), .Q (new_AGEMA_signal_12392) ) ;
    buf_clk new_AGEMA_reg_buffer_6543 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T27), .Q (new_AGEMA_signal_12395) ) ;
    buf_clk new_AGEMA_reg_buffer_6546 ( .C (clk), .D (new_AGEMA_signal_5228), .Q (new_AGEMA_signal_12398) ) ;
    buf_clk new_AGEMA_reg_buffer_6549 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T10), .Q (new_AGEMA_signal_12401) ) ;
    buf_clk new_AGEMA_reg_buffer_6552 ( .C (clk), .D (new_AGEMA_signal_5437), .Q (new_AGEMA_signal_12404) ) ;
    buf_clk new_AGEMA_reg_buffer_6555 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T13), .Q (new_AGEMA_signal_12407) ) ;
    buf_clk new_AGEMA_reg_buffer_6558 ( .C (clk), .D (new_AGEMA_signal_5223), .Q (new_AGEMA_signal_12410) ) ;
    buf_clk new_AGEMA_reg_buffer_6561 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T23), .Q (new_AGEMA_signal_12413) ) ;
    buf_clk new_AGEMA_reg_buffer_6564 ( .C (clk), .D (new_AGEMA_signal_5441), .Q (new_AGEMA_signal_12416) ) ;
    buf_clk new_AGEMA_reg_buffer_6567 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T19), .Q (new_AGEMA_signal_12419) ) ;
    buf_clk new_AGEMA_reg_buffer_6570 ( .C (clk), .D (new_AGEMA_signal_5226), .Q (new_AGEMA_signal_12422) ) ;
    buf_clk new_AGEMA_reg_buffer_6573 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T3), .Q (new_AGEMA_signal_12425) ) ;
    buf_clk new_AGEMA_reg_buffer_6576 ( .C (clk), .D (new_AGEMA_signal_5045), .Q (new_AGEMA_signal_12428) ) ;
    buf_clk new_AGEMA_reg_buffer_6579 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T22), .Q (new_AGEMA_signal_12431) ) ;
    buf_clk new_AGEMA_reg_buffer_6582 ( .C (clk), .D (new_AGEMA_signal_5227), .Q (new_AGEMA_signal_12434) ) ;
    buf_clk new_AGEMA_reg_buffer_6585 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T20), .Q (new_AGEMA_signal_12437) ) ;
    buf_clk new_AGEMA_reg_buffer_6588 ( .C (clk), .D (new_AGEMA_signal_5440), .Q (new_AGEMA_signal_12440) ) ;
    buf_clk new_AGEMA_reg_buffer_6591 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T1), .Q (new_AGEMA_signal_12443) ) ;
    buf_clk new_AGEMA_reg_buffer_6594 ( .C (clk), .D (new_AGEMA_signal_5043), .Q (new_AGEMA_signal_12446) ) ;
    buf_clk new_AGEMA_reg_buffer_6597 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T4), .Q (new_AGEMA_signal_12449) ) ;
    buf_clk new_AGEMA_reg_buffer_6600 ( .C (clk), .D (new_AGEMA_signal_5046), .Q (new_AGEMA_signal_12452) ) ;
    buf_clk new_AGEMA_reg_buffer_6603 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T2), .Q (new_AGEMA_signal_12455) ) ;
    buf_clk new_AGEMA_reg_buffer_6606 ( .C (clk), .D (new_AGEMA_signal_5044), .Q (new_AGEMA_signal_12458) ) ;
    buf_clk new_AGEMA_reg_buffer_6609 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T6), .Q (new_AGEMA_signal_12461) ) ;
    buf_clk new_AGEMA_reg_buffer_6612 ( .C (clk), .D (new_AGEMA_signal_5229), .Q (new_AGEMA_signal_12464) ) ;
    buf_clk new_AGEMA_reg_buffer_6615 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T8), .Q (new_AGEMA_signal_12467) ) ;
    buf_clk new_AGEMA_reg_buffer_6618 ( .C (clk), .D (new_AGEMA_signal_5449), .Q (new_AGEMA_signal_12470) ) ;
    buf_clk new_AGEMA_reg_buffer_6621 ( .C (clk), .D (ciphertext_s0[64]), .Q (new_AGEMA_signal_12473) ) ;
    buf_clk new_AGEMA_reg_buffer_6624 ( .C (clk), .D (ciphertext_s1[64]), .Q (new_AGEMA_signal_12476) ) ;
    buf_clk new_AGEMA_reg_buffer_6627 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T16), .Q (new_AGEMA_signal_12479) ) ;
    buf_clk new_AGEMA_reg_buffer_6630 ( .C (clk), .D (new_AGEMA_signal_5233), .Q (new_AGEMA_signal_12482) ) ;
    buf_clk new_AGEMA_reg_buffer_6633 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T9), .Q (new_AGEMA_signal_12485) ) ;
    buf_clk new_AGEMA_reg_buffer_6636 ( .C (clk), .D (new_AGEMA_signal_5230), .Q (new_AGEMA_signal_12488) ) ;
    buf_clk new_AGEMA_reg_buffer_6639 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T17), .Q (new_AGEMA_signal_12491) ) ;
    buf_clk new_AGEMA_reg_buffer_6642 ( .C (clk), .D (new_AGEMA_signal_5452), .Q (new_AGEMA_signal_12494) ) ;
    buf_clk new_AGEMA_reg_buffer_6645 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T15), .Q (new_AGEMA_signal_12497) ) ;
    buf_clk new_AGEMA_reg_buffer_6648 ( .C (clk), .D (new_AGEMA_signal_5232), .Q (new_AGEMA_signal_12500) ) ;
    buf_clk new_AGEMA_reg_buffer_6651 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T27), .Q (new_AGEMA_signal_12503) ) ;
    buf_clk new_AGEMA_reg_buffer_6654 ( .C (clk), .D (new_AGEMA_signal_5236), .Q (new_AGEMA_signal_12506) ) ;
    buf_clk new_AGEMA_reg_buffer_6657 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T10), .Q (new_AGEMA_signal_12509) ) ;
    buf_clk new_AGEMA_reg_buffer_6660 ( .C (clk), .D (new_AGEMA_signal_5450), .Q (new_AGEMA_signal_12512) ) ;
    buf_clk new_AGEMA_reg_buffer_6663 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T13), .Q (new_AGEMA_signal_12515) ) ;
    buf_clk new_AGEMA_reg_buffer_6666 ( .C (clk), .D (new_AGEMA_signal_5231), .Q (new_AGEMA_signal_12518) ) ;
    buf_clk new_AGEMA_reg_buffer_6669 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T23), .Q (new_AGEMA_signal_12521) ) ;
    buf_clk new_AGEMA_reg_buffer_6672 ( .C (clk), .D (new_AGEMA_signal_5454), .Q (new_AGEMA_signal_12524) ) ;
    buf_clk new_AGEMA_reg_buffer_6675 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T19), .Q (new_AGEMA_signal_12527) ) ;
    buf_clk new_AGEMA_reg_buffer_6678 ( .C (clk), .D (new_AGEMA_signal_5234), .Q (new_AGEMA_signal_12530) ) ;
    buf_clk new_AGEMA_reg_buffer_6681 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T3), .Q (new_AGEMA_signal_12533) ) ;
    buf_clk new_AGEMA_reg_buffer_6684 ( .C (clk), .D (new_AGEMA_signal_5055), .Q (new_AGEMA_signal_12536) ) ;
    buf_clk new_AGEMA_reg_buffer_6687 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T22), .Q (new_AGEMA_signal_12539) ) ;
    buf_clk new_AGEMA_reg_buffer_6690 ( .C (clk), .D (new_AGEMA_signal_5235), .Q (new_AGEMA_signal_12542) ) ;
    buf_clk new_AGEMA_reg_buffer_6693 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T20), .Q (new_AGEMA_signal_12545) ) ;
    buf_clk new_AGEMA_reg_buffer_6696 ( .C (clk), .D (new_AGEMA_signal_5453), .Q (new_AGEMA_signal_12548) ) ;
    buf_clk new_AGEMA_reg_buffer_6699 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T1), .Q (new_AGEMA_signal_12551) ) ;
    buf_clk new_AGEMA_reg_buffer_6702 ( .C (clk), .D (new_AGEMA_signal_5053), .Q (new_AGEMA_signal_12554) ) ;
    buf_clk new_AGEMA_reg_buffer_6705 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T4), .Q (new_AGEMA_signal_12557) ) ;
    buf_clk new_AGEMA_reg_buffer_6708 ( .C (clk), .D (new_AGEMA_signal_5056), .Q (new_AGEMA_signal_12560) ) ;
    buf_clk new_AGEMA_reg_buffer_6711 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T2), .Q (new_AGEMA_signal_12563) ) ;
    buf_clk new_AGEMA_reg_buffer_6714 ( .C (clk), .D (new_AGEMA_signal_5054), .Q (new_AGEMA_signal_12566) ) ;
    buf_clk new_AGEMA_reg_buffer_6717 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T6), .Q (new_AGEMA_signal_12569) ) ;
    buf_clk new_AGEMA_reg_buffer_6720 ( .C (clk), .D (new_AGEMA_signal_5237), .Q (new_AGEMA_signal_12572) ) ;
    buf_clk new_AGEMA_reg_buffer_6723 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T8), .Q (new_AGEMA_signal_12575) ) ;
    buf_clk new_AGEMA_reg_buffer_6726 ( .C (clk), .D (new_AGEMA_signal_5462), .Q (new_AGEMA_signal_12578) ) ;
    buf_clk new_AGEMA_reg_buffer_6729 ( .C (clk), .D (ciphertext_s0[72]), .Q (new_AGEMA_signal_12581) ) ;
    buf_clk new_AGEMA_reg_buffer_6732 ( .C (clk), .D (ciphertext_s1[72]), .Q (new_AGEMA_signal_12584) ) ;
    buf_clk new_AGEMA_reg_buffer_6735 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T16), .Q (new_AGEMA_signal_12587) ) ;
    buf_clk new_AGEMA_reg_buffer_6738 ( .C (clk), .D (new_AGEMA_signal_5241), .Q (new_AGEMA_signal_12590) ) ;
    buf_clk new_AGEMA_reg_buffer_6741 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T9), .Q (new_AGEMA_signal_12593) ) ;
    buf_clk new_AGEMA_reg_buffer_6744 ( .C (clk), .D (new_AGEMA_signal_5238), .Q (new_AGEMA_signal_12596) ) ;
    buf_clk new_AGEMA_reg_buffer_6747 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T17), .Q (new_AGEMA_signal_12599) ) ;
    buf_clk new_AGEMA_reg_buffer_6750 ( .C (clk), .D (new_AGEMA_signal_5465), .Q (new_AGEMA_signal_12602) ) ;
    buf_clk new_AGEMA_reg_buffer_6753 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T15), .Q (new_AGEMA_signal_12605) ) ;
    buf_clk new_AGEMA_reg_buffer_6756 ( .C (clk), .D (new_AGEMA_signal_5240), .Q (new_AGEMA_signal_12608) ) ;
    buf_clk new_AGEMA_reg_buffer_6759 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T27), .Q (new_AGEMA_signal_12611) ) ;
    buf_clk new_AGEMA_reg_buffer_6762 ( .C (clk), .D (new_AGEMA_signal_5244), .Q (new_AGEMA_signal_12614) ) ;
    buf_clk new_AGEMA_reg_buffer_6765 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T10), .Q (new_AGEMA_signal_12617) ) ;
    buf_clk new_AGEMA_reg_buffer_6768 ( .C (clk), .D (new_AGEMA_signal_5463), .Q (new_AGEMA_signal_12620) ) ;
    buf_clk new_AGEMA_reg_buffer_6771 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T13), .Q (new_AGEMA_signal_12623) ) ;
    buf_clk new_AGEMA_reg_buffer_6774 ( .C (clk), .D (new_AGEMA_signal_5239), .Q (new_AGEMA_signal_12626) ) ;
    buf_clk new_AGEMA_reg_buffer_6777 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T23), .Q (new_AGEMA_signal_12629) ) ;
    buf_clk new_AGEMA_reg_buffer_6780 ( .C (clk), .D (new_AGEMA_signal_5467), .Q (new_AGEMA_signal_12632) ) ;
    buf_clk new_AGEMA_reg_buffer_6783 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T19), .Q (new_AGEMA_signal_12635) ) ;
    buf_clk new_AGEMA_reg_buffer_6786 ( .C (clk), .D (new_AGEMA_signal_5242), .Q (new_AGEMA_signal_12638) ) ;
    buf_clk new_AGEMA_reg_buffer_6789 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T3), .Q (new_AGEMA_signal_12641) ) ;
    buf_clk new_AGEMA_reg_buffer_6792 ( .C (clk), .D (new_AGEMA_signal_5065), .Q (new_AGEMA_signal_12644) ) ;
    buf_clk new_AGEMA_reg_buffer_6795 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T22), .Q (new_AGEMA_signal_12647) ) ;
    buf_clk new_AGEMA_reg_buffer_6798 ( .C (clk), .D (new_AGEMA_signal_5243), .Q (new_AGEMA_signal_12650) ) ;
    buf_clk new_AGEMA_reg_buffer_6801 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T20), .Q (new_AGEMA_signal_12653) ) ;
    buf_clk new_AGEMA_reg_buffer_6804 ( .C (clk), .D (new_AGEMA_signal_5466), .Q (new_AGEMA_signal_12656) ) ;
    buf_clk new_AGEMA_reg_buffer_6807 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T1), .Q (new_AGEMA_signal_12659) ) ;
    buf_clk new_AGEMA_reg_buffer_6810 ( .C (clk), .D (new_AGEMA_signal_5063), .Q (new_AGEMA_signal_12662) ) ;
    buf_clk new_AGEMA_reg_buffer_6813 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T4), .Q (new_AGEMA_signal_12665) ) ;
    buf_clk new_AGEMA_reg_buffer_6816 ( .C (clk), .D (new_AGEMA_signal_5066), .Q (new_AGEMA_signal_12668) ) ;
    buf_clk new_AGEMA_reg_buffer_6819 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T2), .Q (new_AGEMA_signal_12671) ) ;
    buf_clk new_AGEMA_reg_buffer_6822 ( .C (clk), .D (new_AGEMA_signal_5064), .Q (new_AGEMA_signal_12674) ) ;
    buf_clk new_AGEMA_reg_buffer_6825 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T6), .Q (new_AGEMA_signal_12677) ) ;
    buf_clk new_AGEMA_reg_buffer_6828 ( .C (clk), .D (new_AGEMA_signal_5245), .Q (new_AGEMA_signal_12680) ) ;
    buf_clk new_AGEMA_reg_buffer_6831 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T8), .Q (new_AGEMA_signal_12683) ) ;
    buf_clk new_AGEMA_reg_buffer_6834 ( .C (clk), .D (new_AGEMA_signal_5475), .Q (new_AGEMA_signal_12686) ) ;
    buf_clk new_AGEMA_reg_buffer_6837 ( .C (clk), .D (ciphertext_s0[80]), .Q (new_AGEMA_signal_12689) ) ;
    buf_clk new_AGEMA_reg_buffer_6840 ( .C (clk), .D (ciphertext_s1[80]), .Q (new_AGEMA_signal_12692) ) ;
    buf_clk new_AGEMA_reg_buffer_6843 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T16), .Q (new_AGEMA_signal_12695) ) ;
    buf_clk new_AGEMA_reg_buffer_6846 ( .C (clk), .D (new_AGEMA_signal_5249), .Q (new_AGEMA_signal_12698) ) ;
    buf_clk new_AGEMA_reg_buffer_6849 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T9), .Q (new_AGEMA_signal_12701) ) ;
    buf_clk new_AGEMA_reg_buffer_6852 ( .C (clk), .D (new_AGEMA_signal_5246), .Q (new_AGEMA_signal_12704) ) ;
    buf_clk new_AGEMA_reg_buffer_6855 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T17), .Q (new_AGEMA_signal_12707) ) ;
    buf_clk new_AGEMA_reg_buffer_6858 ( .C (clk), .D (new_AGEMA_signal_5478), .Q (new_AGEMA_signal_12710) ) ;
    buf_clk new_AGEMA_reg_buffer_6861 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T15), .Q (new_AGEMA_signal_12713) ) ;
    buf_clk new_AGEMA_reg_buffer_6864 ( .C (clk), .D (new_AGEMA_signal_5248), .Q (new_AGEMA_signal_12716) ) ;
    buf_clk new_AGEMA_reg_buffer_6867 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T27), .Q (new_AGEMA_signal_12719) ) ;
    buf_clk new_AGEMA_reg_buffer_6870 ( .C (clk), .D (new_AGEMA_signal_5252), .Q (new_AGEMA_signal_12722) ) ;
    buf_clk new_AGEMA_reg_buffer_6873 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T10), .Q (new_AGEMA_signal_12725) ) ;
    buf_clk new_AGEMA_reg_buffer_6876 ( .C (clk), .D (new_AGEMA_signal_5476), .Q (new_AGEMA_signal_12728) ) ;
    buf_clk new_AGEMA_reg_buffer_6879 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T13), .Q (new_AGEMA_signal_12731) ) ;
    buf_clk new_AGEMA_reg_buffer_6882 ( .C (clk), .D (new_AGEMA_signal_5247), .Q (new_AGEMA_signal_12734) ) ;
    buf_clk new_AGEMA_reg_buffer_6885 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T23), .Q (new_AGEMA_signal_12737) ) ;
    buf_clk new_AGEMA_reg_buffer_6888 ( .C (clk), .D (new_AGEMA_signal_5480), .Q (new_AGEMA_signal_12740) ) ;
    buf_clk new_AGEMA_reg_buffer_6891 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T19), .Q (new_AGEMA_signal_12743) ) ;
    buf_clk new_AGEMA_reg_buffer_6894 ( .C (clk), .D (new_AGEMA_signal_5250), .Q (new_AGEMA_signal_12746) ) ;
    buf_clk new_AGEMA_reg_buffer_6897 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T3), .Q (new_AGEMA_signal_12749) ) ;
    buf_clk new_AGEMA_reg_buffer_6900 ( .C (clk), .D (new_AGEMA_signal_5075), .Q (new_AGEMA_signal_12752) ) ;
    buf_clk new_AGEMA_reg_buffer_6903 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T22), .Q (new_AGEMA_signal_12755) ) ;
    buf_clk new_AGEMA_reg_buffer_6906 ( .C (clk), .D (new_AGEMA_signal_5251), .Q (new_AGEMA_signal_12758) ) ;
    buf_clk new_AGEMA_reg_buffer_6909 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T20), .Q (new_AGEMA_signal_12761) ) ;
    buf_clk new_AGEMA_reg_buffer_6912 ( .C (clk), .D (new_AGEMA_signal_5479), .Q (new_AGEMA_signal_12764) ) ;
    buf_clk new_AGEMA_reg_buffer_6915 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T1), .Q (new_AGEMA_signal_12767) ) ;
    buf_clk new_AGEMA_reg_buffer_6918 ( .C (clk), .D (new_AGEMA_signal_5073), .Q (new_AGEMA_signal_12770) ) ;
    buf_clk new_AGEMA_reg_buffer_6921 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T4), .Q (new_AGEMA_signal_12773) ) ;
    buf_clk new_AGEMA_reg_buffer_6924 ( .C (clk), .D (new_AGEMA_signal_5076), .Q (new_AGEMA_signal_12776) ) ;
    buf_clk new_AGEMA_reg_buffer_6927 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T2), .Q (new_AGEMA_signal_12779) ) ;
    buf_clk new_AGEMA_reg_buffer_6930 ( .C (clk), .D (new_AGEMA_signal_5074), .Q (new_AGEMA_signal_12782) ) ;
    buf_clk new_AGEMA_reg_buffer_6933 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T6), .Q (new_AGEMA_signal_12785) ) ;
    buf_clk new_AGEMA_reg_buffer_6936 ( .C (clk), .D (new_AGEMA_signal_5253), .Q (new_AGEMA_signal_12788) ) ;
    buf_clk new_AGEMA_reg_buffer_6939 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T8), .Q (new_AGEMA_signal_12791) ) ;
    buf_clk new_AGEMA_reg_buffer_6942 ( .C (clk), .D (new_AGEMA_signal_5488), .Q (new_AGEMA_signal_12794) ) ;
    buf_clk new_AGEMA_reg_buffer_6945 ( .C (clk), .D (ciphertext_s0[88]), .Q (new_AGEMA_signal_12797) ) ;
    buf_clk new_AGEMA_reg_buffer_6948 ( .C (clk), .D (ciphertext_s1[88]), .Q (new_AGEMA_signal_12800) ) ;
    buf_clk new_AGEMA_reg_buffer_6951 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T16), .Q (new_AGEMA_signal_12803) ) ;
    buf_clk new_AGEMA_reg_buffer_6954 ( .C (clk), .D (new_AGEMA_signal_5257), .Q (new_AGEMA_signal_12806) ) ;
    buf_clk new_AGEMA_reg_buffer_6957 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T9), .Q (new_AGEMA_signal_12809) ) ;
    buf_clk new_AGEMA_reg_buffer_6960 ( .C (clk), .D (new_AGEMA_signal_5254), .Q (new_AGEMA_signal_12812) ) ;
    buf_clk new_AGEMA_reg_buffer_6963 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T17), .Q (new_AGEMA_signal_12815) ) ;
    buf_clk new_AGEMA_reg_buffer_6966 ( .C (clk), .D (new_AGEMA_signal_5491), .Q (new_AGEMA_signal_12818) ) ;
    buf_clk new_AGEMA_reg_buffer_6969 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T15), .Q (new_AGEMA_signal_12821) ) ;
    buf_clk new_AGEMA_reg_buffer_6972 ( .C (clk), .D (new_AGEMA_signal_5256), .Q (new_AGEMA_signal_12824) ) ;
    buf_clk new_AGEMA_reg_buffer_6975 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T27), .Q (new_AGEMA_signal_12827) ) ;
    buf_clk new_AGEMA_reg_buffer_6978 ( .C (clk), .D (new_AGEMA_signal_5260), .Q (new_AGEMA_signal_12830) ) ;
    buf_clk new_AGEMA_reg_buffer_6981 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T10), .Q (new_AGEMA_signal_12833) ) ;
    buf_clk new_AGEMA_reg_buffer_6984 ( .C (clk), .D (new_AGEMA_signal_5489), .Q (new_AGEMA_signal_12836) ) ;
    buf_clk new_AGEMA_reg_buffer_6987 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T13), .Q (new_AGEMA_signal_12839) ) ;
    buf_clk new_AGEMA_reg_buffer_6990 ( .C (clk), .D (new_AGEMA_signal_5255), .Q (new_AGEMA_signal_12842) ) ;
    buf_clk new_AGEMA_reg_buffer_6993 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T23), .Q (new_AGEMA_signal_12845) ) ;
    buf_clk new_AGEMA_reg_buffer_6996 ( .C (clk), .D (new_AGEMA_signal_5493), .Q (new_AGEMA_signal_12848) ) ;
    buf_clk new_AGEMA_reg_buffer_6999 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T19), .Q (new_AGEMA_signal_12851) ) ;
    buf_clk new_AGEMA_reg_buffer_7002 ( .C (clk), .D (new_AGEMA_signal_5258), .Q (new_AGEMA_signal_12854) ) ;
    buf_clk new_AGEMA_reg_buffer_7005 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T3), .Q (new_AGEMA_signal_12857) ) ;
    buf_clk new_AGEMA_reg_buffer_7008 ( .C (clk), .D (new_AGEMA_signal_5085), .Q (new_AGEMA_signal_12860) ) ;
    buf_clk new_AGEMA_reg_buffer_7011 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T22), .Q (new_AGEMA_signal_12863) ) ;
    buf_clk new_AGEMA_reg_buffer_7014 ( .C (clk), .D (new_AGEMA_signal_5259), .Q (new_AGEMA_signal_12866) ) ;
    buf_clk new_AGEMA_reg_buffer_7017 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T20), .Q (new_AGEMA_signal_12869) ) ;
    buf_clk new_AGEMA_reg_buffer_7020 ( .C (clk), .D (new_AGEMA_signal_5492), .Q (new_AGEMA_signal_12872) ) ;
    buf_clk new_AGEMA_reg_buffer_7023 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T1), .Q (new_AGEMA_signal_12875) ) ;
    buf_clk new_AGEMA_reg_buffer_7026 ( .C (clk), .D (new_AGEMA_signal_5083), .Q (new_AGEMA_signal_12878) ) ;
    buf_clk new_AGEMA_reg_buffer_7029 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T4), .Q (new_AGEMA_signal_12881) ) ;
    buf_clk new_AGEMA_reg_buffer_7032 ( .C (clk), .D (new_AGEMA_signal_5086), .Q (new_AGEMA_signal_12884) ) ;
    buf_clk new_AGEMA_reg_buffer_7035 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T2), .Q (new_AGEMA_signal_12887) ) ;
    buf_clk new_AGEMA_reg_buffer_7038 ( .C (clk), .D (new_AGEMA_signal_5084), .Q (new_AGEMA_signal_12890) ) ;
    buf_clk new_AGEMA_reg_buffer_7041 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T6), .Q (new_AGEMA_signal_12893) ) ;
    buf_clk new_AGEMA_reg_buffer_7044 ( .C (clk), .D (new_AGEMA_signal_5261), .Q (new_AGEMA_signal_12896) ) ;
    buf_clk new_AGEMA_reg_buffer_7047 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T8), .Q (new_AGEMA_signal_12899) ) ;
    buf_clk new_AGEMA_reg_buffer_7050 ( .C (clk), .D (new_AGEMA_signal_5501), .Q (new_AGEMA_signal_12902) ) ;
    buf_clk new_AGEMA_reg_buffer_7053 ( .C (clk), .D (ciphertext_s0[96]), .Q (new_AGEMA_signal_12905) ) ;
    buf_clk new_AGEMA_reg_buffer_7056 ( .C (clk), .D (ciphertext_s1[96]), .Q (new_AGEMA_signal_12908) ) ;
    buf_clk new_AGEMA_reg_buffer_7059 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T16), .Q (new_AGEMA_signal_12911) ) ;
    buf_clk new_AGEMA_reg_buffer_7062 ( .C (clk), .D (new_AGEMA_signal_5265), .Q (new_AGEMA_signal_12914) ) ;
    buf_clk new_AGEMA_reg_buffer_7065 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T9), .Q (new_AGEMA_signal_12917) ) ;
    buf_clk new_AGEMA_reg_buffer_7068 ( .C (clk), .D (new_AGEMA_signal_5262), .Q (new_AGEMA_signal_12920) ) ;
    buf_clk new_AGEMA_reg_buffer_7071 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T17), .Q (new_AGEMA_signal_12923) ) ;
    buf_clk new_AGEMA_reg_buffer_7074 ( .C (clk), .D (new_AGEMA_signal_5504), .Q (new_AGEMA_signal_12926) ) ;
    buf_clk new_AGEMA_reg_buffer_7077 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T15), .Q (new_AGEMA_signal_12929) ) ;
    buf_clk new_AGEMA_reg_buffer_7080 ( .C (clk), .D (new_AGEMA_signal_5264), .Q (new_AGEMA_signal_12932) ) ;
    buf_clk new_AGEMA_reg_buffer_7083 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T27), .Q (new_AGEMA_signal_12935) ) ;
    buf_clk new_AGEMA_reg_buffer_7086 ( .C (clk), .D (new_AGEMA_signal_5268), .Q (new_AGEMA_signal_12938) ) ;
    buf_clk new_AGEMA_reg_buffer_7089 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T10), .Q (new_AGEMA_signal_12941) ) ;
    buf_clk new_AGEMA_reg_buffer_7092 ( .C (clk), .D (new_AGEMA_signal_5502), .Q (new_AGEMA_signal_12944) ) ;
    buf_clk new_AGEMA_reg_buffer_7095 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T13), .Q (new_AGEMA_signal_12947) ) ;
    buf_clk new_AGEMA_reg_buffer_7098 ( .C (clk), .D (new_AGEMA_signal_5263), .Q (new_AGEMA_signal_12950) ) ;
    buf_clk new_AGEMA_reg_buffer_7101 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T23), .Q (new_AGEMA_signal_12953) ) ;
    buf_clk new_AGEMA_reg_buffer_7104 ( .C (clk), .D (new_AGEMA_signal_5506), .Q (new_AGEMA_signal_12956) ) ;
    buf_clk new_AGEMA_reg_buffer_7107 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T19), .Q (new_AGEMA_signal_12959) ) ;
    buf_clk new_AGEMA_reg_buffer_7110 ( .C (clk), .D (new_AGEMA_signal_5266), .Q (new_AGEMA_signal_12962) ) ;
    buf_clk new_AGEMA_reg_buffer_7113 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T3), .Q (new_AGEMA_signal_12965) ) ;
    buf_clk new_AGEMA_reg_buffer_7116 ( .C (clk), .D (new_AGEMA_signal_5095), .Q (new_AGEMA_signal_12968) ) ;
    buf_clk new_AGEMA_reg_buffer_7119 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T22), .Q (new_AGEMA_signal_12971) ) ;
    buf_clk new_AGEMA_reg_buffer_7122 ( .C (clk), .D (new_AGEMA_signal_5267), .Q (new_AGEMA_signal_12974) ) ;
    buf_clk new_AGEMA_reg_buffer_7125 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T20), .Q (new_AGEMA_signal_12977) ) ;
    buf_clk new_AGEMA_reg_buffer_7128 ( .C (clk), .D (new_AGEMA_signal_5505), .Q (new_AGEMA_signal_12980) ) ;
    buf_clk new_AGEMA_reg_buffer_7131 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T1), .Q (new_AGEMA_signal_12983) ) ;
    buf_clk new_AGEMA_reg_buffer_7134 ( .C (clk), .D (new_AGEMA_signal_5093), .Q (new_AGEMA_signal_12986) ) ;
    buf_clk new_AGEMA_reg_buffer_7137 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T4), .Q (new_AGEMA_signal_12989) ) ;
    buf_clk new_AGEMA_reg_buffer_7140 ( .C (clk), .D (new_AGEMA_signal_5096), .Q (new_AGEMA_signal_12992) ) ;
    buf_clk new_AGEMA_reg_buffer_7143 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T2), .Q (new_AGEMA_signal_12995) ) ;
    buf_clk new_AGEMA_reg_buffer_7146 ( .C (clk), .D (new_AGEMA_signal_5094), .Q (new_AGEMA_signal_12998) ) ;
    buf_clk new_AGEMA_reg_buffer_7149 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T6), .Q (new_AGEMA_signal_13001) ) ;
    buf_clk new_AGEMA_reg_buffer_7152 ( .C (clk), .D (new_AGEMA_signal_5269), .Q (new_AGEMA_signal_13004) ) ;
    buf_clk new_AGEMA_reg_buffer_7155 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T8), .Q (new_AGEMA_signal_13007) ) ;
    buf_clk new_AGEMA_reg_buffer_7158 ( .C (clk), .D (new_AGEMA_signal_5514), .Q (new_AGEMA_signal_13010) ) ;
    buf_clk new_AGEMA_reg_buffer_7161 ( .C (clk), .D (ciphertext_s0[104]), .Q (new_AGEMA_signal_13013) ) ;
    buf_clk new_AGEMA_reg_buffer_7164 ( .C (clk), .D (ciphertext_s1[104]), .Q (new_AGEMA_signal_13016) ) ;
    buf_clk new_AGEMA_reg_buffer_7167 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T16), .Q (new_AGEMA_signal_13019) ) ;
    buf_clk new_AGEMA_reg_buffer_7170 ( .C (clk), .D (new_AGEMA_signal_5273), .Q (new_AGEMA_signal_13022) ) ;
    buf_clk new_AGEMA_reg_buffer_7173 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T9), .Q (new_AGEMA_signal_13025) ) ;
    buf_clk new_AGEMA_reg_buffer_7176 ( .C (clk), .D (new_AGEMA_signal_5270), .Q (new_AGEMA_signal_13028) ) ;
    buf_clk new_AGEMA_reg_buffer_7179 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T17), .Q (new_AGEMA_signal_13031) ) ;
    buf_clk new_AGEMA_reg_buffer_7182 ( .C (clk), .D (new_AGEMA_signal_5517), .Q (new_AGEMA_signal_13034) ) ;
    buf_clk new_AGEMA_reg_buffer_7185 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T15), .Q (new_AGEMA_signal_13037) ) ;
    buf_clk new_AGEMA_reg_buffer_7188 ( .C (clk), .D (new_AGEMA_signal_5272), .Q (new_AGEMA_signal_13040) ) ;
    buf_clk new_AGEMA_reg_buffer_7191 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T27), .Q (new_AGEMA_signal_13043) ) ;
    buf_clk new_AGEMA_reg_buffer_7194 ( .C (clk), .D (new_AGEMA_signal_5276), .Q (new_AGEMA_signal_13046) ) ;
    buf_clk new_AGEMA_reg_buffer_7197 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T10), .Q (new_AGEMA_signal_13049) ) ;
    buf_clk new_AGEMA_reg_buffer_7200 ( .C (clk), .D (new_AGEMA_signal_5515), .Q (new_AGEMA_signal_13052) ) ;
    buf_clk new_AGEMA_reg_buffer_7203 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T13), .Q (new_AGEMA_signal_13055) ) ;
    buf_clk new_AGEMA_reg_buffer_7206 ( .C (clk), .D (new_AGEMA_signal_5271), .Q (new_AGEMA_signal_13058) ) ;
    buf_clk new_AGEMA_reg_buffer_7209 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T23), .Q (new_AGEMA_signal_13061) ) ;
    buf_clk new_AGEMA_reg_buffer_7212 ( .C (clk), .D (new_AGEMA_signal_5519), .Q (new_AGEMA_signal_13064) ) ;
    buf_clk new_AGEMA_reg_buffer_7215 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T19), .Q (new_AGEMA_signal_13067) ) ;
    buf_clk new_AGEMA_reg_buffer_7218 ( .C (clk), .D (new_AGEMA_signal_5274), .Q (new_AGEMA_signal_13070) ) ;
    buf_clk new_AGEMA_reg_buffer_7221 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T3), .Q (new_AGEMA_signal_13073) ) ;
    buf_clk new_AGEMA_reg_buffer_7224 ( .C (clk), .D (new_AGEMA_signal_5105), .Q (new_AGEMA_signal_13076) ) ;
    buf_clk new_AGEMA_reg_buffer_7227 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T22), .Q (new_AGEMA_signal_13079) ) ;
    buf_clk new_AGEMA_reg_buffer_7230 ( .C (clk), .D (new_AGEMA_signal_5275), .Q (new_AGEMA_signal_13082) ) ;
    buf_clk new_AGEMA_reg_buffer_7233 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T20), .Q (new_AGEMA_signal_13085) ) ;
    buf_clk new_AGEMA_reg_buffer_7236 ( .C (clk), .D (new_AGEMA_signal_5518), .Q (new_AGEMA_signal_13088) ) ;
    buf_clk new_AGEMA_reg_buffer_7239 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T1), .Q (new_AGEMA_signal_13091) ) ;
    buf_clk new_AGEMA_reg_buffer_7242 ( .C (clk), .D (new_AGEMA_signal_5103), .Q (new_AGEMA_signal_13094) ) ;
    buf_clk new_AGEMA_reg_buffer_7245 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T4), .Q (new_AGEMA_signal_13097) ) ;
    buf_clk new_AGEMA_reg_buffer_7248 ( .C (clk), .D (new_AGEMA_signal_5106), .Q (new_AGEMA_signal_13100) ) ;
    buf_clk new_AGEMA_reg_buffer_7251 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T2), .Q (new_AGEMA_signal_13103) ) ;
    buf_clk new_AGEMA_reg_buffer_7254 ( .C (clk), .D (new_AGEMA_signal_5104), .Q (new_AGEMA_signal_13106) ) ;
    buf_clk new_AGEMA_reg_buffer_7257 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T6), .Q (new_AGEMA_signal_13109) ) ;
    buf_clk new_AGEMA_reg_buffer_7260 ( .C (clk), .D (new_AGEMA_signal_5277), .Q (new_AGEMA_signal_13112) ) ;
    buf_clk new_AGEMA_reg_buffer_7263 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T8), .Q (new_AGEMA_signal_13115) ) ;
    buf_clk new_AGEMA_reg_buffer_7266 ( .C (clk), .D (new_AGEMA_signal_5527), .Q (new_AGEMA_signal_13118) ) ;
    buf_clk new_AGEMA_reg_buffer_7269 ( .C (clk), .D (ciphertext_s0[112]), .Q (new_AGEMA_signal_13121) ) ;
    buf_clk new_AGEMA_reg_buffer_7272 ( .C (clk), .D (ciphertext_s1[112]), .Q (new_AGEMA_signal_13124) ) ;
    buf_clk new_AGEMA_reg_buffer_7275 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T16), .Q (new_AGEMA_signal_13127) ) ;
    buf_clk new_AGEMA_reg_buffer_7278 ( .C (clk), .D (new_AGEMA_signal_5281), .Q (new_AGEMA_signal_13130) ) ;
    buf_clk new_AGEMA_reg_buffer_7281 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T9), .Q (new_AGEMA_signal_13133) ) ;
    buf_clk new_AGEMA_reg_buffer_7284 ( .C (clk), .D (new_AGEMA_signal_5278), .Q (new_AGEMA_signal_13136) ) ;
    buf_clk new_AGEMA_reg_buffer_7287 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T17), .Q (new_AGEMA_signal_13139) ) ;
    buf_clk new_AGEMA_reg_buffer_7290 ( .C (clk), .D (new_AGEMA_signal_5530), .Q (new_AGEMA_signal_13142) ) ;
    buf_clk new_AGEMA_reg_buffer_7293 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T15), .Q (new_AGEMA_signal_13145) ) ;
    buf_clk new_AGEMA_reg_buffer_7296 ( .C (clk), .D (new_AGEMA_signal_5280), .Q (new_AGEMA_signal_13148) ) ;
    buf_clk new_AGEMA_reg_buffer_7299 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T27), .Q (new_AGEMA_signal_13151) ) ;
    buf_clk new_AGEMA_reg_buffer_7302 ( .C (clk), .D (new_AGEMA_signal_5284), .Q (new_AGEMA_signal_13154) ) ;
    buf_clk new_AGEMA_reg_buffer_7305 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T10), .Q (new_AGEMA_signal_13157) ) ;
    buf_clk new_AGEMA_reg_buffer_7308 ( .C (clk), .D (new_AGEMA_signal_5528), .Q (new_AGEMA_signal_13160) ) ;
    buf_clk new_AGEMA_reg_buffer_7311 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T13), .Q (new_AGEMA_signal_13163) ) ;
    buf_clk new_AGEMA_reg_buffer_7314 ( .C (clk), .D (new_AGEMA_signal_5279), .Q (new_AGEMA_signal_13166) ) ;
    buf_clk new_AGEMA_reg_buffer_7317 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T23), .Q (new_AGEMA_signal_13169) ) ;
    buf_clk new_AGEMA_reg_buffer_7320 ( .C (clk), .D (new_AGEMA_signal_5532), .Q (new_AGEMA_signal_13172) ) ;
    buf_clk new_AGEMA_reg_buffer_7323 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T19), .Q (new_AGEMA_signal_13175) ) ;
    buf_clk new_AGEMA_reg_buffer_7326 ( .C (clk), .D (new_AGEMA_signal_5282), .Q (new_AGEMA_signal_13178) ) ;
    buf_clk new_AGEMA_reg_buffer_7329 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T3), .Q (new_AGEMA_signal_13181) ) ;
    buf_clk new_AGEMA_reg_buffer_7332 ( .C (clk), .D (new_AGEMA_signal_5115), .Q (new_AGEMA_signal_13184) ) ;
    buf_clk new_AGEMA_reg_buffer_7335 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T22), .Q (new_AGEMA_signal_13187) ) ;
    buf_clk new_AGEMA_reg_buffer_7338 ( .C (clk), .D (new_AGEMA_signal_5283), .Q (new_AGEMA_signal_13190) ) ;
    buf_clk new_AGEMA_reg_buffer_7341 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T20), .Q (new_AGEMA_signal_13193) ) ;
    buf_clk new_AGEMA_reg_buffer_7344 ( .C (clk), .D (new_AGEMA_signal_5531), .Q (new_AGEMA_signal_13196) ) ;
    buf_clk new_AGEMA_reg_buffer_7347 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T1), .Q (new_AGEMA_signal_13199) ) ;
    buf_clk new_AGEMA_reg_buffer_7350 ( .C (clk), .D (new_AGEMA_signal_5113), .Q (new_AGEMA_signal_13202) ) ;
    buf_clk new_AGEMA_reg_buffer_7353 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T4), .Q (new_AGEMA_signal_13205) ) ;
    buf_clk new_AGEMA_reg_buffer_7356 ( .C (clk), .D (new_AGEMA_signal_5116), .Q (new_AGEMA_signal_13208) ) ;
    buf_clk new_AGEMA_reg_buffer_7359 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T2), .Q (new_AGEMA_signal_13211) ) ;
    buf_clk new_AGEMA_reg_buffer_7362 ( .C (clk), .D (new_AGEMA_signal_5114), .Q (new_AGEMA_signal_13214) ) ;
    buf_clk new_AGEMA_reg_buffer_7365 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T6), .Q (new_AGEMA_signal_13217) ) ;
    buf_clk new_AGEMA_reg_buffer_7368 ( .C (clk), .D (new_AGEMA_signal_5285), .Q (new_AGEMA_signal_13220) ) ;
    buf_clk new_AGEMA_reg_buffer_7371 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T8), .Q (new_AGEMA_signal_13223) ) ;
    buf_clk new_AGEMA_reg_buffer_7374 ( .C (clk), .D (new_AGEMA_signal_5540), .Q (new_AGEMA_signal_13226) ) ;
    buf_clk new_AGEMA_reg_buffer_7377 ( .C (clk), .D (ciphertext_s0[120]), .Q (new_AGEMA_signal_13229) ) ;
    buf_clk new_AGEMA_reg_buffer_7380 ( .C (clk), .D (ciphertext_s1[120]), .Q (new_AGEMA_signal_13232) ) ;
    buf_clk new_AGEMA_reg_buffer_7383 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T16), .Q (new_AGEMA_signal_13235) ) ;
    buf_clk new_AGEMA_reg_buffer_7386 ( .C (clk), .D (new_AGEMA_signal_5289), .Q (new_AGEMA_signal_13238) ) ;
    buf_clk new_AGEMA_reg_buffer_7389 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T9), .Q (new_AGEMA_signal_13241) ) ;
    buf_clk new_AGEMA_reg_buffer_7392 ( .C (clk), .D (new_AGEMA_signal_5286), .Q (new_AGEMA_signal_13244) ) ;
    buf_clk new_AGEMA_reg_buffer_7395 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T17), .Q (new_AGEMA_signal_13247) ) ;
    buf_clk new_AGEMA_reg_buffer_7398 ( .C (clk), .D (new_AGEMA_signal_5543), .Q (new_AGEMA_signal_13250) ) ;
    buf_clk new_AGEMA_reg_buffer_7401 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T15), .Q (new_AGEMA_signal_13253) ) ;
    buf_clk new_AGEMA_reg_buffer_7404 ( .C (clk), .D (new_AGEMA_signal_5288), .Q (new_AGEMA_signal_13256) ) ;
    buf_clk new_AGEMA_reg_buffer_7407 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T27), .Q (new_AGEMA_signal_13259) ) ;
    buf_clk new_AGEMA_reg_buffer_7410 ( .C (clk), .D (new_AGEMA_signal_5292), .Q (new_AGEMA_signal_13262) ) ;
    buf_clk new_AGEMA_reg_buffer_7413 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T10), .Q (new_AGEMA_signal_13265) ) ;
    buf_clk new_AGEMA_reg_buffer_7416 ( .C (clk), .D (new_AGEMA_signal_5541), .Q (new_AGEMA_signal_13268) ) ;
    buf_clk new_AGEMA_reg_buffer_7419 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T13), .Q (new_AGEMA_signal_13271) ) ;
    buf_clk new_AGEMA_reg_buffer_7422 ( .C (clk), .D (new_AGEMA_signal_5287), .Q (new_AGEMA_signal_13274) ) ;
    buf_clk new_AGEMA_reg_buffer_7425 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T23), .Q (new_AGEMA_signal_13277) ) ;
    buf_clk new_AGEMA_reg_buffer_7428 ( .C (clk), .D (new_AGEMA_signal_5545), .Q (new_AGEMA_signal_13280) ) ;
    buf_clk new_AGEMA_reg_buffer_7431 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T19), .Q (new_AGEMA_signal_13283) ) ;
    buf_clk new_AGEMA_reg_buffer_7434 ( .C (clk), .D (new_AGEMA_signal_5290), .Q (new_AGEMA_signal_13286) ) ;
    buf_clk new_AGEMA_reg_buffer_7437 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T3), .Q (new_AGEMA_signal_13289) ) ;
    buf_clk new_AGEMA_reg_buffer_7440 ( .C (clk), .D (new_AGEMA_signal_5125), .Q (new_AGEMA_signal_13292) ) ;
    buf_clk new_AGEMA_reg_buffer_7443 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T22), .Q (new_AGEMA_signal_13295) ) ;
    buf_clk new_AGEMA_reg_buffer_7446 ( .C (clk), .D (new_AGEMA_signal_5291), .Q (new_AGEMA_signal_13298) ) ;
    buf_clk new_AGEMA_reg_buffer_7449 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T20), .Q (new_AGEMA_signal_13301) ) ;
    buf_clk new_AGEMA_reg_buffer_7452 ( .C (clk), .D (new_AGEMA_signal_5544), .Q (new_AGEMA_signal_13304) ) ;
    buf_clk new_AGEMA_reg_buffer_7455 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T1), .Q (new_AGEMA_signal_13307) ) ;
    buf_clk new_AGEMA_reg_buffer_7458 ( .C (clk), .D (new_AGEMA_signal_5123), .Q (new_AGEMA_signal_13310) ) ;
    buf_clk new_AGEMA_reg_buffer_7461 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T4), .Q (new_AGEMA_signal_13313) ) ;
    buf_clk new_AGEMA_reg_buffer_7464 ( .C (clk), .D (new_AGEMA_signal_5126), .Q (new_AGEMA_signal_13316) ) ;
    buf_clk new_AGEMA_reg_buffer_7467 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T2), .Q (new_AGEMA_signal_13319) ) ;
    buf_clk new_AGEMA_reg_buffer_7470 ( .C (clk), .D (new_AGEMA_signal_5124), .Q (new_AGEMA_signal_13322) ) ;
    buf_clk new_AGEMA_reg_buffer_7473 ( .C (clk), .D (key_s0[0]), .Q (new_AGEMA_signal_13325) ) ;
    buf_clk new_AGEMA_reg_buffer_7477 ( .C (clk), .D (key_s1[0]), .Q (new_AGEMA_signal_13329) ) ;
    buf_clk new_AGEMA_reg_buffer_7481 ( .C (clk), .D (key_s0[1]), .Q (new_AGEMA_signal_13333) ) ;
    buf_clk new_AGEMA_reg_buffer_7485 ( .C (clk), .D (key_s1[1]), .Q (new_AGEMA_signal_13337) ) ;
    buf_clk new_AGEMA_reg_buffer_7489 ( .C (clk), .D (key_s0[2]), .Q (new_AGEMA_signal_13341) ) ;
    buf_clk new_AGEMA_reg_buffer_7493 ( .C (clk), .D (key_s1[2]), .Q (new_AGEMA_signal_13345) ) ;
    buf_clk new_AGEMA_reg_buffer_7497 ( .C (clk), .D (key_s0[3]), .Q (new_AGEMA_signal_13349) ) ;
    buf_clk new_AGEMA_reg_buffer_7501 ( .C (clk), .D (key_s1[3]), .Q (new_AGEMA_signal_13353) ) ;
    buf_clk new_AGEMA_reg_buffer_7505 ( .C (clk), .D (key_s0[4]), .Q (new_AGEMA_signal_13357) ) ;
    buf_clk new_AGEMA_reg_buffer_7509 ( .C (clk), .D (key_s1[4]), .Q (new_AGEMA_signal_13361) ) ;
    buf_clk new_AGEMA_reg_buffer_7513 ( .C (clk), .D (key_s0[5]), .Q (new_AGEMA_signal_13365) ) ;
    buf_clk new_AGEMA_reg_buffer_7517 ( .C (clk), .D (key_s1[5]), .Q (new_AGEMA_signal_13369) ) ;
    buf_clk new_AGEMA_reg_buffer_7521 ( .C (clk), .D (key_s0[6]), .Q (new_AGEMA_signal_13373) ) ;
    buf_clk new_AGEMA_reg_buffer_7525 ( .C (clk), .D (key_s1[6]), .Q (new_AGEMA_signal_13377) ) ;
    buf_clk new_AGEMA_reg_buffer_7529 ( .C (clk), .D (key_s0[7]), .Q (new_AGEMA_signal_13381) ) ;
    buf_clk new_AGEMA_reg_buffer_7533 ( .C (clk), .D (key_s1[7]), .Q (new_AGEMA_signal_13385) ) ;
    buf_clk new_AGEMA_reg_buffer_7537 ( .C (clk), .D (key_s0[8]), .Q (new_AGEMA_signal_13389) ) ;
    buf_clk new_AGEMA_reg_buffer_7541 ( .C (clk), .D (key_s1[8]), .Q (new_AGEMA_signal_13393) ) ;
    buf_clk new_AGEMA_reg_buffer_7545 ( .C (clk), .D (key_s0[9]), .Q (new_AGEMA_signal_13397) ) ;
    buf_clk new_AGEMA_reg_buffer_7549 ( .C (clk), .D (key_s1[9]), .Q (new_AGEMA_signal_13401) ) ;
    buf_clk new_AGEMA_reg_buffer_7553 ( .C (clk), .D (key_s0[10]), .Q (new_AGEMA_signal_13405) ) ;
    buf_clk new_AGEMA_reg_buffer_7557 ( .C (clk), .D (key_s1[10]), .Q (new_AGEMA_signal_13409) ) ;
    buf_clk new_AGEMA_reg_buffer_7561 ( .C (clk), .D (key_s0[11]), .Q (new_AGEMA_signal_13413) ) ;
    buf_clk new_AGEMA_reg_buffer_7565 ( .C (clk), .D (key_s1[11]), .Q (new_AGEMA_signal_13417) ) ;
    buf_clk new_AGEMA_reg_buffer_7569 ( .C (clk), .D (key_s0[12]), .Q (new_AGEMA_signal_13421) ) ;
    buf_clk new_AGEMA_reg_buffer_7573 ( .C (clk), .D (key_s1[12]), .Q (new_AGEMA_signal_13425) ) ;
    buf_clk new_AGEMA_reg_buffer_7577 ( .C (clk), .D (key_s0[13]), .Q (new_AGEMA_signal_13429) ) ;
    buf_clk new_AGEMA_reg_buffer_7581 ( .C (clk), .D (key_s1[13]), .Q (new_AGEMA_signal_13433) ) ;
    buf_clk new_AGEMA_reg_buffer_7585 ( .C (clk), .D (key_s0[14]), .Q (new_AGEMA_signal_13437) ) ;
    buf_clk new_AGEMA_reg_buffer_7589 ( .C (clk), .D (key_s1[14]), .Q (new_AGEMA_signal_13441) ) ;
    buf_clk new_AGEMA_reg_buffer_7593 ( .C (clk), .D (key_s0[15]), .Q (new_AGEMA_signal_13445) ) ;
    buf_clk new_AGEMA_reg_buffer_7597 ( .C (clk), .D (key_s1[15]), .Q (new_AGEMA_signal_13449) ) ;
    buf_clk new_AGEMA_reg_buffer_7601 ( .C (clk), .D (key_s0[16]), .Q (new_AGEMA_signal_13453) ) ;
    buf_clk new_AGEMA_reg_buffer_7605 ( .C (clk), .D (key_s1[16]), .Q (new_AGEMA_signal_13457) ) ;
    buf_clk new_AGEMA_reg_buffer_7609 ( .C (clk), .D (key_s0[17]), .Q (new_AGEMA_signal_13461) ) ;
    buf_clk new_AGEMA_reg_buffer_7613 ( .C (clk), .D (key_s1[17]), .Q (new_AGEMA_signal_13465) ) ;
    buf_clk new_AGEMA_reg_buffer_7617 ( .C (clk), .D (key_s0[18]), .Q (new_AGEMA_signal_13469) ) ;
    buf_clk new_AGEMA_reg_buffer_7621 ( .C (clk), .D (key_s1[18]), .Q (new_AGEMA_signal_13473) ) ;
    buf_clk new_AGEMA_reg_buffer_7625 ( .C (clk), .D (key_s0[19]), .Q (new_AGEMA_signal_13477) ) ;
    buf_clk new_AGEMA_reg_buffer_7629 ( .C (clk), .D (key_s1[19]), .Q (new_AGEMA_signal_13481) ) ;
    buf_clk new_AGEMA_reg_buffer_7633 ( .C (clk), .D (key_s0[20]), .Q (new_AGEMA_signal_13485) ) ;
    buf_clk new_AGEMA_reg_buffer_7637 ( .C (clk), .D (key_s1[20]), .Q (new_AGEMA_signal_13489) ) ;
    buf_clk new_AGEMA_reg_buffer_7641 ( .C (clk), .D (key_s0[21]), .Q (new_AGEMA_signal_13493) ) ;
    buf_clk new_AGEMA_reg_buffer_7645 ( .C (clk), .D (key_s1[21]), .Q (new_AGEMA_signal_13497) ) ;
    buf_clk new_AGEMA_reg_buffer_7649 ( .C (clk), .D (key_s0[22]), .Q (new_AGEMA_signal_13501) ) ;
    buf_clk new_AGEMA_reg_buffer_7653 ( .C (clk), .D (key_s1[22]), .Q (new_AGEMA_signal_13505) ) ;
    buf_clk new_AGEMA_reg_buffer_7657 ( .C (clk), .D (key_s0[23]), .Q (new_AGEMA_signal_13509) ) ;
    buf_clk new_AGEMA_reg_buffer_7661 ( .C (clk), .D (key_s1[23]), .Q (new_AGEMA_signal_13513) ) ;
    buf_clk new_AGEMA_reg_buffer_7665 ( .C (clk), .D (key_s0[24]), .Q (new_AGEMA_signal_13517) ) ;
    buf_clk new_AGEMA_reg_buffer_7669 ( .C (clk), .D (key_s1[24]), .Q (new_AGEMA_signal_13521) ) ;
    buf_clk new_AGEMA_reg_buffer_7673 ( .C (clk), .D (key_s0[25]), .Q (new_AGEMA_signal_13525) ) ;
    buf_clk new_AGEMA_reg_buffer_7677 ( .C (clk), .D (key_s1[25]), .Q (new_AGEMA_signal_13529) ) ;
    buf_clk new_AGEMA_reg_buffer_7681 ( .C (clk), .D (key_s0[26]), .Q (new_AGEMA_signal_13533) ) ;
    buf_clk new_AGEMA_reg_buffer_7685 ( .C (clk), .D (key_s1[26]), .Q (new_AGEMA_signal_13537) ) ;
    buf_clk new_AGEMA_reg_buffer_7689 ( .C (clk), .D (key_s0[27]), .Q (new_AGEMA_signal_13541) ) ;
    buf_clk new_AGEMA_reg_buffer_7693 ( .C (clk), .D (key_s1[27]), .Q (new_AGEMA_signal_13545) ) ;
    buf_clk new_AGEMA_reg_buffer_7697 ( .C (clk), .D (key_s0[28]), .Q (new_AGEMA_signal_13549) ) ;
    buf_clk new_AGEMA_reg_buffer_7701 ( .C (clk), .D (key_s1[28]), .Q (new_AGEMA_signal_13553) ) ;
    buf_clk new_AGEMA_reg_buffer_7705 ( .C (clk), .D (key_s0[29]), .Q (new_AGEMA_signal_13557) ) ;
    buf_clk new_AGEMA_reg_buffer_7709 ( .C (clk), .D (key_s1[29]), .Q (new_AGEMA_signal_13561) ) ;
    buf_clk new_AGEMA_reg_buffer_7713 ( .C (clk), .D (key_s0[30]), .Q (new_AGEMA_signal_13565) ) ;
    buf_clk new_AGEMA_reg_buffer_7717 ( .C (clk), .D (key_s1[30]), .Q (new_AGEMA_signal_13569) ) ;
    buf_clk new_AGEMA_reg_buffer_7721 ( .C (clk), .D (key_s0[31]), .Q (new_AGEMA_signal_13573) ) ;
    buf_clk new_AGEMA_reg_buffer_7725 ( .C (clk), .D (key_s1[31]), .Q (new_AGEMA_signal_13577) ) ;
    buf_clk new_AGEMA_reg_buffer_7729 ( .C (clk), .D (key_s0[32]), .Q (new_AGEMA_signal_13581) ) ;
    buf_clk new_AGEMA_reg_buffer_7733 ( .C (clk), .D (key_s1[32]), .Q (new_AGEMA_signal_13585) ) ;
    buf_clk new_AGEMA_reg_buffer_7737 ( .C (clk), .D (key_s0[33]), .Q (new_AGEMA_signal_13589) ) ;
    buf_clk new_AGEMA_reg_buffer_7741 ( .C (clk), .D (key_s1[33]), .Q (new_AGEMA_signal_13593) ) ;
    buf_clk new_AGEMA_reg_buffer_7745 ( .C (clk), .D (key_s0[34]), .Q (new_AGEMA_signal_13597) ) ;
    buf_clk new_AGEMA_reg_buffer_7749 ( .C (clk), .D (key_s1[34]), .Q (new_AGEMA_signal_13601) ) ;
    buf_clk new_AGEMA_reg_buffer_7753 ( .C (clk), .D (key_s0[35]), .Q (new_AGEMA_signal_13605) ) ;
    buf_clk new_AGEMA_reg_buffer_7757 ( .C (clk), .D (key_s1[35]), .Q (new_AGEMA_signal_13609) ) ;
    buf_clk new_AGEMA_reg_buffer_7761 ( .C (clk), .D (key_s0[36]), .Q (new_AGEMA_signal_13613) ) ;
    buf_clk new_AGEMA_reg_buffer_7765 ( .C (clk), .D (key_s1[36]), .Q (new_AGEMA_signal_13617) ) ;
    buf_clk new_AGEMA_reg_buffer_7769 ( .C (clk), .D (key_s0[37]), .Q (new_AGEMA_signal_13621) ) ;
    buf_clk new_AGEMA_reg_buffer_7773 ( .C (clk), .D (key_s1[37]), .Q (new_AGEMA_signal_13625) ) ;
    buf_clk new_AGEMA_reg_buffer_7777 ( .C (clk), .D (key_s0[38]), .Q (new_AGEMA_signal_13629) ) ;
    buf_clk new_AGEMA_reg_buffer_7781 ( .C (clk), .D (key_s1[38]), .Q (new_AGEMA_signal_13633) ) ;
    buf_clk new_AGEMA_reg_buffer_7785 ( .C (clk), .D (key_s0[39]), .Q (new_AGEMA_signal_13637) ) ;
    buf_clk new_AGEMA_reg_buffer_7789 ( .C (clk), .D (key_s1[39]), .Q (new_AGEMA_signal_13641) ) ;
    buf_clk new_AGEMA_reg_buffer_7793 ( .C (clk), .D (key_s0[40]), .Q (new_AGEMA_signal_13645) ) ;
    buf_clk new_AGEMA_reg_buffer_7797 ( .C (clk), .D (key_s1[40]), .Q (new_AGEMA_signal_13649) ) ;
    buf_clk new_AGEMA_reg_buffer_7801 ( .C (clk), .D (key_s0[41]), .Q (new_AGEMA_signal_13653) ) ;
    buf_clk new_AGEMA_reg_buffer_7805 ( .C (clk), .D (key_s1[41]), .Q (new_AGEMA_signal_13657) ) ;
    buf_clk new_AGEMA_reg_buffer_7809 ( .C (clk), .D (key_s0[42]), .Q (new_AGEMA_signal_13661) ) ;
    buf_clk new_AGEMA_reg_buffer_7813 ( .C (clk), .D (key_s1[42]), .Q (new_AGEMA_signal_13665) ) ;
    buf_clk new_AGEMA_reg_buffer_7817 ( .C (clk), .D (key_s0[43]), .Q (new_AGEMA_signal_13669) ) ;
    buf_clk new_AGEMA_reg_buffer_7821 ( .C (clk), .D (key_s1[43]), .Q (new_AGEMA_signal_13673) ) ;
    buf_clk new_AGEMA_reg_buffer_7825 ( .C (clk), .D (key_s0[44]), .Q (new_AGEMA_signal_13677) ) ;
    buf_clk new_AGEMA_reg_buffer_7829 ( .C (clk), .D (key_s1[44]), .Q (new_AGEMA_signal_13681) ) ;
    buf_clk new_AGEMA_reg_buffer_7833 ( .C (clk), .D (key_s0[45]), .Q (new_AGEMA_signal_13685) ) ;
    buf_clk new_AGEMA_reg_buffer_7837 ( .C (clk), .D (key_s1[45]), .Q (new_AGEMA_signal_13689) ) ;
    buf_clk new_AGEMA_reg_buffer_7841 ( .C (clk), .D (key_s0[46]), .Q (new_AGEMA_signal_13693) ) ;
    buf_clk new_AGEMA_reg_buffer_7845 ( .C (clk), .D (key_s1[46]), .Q (new_AGEMA_signal_13697) ) ;
    buf_clk new_AGEMA_reg_buffer_7849 ( .C (clk), .D (key_s0[47]), .Q (new_AGEMA_signal_13701) ) ;
    buf_clk new_AGEMA_reg_buffer_7853 ( .C (clk), .D (key_s1[47]), .Q (new_AGEMA_signal_13705) ) ;
    buf_clk new_AGEMA_reg_buffer_7857 ( .C (clk), .D (key_s0[48]), .Q (new_AGEMA_signal_13709) ) ;
    buf_clk new_AGEMA_reg_buffer_7861 ( .C (clk), .D (key_s1[48]), .Q (new_AGEMA_signal_13713) ) ;
    buf_clk new_AGEMA_reg_buffer_7865 ( .C (clk), .D (key_s0[49]), .Q (new_AGEMA_signal_13717) ) ;
    buf_clk new_AGEMA_reg_buffer_7869 ( .C (clk), .D (key_s1[49]), .Q (new_AGEMA_signal_13721) ) ;
    buf_clk new_AGEMA_reg_buffer_7873 ( .C (clk), .D (key_s0[50]), .Q (new_AGEMA_signal_13725) ) ;
    buf_clk new_AGEMA_reg_buffer_7877 ( .C (clk), .D (key_s1[50]), .Q (new_AGEMA_signal_13729) ) ;
    buf_clk new_AGEMA_reg_buffer_7881 ( .C (clk), .D (key_s0[51]), .Q (new_AGEMA_signal_13733) ) ;
    buf_clk new_AGEMA_reg_buffer_7885 ( .C (clk), .D (key_s1[51]), .Q (new_AGEMA_signal_13737) ) ;
    buf_clk new_AGEMA_reg_buffer_7889 ( .C (clk), .D (key_s0[52]), .Q (new_AGEMA_signal_13741) ) ;
    buf_clk new_AGEMA_reg_buffer_7893 ( .C (clk), .D (key_s1[52]), .Q (new_AGEMA_signal_13745) ) ;
    buf_clk new_AGEMA_reg_buffer_7897 ( .C (clk), .D (key_s0[53]), .Q (new_AGEMA_signal_13749) ) ;
    buf_clk new_AGEMA_reg_buffer_7901 ( .C (clk), .D (key_s1[53]), .Q (new_AGEMA_signal_13753) ) ;
    buf_clk new_AGEMA_reg_buffer_7905 ( .C (clk), .D (key_s0[54]), .Q (new_AGEMA_signal_13757) ) ;
    buf_clk new_AGEMA_reg_buffer_7909 ( .C (clk), .D (key_s1[54]), .Q (new_AGEMA_signal_13761) ) ;
    buf_clk new_AGEMA_reg_buffer_7913 ( .C (clk), .D (key_s0[55]), .Q (new_AGEMA_signal_13765) ) ;
    buf_clk new_AGEMA_reg_buffer_7917 ( .C (clk), .D (key_s1[55]), .Q (new_AGEMA_signal_13769) ) ;
    buf_clk new_AGEMA_reg_buffer_7921 ( .C (clk), .D (key_s0[56]), .Q (new_AGEMA_signal_13773) ) ;
    buf_clk new_AGEMA_reg_buffer_7925 ( .C (clk), .D (key_s1[56]), .Q (new_AGEMA_signal_13777) ) ;
    buf_clk new_AGEMA_reg_buffer_7929 ( .C (clk), .D (key_s0[57]), .Q (new_AGEMA_signal_13781) ) ;
    buf_clk new_AGEMA_reg_buffer_7933 ( .C (clk), .D (key_s1[57]), .Q (new_AGEMA_signal_13785) ) ;
    buf_clk new_AGEMA_reg_buffer_7937 ( .C (clk), .D (key_s0[58]), .Q (new_AGEMA_signal_13789) ) ;
    buf_clk new_AGEMA_reg_buffer_7941 ( .C (clk), .D (key_s1[58]), .Q (new_AGEMA_signal_13793) ) ;
    buf_clk new_AGEMA_reg_buffer_7945 ( .C (clk), .D (key_s0[59]), .Q (new_AGEMA_signal_13797) ) ;
    buf_clk new_AGEMA_reg_buffer_7949 ( .C (clk), .D (key_s1[59]), .Q (new_AGEMA_signal_13801) ) ;
    buf_clk new_AGEMA_reg_buffer_7953 ( .C (clk), .D (key_s0[60]), .Q (new_AGEMA_signal_13805) ) ;
    buf_clk new_AGEMA_reg_buffer_7957 ( .C (clk), .D (key_s1[60]), .Q (new_AGEMA_signal_13809) ) ;
    buf_clk new_AGEMA_reg_buffer_7961 ( .C (clk), .D (key_s0[61]), .Q (new_AGEMA_signal_13813) ) ;
    buf_clk new_AGEMA_reg_buffer_7965 ( .C (clk), .D (key_s1[61]), .Q (new_AGEMA_signal_13817) ) ;
    buf_clk new_AGEMA_reg_buffer_7969 ( .C (clk), .D (key_s0[62]), .Q (new_AGEMA_signal_13821) ) ;
    buf_clk new_AGEMA_reg_buffer_7973 ( .C (clk), .D (key_s1[62]), .Q (new_AGEMA_signal_13825) ) ;
    buf_clk new_AGEMA_reg_buffer_7977 ( .C (clk), .D (key_s0[63]), .Q (new_AGEMA_signal_13829) ) ;
    buf_clk new_AGEMA_reg_buffer_7981 ( .C (clk), .D (key_s1[63]), .Q (new_AGEMA_signal_13833) ) ;
    buf_clk new_AGEMA_reg_buffer_7985 ( .C (clk), .D (key_s0[64]), .Q (new_AGEMA_signal_13837) ) ;
    buf_clk new_AGEMA_reg_buffer_7989 ( .C (clk), .D (key_s1[64]), .Q (new_AGEMA_signal_13841) ) ;
    buf_clk new_AGEMA_reg_buffer_7993 ( .C (clk), .D (key_s0[65]), .Q (new_AGEMA_signal_13845) ) ;
    buf_clk new_AGEMA_reg_buffer_7997 ( .C (clk), .D (key_s1[65]), .Q (new_AGEMA_signal_13849) ) ;
    buf_clk new_AGEMA_reg_buffer_8001 ( .C (clk), .D (key_s0[66]), .Q (new_AGEMA_signal_13853) ) ;
    buf_clk new_AGEMA_reg_buffer_8005 ( .C (clk), .D (key_s1[66]), .Q (new_AGEMA_signal_13857) ) ;
    buf_clk new_AGEMA_reg_buffer_8009 ( .C (clk), .D (key_s0[67]), .Q (new_AGEMA_signal_13861) ) ;
    buf_clk new_AGEMA_reg_buffer_8013 ( .C (clk), .D (key_s1[67]), .Q (new_AGEMA_signal_13865) ) ;
    buf_clk new_AGEMA_reg_buffer_8017 ( .C (clk), .D (key_s0[68]), .Q (new_AGEMA_signal_13869) ) ;
    buf_clk new_AGEMA_reg_buffer_8021 ( .C (clk), .D (key_s1[68]), .Q (new_AGEMA_signal_13873) ) ;
    buf_clk new_AGEMA_reg_buffer_8025 ( .C (clk), .D (key_s0[69]), .Q (new_AGEMA_signal_13877) ) ;
    buf_clk new_AGEMA_reg_buffer_8029 ( .C (clk), .D (key_s1[69]), .Q (new_AGEMA_signal_13881) ) ;
    buf_clk new_AGEMA_reg_buffer_8033 ( .C (clk), .D (key_s0[70]), .Q (new_AGEMA_signal_13885) ) ;
    buf_clk new_AGEMA_reg_buffer_8037 ( .C (clk), .D (key_s1[70]), .Q (new_AGEMA_signal_13889) ) ;
    buf_clk new_AGEMA_reg_buffer_8041 ( .C (clk), .D (key_s0[71]), .Q (new_AGEMA_signal_13893) ) ;
    buf_clk new_AGEMA_reg_buffer_8045 ( .C (clk), .D (key_s1[71]), .Q (new_AGEMA_signal_13897) ) ;
    buf_clk new_AGEMA_reg_buffer_8049 ( .C (clk), .D (key_s0[72]), .Q (new_AGEMA_signal_13901) ) ;
    buf_clk new_AGEMA_reg_buffer_8053 ( .C (clk), .D (key_s1[72]), .Q (new_AGEMA_signal_13905) ) ;
    buf_clk new_AGEMA_reg_buffer_8057 ( .C (clk), .D (key_s0[73]), .Q (new_AGEMA_signal_13909) ) ;
    buf_clk new_AGEMA_reg_buffer_8061 ( .C (clk), .D (key_s1[73]), .Q (new_AGEMA_signal_13913) ) ;
    buf_clk new_AGEMA_reg_buffer_8065 ( .C (clk), .D (key_s0[74]), .Q (new_AGEMA_signal_13917) ) ;
    buf_clk new_AGEMA_reg_buffer_8069 ( .C (clk), .D (key_s1[74]), .Q (new_AGEMA_signal_13921) ) ;
    buf_clk new_AGEMA_reg_buffer_8073 ( .C (clk), .D (key_s0[75]), .Q (new_AGEMA_signal_13925) ) ;
    buf_clk new_AGEMA_reg_buffer_8077 ( .C (clk), .D (key_s1[75]), .Q (new_AGEMA_signal_13929) ) ;
    buf_clk new_AGEMA_reg_buffer_8081 ( .C (clk), .D (key_s0[76]), .Q (new_AGEMA_signal_13933) ) ;
    buf_clk new_AGEMA_reg_buffer_8085 ( .C (clk), .D (key_s1[76]), .Q (new_AGEMA_signal_13937) ) ;
    buf_clk new_AGEMA_reg_buffer_8089 ( .C (clk), .D (key_s0[77]), .Q (new_AGEMA_signal_13941) ) ;
    buf_clk new_AGEMA_reg_buffer_8093 ( .C (clk), .D (key_s1[77]), .Q (new_AGEMA_signal_13945) ) ;
    buf_clk new_AGEMA_reg_buffer_8097 ( .C (clk), .D (key_s0[78]), .Q (new_AGEMA_signal_13949) ) ;
    buf_clk new_AGEMA_reg_buffer_8101 ( .C (clk), .D (key_s1[78]), .Q (new_AGEMA_signal_13953) ) ;
    buf_clk new_AGEMA_reg_buffer_8105 ( .C (clk), .D (key_s0[79]), .Q (new_AGEMA_signal_13957) ) ;
    buf_clk new_AGEMA_reg_buffer_8109 ( .C (clk), .D (key_s1[79]), .Q (new_AGEMA_signal_13961) ) ;
    buf_clk new_AGEMA_reg_buffer_8113 ( .C (clk), .D (key_s0[80]), .Q (new_AGEMA_signal_13965) ) ;
    buf_clk new_AGEMA_reg_buffer_8117 ( .C (clk), .D (key_s1[80]), .Q (new_AGEMA_signal_13969) ) ;
    buf_clk new_AGEMA_reg_buffer_8121 ( .C (clk), .D (key_s0[81]), .Q (new_AGEMA_signal_13973) ) ;
    buf_clk new_AGEMA_reg_buffer_8125 ( .C (clk), .D (key_s1[81]), .Q (new_AGEMA_signal_13977) ) ;
    buf_clk new_AGEMA_reg_buffer_8129 ( .C (clk), .D (key_s0[82]), .Q (new_AGEMA_signal_13981) ) ;
    buf_clk new_AGEMA_reg_buffer_8133 ( .C (clk), .D (key_s1[82]), .Q (new_AGEMA_signal_13985) ) ;
    buf_clk new_AGEMA_reg_buffer_8137 ( .C (clk), .D (key_s0[83]), .Q (new_AGEMA_signal_13989) ) ;
    buf_clk new_AGEMA_reg_buffer_8141 ( .C (clk), .D (key_s1[83]), .Q (new_AGEMA_signal_13993) ) ;
    buf_clk new_AGEMA_reg_buffer_8145 ( .C (clk), .D (key_s0[84]), .Q (new_AGEMA_signal_13997) ) ;
    buf_clk new_AGEMA_reg_buffer_8149 ( .C (clk), .D (key_s1[84]), .Q (new_AGEMA_signal_14001) ) ;
    buf_clk new_AGEMA_reg_buffer_8153 ( .C (clk), .D (key_s0[85]), .Q (new_AGEMA_signal_14005) ) ;
    buf_clk new_AGEMA_reg_buffer_8157 ( .C (clk), .D (key_s1[85]), .Q (new_AGEMA_signal_14009) ) ;
    buf_clk new_AGEMA_reg_buffer_8161 ( .C (clk), .D (key_s0[86]), .Q (new_AGEMA_signal_14013) ) ;
    buf_clk new_AGEMA_reg_buffer_8165 ( .C (clk), .D (key_s1[86]), .Q (new_AGEMA_signal_14017) ) ;
    buf_clk new_AGEMA_reg_buffer_8169 ( .C (clk), .D (key_s0[87]), .Q (new_AGEMA_signal_14021) ) ;
    buf_clk new_AGEMA_reg_buffer_8173 ( .C (clk), .D (key_s1[87]), .Q (new_AGEMA_signal_14025) ) ;
    buf_clk new_AGEMA_reg_buffer_8177 ( .C (clk), .D (key_s0[88]), .Q (new_AGEMA_signal_14029) ) ;
    buf_clk new_AGEMA_reg_buffer_8181 ( .C (clk), .D (key_s1[88]), .Q (new_AGEMA_signal_14033) ) ;
    buf_clk new_AGEMA_reg_buffer_8185 ( .C (clk), .D (key_s0[89]), .Q (new_AGEMA_signal_14037) ) ;
    buf_clk new_AGEMA_reg_buffer_8189 ( .C (clk), .D (key_s1[89]), .Q (new_AGEMA_signal_14041) ) ;
    buf_clk new_AGEMA_reg_buffer_8193 ( .C (clk), .D (key_s0[90]), .Q (new_AGEMA_signal_14045) ) ;
    buf_clk new_AGEMA_reg_buffer_8197 ( .C (clk), .D (key_s1[90]), .Q (new_AGEMA_signal_14049) ) ;
    buf_clk new_AGEMA_reg_buffer_8201 ( .C (clk), .D (key_s0[91]), .Q (new_AGEMA_signal_14053) ) ;
    buf_clk new_AGEMA_reg_buffer_8205 ( .C (clk), .D (key_s1[91]), .Q (new_AGEMA_signal_14057) ) ;
    buf_clk new_AGEMA_reg_buffer_8209 ( .C (clk), .D (key_s0[92]), .Q (new_AGEMA_signal_14061) ) ;
    buf_clk new_AGEMA_reg_buffer_8213 ( .C (clk), .D (key_s1[92]), .Q (new_AGEMA_signal_14065) ) ;
    buf_clk new_AGEMA_reg_buffer_8217 ( .C (clk), .D (key_s0[93]), .Q (new_AGEMA_signal_14069) ) ;
    buf_clk new_AGEMA_reg_buffer_8221 ( .C (clk), .D (key_s1[93]), .Q (new_AGEMA_signal_14073) ) ;
    buf_clk new_AGEMA_reg_buffer_8225 ( .C (clk), .D (key_s0[94]), .Q (new_AGEMA_signal_14077) ) ;
    buf_clk new_AGEMA_reg_buffer_8229 ( .C (clk), .D (key_s1[94]), .Q (new_AGEMA_signal_14081) ) ;
    buf_clk new_AGEMA_reg_buffer_8233 ( .C (clk), .D (key_s0[95]), .Q (new_AGEMA_signal_14085) ) ;
    buf_clk new_AGEMA_reg_buffer_8237 ( .C (clk), .D (key_s1[95]), .Q (new_AGEMA_signal_14089) ) ;
    buf_clk new_AGEMA_reg_buffer_8241 ( .C (clk), .D (key_s0[96]), .Q (new_AGEMA_signal_14093) ) ;
    buf_clk new_AGEMA_reg_buffer_8245 ( .C (clk), .D (key_s1[96]), .Q (new_AGEMA_signal_14097) ) ;
    buf_clk new_AGEMA_reg_buffer_8249 ( .C (clk), .D (key_s0[97]), .Q (new_AGEMA_signal_14101) ) ;
    buf_clk new_AGEMA_reg_buffer_8253 ( .C (clk), .D (key_s1[97]), .Q (new_AGEMA_signal_14105) ) ;
    buf_clk new_AGEMA_reg_buffer_8257 ( .C (clk), .D (key_s0[98]), .Q (new_AGEMA_signal_14109) ) ;
    buf_clk new_AGEMA_reg_buffer_8261 ( .C (clk), .D (key_s1[98]), .Q (new_AGEMA_signal_14113) ) ;
    buf_clk new_AGEMA_reg_buffer_8265 ( .C (clk), .D (key_s0[99]), .Q (new_AGEMA_signal_14117) ) ;
    buf_clk new_AGEMA_reg_buffer_8269 ( .C (clk), .D (key_s1[99]), .Q (new_AGEMA_signal_14121) ) ;
    buf_clk new_AGEMA_reg_buffer_8273 ( .C (clk), .D (key_s0[100]), .Q (new_AGEMA_signal_14125) ) ;
    buf_clk new_AGEMA_reg_buffer_8277 ( .C (clk), .D (key_s1[100]), .Q (new_AGEMA_signal_14129) ) ;
    buf_clk new_AGEMA_reg_buffer_8281 ( .C (clk), .D (key_s0[101]), .Q (new_AGEMA_signal_14133) ) ;
    buf_clk new_AGEMA_reg_buffer_8285 ( .C (clk), .D (key_s1[101]), .Q (new_AGEMA_signal_14137) ) ;
    buf_clk new_AGEMA_reg_buffer_8289 ( .C (clk), .D (key_s0[102]), .Q (new_AGEMA_signal_14141) ) ;
    buf_clk new_AGEMA_reg_buffer_8293 ( .C (clk), .D (key_s1[102]), .Q (new_AGEMA_signal_14145) ) ;
    buf_clk new_AGEMA_reg_buffer_8297 ( .C (clk), .D (key_s0[103]), .Q (new_AGEMA_signal_14149) ) ;
    buf_clk new_AGEMA_reg_buffer_8301 ( .C (clk), .D (key_s1[103]), .Q (new_AGEMA_signal_14153) ) ;
    buf_clk new_AGEMA_reg_buffer_8305 ( .C (clk), .D (key_s0[104]), .Q (new_AGEMA_signal_14157) ) ;
    buf_clk new_AGEMA_reg_buffer_8309 ( .C (clk), .D (key_s1[104]), .Q (new_AGEMA_signal_14161) ) ;
    buf_clk new_AGEMA_reg_buffer_8313 ( .C (clk), .D (key_s0[105]), .Q (new_AGEMA_signal_14165) ) ;
    buf_clk new_AGEMA_reg_buffer_8317 ( .C (clk), .D (key_s1[105]), .Q (new_AGEMA_signal_14169) ) ;
    buf_clk new_AGEMA_reg_buffer_8321 ( .C (clk), .D (key_s0[106]), .Q (new_AGEMA_signal_14173) ) ;
    buf_clk new_AGEMA_reg_buffer_8325 ( .C (clk), .D (key_s1[106]), .Q (new_AGEMA_signal_14177) ) ;
    buf_clk new_AGEMA_reg_buffer_8329 ( .C (clk), .D (key_s0[107]), .Q (new_AGEMA_signal_14181) ) ;
    buf_clk new_AGEMA_reg_buffer_8333 ( .C (clk), .D (key_s1[107]), .Q (new_AGEMA_signal_14185) ) ;
    buf_clk new_AGEMA_reg_buffer_8337 ( .C (clk), .D (key_s0[108]), .Q (new_AGEMA_signal_14189) ) ;
    buf_clk new_AGEMA_reg_buffer_8341 ( .C (clk), .D (key_s1[108]), .Q (new_AGEMA_signal_14193) ) ;
    buf_clk new_AGEMA_reg_buffer_8345 ( .C (clk), .D (key_s0[109]), .Q (new_AGEMA_signal_14197) ) ;
    buf_clk new_AGEMA_reg_buffer_8349 ( .C (clk), .D (key_s1[109]), .Q (new_AGEMA_signal_14201) ) ;
    buf_clk new_AGEMA_reg_buffer_8353 ( .C (clk), .D (key_s0[110]), .Q (new_AGEMA_signal_14205) ) ;
    buf_clk new_AGEMA_reg_buffer_8357 ( .C (clk), .D (key_s1[110]), .Q (new_AGEMA_signal_14209) ) ;
    buf_clk new_AGEMA_reg_buffer_8361 ( .C (clk), .D (key_s0[111]), .Q (new_AGEMA_signal_14213) ) ;
    buf_clk new_AGEMA_reg_buffer_8365 ( .C (clk), .D (key_s1[111]), .Q (new_AGEMA_signal_14217) ) ;
    buf_clk new_AGEMA_reg_buffer_8369 ( .C (clk), .D (key_s0[112]), .Q (new_AGEMA_signal_14221) ) ;
    buf_clk new_AGEMA_reg_buffer_8373 ( .C (clk), .D (key_s1[112]), .Q (new_AGEMA_signal_14225) ) ;
    buf_clk new_AGEMA_reg_buffer_8377 ( .C (clk), .D (key_s0[113]), .Q (new_AGEMA_signal_14229) ) ;
    buf_clk new_AGEMA_reg_buffer_8381 ( .C (clk), .D (key_s1[113]), .Q (new_AGEMA_signal_14233) ) ;
    buf_clk new_AGEMA_reg_buffer_8385 ( .C (clk), .D (key_s0[114]), .Q (new_AGEMA_signal_14237) ) ;
    buf_clk new_AGEMA_reg_buffer_8389 ( .C (clk), .D (key_s1[114]), .Q (new_AGEMA_signal_14241) ) ;
    buf_clk new_AGEMA_reg_buffer_8393 ( .C (clk), .D (key_s0[115]), .Q (new_AGEMA_signal_14245) ) ;
    buf_clk new_AGEMA_reg_buffer_8397 ( .C (clk), .D (key_s1[115]), .Q (new_AGEMA_signal_14249) ) ;
    buf_clk new_AGEMA_reg_buffer_8401 ( .C (clk), .D (key_s0[116]), .Q (new_AGEMA_signal_14253) ) ;
    buf_clk new_AGEMA_reg_buffer_8405 ( .C (clk), .D (key_s1[116]), .Q (new_AGEMA_signal_14257) ) ;
    buf_clk new_AGEMA_reg_buffer_8409 ( .C (clk), .D (key_s0[117]), .Q (new_AGEMA_signal_14261) ) ;
    buf_clk new_AGEMA_reg_buffer_8413 ( .C (clk), .D (key_s1[117]), .Q (new_AGEMA_signal_14265) ) ;
    buf_clk new_AGEMA_reg_buffer_8417 ( .C (clk), .D (key_s0[118]), .Q (new_AGEMA_signal_14269) ) ;
    buf_clk new_AGEMA_reg_buffer_8421 ( .C (clk), .D (key_s1[118]), .Q (new_AGEMA_signal_14273) ) ;
    buf_clk new_AGEMA_reg_buffer_8425 ( .C (clk), .D (key_s0[119]), .Q (new_AGEMA_signal_14277) ) ;
    buf_clk new_AGEMA_reg_buffer_8429 ( .C (clk), .D (key_s1[119]), .Q (new_AGEMA_signal_14281) ) ;
    buf_clk new_AGEMA_reg_buffer_8433 ( .C (clk), .D (key_s0[120]), .Q (new_AGEMA_signal_14285) ) ;
    buf_clk new_AGEMA_reg_buffer_8437 ( .C (clk), .D (key_s1[120]), .Q (new_AGEMA_signal_14289) ) ;
    buf_clk new_AGEMA_reg_buffer_8441 ( .C (clk), .D (key_s0[121]), .Q (new_AGEMA_signal_14293) ) ;
    buf_clk new_AGEMA_reg_buffer_8445 ( .C (clk), .D (key_s1[121]), .Q (new_AGEMA_signal_14297) ) ;
    buf_clk new_AGEMA_reg_buffer_8449 ( .C (clk), .D (key_s0[122]), .Q (new_AGEMA_signal_14301) ) ;
    buf_clk new_AGEMA_reg_buffer_8453 ( .C (clk), .D (key_s1[122]), .Q (new_AGEMA_signal_14305) ) ;
    buf_clk new_AGEMA_reg_buffer_8457 ( .C (clk), .D (key_s0[123]), .Q (new_AGEMA_signal_14309) ) ;
    buf_clk new_AGEMA_reg_buffer_8461 ( .C (clk), .D (key_s1[123]), .Q (new_AGEMA_signal_14313) ) ;
    buf_clk new_AGEMA_reg_buffer_8465 ( .C (clk), .D (key_s0[124]), .Q (new_AGEMA_signal_14317) ) ;
    buf_clk new_AGEMA_reg_buffer_8469 ( .C (clk), .D (key_s1[124]), .Q (new_AGEMA_signal_14321) ) ;
    buf_clk new_AGEMA_reg_buffer_8473 ( .C (clk), .D (key_s0[125]), .Q (new_AGEMA_signal_14325) ) ;
    buf_clk new_AGEMA_reg_buffer_8477 ( .C (clk), .D (key_s1[125]), .Q (new_AGEMA_signal_14329) ) ;
    buf_clk new_AGEMA_reg_buffer_8481 ( .C (clk), .D (key_s0[126]), .Q (new_AGEMA_signal_14333) ) ;
    buf_clk new_AGEMA_reg_buffer_8485 ( .C (clk), .D (key_s1[126]), .Q (new_AGEMA_signal_14337) ) ;
    buf_clk new_AGEMA_reg_buffer_8489 ( .C (clk), .D (key_s0[127]), .Q (new_AGEMA_signal_14341) ) ;
    buf_clk new_AGEMA_reg_buffer_8493 ( .C (clk), .D (key_s1[127]), .Q (new_AGEMA_signal_14345) ) ;
    buf_clk new_AGEMA_reg_buffer_8497 ( .C (clk), .D (RoundKey[9]), .Q (new_AGEMA_signal_14349) ) ;
    buf_clk new_AGEMA_reg_buffer_8501 ( .C (clk), .D (new_AGEMA_signal_4931), .Q (new_AGEMA_signal_14353) ) ;
    buf_clk new_AGEMA_reg_buffer_8505 ( .C (clk), .D (RoundKey[8]), .Q (new_AGEMA_signal_14357) ) ;
    buf_clk new_AGEMA_reg_buffer_8509 ( .C (clk), .D (new_AGEMA_signal_4898), .Q (new_AGEMA_signal_14361) ) ;
    buf_clk new_AGEMA_reg_buffer_8513 ( .C (clk), .D (RoundKey[7]), .Q (new_AGEMA_signal_14365) ) ;
    buf_clk new_AGEMA_reg_buffer_8517 ( .C (clk), .D (new_AGEMA_signal_4865), .Q (new_AGEMA_signal_14369) ) ;
    buf_clk new_AGEMA_reg_buffer_8521 ( .C (clk), .D (RoundKey[6]), .Q (new_AGEMA_signal_14373) ) ;
    buf_clk new_AGEMA_reg_buffer_8525 ( .C (clk), .D (new_AGEMA_signal_4832), .Q (new_AGEMA_signal_14377) ) ;
    buf_clk new_AGEMA_reg_buffer_8529 ( .C (clk), .D (RoundKey[5]), .Q (new_AGEMA_signal_14381) ) ;
    buf_clk new_AGEMA_reg_buffer_8533 ( .C (clk), .D (new_AGEMA_signal_4799), .Q (new_AGEMA_signal_14385) ) ;
    buf_clk new_AGEMA_reg_buffer_8537 ( .C (clk), .D (RoundKey[4]), .Q (new_AGEMA_signal_14389) ) ;
    buf_clk new_AGEMA_reg_buffer_8541 ( .C (clk), .D (new_AGEMA_signal_4766), .Q (new_AGEMA_signal_14393) ) ;
    buf_clk new_AGEMA_reg_buffer_8545 ( .C (clk), .D (RoundKey[41]), .Q (new_AGEMA_signal_14397) ) ;
    buf_clk new_AGEMA_reg_buffer_8549 ( .C (clk), .D (new_AGEMA_signal_4739), .Q (new_AGEMA_signal_14401) ) ;
    buf_clk new_AGEMA_reg_buffer_8553 ( .C (clk), .D (RoundKey[73]), .Q (new_AGEMA_signal_14405) ) ;
    buf_clk new_AGEMA_reg_buffer_8557 ( .C (clk), .D (new_AGEMA_signal_4844), .Q (new_AGEMA_signal_14409) ) ;
    buf_clk new_AGEMA_reg_buffer_8561 ( .C (clk), .D (RoundKey[40]), .Q (new_AGEMA_signal_14413) ) ;
    buf_clk new_AGEMA_reg_buffer_8565 ( .C (clk), .D (new_AGEMA_signal_4736), .Q (new_AGEMA_signal_14417) ) ;
    buf_clk new_AGEMA_reg_buffer_8569 ( .C (clk), .D (RoundKey[72]), .Q (new_AGEMA_signal_14421) ) ;
    buf_clk new_AGEMA_reg_buffer_8573 ( .C (clk), .D (new_AGEMA_signal_4841), .Q (new_AGEMA_signal_14425) ) ;
    buf_clk new_AGEMA_reg_buffer_8577 ( .C (clk), .D (RoundKey[3]), .Q (new_AGEMA_signal_14429) ) ;
    buf_clk new_AGEMA_reg_buffer_8581 ( .C (clk), .D (new_AGEMA_signal_4733), .Q (new_AGEMA_signal_14433) ) ;
    buf_clk new_AGEMA_reg_buffer_8585 ( .C (clk), .D (RoundKey[39]), .Q (new_AGEMA_signal_14437) ) ;
    buf_clk new_AGEMA_reg_buffer_8589 ( .C (clk), .D (new_AGEMA_signal_4730), .Q (new_AGEMA_signal_14441) ) ;
    buf_clk new_AGEMA_reg_buffer_8593 ( .C (clk), .D (RoundKey[71]), .Q (new_AGEMA_signal_14445) ) ;
    buf_clk new_AGEMA_reg_buffer_8597 ( .C (clk), .D (new_AGEMA_signal_4838), .Q (new_AGEMA_signal_14449) ) ;
    buf_clk new_AGEMA_reg_buffer_8601 ( .C (clk), .D (RoundKey[38]), .Q (new_AGEMA_signal_14453) ) ;
    buf_clk new_AGEMA_reg_buffer_8605 ( .C (clk), .D (new_AGEMA_signal_4727), .Q (new_AGEMA_signal_14457) ) ;
    buf_clk new_AGEMA_reg_buffer_8609 ( .C (clk), .D (RoundKey[70]), .Q (new_AGEMA_signal_14461) ) ;
    buf_clk new_AGEMA_reg_buffer_8613 ( .C (clk), .D (new_AGEMA_signal_4835), .Q (new_AGEMA_signal_14465) ) ;
    buf_clk new_AGEMA_reg_buffer_8617 ( .C (clk), .D (RoundKey[37]), .Q (new_AGEMA_signal_14469) ) ;
    buf_clk new_AGEMA_reg_buffer_8621 ( .C (clk), .D (new_AGEMA_signal_4724), .Q (new_AGEMA_signal_14473) ) ;
    buf_clk new_AGEMA_reg_buffer_8625 ( .C (clk), .D (RoundKey[69]), .Q (new_AGEMA_signal_14477) ) ;
    buf_clk new_AGEMA_reg_buffer_8629 ( .C (clk), .D (new_AGEMA_signal_4829), .Q (new_AGEMA_signal_14481) ) ;
    buf_clk new_AGEMA_reg_buffer_8633 ( .C (clk), .D (RoundKey[36]), .Q (new_AGEMA_signal_14485) ) ;
    buf_clk new_AGEMA_reg_buffer_8637 ( .C (clk), .D (new_AGEMA_signal_4721), .Q (new_AGEMA_signal_14489) ) ;
    buf_clk new_AGEMA_reg_buffer_8641 ( .C (clk), .D (RoundKey[68]), .Q (new_AGEMA_signal_14493) ) ;
    buf_clk new_AGEMA_reg_buffer_8645 ( .C (clk), .D (new_AGEMA_signal_4826), .Q (new_AGEMA_signal_14497) ) ;
    buf_clk new_AGEMA_reg_buffer_8649 ( .C (clk), .D (RoundKey[35]), .Q (new_AGEMA_signal_14501) ) ;
    buf_clk new_AGEMA_reg_buffer_8653 ( .C (clk), .D (new_AGEMA_signal_4718), .Q (new_AGEMA_signal_14505) ) ;
    buf_clk new_AGEMA_reg_buffer_8657 ( .C (clk), .D (RoundKey[67]), .Q (new_AGEMA_signal_14509) ) ;
    buf_clk new_AGEMA_reg_buffer_8661 ( .C (clk), .D (new_AGEMA_signal_4823), .Q (new_AGEMA_signal_14513) ) ;
    buf_clk new_AGEMA_reg_buffer_8665 ( .C (clk), .D (RoundKey[99]), .Q (new_AGEMA_signal_14517) ) ;
    buf_clk new_AGEMA_reg_buffer_8669 ( .C (clk), .D (new_AGEMA_signal_4928), .Q (new_AGEMA_signal_14521) ) ;
    buf_clk new_AGEMA_reg_buffer_8673 ( .C (clk), .D (RoundKey[31]), .Q (new_AGEMA_signal_14525) ) ;
    buf_clk new_AGEMA_reg_buffer_8677 ( .C (clk), .D (new_AGEMA_signal_4706), .Q (new_AGEMA_signal_14529) ) ;
    buf_clk new_AGEMA_reg_buffer_8681 ( .C (clk), .D (RoundKey[63]), .Q (new_AGEMA_signal_14533) ) ;
    buf_clk new_AGEMA_reg_buffer_8685 ( .C (clk), .D (new_AGEMA_signal_4811), .Q (new_AGEMA_signal_14537) ) ;
    buf_clk new_AGEMA_reg_buffer_8689 ( .C (clk), .D (RoundKey[95]), .Q (new_AGEMA_signal_14541) ) ;
    buf_clk new_AGEMA_reg_buffer_8693 ( .C (clk), .D (new_AGEMA_signal_4916), .Q (new_AGEMA_signal_14545) ) ;
    buf_clk new_AGEMA_reg_buffer_8697 ( .C (clk), .D (RoundKey[30]), .Q (new_AGEMA_signal_14549) ) ;
    buf_clk new_AGEMA_reg_buffer_8701 ( .C (clk), .D (new_AGEMA_signal_4703), .Q (new_AGEMA_signal_14553) ) ;
    buf_clk new_AGEMA_reg_buffer_8705 ( .C (clk), .D (RoundKey[62]), .Q (new_AGEMA_signal_14557) ) ;
    buf_clk new_AGEMA_reg_buffer_8709 ( .C (clk), .D (new_AGEMA_signal_4808), .Q (new_AGEMA_signal_14561) ) ;
    buf_clk new_AGEMA_reg_buffer_8713 ( .C (clk), .D (RoundKey[94]), .Q (new_AGEMA_signal_14565) ) ;
    buf_clk new_AGEMA_reg_buffer_8717 ( .C (clk), .D (new_AGEMA_signal_4913), .Q (new_AGEMA_signal_14569) ) ;
    buf_clk new_AGEMA_reg_buffer_8721 ( .C (clk), .D (RoundKey[2]), .Q (new_AGEMA_signal_14573) ) ;
    buf_clk new_AGEMA_reg_buffer_8725 ( .C (clk), .D (new_AGEMA_signal_4700), .Q (new_AGEMA_signal_14577) ) ;
    buf_clk new_AGEMA_reg_buffer_8729 ( .C (clk), .D (RoundKey[34]), .Q (new_AGEMA_signal_14581) ) ;
    buf_clk new_AGEMA_reg_buffer_8733 ( .C (clk), .D (new_AGEMA_signal_4715), .Q (new_AGEMA_signal_14585) ) ;
    buf_clk new_AGEMA_reg_buffer_8737 ( .C (clk), .D (RoundKey[66]), .Q (new_AGEMA_signal_14589) ) ;
    buf_clk new_AGEMA_reg_buffer_8741 ( .C (clk), .D (new_AGEMA_signal_4820), .Q (new_AGEMA_signal_14593) ) ;
    buf_clk new_AGEMA_reg_buffer_8745 ( .C (clk), .D (RoundKey[98]), .Q (new_AGEMA_signal_14597) ) ;
    buf_clk new_AGEMA_reg_buffer_8749 ( .C (clk), .D (new_AGEMA_signal_4925), .Q (new_AGEMA_signal_14601) ) ;
    buf_clk new_AGEMA_reg_buffer_8753 ( .C (clk), .D (RoundKey[29]), .Q (new_AGEMA_signal_14605) ) ;
    buf_clk new_AGEMA_reg_buffer_8757 ( .C (clk), .D (new_AGEMA_signal_4697), .Q (new_AGEMA_signal_14609) ) ;
    buf_clk new_AGEMA_reg_buffer_8761 ( .C (clk), .D (RoundKey[61]), .Q (new_AGEMA_signal_14613) ) ;
    buf_clk new_AGEMA_reg_buffer_8765 ( .C (clk), .D (new_AGEMA_signal_4805), .Q (new_AGEMA_signal_14617) ) ;
    buf_clk new_AGEMA_reg_buffer_8769 ( .C (clk), .D (RoundKey[93]), .Q (new_AGEMA_signal_14621) ) ;
    buf_clk new_AGEMA_reg_buffer_8773 ( .C (clk), .D (new_AGEMA_signal_4910), .Q (new_AGEMA_signal_14625) ) ;
    buf_clk new_AGEMA_reg_buffer_8777 ( .C (clk), .D (RoundKey[28]), .Q (new_AGEMA_signal_14629) ) ;
    buf_clk new_AGEMA_reg_buffer_8781 ( .C (clk), .D (new_AGEMA_signal_4694), .Q (new_AGEMA_signal_14633) ) ;
    buf_clk new_AGEMA_reg_buffer_8785 ( .C (clk), .D (RoundKey[60]), .Q (new_AGEMA_signal_14637) ) ;
    buf_clk new_AGEMA_reg_buffer_8789 ( .C (clk), .D (new_AGEMA_signal_4802), .Q (new_AGEMA_signal_14641) ) ;
    buf_clk new_AGEMA_reg_buffer_8793 ( .C (clk), .D (RoundKey[92]), .Q (new_AGEMA_signal_14645) ) ;
    buf_clk new_AGEMA_reg_buffer_8797 ( .C (clk), .D (new_AGEMA_signal_4907), .Q (new_AGEMA_signal_14649) ) ;
    buf_clk new_AGEMA_reg_buffer_8801 ( .C (clk), .D (RoundKey[27]), .Q (new_AGEMA_signal_14653) ) ;
    buf_clk new_AGEMA_reg_buffer_8805 ( .C (clk), .D (new_AGEMA_signal_4691), .Q (new_AGEMA_signal_14657) ) ;
    buf_clk new_AGEMA_reg_buffer_8809 ( .C (clk), .D (RoundKey[59]), .Q (new_AGEMA_signal_14661) ) ;
    buf_clk new_AGEMA_reg_buffer_8813 ( .C (clk), .D (new_AGEMA_signal_4796), .Q (new_AGEMA_signal_14665) ) ;
    buf_clk new_AGEMA_reg_buffer_8817 ( .C (clk), .D (RoundKey[91]), .Q (new_AGEMA_signal_14669) ) ;
    buf_clk new_AGEMA_reg_buffer_8821 ( .C (clk), .D (new_AGEMA_signal_4904), .Q (new_AGEMA_signal_14673) ) ;
    buf_clk new_AGEMA_reg_buffer_8825 ( .C (clk), .D (RoundKey[26]), .Q (new_AGEMA_signal_14677) ) ;
    buf_clk new_AGEMA_reg_buffer_8829 ( .C (clk), .D (new_AGEMA_signal_4688), .Q (new_AGEMA_signal_14681) ) ;
    buf_clk new_AGEMA_reg_buffer_8833 ( .C (clk), .D (RoundKey[58]), .Q (new_AGEMA_signal_14685) ) ;
    buf_clk new_AGEMA_reg_buffer_8837 ( .C (clk), .D (new_AGEMA_signal_4793), .Q (new_AGEMA_signal_14689) ) ;
    buf_clk new_AGEMA_reg_buffer_8841 ( .C (clk), .D (RoundKey[90]), .Q (new_AGEMA_signal_14693) ) ;
    buf_clk new_AGEMA_reg_buffer_8845 ( .C (clk), .D (new_AGEMA_signal_4901), .Q (new_AGEMA_signal_14697) ) ;
    buf_clk new_AGEMA_reg_buffer_8849 ( .C (clk), .D (RoundKey[25]), .Q (new_AGEMA_signal_14701) ) ;
    buf_clk new_AGEMA_reg_buffer_8853 ( .C (clk), .D (new_AGEMA_signal_4685), .Q (new_AGEMA_signal_14705) ) ;
    buf_clk new_AGEMA_reg_buffer_8857 ( .C (clk), .D (RoundKey[57]), .Q (new_AGEMA_signal_14709) ) ;
    buf_clk new_AGEMA_reg_buffer_8861 ( .C (clk), .D (new_AGEMA_signal_4790), .Q (new_AGEMA_signal_14713) ) ;
    buf_clk new_AGEMA_reg_buffer_8865 ( .C (clk), .D (RoundKey[89]), .Q (new_AGEMA_signal_14717) ) ;
    buf_clk new_AGEMA_reg_buffer_8869 ( .C (clk), .D (new_AGEMA_signal_4895), .Q (new_AGEMA_signal_14721) ) ;
    buf_clk new_AGEMA_reg_buffer_8873 ( .C (clk), .D (RoundKey[24]), .Q (new_AGEMA_signal_14725) ) ;
    buf_clk new_AGEMA_reg_buffer_8877 ( .C (clk), .D (new_AGEMA_signal_4682), .Q (new_AGEMA_signal_14729) ) ;
    buf_clk new_AGEMA_reg_buffer_8881 ( .C (clk), .D (RoundKey[56]), .Q (new_AGEMA_signal_14733) ) ;
    buf_clk new_AGEMA_reg_buffer_8885 ( .C (clk), .D (new_AGEMA_signal_4787), .Q (new_AGEMA_signal_14737) ) ;
    buf_clk new_AGEMA_reg_buffer_8889 ( .C (clk), .D (RoundKey[88]), .Q (new_AGEMA_signal_14741) ) ;
    buf_clk new_AGEMA_reg_buffer_8893 ( .C (clk), .D (new_AGEMA_signal_4892), .Q (new_AGEMA_signal_14745) ) ;
    buf_clk new_AGEMA_reg_buffer_8897 ( .C (clk), .D (RoundKey[23]), .Q (new_AGEMA_signal_14749) ) ;
    buf_clk new_AGEMA_reg_buffer_8901 ( .C (clk), .D (new_AGEMA_signal_4679), .Q (new_AGEMA_signal_14753) ) ;
    buf_clk new_AGEMA_reg_buffer_8905 ( .C (clk), .D (RoundKey[55]), .Q (new_AGEMA_signal_14757) ) ;
    buf_clk new_AGEMA_reg_buffer_8909 ( .C (clk), .D (new_AGEMA_signal_4784), .Q (new_AGEMA_signal_14761) ) ;
    buf_clk new_AGEMA_reg_buffer_8913 ( .C (clk), .D (RoundKey[87]), .Q (new_AGEMA_signal_14765) ) ;
    buf_clk new_AGEMA_reg_buffer_8917 ( .C (clk), .D (new_AGEMA_signal_4889), .Q (new_AGEMA_signal_14769) ) ;
    buf_clk new_AGEMA_reg_buffer_8921 ( .C (clk), .D (RoundKey[22]), .Q (new_AGEMA_signal_14773) ) ;
    buf_clk new_AGEMA_reg_buffer_8925 ( .C (clk), .D (new_AGEMA_signal_4676), .Q (new_AGEMA_signal_14777) ) ;
    buf_clk new_AGEMA_reg_buffer_8929 ( .C (clk), .D (RoundKey[54]), .Q (new_AGEMA_signal_14781) ) ;
    buf_clk new_AGEMA_reg_buffer_8933 ( .C (clk), .D (new_AGEMA_signal_4781), .Q (new_AGEMA_signal_14785) ) ;
    buf_clk new_AGEMA_reg_buffer_8937 ( .C (clk), .D (RoundKey[86]), .Q (new_AGEMA_signal_14789) ) ;
    buf_clk new_AGEMA_reg_buffer_8941 ( .C (clk), .D (new_AGEMA_signal_4886), .Q (new_AGEMA_signal_14793) ) ;
    buf_clk new_AGEMA_reg_buffer_8945 ( .C (clk), .D (RoundKey[21]), .Q (new_AGEMA_signal_14797) ) ;
    buf_clk new_AGEMA_reg_buffer_8949 ( .C (clk), .D (new_AGEMA_signal_4673), .Q (new_AGEMA_signal_14801) ) ;
    buf_clk new_AGEMA_reg_buffer_8953 ( .C (clk), .D (RoundKey[53]), .Q (new_AGEMA_signal_14805) ) ;
    buf_clk new_AGEMA_reg_buffer_8957 ( .C (clk), .D (new_AGEMA_signal_4778), .Q (new_AGEMA_signal_14809) ) ;
    buf_clk new_AGEMA_reg_buffer_8961 ( .C (clk), .D (RoundKey[85]), .Q (new_AGEMA_signal_14813) ) ;
    buf_clk new_AGEMA_reg_buffer_8965 ( .C (clk), .D (new_AGEMA_signal_4883), .Q (new_AGEMA_signal_14817) ) ;
    buf_clk new_AGEMA_reg_buffer_8969 ( .C (clk), .D (RoundKey[20]), .Q (new_AGEMA_signal_14821) ) ;
    buf_clk new_AGEMA_reg_buffer_8973 ( .C (clk), .D (new_AGEMA_signal_4670), .Q (new_AGEMA_signal_14825) ) ;
    buf_clk new_AGEMA_reg_buffer_8977 ( .C (clk), .D (RoundKey[52]), .Q (new_AGEMA_signal_14829) ) ;
    buf_clk new_AGEMA_reg_buffer_8981 ( .C (clk), .D (new_AGEMA_signal_4775), .Q (new_AGEMA_signal_14833) ) ;
    buf_clk new_AGEMA_reg_buffer_8985 ( .C (clk), .D (RoundKey[84]), .Q (new_AGEMA_signal_14837) ) ;
    buf_clk new_AGEMA_reg_buffer_8989 ( .C (clk), .D (new_AGEMA_signal_4880), .Q (new_AGEMA_signal_14841) ) ;
    buf_clk new_AGEMA_reg_buffer_8993 ( .C (clk), .D (RoundKey[1]), .Q (new_AGEMA_signal_14845) ) ;
    buf_clk new_AGEMA_reg_buffer_8997 ( .C (clk), .D (new_AGEMA_signal_4667), .Q (new_AGEMA_signal_14849) ) ;
    buf_clk new_AGEMA_reg_buffer_9001 ( .C (clk), .D (RoundKey[33]), .Q (new_AGEMA_signal_14853) ) ;
    buf_clk new_AGEMA_reg_buffer_9005 ( .C (clk), .D (new_AGEMA_signal_4712), .Q (new_AGEMA_signal_14857) ) ;
    buf_clk new_AGEMA_reg_buffer_9009 ( .C (clk), .D (RoundKey[65]), .Q (new_AGEMA_signal_14861) ) ;
    buf_clk new_AGEMA_reg_buffer_9013 ( .C (clk), .D (new_AGEMA_signal_4817), .Q (new_AGEMA_signal_14865) ) ;
    buf_clk new_AGEMA_reg_buffer_9017 ( .C (clk), .D (RoundKey[97]), .Q (new_AGEMA_signal_14869) ) ;
    buf_clk new_AGEMA_reg_buffer_9021 ( .C (clk), .D (new_AGEMA_signal_4922), .Q (new_AGEMA_signal_14873) ) ;
    buf_clk new_AGEMA_reg_buffer_9025 ( .C (clk), .D (RoundKey[19]), .Q (new_AGEMA_signal_14877) ) ;
    buf_clk new_AGEMA_reg_buffer_9029 ( .C (clk), .D (new_AGEMA_signal_4664), .Q (new_AGEMA_signal_14881) ) ;
    buf_clk new_AGEMA_reg_buffer_9033 ( .C (clk), .D (RoundKey[51]), .Q (new_AGEMA_signal_14885) ) ;
    buf_clk new_AGEMA_reg_buffer_9037 ( .C (clk), .D (new_AGEMA_signal_4772), .Q (new_AGEMA_signal_14889) ) ;
    buf_clk new_AGEMA_reg_buffer_9041 ( .C (clk), .D (RoundKey[83]), .Q (new_AGEMA_signal_14893) ) ;
    buf_clk new_AGEMA_reg_buffer_9045 ( .C (clk), .D (new_AGEMA_signal_4877), .Q (new_AGEMA_signal_14897) ) ;
    buf_clk new_AGEMA_reg_buffer_9049 ( .C (clk), .D (RoundKey[18]), .Q (new_AGEMA_signal_14901) ) ;
    buf_clk new_AGEMA_reg_buffer_9053 ( .C (clk), .D (new_AGEMA_signal_4661), .Q (new_AGEMA_signal_14905) ) ;
    buf_clk new_AGEMA_reg_buffer_9057 ( .C (clk), .D (RoundKey[50]), .Q (new_AGEMA_signal_14909) ) ;
    buf_clk new_AGEMA_reg_buffer_9061 ( .C (clk), .D (new_AGEMA_signal_4769), .Q (new_AGEMA_signal_14913) ) ;
    buf_clk new_AGEMA_reg_buffer_9065 ( .C (clk), .D (RoundKey[82]), .Q (new_AGEMA_signal_14917) ) ;
    buf_clk new_AGEMA_reg_buffer_9069 ( .C (clk), .D (new_AGEMA_signal_4874), .Q (new_AGEMA_signal_14921) ) ;
    buf_clk new_AGEMA_reg_buffer_9073 ( .C (clk), .D (RoundKey[17]), .Q (new_AGEMA_signal_14925) ) ;
    buf_clk new_AGEMA_reg_buffer_9077 ( .C (clk), .D (new_AGEMA_signal_4658), .Q (new_AGEMA_signal_14929) ) ;
    buf_clk new_AGEMA_reg_buffer_9081 ( .C (clk), .D (RoundKey[49]), .Q (new_AGEMA_signal_14933) ) ;
    buf_clk new_AGEMA_reg_buffer_9085 ( .C (clk), .D (new_AGEMA_signal_4763), .Q (new_AGEMA_signal_14937) ) ;
    buf_clk new_AGEMA_reg_buffer_9089 ( .C (clk), .D (RoundKey[81]), .Q (new_AGEMA_signal_14941) ) ;
    buf_clk new_AGEMA_reg_buffer_9093 ( .C (clk), .D (new_AGEMA_signal_4871), .Q (new_AGEMA_signal_14945) ) ;
    buf_clk new_AGEMA_reg_buffer_9097 ( .C (clk), .D (RoundKey[16]), .Q (new_AGEMA_signal_14949) ) ;
    buf_clk new_AGEMA_reg_buffer_9101 ( .C (clk), .D (new_AGEMA_signal_4655), .Q (new_AGEMA_signal_14953) ) ;
    buf_clk new_AGEMA_reg_buffer_9105 ( .C (clk), .D (RoundKey[48]), .Q (new_AGEMA_signal_14957) ) ;
    buf_clk new_AGEMA_reg_buffer_9109 ( .C (clk), .D (new_AGEMA_signal_4760), .Q (new_AGEMA_signal_14961) ) ;
    buf_clk new_AGEMA_reg_buffer_9113 ( .C (clk), .D (RoundKey[80]), .Q (new_AGEMA_signal_14965) ) ;
    buf_clk new_AGEMA_reg_buffer_9117 ( .C (clk), .D (new_AGEMA_signal_4868), .Q (new_AGEMA_signal_14969) ) ;
    buf_clk new_AGEMA_reg_buffer_9121 ( .C (clk), .D (RoundKey[15]), .Q (new_AGEMA_signal_14973) ) ;
    buf_clk new_AGEMA_reg_buffer_9125 ( .C (clk), .D (new_AGEMA_signal_4652), .Q (new_AGEMA_signal_14977) ) ;
    buf_clk new_AGEMA_reg_buffer_9129 ( .C (clk), .D (RoundKey[47]), .Q (new_AGEMA_signal_14981) ) ;
    buf_clk new_AGEMA_reg_buffer_9133 ( .C (clk), .D (new_AGEMA_signal_4757), .Q (new_AGEMA_signal_14985) ) ;
    buf_clk new_AGEMA_reg_buffer_9137 ( .C (clk), .D (RoundKey[79]), .Q (new_AGEMA_signal_14989) ) ;
    buf_clk new_AGEMA_reg_buffer_9141 ( .C (clk), .D (new_AGEMA_signal_4862), .Q (new_AGEMA_signal_14993) ) ;
    buf_clk new_AGEMA_reg_buffer_9145 ( .C (clk), .D (RoundKey[14]), .Q (new_AGEMA_signal_14997) ) ;
    buf_clk new_AGEMA_reg_buffer_9149 ( .C (clk), .D (new_AGEMA_signal_4649), .Q (new_AGEMA_signal_15001) ) ;
    buf_clk new_AGEMA_reg_buffer_9153 ( .C (clk), .D (RoundKey[46]), .Q (new_AGEMA_signal_15005) ) ;
    buf_clk new_AGEMA_reg_buffer_9157 ( .C (clk), .D (new_AGEMA_signal_4754), .Q (new_AGEMA_signal_15009) ) ;
    buf_clk new_AGEMA_reg_buffer_9161 ( .C (clk), .D (RoundKey[78]), .Q (new_AGEMA_signal_15013) ) ;
    buf_clk new_AGEMA_reg_buffer_9165 ( .C (clk), .D (new_AGEMA_signal_4859), .Q (new_AGEMA_signal_15017) ) ;
    buf_clk new_AGEMA_reg_buffer_9169 ( .C (clk), .D (RoundKey[13]), .Q (new_AGEMA_signal_15021) ) ;
    buf_clk new_AGEMA_reg_buffer_9173 ( .C (clk), .D (new_AGEMA_signal_4646), .Q (new_AGEMA_signal_15025) ) ;
    buf_clk new_AGEMA_reg_buffer_9177 ( .C (clk), .D (RoundKey[45]), .Q (new_AGEMA_signal_15029) ) ;
    buf_clk new_AGEMA_reg_buffer_9181 ( .C (clk), .D (new_AGEMA_signal_4751), .Q (new_AGEMA_signal_15033) ) ;
    buf_clk new_AGEMA_reg_buffer_9185 ( .C (clk), .D (RoundKey[77]), .Q (new_AGEMA_signal_15037) ) ;
    buf_clk new_AGEMA_reg_buffer_9189 ( .C (clk), .D (new_AGEMA_signal_4856), .Q (new_AGEMA_signal_15041) ) ;
    buf_clk new_AGEMA_reg_buffer_9193 ( .C (clk), .D (RoundKey[12]), .Q (new_AGEMA_signal_15045) ) ;
    buf_clk new_AGEMA_reg_buffer_9197 ( .C (clk), .D (new_AGEMA_signal_4643), .Q (new_AGEMA_signal_15049) ) ;
    buf_clk new_AGEMA_reg_buffer_9201 ( .C (clk), .D (RoundKey[44]), .Q (new_AGEMA_signal_15053) ) ;
    buf_clk new_AGEMA_reg_buffer_9205 ( .C (clk), .D (new_AGEMA_signal_4748), .Q (new_AGEMA_signal_15057) ) ;
    buf_clk new_AGEMA_reg_buffer_9209 ( .C (clk), .D (RoundKey[76]), .Q (new_AGEMA_signal_15061) ) ;
    buf_clk new_AGEMA_reg_buffer_9213 ( .C (clk), .D (new_AGEMA_signal_4853), .Q (new_AGEMA_signal_15065) ) ;
    buf_clk new_AGEMA_reg_buffer_9217 ( .C (clk), .D (RoundKey[127]), .Q (new_AGEMA_signal_15069) ) ;
    buf_clk new_AGEMA_reg_buffer_9221 ( .C (clk), .D (new_AGEMA_signal_4640), .Q (new_AGEMA_signal_15073) ) ;
    buf_clk new_AGEMA_reg_buffer_9225 ( .C (clk), .D (RoundKey[126]), .Q (new_AGEMA_signal_15077) ) ;
    buf_clk new_AGEMA_reg_buffer_9229 ( .C (clk), .D (new_AGEMA_signal_4637), .Q (new_AGEMA_signal_15081) ) ;
    buf_clk new_AGEMA_reg_buffer_9233 ( .C (clk), .D (RoundKey[125]), .Q (new_AGEMA_signal_15085) ) ;
    buf_clk new_AGEMA_reg_buffer_9237 ( .C (clk), .D (new_AGEMA_signal_4634), .Q (new_AGEMA_signal_15089) ) ;
    buf_clk new_AGEMA_reg_buffer_9241 ( .C (clk), .D (RoundKey[124]), .Q (new_AGEMA_signal_15093) ) ;
    buf_clk new_AGEMA_reg_buffer_9245 ( .C (clk), .D (new_AGEMA_signal_4631), .Q (new_AGEMA_signal_15097) ) ;
    buf_clk new_AGEMA_reg_buffer_9249 ( .C (clk), .D (RoundKey[123]), .Q (new_AGEMA_signal_15101) ) ;
    buf_clk new_AGEMA_reg_buffer_9253 ( .C (clk), .D (new_AGEMA_signal_4628), .Q (new_AGEMA_signal_15105) ) ;
    buf_clk new_AGEMA_reg_buffer_9257 ( .C (clk), .D (RoundKey[122]), .Q (new_AGEMA_signal_15109) ) ;
    buf_clk new_AGEMA_reg_buffer_9261 ( .C (clk), .D (new_AGEMA_signal_4625), .Q (new_AGEMA_signal_15113) ) ;
    buf_clk new_AGEMA_reg_buffer_9265 ( .C (clk), .D (RoundKey[121]), .Q (new_AGEMA_signal_15117) ) ;
    buf_clk new_AGEMA_reg_buffer_9269 ( .C (clk), .D (new_AGEMA_signal_4622), .Q (new_AGEMA_signal_15121) ) ;
    buf_clk new_AGEMA_reg_buffer_9273 ( .C (clk), .D (RoundKey[120]), .Q (new_AGEMA_signal_15125) ) ;
    buf_clk new_AGEMA_reg_buffer_9277 ( .C (clk), .D (new_AGEMA_signal_4619), .Q (new_AGEMA_signal_15129) ) ;
    buf_clk new_AGEMA_reg_buffer_9281 ( .C (clk), .D (RoundKey[11]), .Q (new_AGEMA_signal_15133) ) ;
    buf_clk new_AGEMA_reg_buffer_9285 ( .C (clk), .D (new_AGEMA_signal_4616), .Q (new_AGEMA_signal_15137) ) ;
    buf_clk new_AGEMA_reg_buffer_9289 ( .C (clk), .D (RoundKey[43]), .Q (new_AGEMA_signal_15141) ) ;
    buf_clk new_AGEMA_reg_buffer_9293 ( .C (clk), .D (new_AGEMA_signal_4745), .Q (new_AGEMA_signal_15145) ) ;
    buf_clk new_AGEMA_reg_buffer_9297 ( .C (clk), .D (RoundKey[75]), .Q (new_AGEMA_signal_15149) ) ;
    buf_clk new_AGEMA_reg_buffer_9301 ( .C (clk), .D (new_AGEMA_signal_4850), .Q (new_AGEMA_signal_15153) ) ;
    buf_clk new_AGEMA_reg_buffer_9305 ( .C (clk), .D (RoundKey[119]), .Q (new_AGEMA_signal_15157) ) ;
    buf_clk new_AGEMA_reg_buffer_9309 ( .C (clk), .D (new_AGEMA_signal_4613), .Q (new_AGEMA_signal_15161) ) ;
    buf_clk new_AGEMA_reg_buffer_9313 ( .C (clk), .D (RoundKey[118]), .Q (new_AGEMA_signal_15165) ) ;
    buf_clk new_AGEMA_reg_buffer_9317 ( .C (clk), .D (new_AGEMA_signal_4610), .Q (new_AGEMA_signal_15169) ) ;
    buf_clk new_AGEMA_reg_buffer_9321 ( .C (clk), .D (RoundKey[117]), .Q (new_AGEMA_signal_15173) ) ;
    buf_clk new_AGEMA_reg_buffer_9325 ( .C (clk), .D (new_AGEMA_signal_4607), .Q (new_AGEMA_signal_15177) ) ;
    buf_clk new_AGEMA_reg_buffer_9329 ( .C (clk), .D (RoundKey[116]), .Q (new_AGEMA_signal_15181) ) ;
    buf_clk new_AGEMA_reg_buffer_9333 ( .C (clk), .D (new_AGEMA_signal_4604), .Q (new_AGEMA_signal_15185) ) ;
    buf_clk new_AGEMA_reg_buffer_9337 ( .C (clk), .D (RoundKey[115]), .Q (new_AGEMA_signal_15189) ) ;
    buf_clk new_AGEMA_reg_buffer_9341 ( .C (clk), .D (new_AGEMA_signal_4601), .Q (new_AGEMA_signal_15193) ) ;
    buf_clk new_AGEMA_reg_buffer_9345 ( .C (clk), .D (RoundKey[114]), .Q (new_AGEMA_signal_15197) ) ;
    buf_clk new_AGEMA_reg_buffer_9349 ( .C (clk), .D (new_AGEMA_signal_4598), .Q (new_AGEMA_signal_15201) ) ;
    buf_clk new_AGEMA_reg_buffer_9353 ( .C (clk), .D (RoundKey[113]), .Q (new_AGEMA_signal_15205) ) ;
    buf_clk new_AGEMA_reg_buffer_9357 ( .C (clk), .D (new_AGEMA_signal_4595), .Q (new_AGEMA_signal_15209) ) ;
    buf_clk new_AGEMA_reg_buffer_9361 ( .C (clk), .D (RoundKey[112]), .Q (new_AGEMA_signal_15213) ) ;
    buf_clk new_AGEMA_reg_buffer_9365 ( .C (clk), .D (new_AGEMA_signal_4592), .Q (new_AGEMA_signal_15217) ) ;
    buf_clk new_AGEMA_reg_buffer_9369 ( .C (clk), .D (RoundKey[111]), .Q (new_AGEMA_signal_15221) ) ;
    buf_clk new_AGEMA_reg_buffer_9373 ( .C (clk), .D (new_AGEMA_signal_4589), .Q (new_AGEMA_signal_15225) ) ;
    buf_clk new_AGEMA_reg_buffer_9377 ( .C (clk), .D (RoundKey[110]), .Q (new_AGEMA_signal_15229) ) ;
    buf_clk new_AGEMA_reg_buffer_9381 ( .C (clk), .D (new_AGEMA_signal_4586), .Q (new_AGEMA_signal_15233) ) ;
    buf_clk new_AGEMA_reg_buffer_9385 ( .C (clk), .D (RoundKey[10]), .Q (new_AGEMA_signal_15237) ) ;
    buf_clk new_AGEMA_reg_buffer_9389 ( .C (clk), .D (new_AGEMA_signal_4583), .Q (new_AGEMA_signal_15241) ) ;
    buf_clk new_AGEMA_reg_buffer_9393 ( .C (clk), .D (RoundKey[42]), .Q (new_AGEMA_signal_15245) ) ;
    buf_clk new_AGEMA_reg_buffer_9397 ( .C (clk), .D (new_AGEMA_signal_4742), .Q (new_AGEMA_signal_15249) ) ;
    buf_clk new_AGEMA_reg_buffer_9401 ( .C (clk), .D (RoundKey[74]), .Q (new_AGEMA_signal_15253) ) ;
    buf_clk new_AGEMA_reg_buffer_9405 ( .C (clk), .D (new_AGEMA_signal_4847), .Q (new_AGEMA_signal_15257) ) ;
    buf_clk new_AGEMA_reg_buffer_9409 ( .C (clk), .D (RoundKey[109]), .Q (new_AGEMA_signal_15261) ) ;
    buf_clk new_AGEMA_reg_buffer_9413 ( .C (clk), .D (new_AGEMA_signal_4580), .Q (new_AGEMA_signal_15265) ) ;
    buf_clk new_AGEMA_reg_buffer_9417 ( .C (clk), .D (RoundKey[108]), .Q (new_AGEMA_signal_15269) ) ;
    buf_clk new_AGEMA_reg_buffer_9421 ( .C (clk), .D (new_AGEMA_signal_4577), .Q (new_AGEMA_signal_15273) ) ;
    buf_clk new_AGEMA_reg_buffer_9425 ( .C (clk), .D (RoundKey[107]), .Q (new_AGEMA_signal_15277) ) ;
    buf_clk new_AGEMA_reg_buffer_9429 ( .C (clk), .D (new_AGEMA_signal_4574), .Q (new_AGEMA_signal_15281) ) ;
    buf_clk new_AGEMA_reg_buffer_9433 ( .C (clk), .D (RoundKey[106]), .Q (new_AGEMA_signal_15285) ) ;
    buf_clk new_AGEMA_reg_buffer_9437 ( .C (clk), .D (new_AGEMA_signal_4571), .Q (new_AGEMA_signal_15289) ) ;
    buf_clk new_AGEMA_reg_buffer_9441 ( .C (clk), .D (RoundKey[105]), .Q (new_AGEMA_signal_15293) ) ;
    buf_clk new_AGEMA_reg_buffer_9445 ( .C (clk), .D (new_AGEMA_signal_4568), .Q (new_AGEMA_signal_15297) ) ;
    buf_clk new_AGEMA_reg_buffer_9449 ( .C (clk), .D (RoundKey[104]), .Q (new_AGEMA_signal_15301) ) ;
    buf_clk new_AGEMA_reg_buffer_9453 ( .C (clk), .D (new_AGEMA_signal_4565), .Q (new_AGEMA_signal_15305) ) ;
    buf_clk new_AGEMA_reg_buffer_9457 ( .C (clk), .D (RoundKey[103]), .Q (new_AGEMA_signal_15309) ) ;
    buf_clk new_AGEMA_reg_buffer_9461 ( .C (clk), .D (new_AGEMA_signal_4562), .Q (new_AGEMA_signal_15313) ) ;
    buf_clk new_AGEMA_reg_buffer_9465 ( .C (clk), .D (RoundKey[102]), .Q (new_AGEMA_signal_15317) ) ;
    buf_clk new_AGEMA_reg_buffer_9469 ( .C (clk), .D (new_AGEMA_signal_4559), .Q (new_AGEMA_signal_15321) ) ;
    buf_clk new_AGEMA_reg_buffer_9473 ( .C (clk), .D (RoundKey[101]), .Q (new_AGEMA_signal_15325) ) ;
    buf_clk new_AGEMA_reg_buffer_9477 ( .C (clk), .D (new_AGEMA_signal_4556), .Q (new_AGEMA_signal_15329) ) ;
    buf_clk new_AGEMA_reg_buffer_9481 ( .C (clk), .D (RoundKey[100]), .Q (new_AGEMA_signal_15333) ) ;
    buf_clk new_AGEMA_reg_buffer_9485 ( .C (clk), .D (new_AGEMA_signal_4553), .Q (new_AGEMA_signal_15337) ) ;
    buf_clk new_AGEMA_reg_buffer_9489 ( .C (clk), .D (RoundKey[0]), .Q (new_AGEMA_signal_15341) ) ;
    buf_clk new_AGEMA_reg_buffer_9493 ( .C (clk), .D (new_AGEMA_signal_4550), .Q (new_AGEMA_signal_15345) ) ;
    buf_clk new_AGEMA_reg_buffer_9497 ( .C (clk), .D (RoundKey[32]), .Q (new_AGEMA_signal_15349) ) ;
    buf_clk new_AGEMA_reg_buffer_9501 ( .C (clk), .D (new_AGEMA_signal_4709), .Q (new_AGEMA_signal_15353) ) ;
    buf_clk new_AGEMA_reg_buffer_9505 ( .C (clk), .D (RoundKey[64]), .Q (new_AGEMA_signal_15357) ) ;
    buf_clk new_AGEMA_reg_buffer_9509 ( .C (clk), .D (new_AGEMA_signal_4814), .Q (new_AGEMA_signal_15361) ) ;
    buf_clk new_AGEMA_reg_buffer_9513 ( .C (clk), .D (RoundKey[96]), .Q (new_AGEMA_signal_15365) ) ;
    buf_clk new_AGEMA_reg_buffer_9517 ( .C (clk), .D (new_AGEMA_signal_4919), .Q (new_AGEMA_signal_15369) ) ;
    buf_clk new_AGEMA_reg_buffer_9521 ( .C (clk), .D (n283), .Q (new_AGEMA_signal_15373) ) ;
    buf_clk new_AGEMA_reg_buffer_9525 ( .C (clk), .D (n285), .Q (new_AGEMA_signal_15377) ) ;
    buf_clk new_AGEMA_reg_buffer_9529 ( .C (clk), .D (Rcon[5]), .Q (new_AGEMA_signal_15381) ) ;
    buf_clk new_AGEMA_reg_buffer_9533 ( .C (clk), .D (Rcon[4]), .Q (new_AGEMA_signal_15385) ) ;
    buf_clk new_AGEMA_reg_buffer_9537 ( .C (clk), .D (Rcon[3]), .Q (new_AGEMA_signal_15389) ) ;
    buf_clk new_AGEMA_reg_buffer_9541 ( .C (clk), .D (Rcon[2]), .Q (new_AGEMA_signal_15393) ) ;
    buf_clk new_AGEMA_reg_buffer_9545 ( .C (clk), .D (Rcon[1]), .Q (new_AGEMA_signal_15397) ) ;
    buf_clk new_AGEMA_reg_buffer_9549 ( .C (clk), .D (Rcon[0]), .Q (new_AGEMA_signal_15401) ) ;
    buf_clk new_AGEMA_reg_buffer_9553 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6), .Q (new_AGEMA_signal_15405) ) ;
    buf_clk new_AGEMA_reg_buffer_9556 ( .C (clk), .D (new_AGEMA_signal_5133), .Q (new_AGEMA_signal_15408) ) ;
    buf_clk new_AGEMA_reg_buffer_9559 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8), .Q (new_AGEMA_signal_15411) ) ;
    buf_clk new_AGEMA_reg_buffer_9562 ( .C (clk), .D (new_AGEMA_signal_5293), .Q (new_AGEMA_signal_15414) ) ;
    buf_clk new_AGEMA_reg_buffer_9565 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16), .Q (new_AGEMA_signal_15417) ) ;
    buf_clk new_AGEMA_reg_buffer_9568 ( .C (clk), .D (new_AGEMA_signal_5137), .Q (new_AGEMA_signal_15420) ) ;
    buf_clk new_AGEMA_reg_buffer_9571 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9), .Q (new_AGEMA_signal_15423) ) ;
    buf_clk new_AGEMA_reg_buffer_9574 ( .C (clk), .D (new_AGEMA_signal_5134), .Q (new_AGEMA_signal_15426) ) ;
    buf_clk new_AGEMA_reg_buffer_9577 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17), .Q (new_AGEMA_signal_15429) ) ;
    buf_clk new_AGEMA_reg_buffer_9580 ( .C (clk), .D (new_AGEMA_signal_5296), .Q (new_AGEMA_signal_15432) ) ;
    buf_clk new_AGEMA_reg_buffer_9583 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15), .Q (new_AGEMA_signal_15435) ) ;
    buf_clk new_AGEMA_reg_buffer_9586 ( .C (clk), .D (new_AGEMA_signal_5136), .Q (new_AGEMA_signal_15438) ) ;
    buf_clk new_AGEMA_reg_buffer_9589 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27), .Q (new_AGEMA_signal_15441) ) ;
    buf_clk new_AGEMA_reg_buffer_9592 ( .C (clk), .D (new_AGEMA_signal_5140), .Q (new_AGEMA_signal_15444) ) ;
    buf_clk new_AGEMA_reg_buffer_9595 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10), .Q (new_AGEMA_signal_15447) ) ;
    buf_clk new_AGEMA_reg_buffer_9598 ( .C (clk), .D (new_AGEMA_signal_5294), .Q (new_AGEMA_signal_15450) ) ;
    buf_clk new_AGEMA_reg_buffer_9601 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13), .Q (new_AGEMA_signal_15453) ) ;
    buf_clk new_AGEMA_reg_buffer_9604 ( .C (clk), .D (new_AGEMA_signal_5135), .Q (new_AGEMA_signal_15456) ) ;
    buf_clk new_AGEMA_reg_buffer_9607 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23), .Q (new_AGEMA_signal_15459) ) ;
    buf_clk new_AGEMA_reg_buffer_9610 ( .C (clk), .D (new_AGEMA_signal_5298), .Q (new_AGEMA_signal_15462) ) ;
    buf_clk new_AGEMA_reg_buffer_9613 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19), .Q (new_AGEMA_signal_15465) ) ;
    buf_clk new_AGEMA_reg_buffer_9616 ( .C (clk), .D (new_AGEMA_signal_5138), .Q (new_AGEMA_signal_15468) ) ;
    buf_clk new_AGEMA_reg_buffer_9619 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3), .Q (new_AGEMA_signal_15471) ) ;
    buf_clk new_AGEMA_reg_buffer_9622 ( .C (clk), .D (new_AGEMA_signal_4935), .Q (new_AGEMA_signal_15474) ) ;
    buf_clk new_AGEMA_reg_buffer_9625 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22), .Q (new_AGEMA_signal_15477) ) ;
    buf_clk new_AGEMA_reg_buffer_9628 ( .C (clk), .D (new_AGEMA_signal_5139), .Q (new_AGEMA_signal_15480) ) ;
    buf_clk new_AGEMA_reg_buffer_9631 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20), .Q (new_AGEMA_signal_15483) ) ;
    buf_clk new_AGEMA_reg_buffer_9634 ( .C (clk), .D (new_AGEMA_signal_5297), .Q (new_AGEMA_signal_15486) ) ;
    buf_clk new_AGEMA_reg_buffer_9637 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1), .Q (new_AGEMA_signal_15489) ) ;
    buf_clk new_AGEMA_reg_buffer_9640 ( .C (clk), .D (new_AGEMA_signal_4933), .Q (new_AGEMA_signal_15492) ) ;
    buf_clk new_AGEMA_reg_buffer_9643 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4), .Q (new_AGEMA_signal_15495) ) ;
    buf_clk new_AGEMA_reg_buffer_9646 ( .C (clk), .D (new_AGEMA_signal_4936), .Q (new_AGEMA_signal_15498) ) ;
    buf_clk new_AGEMA_reg_buffer_9649 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2), .Q (new_AGEMA_signal_15501) ) ;
    buf_clk new_AGEMA_reg_buffer_9652 ( .C (clk), .D (new_AGEMA_signal_4934), .Q (new_AGEMA_signal_15504) ) ;
    buf_clk new_AGEMA_reg_buffer_9655 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6), .Q (new_AGEMA_signal_15507) ) ;
    buf_clk new_AGEMA_reg_buffer_9658 ( .C (clk), .D (new_AGEMA_signal_5141), .Q (new_AGEMA_signal_15510) ) ;
    buf_clk new_AGEMA_reg_buffer_9661 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8), .Q (new_AGEMA_signal_15513) ) ;
    buf_clk new_AGEMA_reg_buffer_9664 ( .C (clk), .D (new_AGEMA_signal_5306), .Q (new_AGEMA_signal_15516) ) ;
    buf_clk new_AGEMA_reg_buffer_9667 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16), .Q (new_AGEMA_signal_15519) ) ;
    buf_clk new_AGEMA_reg_buffer_9670 ( .C (clk), .D (new_AGEMA_signal_5145), .Q (new_AGEMA_signal_15522) ) ;
    buf_clk new_AGEMA_reg_buffer_9673 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9), .Q (new_AGEMA_signal_15525) ) ;
    buf_clk new_AGEMA_reg_buffer_9676 ( .C (clk), .D (new_AGEMA_signal_5142), .Q (new_AGEMA_signal_15528) ) ;
    buf_clk new_AGEMA_reg_buffer_9679 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17), .Q (new_AGEMA_signal_15531) ) ;
    buf_clk new_AGEMA_reg_buffer_9682 ( .C (clk), .D (new_AGEMA_signal_5309), .Q (new_AGEMA_signal_15534) ) ;
    buf_clk new_AGEMA_reg_buffer_9685 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15), .Q (new_AGEMA_signal_15537) ) ;
    buf_clk new_AGEMA_reg_buffer_9688 ( .C (clk), .D (new_AGEMA_signal_5144), .Q (new_AGEMA_signal_15540) ) ;
    buf_clk new_AGEMA_reg_buffer_9691 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27), .Q (new_AGEMA_signal_15543) ) ;
    buf_clk new_AGEMA_reg_buffer_9694 ( .C (clk), .D (new_AGEMA_signal_5148), .Q (new_AGEMA_signal_15546) ) ;
    buf_clk new_AGEMA_reg_buffer_9697 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10), .Q (new_AGEMA_signal_15549) ) ;
    buf_clk new_AGEMA_reg_buffer_9700 ( .C (clk), .D (new_AGEMA_signal_5307), .Q (new_AGEMA_signal_15552) ) ;
    buf_clk new_AGEMA_reg_buffer_9703 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13), .Q (new_AGEMA_signal_15555) ) ;
    buf_clk new_AGEMA_reg_buffer_9706 ( .C (clk), .D (new_AGEMA_signal_5143), .Q (new_AGEMA_signal_15558) ) ;
    buf_clk new_AGEMA_reg_buffer_9709 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23), .Q (new_AGEMA_signal_15561) ) ;
    buf_clk new_AGEMA_reg_buffer_9712 ( .C (clk), .D (new_AGEMA_signal_5311), .Q (new_AGEMA_signal_15564) ) ;
    buf_clk new_AGEMA_reg_buffer_9715 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19), .Q (new_AGEMA_signal_15567) ) ;
    buf_clk new_AGEMA_reg_buffer_9718 ( .C (clk), .D (new_AGEMA_signal_5146), .Q (new_AGEMA_signal_15570) ) ;
    buf_clk new_AGEMA_reg_buffer_9721 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3), .Q (new_AGEMA_signal_15573) ) ;
    buf_clk new_AGEMA_reg_buffer_9724 ( .C (clk), .D (new_AGEMA_signal_4945), .Q (new_AGEMA_signal_15576) ) ;
    buf_clk new_AGEMA_reg_buffer_9727 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22), .Q (new_AGEMA_signal_15579) ) ;
    buf_clk new_AGEMA_reg_buffer_9730 ( .C (clk), .D (new_AGEMA_signal_5147), .Q (new_AGEMA_signal_15582) ) ;
    buf_clk new_AGEMA_reg_buffer_9733 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20), .Q (new_AGEMA_signal_15585) ) ;
    buf_clk new_AGEMA_reg_buffer_9736 ( .C (clk), .D (new_AGEMA_signal_5310), .Q (new_AGEMA_signal_15588) ) ;
    buf_clk new_AGEMA_reg_buffer_9739 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1), .Q (new_AGEMA_signal_15591) ) ;
    buf_clk new_AGEMA_reg_buffer_9742 ( .C (clk), .D (new_AGEMA_signal_4943), .Q (new_AGEMA_signal_15594) ) ;
    buf_clk new_AGEMA_reg_buffer_9745 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4), .Q (new_AGEMA_signal_15597) ) ;
    buf_clk new_AGEMA_reg_buffer_9748 ( .C (clk), .D (new_AGEMA_signal_4946), .Q (new_AGEMA_signal_15600) ) ;
    buf_clk new_AGEMA_reg_buffer_9751 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2), .Q (new_AGEMA_signal_15603) ) ;
    buf_clk new_AGEMA_reg_buffer_9754 ( .C (clk), .D (new_AGEMA_signal_4944), .Q (new_AGEMA_signal_15606) ) ;
    buf_clk new_AGEMA_reg_buffer_9757 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6), .Q (new_AGEMA_signal_15609) ) ;
    buf_clk new_AGEMA_reg_buffer_9760 ( .C (clk), .D (new_AGEMA_signal_5149), .Q (new_AGEMA_signal_15612) ) ;
    buf_clk new_AGEMA_reg_buffer_9763 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8), .Q (new_AGEMA_signal_15615) ) ;
    buf_clk new_AGEMA_reg_buffer_9766 ( .C (clk), .D (new_AGEMA_signal_5319), .Q (new_AGEMA_signal_15618) ) ;
    buf_clk new_AGEMA_reg_buffer_9769 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16), .Q (new_AGEMA_signal_15621) ) ;
    buf_clk new_AGEMA_reg_buffer_9772 ( .C (clk), .D (new_AGEMA_signal_5153), .Q (new_AGEMA_signal_15624) ) ;
    buf_clk new_AGEMA_reg_buffer_9775 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9), .Q (new_AGEMA_signal_15627) ) ;
    buf_clk new_AGEMA_reg_buffer_9778 ( .C (clk), .D (new_AGEMA_signal_5150), .Q (new_AGEMA_signal_15630) ) ;
    buf_clk new_AGEMA_reg_buffer_9781 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17), .Q (new_AGEMA_signal_15633) ) ;
    buf_clk new_AGEMA_reg_buffer_9784 ( .C (clk), .D (new_AGEMA_signal_5322), .Q (new_AGEMA_signal_15636) ) ;
    buf_clk new_AGEMA_reg_buffer_9787 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15), .Q (new_AGEMA_signal_15639) ) ;
    buf_clk new_AGEMA_reg_buffer_9790 ( .C (clk), .D (new_AGEMA_signal_5152), .Q (new_AGEMA_signal_15642) ) ;
    buf_clk new_AGEMA_reg_buffer_9793 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27), .Q (new_AGEMA_signal_15645) ) ;
    buf_clk new_AGEMA_reg_buffer_9796 ( .C (clk), .D (new_AGEMA_signal_5156), .Q (new_AGEMA_signal_15648) ) ;
    buf_clk new_AGEMA_reg_buffer_9799 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10), .Q (new_AGEMA_signal_15651) ) ;
    buf_clk new_AGEMA_reg_buffer_9802 ( .C (clk), .D (new_AGEMA_signal_5320), .Q (new_AGEMA_signal_15654) ) ;
    buf_clk new_AGEMA_reg_buffer_9805 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13), .Q (new_AGEMA_signal_15657) ) ;
    buf_clk new_AGEMA_reg_buffer_9808 ( .C (clk), .D (new_AGEMA_signal_5151), .Q (new_AGEMA_signal_15660) ) ;
    buf_clk new_AGEMA_reg_buffer_9811 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23), .Q (new_AGEMA_signal_15663) ) ;
    buf_clk new_AGEMA_reg_buffer_9814 ( .C (clk), .D (new_AGEMA_signal_5324), .Q (new_AGEMA_signal_15666) ) ;
    buf_clk new_AGEMA_reg_buffer_9817 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19), .Q (new_AGEMA_signal_15669) ) ;
    buf_clk new_AGEMA_reg_buffer_9820 ( .C (clk), .D (new_AGEMA_signal_5154), .Q (new_AGEMA_signal_15672) ) ;
    buf_clk new_AGEMA_reg_buffer_9823 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3), .Q (new_AGEMA_signal_15675) ) ;
    buf_clk new_AGEMA_reg_buffer_9826 ( .C (clk), .D (new_AGEMA_signal_4955), .Q (new_AGEMA_signal_15678) ) ;
    buf_clk new_AGEMA_reg_buffer_9829 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22), .Q (new_AGEMA_signal_15681) ) ;
    buf_clk new_AGEMA_reg_buffer_9832 ( .C (clk), .D (new_AGEMA_signal_5155), .Q (new_AGEMA_signal_15684) ) ;
    buf_clk new_AGEMA_reg_buffer_9835 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20), .Q (new_AGEMA_signal_15687) ) ;
    buf_clk new_AGEMA_reg_buffer_9838 ( .C (clk), .D (new_AGEMA_signal_5323), .Q (new_AGEMA_signal_15690) ) ;
    buf_clk new_AGEMA_reg_buffer_9841 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1), .Q (new_AGEMA_signal_15693) ) ;
    buf_clk new_AGEMA_reg_buffer_9844 ( .C (clk), .D (new_AGEMA_signal_4953), .Q (new_AGEMA_signal_15696) ) ;
    buf_clk new_AGEMA_reg_buffer_9847 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4), .Q (new_AGEMA_signal_15699) ) ;
    buf_clk new_AGEMA_reg_buffer_9850 ( .C (clk), .D (new_AGEMA_signal_4956), .Q (new_AGEMA_signal_15702) ) ;
    buf_clk new_AGEMA_reg_buffer_9853 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2), .Q (new_AGEMA_signal_15705) ) ;
    buf_clk new_AGEMA_reg_buffer_9856 ( .C (clk), .D (new_AGEMA_signal_4954), .Q (new_AGEMA_signal_15708) ) ;
    buf_clk new_AGEMA_reg_buffer_9859 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6), .Q (new_AGEMA_signal_15711) ) ;
    buf_clk new_AGEMA_reg_buffer_9862 ( .C (clk), .D (new_AGEMA_signal_5157), .Q (new_AGEMA_signal_15714) ) ;
    buf_clk new_AGEMA_reg_buffer_9865 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8), .Q (new_AGEMA_signal_15717) ) ;
    buf_clk new_AGEMA_reg_buffer_9868 ( .C (clk), .D (new_AGEMA_signal_5332), .Q (new_AGEMA_signal_15720) ) ;
    buf_clk new_AGEMA_reg_buffer_9871 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16), .Q (new_AGEMA_signal_15723) ) ;
    buf_clk new_AGEMA_reg_buffer_9874 ( .C (clk), .D (new_AGEMA_signal_5161), .Q (new_AGEMA_signal_15726) ) ;
    buf_clk new_AGEMA_reg_buffer_9877 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9), .Q (new_AGEMA_signal_15729) ) ;
    buf_clk new_AGEMA_reg_buffer_9880 ( .C (clk), .D (new_AGEMA_signal_5158), .Q (new_AGEMA_signal_15732) ) ;
    buf_clk new_AGEMA_reg_buffer_9883 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17), .Q (new_AGEMA_signal_15735) ) ;
    buf_clk new_AGEMA_reg_buffer_9886 ( .C (clk), .D (new_AGEMA_signal_5335), .Q (new_AGEMA_signal_15738) ) ;
    buf_clk new_AGEMA_reg_buffer_9889 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15), .Q (new_AGEMA_signal_15741) ) ;
    buf_clk new_AGEMA_reg_buffer_9892 ( .C (clk), .D (new_AGEMA_signal_5160), .Q (new_AGEMA_signal_15744) ) ;
    buf_clk new_AGEMA_reg_buffer_9895 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27), .Q (new_AGEMA_signal_15747) ) ;
    buf_clk new_AGEMA_reg_buffer_9898 ( .C (clk), .D (new_AGEMA_signal_5164), .Q (new_AGEMA_signal_15750) ) ;
    buf_clk new_AGEMA_reg_buffer_9901 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10), .Q (new_AGEMA_signal_15753) ) ;
    buf_clk new_AGEMA_reg_buffer_9904 ( .C (clk), .D (new_AGEMA_signal_5333), .Q (new_AGEMA_signal_15756) ) ;
    buf_clk new_AGEMA_reg_buffer_9907 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13), .Q (new_AGEMA_signal_15759) ) ;
    buf_clk new_AGEMA_reg_buffer_9910 ( .C (clk), .D (new_AGEMA_signal_5159), .Q (new_AGEMA_signal_15762) ) ;
    buf_clk new_AGEMA_reg_buffer_9913 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23), .Q (new_AGEMA_signal_15765) ) ;
    buf_clk new_AGEMA_reg_buffer_9916 ( .C (clk), .D (new_AGEMA_signal_5337), .Q (new_AGEMA_signal_15768) ) ;
    buf_clk new_AGEMA_reg_buffer_9919 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19), .Q (new_AGEMA_signal_15771) ) ;
    buf_clk new_AGEMA_reg_buffer_9922 ( .C (clk), .D (new_AGEMA_signal_5162), .Q (new_AGEMA_signal_15774) ) ;
    buf_clk new_AGEMA_reg_buffer_9925 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3), .Q (new_AGEMA_signal_15777) ) ;
    buf_clk new_AGEMA_reg_buffer_9928 ( .C (clk), .D (new_AGEMA_signal_4965), .Q (new_AGEMA_signal_15780) ) ;
    buf_clk new_AGEMA_reg_buffer_9931 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22), .Q (new_AGEMA_signal_15783) ) ;
    buf_clk new_AGEMA_reg_buffer_9934 ( .C (clk), .D (new_AGEMA_signal_5163), .Q (new_AGEMA_signal_15786) ) ;
    buf_clk new_AGEMA_reg_buffer_9937 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20), .Q (new_AGEMA_signal_15789) ) ;
    buf_clk new_AGEMA_reg_buffer_9940 ( .C (clk), .D (new_AGEMA_signal_5336), .Q (new_AGEMA_signal_15792) ) ;
    buf_clk new_AGEMA_reg_buffer_9943 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1), .Q (new_AGEMA_signal_15795) ) ;
    buf_clk new_AGEMA_reg_buffer_9946 ( .C (clk), .D (new_AGEMA_signal_4963), .Q (new_AGEMA_signal_15798) ) ;
    buf_clk new_AGEMA_reg_buffer_9949 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4), .Q (new_AGEMA_signal_15801) ) ;
    buf_clk new_AGEMA_reg_buffer_9952 ( .C (clk), .D (new_AGEMA_signal_4966), .Q (new_AGEMA_signal_15804) ) ;
    buf_clk new_AGEMA_reg_buffer_9955 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2), .Q (new_AGEMA_signal_15807) ) ;
    buf_clk new_AGEMA_reg_buffer_9958 ( .C (clk), .D (new_AGEMA_signal_4964), .Q (new_AGEMA_signal_15810) ) ;
    buf_clk new_AGEMA_reg_buffer_9961 ( .C (clk), .D (RoundCounterIns_N7), .Q (new_AGEMA_signal_15813) ) ;
    buf_clk new_AGEMA_reg_buffer_9965 ( .C (clk), .D (RoundCounterIns_N8), .Q (new_AGEMA_signal_15817) ) ;
    buf_clk new_AGEMA_reg_buffer_9969 ( .C (clk), .D (RoundCounterIns_n1), .Q (new_AGEMA_signal_15821) ) ;
    buf_clk new_AGEMA_reg_buffer_9973 ( .C (clk), .D (RoundCounterIns_N10), .Q (new_AGEMA_signal_15825) ) ;

    /* cells in depth 2 */
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M25_U1 ( .a ({new_AGEMA_signal_5852, SubBytesIns_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_5850, SubBytesIns_Inst_Sbox_0_M20}), .clk (clk), .r ({Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_5930, SubBytesIns_Inst_Sbox_0_M25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M26_U1 ( .a ({new_AGEMA_signal_10222, new_AGEMA_signal_10221}), .b ({new_AGEMA_signal_5930, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_6014, SubBytesIns_Inst_Sbox_0_M26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M28_U1 ( .a ({new_AGEMA_signal_10224, new_AGEMA_signal_10223}), .b ({new_AGEMA_signal_5930, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_6015, SubBytesIns_Inst_Sbox_0_M28}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M31_U1 ( .a ({new_AGEMA_signal_5850, SubBytesIns_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_5929, SubBytesIns_Inst_Sbox_0_M23}), .clk (clk), .r ({Fresh[363], Fresh[362]}), .c ({new_AGEMA_signal_6016, SubBytesIns_Inst_Sbox_0_M31}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M33_U1 ( .a ({new_AGEMA_signal_10226, new_AGEMA_signal_10225}), .b ({new_AGEMA_signal_5930, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_6017, SubBytesIns_Inst_Sbox_0_M33}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M34_U1 ( .a ({new_AGEMA_signal_5851, SubBytesIns_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_5852, SubBytesIns_Inst_Sbox_0_M22}), .clk (clk), .r ({Fresh[365], Fresh[364]}), .c ({new_AGEMA_signal_5932, SubBytesIns_Inst_Sbox_0_M34}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M36_U1 ( .a ({new_AGEMA_signal_10228, new_AGEMA_signal_10227}), .b ({new_AGEMA_signal_5930, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_6117, SubBytesIns_Inst_Sbox_0_M36}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M25_U1 ( .a ({new_AGEMA_signal_5856, SubBytesIns_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_5854, SubBytesIns_Inst_Sbox_1_M20}), .clk (clk), .r ({Fresh[367], Fresh[366]}), .c ({new_AGEMA_signal_5934, SubBytesIns_Inst_Sbox_1_M25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M26_U1 ( .a ({new_AGEMA_signal_10230, new_AGEMA_signal_10229}), .b ({new_AGEMA_signal_5934, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_6019, SubBytesIns_Inst_Sbox_1_M26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M28_U1 ( .a ({new_AGEMA_signal_10232, new_AGEMA_signal_10231}), .b ({new_AGEMA_signal_5934, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_6020, SubBytesIns_Inst_Sbox_1_M28}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M31_U1 ( .a ({new_AGEMA_signal_5854, SubBytesIns_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_5933, SubBytesIns_Inst_Sbox_1_M23}), .clk (clk), .r ({Fresh[369], Fresh[368]}), .c ({new_AGEMA_signal_6021, SubBytesIns_Inst_Sbox_1_M31}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M33_U1 ( .a ({new_AGEMA_signal_10234, new_AGEMA_signal_10233}), .b ({new_AGEMA_signal_5934, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_6022, SubBytesIns_Inst_Sbox_1_M33}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M34_U1 ( .a ({new_AGEMA_signal_5855, SubBytesIns_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_5856, SubBytesIns_Inst_Sbox_1_M22}), .clk (clk), .r ({Fresh[371], Fresh[370]}), .c ({new_AGEMA_signal_5936, SubBytesIns_Inst_Sbox_1_M34}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M36_U1 ( .a ({new_AGEMA_signal_10236, new_AGEMA_signal_10235}), .b ({new_AGEMA_signal_5934, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_6122, SubBytesIns_Inst_Sbox_1_M36}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M25_U1 ( .a ({new_AGEMA_signal_5860, SubBytesIns_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_5858, SubBytesIns_Inst_Sbox_2_M20}), .clk (clk), .r ({Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_5938, SubBytesIns_Inst_Sbox_2_M25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M26_U1 ( .a ({new_AGEMA_signal_10238, new_AGEMA_signal_10237}), .b ({new_AGEMA_signal_5938, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_6024, SubBytesIns_Inst_Sbox_2_M26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M28_U1 ( .a ({new_AGEMA_signal_10240, new_AGEMA_signal_10239}), .b ({new_AGEMA_signal_5938, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_6025, SubBytesIns_Inst_Sbox_2_M28}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M31_U1 ( .a ({new_AGEMA_signal_5858, SubBytesIns_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_5937, SubBytesIns_Inst_Sbox_2_M23}), .clk (clk), .r ({Fresh[375], Fresh[374]}), .c ({new_AGEMA_signal_6026, SubBytesIns_Inst_Sbox_2_M31}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M33_U1 ( .a ({new_AGEMA_signal_10242, new_AGEMA_signal_10241}), .b ({new_AGEMA_signal_5938, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_6027, SubBytesIns_Inst_Sbox_2_M33}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M34_U1 ( .a ({new_AGEMA_signal_5859, SubBytesIns_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_5860, SubBytesIns_Inst_Sbox_2_M22}), .clk (clk), .r ({Fresh[377], Fresh[376]}), .c ({new_AGEMA_signal_5940, SubBytesIns_Inst_Sbox_2_M34}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M36_U1 ( .a ({new_AGEMA_signal_10244, new_AGEMA_signal_10243}), .b ({new_AGEMA_signal_5938, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_6127, SubBytesIns_Inst_Sbox_2_M36}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M25_U1 ( .a ({new_AGEMA_signal_5864, SubBytesIns_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_5862, SubBytesIns_Inst_Sbox_3_M20}), .clk (clk), .r ({Fresh[379], Fresh[378]}), .c ({new_AGEMA_signal_5942, SubBytesIns_Inst_Sbox_3_M25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M26_U1 ( .a ({new_AGEMA_signal_10246, new_AGEMA_signal_10245}), .b ({new_AGEMA_signal_5942, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_6029, SubBytesIns_Inst_Sbox_3_M26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M28_U1 ( .a ({new_AGEMA_signal_10248, new_AGEMA_signal_10247}), .b ({new_AGEMA_signal_5942, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_6030, SubBytesIns_Inst_Sbox_3_M28}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M31_U1 ( .a ({new_AGEMA_signal_5862, SubBytesIns_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_5941, SubBytesIns_Inst_Sbox_3_M23}), .clk (clk), .r ({Fresh[381], Fresh[380]}), .c ({new_AGEMA_signal_6031, SubBytesIns_Inst_Sbox_3_M31}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M33_U1 ( .a ({new_AGEMA_signal_10250, new_AGEMA_signal_10249}), .b ({new_AGEMA_signal_5942, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_6032, SubBytesIns_Inst_Sbox_3_M33}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M34_U1 ( .a ({new_AGEMA_signal_5863, SubBytesIns_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_5864, SubBytesIns_Inst_Sbox_3_M22}), .clk (clk), .r ({Fresh[383], Fresh[382]}), .c ({new_AGEMA_signal_5944, SubBytesIns_Inst_Sbox_3_M34}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M36_U1 ( .a ({new_AGEMA_signal_10252, new_AGEMA_signal_10251}), .b ({new_AGEMA_signal_5942, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_6132, SubBytesIns_Inst_Sbox_3_M36}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M25_U1 ( .a ({new_AGEMA_signal_5868, SubBytesIns_Inst_Sbox_4_M22}), .b ({new_AGEMA_signal_5866, SubBytesIns_Inst_Sbox_4_M20}), .clk (clk), .r ({Fresh[385], Fresh[384]}), .c ({new_AGEMA_signal_5946, SubBytesIns_Inst_Sbox_4_M25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M26_U1 ( .a ({new_AGEMA_signal_10254, new_AGEMA_signal_10253}), .b ({new_AGEMA_signal_5946, SubBytesIns_Inst_Sbox_4_M25}), .c ({new_AGEMA_signal_6034, SubBytesIns_Inst_Sbox_4_M26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M28_U1 ( .a ({new_AGEMA_signal_10256, new_AGEMA_signal_10255}), .b ({new_AGEMA_signal_5946, SubBytesIns_Inst_Sbox_4_M25}), .c ({new_AGEMA_signal_6035, SubBytesIns_Inst_Sbox_4_M28}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M31_U1 ( .a ({new_AGEMA_signal_5866, SubBytesIns_Inst_Sbox_4_M20}), .b ({new_AGEMA_signal_5945, SubBytesIns_Inst_Sbox_4_M23}), .clk (clk), .r ({Fresh[387], Fresh[386]}), .c ({new_AGEMA_signal_6036, SubBytesIns_Inst_Sbox_4_M31}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M33_U1 ( .a ({new_AGEMA_signal_10258, new_AGEMA_signal_10257}), .b ({new_AGEMA_signal_5946, SubBytesIns_Inst_Sbox_4_M25}), .c ({new_AGEMA_signal_6037, SubBytesIns_Inst_Sbox_4_M33}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M34_U1 ( .a ({new_AGEMA_signal_5867, SubBytesIns_Inst_Sbox_4_M21}), .b ({new_AGEMA_signal_5868, SubBytesIns_Inst_Sbox_4_M22}), .clk (clk), .r ({Fresh[389], Fresh[388]}), .c ({new_AGEMA_signal_5948, SubBytesIns_Inst_Sbox_4_M34}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M36_U1 ( .a ({new_AGEMA_signal_10260, new_AGEMA_signal_10259}), .b ({new_AGEMA_signal_5946, SubBytesIns_Inst_Sbox_4_M25}), .c ({new_AGEMA_signal_6137, SubBytesIns_Inst_Sbox_4_M36}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M25_U1 ( .a ({new_AGEMA_signal_5872, SubBytesIns_Inst_Sbox_5_M22}), .b ({new_AGEMA_signal_5870, SubBytesIns_Inst_Sbox_5_M20}), .clk (clk), .r ({Fresh[391], Fresh[390]}), .c ({new_AGEMA_signal_5950, SubBytesIns_Inst_Sbox_5_M25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M26_U1 ( .a ({new_AGEMA_signal_10262, new_AGEMA_signal_10261}), .b ({new_AGEMA_signal_5950, SubBytesIns_Inst_Sbox_5_M25}), .c ({new_AGEMA_signal_6039, SubBytesIns_Inst_Sbox_5_M26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M28_U1 ( .a ({new_AGEMA_signal_10264, new_AGEMA_signal_10263}), .b ({new_AGEMA_signal_5950, SubBytesIns_Inst_Sbox_5_M25}), .c ({new_AGEMA_signal_6040, SubBytesIns_Inst_Sbox_5_M28}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M31_U1 ( .a ({new_AGEMA_signal_5870, SubBytesIns_Inst_Sbox_5_M20}), .b ({new_AGEMA_signal_5949, SubBytesIns_Inst_Sbox_5_M23}), .clk (clk), .r ({Fresh[393], Fresh[392]}), .c ({new_AGEMA_signal_6041, SubBytesIns_Inst_Sbox_5_M31}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M33_U1 ( .a ({new_AGEMA_signal_10266, new_AGEMA_signal_10265}), .b ({new_AGEMA_signal_5950, SubBytesIns_Inst_Sbox_5_M25}), .c ({new_AGEMA_signal_6042, SubBytesIns_Inst_Sbox_5_M33}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M34_U1 ( .a ({new_AGEMA_signal_5871, SubBytesIns_Inst_Sbox_5_M21}), .b ({new_AGEMA_signal_5872, SubBytesIns_Inst_Sbox_5_M22}), .clk (clk), .r ({Fresh[395], Fresh[394]}), .c ({new_AGEMA_signal_5952, SubBytesIns_Inst_Sbox_5_M34}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M36_U1 ( .a ({new_AGEMA_signal_10268, new_AGEMA_signal_10267}), .b ({new_AGEMA_signal_5950, SubBytesIns_Inst_Sbox_5_M25}), .c ({new_AGEMA_signal_6142, SubBytesIns_Inst_Sbox_5_M36}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M25_U1 ( .a ({new_AGEMA_signal_5876, SubBytesIns_Inst_Sbox_6_M22}), .b ({new_AGEMA_signal_5874, SubBytesIns_Inst_Sbox_6_M20}), .clk (clk), .r ({Fresh[397], Fresh[396]}), .c ({new_AGEMA_signal_5954, SubBytesIns_Inst_Sbox_6_M25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M26_U1 ( .a ({new_AGEMA_signal_10270, new_AGEMA_signal_10269}), .b ({new_AGEMA_signal_5954, SubBytesIns_Inst_Sbox_6_M25}), .c ({new_AGEMA_signal_6044, SubBytesIns_Inst_Sbox_6_M26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M28_U1 ( .a ({new_AGEMA_signal_10272, new_AGEMA_signal_10271}), .b ({new_AGEMA_signal_5954, SubBytesIns_Inst_Sbox_6_M25}), .c ({new_AGEMA_signal_6045, SubBytesIns_Inst_Sbox_6_M28}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M31_U1 ( .a ({new_AGEMA_signal_5874, SubBytesIns_Inst_Sbox_6_M20}), .b ({new_AGEMA_signal_5953, SubBytesIns_Inst_Sbox_6_M23}), .clk (clk), .r ({Fresh[399], Fresh[398]}), .c ({new_AGEMA_signal_6046, SubBytesIns_Inst_Sbox_6_M31}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M33_U1 ( .a ({new_AGEMA_signal_10274, new_AGEMA_signal_10273}), .b ({new_AGEMA_signal_5954, SubBytesIns_Inst_Sbox_6_M25}), .c ({new_AGEMA_signal_6047, SubBytesIns_Inst_Sbox_6_M33}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M34_U1 ( .a ({new_AGEMA_signal_5875, SubBytesIns_Inst_Sbox_6_M21}), .b ({new_AGEMA_signal_5876, SubBytesIns_Inst_Sbox_6_M22}), .clk (clk), .r ({Fresh[401], Fresh[400]}), .c ({new_AGEMA_signal_5956, SubBytesIns_Inst_Sbox_6_M34}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M36_U1 ( .a ({new_AGEMA_signal_10276, new_AGEMA_signal_10275}), .b ({new_AGEMA_signal_5954, SubBytesIns_Inst_Sbox_6_M25}), .c ({new_AGEMA_signal_6147, SubBytesIns_Inst_Sbox_6_M36}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M25_U1 ( .a ({new_AGEMA_signal_5880, SubBytesIns_Inst_Sbox_7_M22}), .b ({new_AGEMA_signal_5878, SubBytesIns_Inst_Sbox_7_M20}), .clk (clk), .r ({Fresh[403], Fresh[402]}), .c ({new_AGEMA_signal_5958, SubBytesIns_Inst_Sbox_7_M25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M26_U1 ( .a ({new_AGEMA_signal_10278, new_AGEMA_signal_10277}), .b ({new_AGEMA_signal_5958, SubBytesIns_Inst_Sbox_7_M25}), .c ({new_AGEMA_signal_6049, SubBytesIns_Inst_Sbox_7_M26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M28_U1 ( .a ({new_AGEMA_signal_10280, new_AGEMA_signal_10279}), .b ({new_AGEMA_signal_5958, SubBytesIns_Inst_Sbox_7_M25}), .c ({new_AGEMA_signal_6050, SubBytesIns_Inst_Sbox_7_M28}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M31_U1 ( .a ({new_AGEMA_signal_5878, SubBytesIns_Inst_Sbox_7_M20}), .b ({new_AGEMA_signal_5957, SubBytesIns_Inst_Sbox_7_M23}), .clk (clk), .r ({Fresh[405], Fresh[404]}), .c ({new_AGEMA_signal_6051, SubBytesIns_Inst_Sbox_7_M31}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M33_U1 ( .a ({new_AGEMA_signal_10282, new_AGEMA_signal_10281}), .b ({new_AGEMA_signal_5958, SubBytesIns_Inst_Sbox_7_M25}), .c ({new_AGEMA_signal_6052, SubBytesIns_Inst_Sbox_7_M33}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M34_U1 ( .a ({new_AGEMA_signal_5879, SubBytesIns_Inst_Sbox_7_M21}), .b ({new_AGEMA_signal_5880, SubBytesIns_Inst_Sbox_7_M22}), .clk (clk), .r ({Fresh[407], Fresh[406]}), .c ({new_AGEMA_signal_5960, SubBytesIns_Inst_Sbox_7_M34}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M36_U1 ( .a ({new_AGEMA_signal_10284, new_AGEMA_signal_10283}), .b ({new_AGEMA_signal_5958, SubBytesIns_Inst_Sbox_7_M25}), .c ({new_AGEMA_signal_6152, SubBytesIns_Inst_Sbox_7_M36}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M25_U1 ( .a ({new_AGEMA_signal_5884, SubBytesIns_Inst_Sbox_8_M22}), .b ({new_AGEMA_signal_5882, SubBytesIns_Inst_Sbox_8_M20}), .clk (clk), .r ({Fresh[409], Fresh[408]}), .c ({new_AGEMA_signal_5962, SubBytesIns_Inst_Sbox_8_M25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M26_U1 ( .a ({new_AGEMA_signal_10286, new_AGEMA_signal_10285}), .b ({new_AGEMA_signal_5962, SubBytesIns_Inst_Sbox_8_M25}), .c ({new_AGEMA_signal_6054, SubBytesIns_Inst_Sbox_8_M26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M28_U1 ( .a ({new_AGEMA_signal_10288, new_AGEMA_signal_10287}), .b ({new_AGEMA_signal_5962, SubBytesIns_Inst_Sbox_8_M25}), .c ({new_AGEMA_signal_6055, SubBytesIns_Inst_Sbox_8_M28}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M31_U1 ( .a ({new_AGEMA_signal_5882, SubBytesIns_Inst_Sbox_8_M20}), .b ({new_AGEMA_signal_5961, SubBytesIns_Inst_Sbox_8_M23}), .clk (clk), .r ({Fresh[411], Fresh[410]}), .c ({new_AGEMA_signal_6056, SubBytesIns_Inst_Sbox_8_M31}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M33_U1 ( .a ({new_AGEMA_signal_10290, new_AGEMA_signal_10289}), .b ({new_AGEMA_signal_5962, SubBytesIns_Inst_Sbox_8_M25}), .c ({new_AGEMA_signal_6057, SubBytesIns_Inst_Sbox_8_M33}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M34_U1 ( .a ({new_AGEMA_signal_5883, SubBytesIns_Inst_Sbox_8_M21}), .b ({new_AGEMA_signal_5884, SubBytesIns_Inst_Sbox_8_M22}), .clk (clk), .r ({Fresh[413], Fresh[412]}), .c ({new_AGEMA_signal_5964, SubBytesIns_Inst_Sbox_8_M34}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M36_U1 ( .a ({new_AGEMA_signal_10292, new_AGEMA_signal_10291}), .b ({new_AGEMA_signal_5962, SubBytesIns_Inst_Sbox_8_M25}), .c ({new_AGEMA_signal_6157, SubBytesIns_Inst_Sbox_8_M36}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M25_U1 ( .a ({new_AGEMA_signal_5888, SubBytesIns_Inst_Sbox_9_M22}), .b ({new_AGEMA_signal_5886, SubBytesIns_Inst_Sbox_9_M20}), .clk (clk), .r ({Fresh[415], Fresh[414]}), .c ({new_AGEMA_signal_5966, SubBytesIns_Inst_Sbox_9_M25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M26_U1 ( .a ({new_AGEMA_signal_10294, new_AGEMA_signal_10293}), .b ({new_AGEMA_signal_5966, SubBytesIns_Inst_Sbox_9_M25}), .c ({new_AGEMA_signal_6059, SubBytesIns_Inst_Sbox_9_M26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M28_U1 ( .a ({new_AGEMA_signal_10296, new_AGEMA_signal_10295}), .b ({new_AGEMA_signal_5966, SubBytesIns_Inst_Sbox_9_M25}), .c ({new_AGEMA_signal_6060, SubBytesIns_Inst_Sbox_9_M28}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M31_U1 ( .a ({new_AGEMA_signal_5886, SubBytesIns_Inst_Sbox_9_M20}), .b ({new_AGEMA_signal_5965, SubBytesIns_Inst_Sbox_9_M23}), .clk (clk), .r ({Fresh[417], Fresh[416]}), .c ({new_AGEMA_signal_6061, SubBytesIns_Inst_Sbox_9_M31}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M33_U1 ( .a ({new_AGEMA_signal_10298, new_AGEMA_signal_10297}), .b ({new_AGEMA_signal_5966, SubBytesIns_Inst_Sbox_9_M25}), .c ({new_AGEMA_signal_6062, SubBytesIns_Inst_Sbox_9_M33}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M34_U1 ( .a ({new_AGEMA_signal_5887, SubBytesIns_Inst_Sbox_9_M21}), .b ({new_AGEMA_signal_5888, SubBytesIns_Inst_Sbox_9_M22}), .clk (clk), .r ({Fresh[419], Fresh[418]}), .c ({new_AGEMA_signal_5968, SubBytesIns_Inst_Sbox_9_M34}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M36_U1 ( .a ({new_AGEMA_signal_10300, new_AGEMA_signal_10299}), .b ({new_AGEMA_signal_5966, SubBytesIns_Inst_Sbox_9_M25}), .c ({new_AGEMA_signal_6162, SubBytesIns_Inst_Sbox_9_M36}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M25_U1 ( .a ({new_AGEMA_signal_5892, SubBytesIns_Inst_Sbox_10_M22}), .b ({new_AGEMA_signal_5890, SubBytesIns_Inst_Sbox_10_M20}), .clk (clk), .r ({Fresh[421], Fresh[420]}), .c ({new_AGEMA_signal_5970, SubBytesIns_Inst_Sbox_10_M25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M26_U1 ( .a ({new_AGEMA_signal_10302, new_AGEMA_signal_10301}), .b ({new_AGEMA_signal_5970, SubBytesIns_Inst_Sbox_10_M25}), .c ({new_AGEMA_signal_6064, SubBytesIns_Inst_Sbox_10_M26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M28_U1 ( .a ({new_AGEMA_signal_10304, new_AGEMA_signal_10303}), .b ({new_AGEMA_signal_5970, SubBytesIns_Inst_Sbox_10_M25}), .c ({new_AGEMA_signal_6065, SubBytesIns_Inst_Sbox_10_M28}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M31_U1 ( .a ({new_AGEMA_signal_5890, SubBytesIns_Inst_Sbox_10_M20}), .b ({new_AGEMA_signal_5969, SubBytesIns_Inst_Sbox_10_M23}), .clk (clk), .r ({Fresh[423], Fresh[422]}), .c ({new_AGEMA_signal_6066, SubBytesIns_Inst_Sbox_10_M31}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M33_U1 ( .a ({new_AGEMA_signal_10306, new_AGEMA_signal_10305}), .b ({new_AGEMA_signal_5970, SubBytesIns_Inst_Sbox_10_M25}), .c ({new_AGEMA_signal_6067, SubBytesIns_Inst_Sbox_10_M33}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M34_U1 ( .a ({new_AGEMA_signal_5891, SubBytesIns_Inst_Sbox_10_M21}), .b ({new_AGEMA_signal_5892, SubBytesIns_Inst_Sbox_10_M22}), .clk (clk), .r ({Fresh[425], Fresh[424]}), .c ({new_AGEMA_signal_5972, SubBytesIns_Inst_Sbox_10_M34}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M36_U1 ( .a ({new_AGEMA_signal_10308, new_AGEMA_signal_10307}), .b ({new_AGEMA_signal_5970, SubBytesIns_Inst_Sbox_10_M25}), .c ({new_AGEMA_signal_6167, SubBytesIns_Inst_Sbox_10_M36}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M25_U1 ( .a ({new_AGEMA_signal_5896, SubBytesIns_Inst_Sbox_11_M22}), .b ({new_AGEMA_signal_5894, SubBytesIns_Inst_Sbox_11_M20}), .clk (clk), .r ({Fresh[427], Fresh[426]}), .c ({new_AGEMA_signal_5974, SubBytesIns_Inst_Sbox_11_M25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M26_U1 ( .a ({new_AGEMA_signal_10310, new_AGEMA_signal_10309}), .b ({new_AGEMA_signal_5974, SubBytesIns_Inst_Sbox_11_M25}), .c ({new_AGEMA_signal_6069, SubBytesIns_Inst_Sbox_11_M26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M28_U1 ( .a ({new_AGEMA_signal_10312, new_AGEMA_signal_10311}), .b ({new_AGEMA_signal_5974, SubBytesIns_Inst_Sbox_11_M25}), .c ({new_AGEMA_signal_6070, SubBytesIns_Inst_Sbox_11_M28}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M31_U1 ( .a ({new_AGEMA_signal_5894, SubBytesIns_Inst_Sbox_11_M20}), .b ({new_AGEMA_signal_5973, SubBytesIns_Inst_Sbox_11_M23}), .clk (clk), .r ({Fresh[429], Fresh[428]}), .c ({new_AGEMA_signal_6071, SubBytesIns_Inst_Sbox_11_M31}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M33_U1 ( .a ({new_AGEMA_signal_10314, new_AGEMA_signal_10313}), .b ({new_AGEMA_signal_5974, SubBytesIns_Inst_Sbox_11_M25}), .c ({new_AGEMA_signal_6072, SubBytesIns_Inst_Sbox_11_M33}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M34_U1 ( .a ({new_AGEMA_signal_5895, SubBytesIns_Inst_Sbox_11_M21}), .b ({new_AGEMA_signal_5896, SubBytesIns_Inst_Sbox_11_M22}), .clk (clk), .r ({Fresh[431], Fresh[430]}), .c ({new_AGEMA_signal_5976, SubBytesIns_Inst_Sbox_11_M34}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M36_U1 ( .a ({new_AGEMA_signal_10316, new_AGEMA_signal_10315}), .b ({new_AGEMA_signal_5974, SubBytesIns_Inst_Sbox_11_M25}), .c ({new_AGEMA_signal_6172, SubBytesIns_Inst_Sbox_11_M36}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M25_U1 ( .a ({new_AGEMA_signal_5900, SubBytesIns_Inst_Sbox_12_M22}), .b ({new_AGEMA_signal_5898, SubBytesIns_Inst_Sbox_12_M20}), .clk (clk), .r ({Fresh[433], Fresh[432]}), .c ({new_AGEMA_signal_5978, SubBytesIns_Inst_Sbox_12_M25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M26_U1 ( .a ({new_AGEMA_signal_10318, new_AGEMA_signal_10317}), .b ({new_AGEMA_signal_5978, SubBytesIns_Inst_Sbox_12_M25}), .c ({new_AGEMA_signal_6074, SubBytesIns_Inst_Sbox_12_M26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M28_U1 ( .a ({new_AGEMA_signal_10320, new_AGEMA_signal_10319}), .b ({new_AGEMA_signal_5978, SubBytesIns_Inst_Sbox_12_M25}), .c ({new_AGEMA_signal_6075, SubBytesIns_Inst_Sbox_12_M28}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M31_U1 ( .a ({new_AGEMA_signal_5898, SubBytesIns_Inst_Sbox_12_M20}), .b ({new_AGEMA_signal_5977, SubBytesIns_Inst_Sbox_12_M23}), .clk (clk), .r ({Fresh[435], Fresh[434]}), .c ({new_AGEMA_signal_6076, SubBytesIns_Inst_Sbox_12_M31}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M33_U1 ( .a ({new_AGEMA_signal_10322, new_AGEMA_signal_10321}), .b ({new_AGEMA_signal_5978, SubBytesIns_Inst_Sbox_12_M25}), .c ({new_AGEMA_signal_6077, SubBytesIns_Inst_Sbox_12_M33}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M34_U1 ( .a ({new_AGEMA_signal_5899, SubBytesIns_Inst_Sbox_12_M21}), .b ({new_AGEMA_signal_5900, SubBytesIns_Inst_Sbox_12_M22}), .clk (clk), .r ({Fresh[437], Fresh[436]}), .c ({new_AGEMA_signal_5980, SubBytesIns_Inst_Sbox_12_M34}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M36_U1 ( .a ({new_AGEMA_signal_10324, new_AGEMA_signal_10323}), .b ({new_AGEMA_signal_5978, SubBytesIns_Inst_Sbox_12_M25}), .c ({new_AGEMA_signal_6177, SubBytesIns_Inst_Sbox_12_M36}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M25_U1 ( .a ({new_AGEMA_signal_5904, SubBytesIns_Inst_Sbox_13_M22}), .b ({new_AGEMA_signal_5902, SubBytesIns_Inst_Sbox_13_M20}), .clk (clk), .r ({Fresh[439], Fresh[438]}), .c ({new_AGEMA_signal_5982, SubBytesIns_Inst_Sbox_13_M25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M26_U1 ( .a ({new_AGEMA_signal_10326, new_AGEMA_signal_10325}), .b ({new_AGEMA_signal_5982, SubBytesIns_Inst_Sbox_13_M25}), .c ({new_AGEMA_signal_6079, SubBytesIns_Inst_Sbox_13_M26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M28_U1 ( .a ({new_AGEMA_signal_10328, new_AGEMA_signal_10327}), .b ({new_AGEMA_signal_5982, SubBytesIns_Inst_Sbox_13_M25}), .c ({new_AGEMA_signal_6080, SubBytesIns_Inst_Sbox_13_M28}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M31_U1 ( .a ({new_AGEMA_signal_5902, SubBytesIns_Inst_Sbox_13_M20}), .b ({new_AGEMA_signal_5981, SubBytesIns_Inst_Sbox_13_M23}), .clk (clk), .r ({Fresh[441], Fresh[440]}), .c ({new_AGEMA_signal_6081, SubBytesIns_Inst_Sbox_13_M31}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M33_U1 ( .a ({new_AGEMA_signal_10330, new_AGEMA_signal_10329}), .b ({new_AGEMA_signal_5982, SubBytesIns_Inst_Sbox_13_M25}), .c ({new_AGEMA_signal_6082, SubBytesIns_Inst_Sbox_13_M33}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M34_U1 ( .a ({new_AGEMA_signal_5903, SubBytesIns_Inst_Sbox_13_M21}), .b ({new_AGEMA_signal_5904, SubBytesIns_Inst_Sbox_13_M22}), .clk (clk), .r ({Fresh[443], Fresh[442]}), .c ({new_AGEMA_signal_5984, SubBytesIns_Inst_Sbox_13_M34}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M36_U1 ( .a ({new_AGEMA_signal_10332, new_AGEMA_signal_10331}), .b ({new_AGEMA_signal_5982, SubBytesIns_Inst_Sbox_13_M25}), .c ({new_AGEMA_signal_6182, SubBytesIns_Inst_Sbox_13_M36}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M25_U1 ( .a ({new_AGEMA_signal_5908, SubBytesIns_Inst_Sbox_14_M22}), .b ({new_AGEMA_signal_5906, SubBytesIns_Inst_Sbox_14_M20}), .clk (clk), .r ({Fresh[445], Fresh[444]}), .c ({new_AGEMA_signal_5986, SubBytesIns_Inst_Sbox_14_M25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M26_U1 ( .a ({new_AGEMA_signal_10334, new_AGEMA_signal_10333}), .b ({new_AGEMA_signal_5986, SubBytesIns_Inst_Sbox_14_M25}), .c ({new_AGEMA_signal_6084, SubBytesIns_Inst_Sbox_14_M26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M28_U1 ( .a ({new_AGEMA_signal_10336, new_AGEMA_signal_10335}), .b ({new_AGEMA_signal_5986, SubBytesIns_Inst_Sbox_14_M25}), .c ({new_AGEMA_signal_6085, SubBytesIns_Inst_Sbox_14_M28}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M31_U1 ( .a ({new_AGEMA_signal_5906, SubBytesIns_Inst_Sbox_14_M20}), .b ({new_AGEMA_signal_5985, SubBytesIns_Inst_Sbox_14_M23}), .clk (clk), .r ({Fresh[447], Fresh[446]}), .c ({new_AGEMA_signal_6086, SubBytesIns_Inst_Sbox_14_M31}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M33_U1 ( .a ({new_AGEMA_signal_10338, new_AGEMA_signal_10337}), .b ({new_AGEMA_signal_5986, SubBytesIns_Inst_Sbox_14_M25}), .c ({new_AGEMA_signal_6087, SubBytesIns_Inst_Sbox_14_M33}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M34_U1 ( .a ({new_AGEMA_signal_5907, SubBytesIns_Inst_Sbox_14_M21}), .b ({new_AGEMA_signal_5908, SubBytesIns_Inst_Sbox_14_M22}), .clk (clk), .r ({Fresh[449], Fresh[448]}), .c ({new_AGEMA_signal_5988, SubBytesIns_Inst_Sbox_14_M34}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M36_U1 ( .a ({new_AGEMA_signal_10340, new_AGEMA_signal_10339}), .b ({new_AGEMA_signal_5986, SubBytesIns_Inst_Sbox_14_M25}), .c ({new_AGEMA_signal_6187, SubBytesIns_Inst_Sbox_14_M36}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M25_U1 ( .a ({new_AGEMA_signal_5912, SubBytesIns_Inst_Sbox_15_M22}), .b ({new_AGEMA_signal_5910, SubBytesIns_Inst_Sbox_15_M20}), .clk (clk), .r ({Fresh[451], Fresh[450]}), .c ({new_AGEMA_signal_5990, SubBytesIns_Inst_Sbox_15_M25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M26_U1 ( .a ({new_AGEMA_signal_10342, new_AGEMA_signal_10341}), .b ({new_AGEMA_signal_5990, SubBytesIns_Inst_Sbox_15_M25}), .c ({new_AGEMA_signal_6089, SubBytesIns_Inst_Sbox_15_M26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M28_U1 ( .a ({new_AGEMA_signal_10344, new_AGEMA_signal_10343}), .b ({new_AGEMA_signal_5990, SubBytesIns_Inst_Sbox_15_M25}), .c ({new_AGEMA_signal_6090, SubBytesIns_Inst_Sbox_15_M28}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M31_U1 ( .a ({new_AGEMA_signal_5910, SubBytesIns_Inst_Sbox_15_M20}), .b ({new_AGEMA_signal_5989, SubBytesIns_Inst_Sbox_15_M23}), .clk (clk), .r ({Fresh[453], Fresh[452]}), .c ({new_AGEMA_signal_6091, SubBytesIns_Inst_Sbox_15_M31}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M33_U1 ( .a ({new_AGEMA_signal_10346, new_AGEMA_signal_10345}), .b ({new_AGEMA_signal_5990, SubBytesIns_Inst_Sbox_15_M25}), .c ({new_AGEMA_signal_6092, SubBytesIns_Inst_Sbox_15_M33}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M34_U1 ( .a ({new_AGEMA_signal_5911, SubBytesIns_Inst_Sbox_15_M21}), .b ({new_AGEMA_signal_5912, SubBytesIns_Inst_Sbox_15_M22}), .clk (clk), .r ({Fresh[455], Fresh[454]}), .c ({new_AGEMA_signal_5992, SubBytesIns_Inst_Sbox_15_M34}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M36_U1 ( .a ({new_AGEMA_signal_10348, new_AGEMA_signal_10347}), .b ({new_AGEMA_signal_5990, SubBytesIns_Inst_Sbox_15_M25}), .c ({new_AGEMA_signal_6192, SubBytesIns_Inst_Sbox_15_M36}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M25_U1 ( .a ({new_AGEMA_signal_5836, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_5834, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20}), .clk (clk), .r ({Fresh[457], Fresh[456]}), .c ({new_AGEMA_signal_5914, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M26_U1 ( .a ({new_AGEMA_signal_10350, new_AGEMA_signal_10349}), .b ({new_AGEMA_signal_5914, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_5994, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M28_U1 ( .a ({new_AGEMA_signal_10352, new_AGEMA_signal_10351}), .b ({new_AGEMA_signal_5914, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_5995, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M28}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M31_U1 ( .a ({new_AGEMA_signal_5834, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_5913, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23}), .clk (clk), .r ({Fresh[459], Fresh[458]}), .c ({new_AGEMA_signal_5996, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M31}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M33_U1 ( .a ({new_AGEMA_signal_10354, new_AGEMA_signal_10353}), .b ({new_AGEMA_signal_5914, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_5997, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M33}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M34_U1 ( .a ({new_AGEMA_signal_5835, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_5836, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22}), .clk (clk), .r ({Fresh[461], Fresh[460]}), .c ({new_AGEMA_signal_5916, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M34}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M36_U1 ( .a ({new_AGEMA_signal_10356, new_AGEMA_signal_10355}), .b ({new_AGEMA_signal_5914, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_6097, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M36}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M25_U1 ( .a ({new_AGEMA_signal_5840, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_5838, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20}), .clk (clk), .r ({Fresh[463], Fresh[462]}), .c ({new_AGEMA_signal_5918, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M26_U1 ( .a ({new_AGEMA_signal_10358, new_AGEMA_signal_10357}), .b ({new_AGEMA_signal_5918, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_5999, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M28_U1 ( .a ({new_AGEMA_signal_10360, new_AGEMA_signal_10359}), .b ({new_AGEMA_signal_5918, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_6000, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M28}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M31_U1 ( .a ({new_AGEMA_signal_5838, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_5917, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23}), .clk (clk), .r ({Fresh[465], Fresh[464]}), .c ({new_AGEMA_signal_6001, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M31}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M33_U1 ( .a ({new_AGEMA_signal_10362, new_AGEMA_signal_10361}), .b ({new_AGEMA_signal_5918, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_6002, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M33}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M34_U1 ( .a ({new_AGEMA_signal_5839, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_5840, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22}), .clk (clk), .r ({Fresh[467], Fresh[466]}), .c ({new_AGEMA_signal_5920, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M34}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M36_U1 ( .a ({new_AGEMA_signal_10364, new_AGEMA_signal_10363}), .b ({new_AGEMA_signal_5918, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_6102, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M36}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M25_U1 ( .a ({new_AGEMA_signal_5844, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_5842, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20}), .clk (clk), .r ({Fresh[469], Fresh[468]}), .c ({new_AGEMA_signal_5922, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M26_U1 ( .a ({new_AGEMA_signal_10366, new_AGEMA_signal_10365}), .b ({new_AGEMA_signal_5922, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_6004, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M28_U1 ( .a ({new_AGEMA_signal_10368, new_AGEMA_signal_10367}), .b ({new_AGEMA_signal_5922, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_6005, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M28}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M31_U1 ( .a ({new_AGEMA_signal_5842, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_5921, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23}), .clk (clk), .r ({Fresh[471], Fresh[470]}), .c ({new_AGEMA_signal_6006, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M31}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M33_U1 ( .a ({new_AGEMA_signal_10370, new_AGEMA_signal_10369}), .b ({new_AGEMA_signal_5922, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_6007, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M33}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M34_U1 ( .a ({new_AGEMA_signal_5843, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_5844, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22}), .clk (clk), .r ({Fresh[473], Fresh[472]}), .c ({new_AGEMA_signal_5924, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M34}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M36_U1 ( .a ({new_AGEMA_signal_10372, new_AGEMA_signal_10371}), .b ({new_AGEMA_signal_5922, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_6107, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M36}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M25_U1 ( .a ({new_AGEMA_signal_5848, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_5846, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20}), .clk (clk), .r ({Fresh[475], Fresh[474]}), .c ({new_AGEMA_signal_5926, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M26_U1 ( .a ({new_AGEMA_signal_10374, new_AGEMA_signal_10373}), .b ({new_AGEMA_signal_5926, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_6009, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M28_U1 ( .a ({new_AGEMA_signal_10376, new_AGEMA_signal_10375}), .b ({new_AGEMA_signal_5926, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_6010, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M28}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M31_U1 ( .a ({new_AGEMA_signal_5846, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_5925, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23}), .clk (clk), .r ({Fresh[477], Fresh[476]}), .c ({new_AGEMA_signal_6011, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M31}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M33_U1 ( .a ({new_AGEMA_signal_10378, new_AGEMA_signal_10377}), .b ({new_AGEMA_signal_5926, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_6012, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M33}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M34_U1 ( .a ({new_AGEMA_signal_5847, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_5848, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22}), .clk (clk), .r ({Fresh[479], Fresh[478]}), .c ({new_AGEMA_signal_5928, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M34}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M36_U1 ( .a ({new_AGEMA_signal_10380, new_AGEMA_signal_10379}), .b ({new_AGEMA_signal_5926, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_6112, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M36}) ) ;
    buf_clk new_AGEMA_reg_buffer_4369 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M21), .Q (new_AGEMA_signal_10221) ) ;
    buf_clk new_AGEMA_reg_buffer_4370 ( .C (clk), .D (new_AGEMA_signal_5851), .Q (new_AGEMA_signal_10222) ) ;
    buf_clk new_AGEMA_reg_buffer_4371 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M23), .Q (new_AGEMA_signal_10223) ) ;
    buf_clk new_AGEMA_reg_buffer_4372 ( .C (clk), .D (new_AGEMA_signal_5929), .Q (new_AGEMA_signal_10224) ) ;
    buf_clk new_AGEMA_reg_buffer_4373 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M27), .Q (new_AGEMA_signal_10225) ) ;
    buf_clk new_AGEMA_reg_buffer_4374 ( .C (clk), .D (new_AGEMA_signal_5931), .Q (new_AGEMA_signal_10226) ) ;
    buf_clk new_AGEMA_reg_buffer_4375 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M24), .Q (new_AGEMA_signal_10227) ) ;
    buf_clk new_AGEMA_reg_buffer_4376 ( .C (clk), .D (new_AGEMA_signal_6013), .Q (new_AGEMA_signal_10228) ) ;
    buf_clk new_AGEMA_reg_buffer_4377 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M21), .Q (new_AGEMA_signal_10229) ) ;
    buf_clk new_AGEMA_reg_buffer_4378 ( .C (clk), .D (new_AGEMA_signal_5855), .Q (new_AGEMA_signal_10230) ) ;
    buf_clk new_AGEMA_reg_buffer_4379 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M23), .Q (new_AGEMA_signal_10231) ) ;
    buf_clk new_AGEMA_reg_buffer_4380 ( .C (clk), .D (new_AGEMA_signal_5933), .Q (new_AGEMA_signal_10232) ) ;
    buf_clk new_AGEMA_reg_buffer_4381 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M27), .Q (new_AGEMA_signal_10233) ) ;
    buf_clk new_AGEMA_reg_buffer_4382 ( .C (clk), .D (new_AGEMA_signal_5935), .Q (new_AGEMA_signal_10234) ) ;
    buf_clk new_AGEMA_reg_buffer_4383 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M24), .Q (new_AGEMA_signal_10235) ) ;
    buf_clk new_AGEMA_reg_buffer_4384 ( .C (clk), .D (new_AGEMA_signal_6018), .Q (new_AGEMA_signal_10236) ) ;
    buf_clk new_AGEMA_reg_buffer_4385 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M21), .Q (new_AGEMA_signal_10237) ) ;
    buf_clk new_AGEMA_reg_buffer_4386 ( .C (clk), .D (new_AGEMA_signal_5859), .Q (new_AGEMA_signal_10238) ) ;
    buf_clk new_AGEMA_reg_buffer_4387 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M23), .Q (new_AGEMA_signal_10239) ) ;
    buf_clk new_AGEMA_reg_buffer_4388 ( .C (clk), .D (new_AGEMA_signal_5937), .Q (new_AGEMA_signal_10240) ) ;
    buf_clk new_AGEMA_reg_buffer_4389 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M27), .Q (new_AGEMA_signal_10241) ) ;
    buf_clk new_AGEMA_reg_buffer_4390 ( .C (clk), .D (new_AGEMA_signal_5939), .Q (new_AGEMA_signal_10242) ) ;
    buf_clk new_AGEMA_reg_buffer_4391 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M24), .Q (new_AGEMA_signal_10243) ) ;
    buf_clk new_AGEMA_reg_buffer_4392 ( .C (clk), .D (new_AGEMA_signal_6023), .Q (new_AGEMA_signal_10244) ) ;
    buf_clk new_AGEMA_reg_buffer_4393 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M21), .Q (new_AGEMA_signal_10245) ) ;
    buf_clk new_AGEMA_reg_buffer_4394 ( .C (clk), .D (new_AGEMA_signal_5863), .Q (new_AGEMA_signal_10246) ) ;
    buf_clk new_AGEMA_reg_buffer_4395 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M23), .Q (new_AGEMA_signal_10247) ) ;
    buf_clk new_AGEMA_reg_buffer_4396 ( .C (clk), .D (new_AGEMA_signal_5941), .Q (new_AGEMA_signal_10248) ) ;
    buf_clk new_AGEMA_reg_buffer_4397 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M27), .Q (new_AGEMA_signal_10249) ) ;
    buf_clk new_AGEMA_reg_buffer_4398 ( .C (clk), .D (new_AGEMA_signal_5943), .Q (new_AGEMA_signal_10250) ) ;
    buf_clk new_AGEMA_reg_buffer_4399 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M24), .Q (new_AGEMA_signal_10251) ) ;
    buf_clk new_AGEMA_reg_buffer_4400 ( .C (clk), .D (new_AGEMA_signal_6028), .Q (new_AGEMA_signal_10252) ) ;
    buf_clk new_AGEMA_reg_buffer_4401 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_M21), .Q (new_AGEMA_signal_10253) ) ;
    buf_clk new_AGEMA_reg_buffer_4402 ( .C (clk), .D (new_AGEMA_signal_5867), .Q (new_AGEMA_signal_10254) ) ;
    buf_clk new_AGEMA_reg_buffer_4403 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_M23), .Q (new_AGEMA_signal_10255) ) ;
    buf_clk new_AGEMA_reg_buffer_4404 ( .C (clk), .D (new_AGEMA_signal_5945), .Q (new_AGEMA_signal_10256) ) ;
    buf_clk new_AGEMA_reg_buffer_4405 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_M27), .Q (new_AGEMA_signal_10257) ) ;
    buf_clk new_AGEMA_reg_buffer_4406 ( .C (clk), .D (new_AGEMA_signal_5947), .Q (new_AGEMA_signal_10258) ) ;
    buf_clk new_AGEMA_reg_buffer_4407 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_M24), .Q (new_AGEMA_signal_10259) ) ;
    buf_clk new_AGEMA_reg_buffer_4408 ( .C (clk), .D (new_AGEMA_signal_6033), .Q (new_AGEMA_signal_10260) ) ;
    buf_clk new_AGEMA_reg_buffer_4409 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_M21), .Q (new_AGEMA_signal_10261) ) ;
    buf_clk new_AGEMA_reg_buffer_4410 ( .C (clk), .D (new_AGEMA_signal_5871), .Q (new_AGEMA_signal_10262) ) ;
    buf_clk new_AGEMA_reg_buffer_4411 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_M23), .Q (new_AGEMA_signal_10263) ) ;
    buf_clk new_AGEMA_reg_buffer_4412 ( .C (clk), .D (new_AGEMA_signal_5949), .Q (new_AGEMA_signal_10264) ) ;
    buf_clk new_AGEMA_reg_buffer_4413 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_M27), .Q (new_AGEMA_signal_10265) ) ;
    buf_clk new_AGEMA_reg_buffer_4414 ( .C (clk), .D (new_AGEMA_signal_5951), .Q (new_AGEMA_signal_10266) ) ;
    buf_clk new_AGEMA_reg_buffer_4415 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_M24), .Q (new_AGEMA_signal_10267) ) ;
    buf_clk new_AGEMA_reg_buffer_4416 ( .C (clk), .D (new_AGEMA_signal_6038), .Q (new_AGEMA_signal_10268) ) ;
    buf_clk new_AGEMA_reg_buffer_4417 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_M21), .Q (new_AGEMA_signal_10269) ) ;
    buf_clk new_AGEMA_reg_buffer_4418 ( .C (clk), .D (new_AGEMA_signal_5875), .Q (new_AGEMA_signal_10270) ) ;
    buf_clk new_AGEMA_reg_buffer_4419 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_M23), .Q (new_AGEMA_signal_10271) ) ;
    buf_clk new_AGEMA_reg_buffer_4420 ( .C (clk), .D (new_AGEMA_signal_5953), .Q (new_AGEMA_signal_10272) ) ;
    buf_clk new_AGEMA_reg_buffer_4421 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_M27), .Q (new_AGEMA_signal_10273) ) ;
    buf_clk new_AGEMA_reg_buffer_4422 ( .C (clk), .D (new_AGEMA_signal_5955), .Q (new_AGEMA_signal_10274) ) ;
    buf_clk new_AGEMA_reg_buffer_4423 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_M24), .Q (new_AGEMA_signal_10275) ) ;
    buf_clk new_AGEMA_reg_buffer_4424 ( .C (clk), .D (new_AGEMA_signal_6043), .Q (new_AGEMA_signal_10276) ) ;
    buf_clk new_AGEMA_reg_buffer_4425 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_M21), .Q (new_AGEMA_signal_10277) ) ;
    buf_clk new_AGEMA_reg_buffer_4426 ( .C (clk), .D (new_AGEMA_signal_5879), .Q (new_AGEMA_signal_10278) ) ;
    buf_clk new_AGEMA_reg_buffer_4427 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_M23), .Q (new_AGEMA_signal_10279) ) ;
    buf_clk new_AGEMA_reg_buffer_4428 ( .C (clk), .D (new_AGEMA_signal_5957), .Q (new_AGEMA_signal_10280) ) ;
    buf_clk new_AGEMA_reg_buffer_4429 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_M27), .Q (new_AGEMA_signal_10281) ) ;
    buf_clk new_AGEMA_reg_buffer_4430 ( .C (clk), .D (new_AGEMA_signal_5959), .Q (new_AGEMA_signal_10282) ) ;
    buf_clk new_AGEMA_reg_buffer_4431 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_M24), .Q (new_AGEMA_signal_10283) ) ;
    buf_clk new_AGEMA_reg_buffer_4432 ( .C (clk), .D (new_AGEMA_signal_6048), .Q (new_AGEMA_signal_10284) ) ;
    buf_clk new_AGEMA_reg_buffer_4433 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_M21), .Q (new_AGEMA_signal_10285) ) ;
    buf_clk new_AGEMA_reg_buffer_4434 ( .C (clk), .D (new_AGEMA_signal_5883), .Q (new_AGEMA_signal_10286) ) ;
    buf_clk new_AGEMA_reg_buffer_4435 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_M23), .Q (new_AGEMA_signal_10287) ) ;
    buf_clk new_AGEMA_reg_buffer_4436 ( .C (clk), .D (new_AGEMA_signal_5961), .Q (new_AGEMA_signal_10288) ) ;
    buf_clk new_AGEMA_reg_buffer_4437 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_M27), .Q (new_AGEMA_signal_10289) ) ;
    buf_clk new_AGEMA_reg_buffer_4438 ( .C (clk), .D (new_AGEMA_signal_5963), .Q (new_AGEMA_signal_10290) ) ;
    buf_clk new_AGEMA_reg_buffer_4439 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_M24), .Q (new_AGEMA_signal_10291) ) ;
    buf_clk new_AGEMA_reg_buffer_4440 ( .C (clk), .D (new_AGEMA_signal_6053), .Q (new_AGEMA_signal_10292) ) ;
    buf_clk new_AGEMA_reg_buffer_4441 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_M21), .Q (new_AGEMA_signal_10293) ) ;
    buf_clk new_AGEMA_reg_buffer_4442 ( .C (clk), .D (new_AGEMA_signal_5887), .Q (new_AGEMA_signal_10294) ) ;
    buf_clk new_AGEMA_reg_buffer_4443 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_M23), .Q (new_AGEMA_signal_10295) ) ;
    buf_clk new_AGEMA_reg_buffer_4444 ( .C (clk), .D (new_AGEMA_signal_5965), .Q (new_AGEMA_signal_10296) ) ;
    buf_clk new_AGEMA_reg_buffer_4445 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_M27), .Q (new_AGEMA_signal_10297) ) ;
    buf_clk new_AGEMA_reg_buffer_4446 ( .C (clk), .D (new_AGEMA_signal_5967), .Q (new_AGEMA_signal_10298) ) ;
    buf_clk new_AGEMA_reg_buffer_4447 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_M24), .Q (new_AGEMA_signal_10299) ) ;
    buf_clk new_AGEMA_reg_buffer_4448 ( .C (clk), .D (new_AGEMA_signal_6058), .Q (new_AGEMA_signal_10300) ) ;
    buf_clk new_AGEMA_reg_buffer_4449 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_M21), .Q (new_AGEMA_signal_10301) ) ;
    buf_clk new_AGEMA_reg_buffer_4450 ( .C (clk), .D (new_AGEMA_signal_5891), .Q (new_AGEMA_signal_10302) ) ;
    buf_clk new_AGEMA_reg_buffer_4451 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_M23), .Q (new_AGEMA_signal_10303) ) ;
    buf_clk new_AGEMA_reg_buffer_4452 ( .C (clk), .D (new_AGEMA_signal_5969), .Q (new_AGEMA_signal_10304) ) ;
    buf_clk new_AGEMA_reg_buffer_4453 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_M27), .Q (new_AGEMA_signal_10305) ) ;
    buf_clk new_AGEMA_reg_buffer_4454 ( .C (clk), .D (new_AGEMA_signal_5971), .Q (new_AGEMA_signal_10306) ) ;
    buf_clk new_AGEMA_reg_buffer_4455 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_M24), .Q (new_AGEMA_signal_10307) ) ;
    buf_clk new_AGEMA_reg_buffer_4456 ( .C (clk), .D (new_AGEMA_signal_6063), .Q (new_AGEMA_signal_10308) ) ;
    buf_clk new_AGEMA_reg_buffer_4457 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_M21), .Q (new_AGEMA_signal_10309) ) ;
    buf_clk new_AGEMA_reg_buffer_4458 ( .C (clk), .D (new_AGEMA_signal_5895), .Q (new_AGEMA_signal_10310) ) ;
    buf_clk new_AGEMA_reg_buffer_4459 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_M23), .Q (new_AGEMA_signal_10311) ) ;
    buf_clk new_AGEMA_reg_buffer_4460 ( .C (clk), .D (new_AGEMA_signal_5973), .Q (new_AGEMA_signal_10312) ) ;
    buf_clk new_AGEMA_reg_buffer_4461 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_M27), .Q (new_AGEMA_signal_10313) ) ;
    buf_clk new_AGEMA_reg_buffer_4462 ( .C (clk), .D (new_AGEMA_signal_5975), .Q (new_AGEMA_signal_10314) ) ;
    buf_clk new_AGEMA_reg_buffer_4463 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_M24), .Q (new_AGEMA_signal_10315) ) ;
    buf_clk new_AGEMA_reg_buffer_4464 ( .C (clk), .D (new_AGEMA_signal_6068), .Q (new_AGEMA_signal_10316) ) ;
    buf_clk new_AGEMA_reg_buffer_4465 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_M21), .Q (new_AGEMA_signal_10317) ) ;
    buf_clk new_AGEMA_reg_buffer_4466 ( .C (clk), .D (new_AGEMA_signal_5899), .Q (new_AGEMA_signal_10318) ) ;
    buf_clk new_AGEMA_reg_buffer_4467 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_M23), .Q (new_AGEMA_signal_10319) ) ;
    buf_clk new_AGEMA_reg_buffer_4468 ( .C (clk), .D (new_AGEMA_signal_5977), .Q (new_AGEMA_signal_10320) ) ;
    buf_clk new_AGEMA_reg_buffer_4469 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_M27), .Q (new_AGEMA_signal_10321) ) ;
    buf_clk new_AGEMA_reg_buffer_4470 ( .C (clk), .D (new_AGEMA_signal_5979), .Q (new_AGEMA_signal_10322) ) ;
    buf_clk new_AGEMA_reg_buffer_4471 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_M24), .Q (new_AGEMA_signal_10323) ) ;
    buf_clk new_AGEMA_reg_buffer_4472 ( .C (clk), .D (new_AGEMA_signal_6073), .Q (new_AGEMA_signal_10324) ) ;
    buf_clk new_AGEMA_reg_buffer_4473 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_M21), .Q (new_AGEMA_signal_10325) ) ;
    buf_clk new_AGEMA_reg_buffer_4474 ( .C (clk), .D (new_AGEMA_signal_5903), .Q (new_AGEMA_signal_10326) ) ;
    buf_clk new_AGEMA_reg_buffer_4475 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_M23), .Q (new_AGEMA_signal_10327) ) ;
    buf_clk new_AGEMA_reg_buffer_4476 ( .C (clk), .D (new_AGEMA_signal_5981), .Q (new_AGEMA_signal_10328) ) ;
    buf_clk new_AGEMA_reg_buffer_4477 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_M27), .Q (new_AGEMA_signal_10329) ) ;
    buf_clk new_AGEMA_reg_buffer_4478 ( .C (clk), .D (new_AGEMA_signal_5983), .Q (new_AGEMA_signal_10330) ) ;
    buf_clk new_AGEMA_reg_buffer_4479 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_M24), .Q (new_AGEMA_signal_10331) ) ;
    buf_clk new_AGEMA_reg_buffer_4480 ( .C (clk), .D (new_AGEMA_signal_6078), .Q (new_AGEMA_signal_10332) ) ;
    buf_clk new_AGEMA_reg_buffer_4481 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_M21), .Q (new_AGEMA_signal_10333) ) ;
    buf_clk new_AGEMA_reg_buffer_4482 ( .C (clk), .D (new_AGEMA_signal_5907), .Q (new_AGEMA_signal_10334) ) ;
    buf_clk new_AGEMA_reg_buffer_4483 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_M23), .Q (new_AGEMA_signal_10335) ) ;
    buf_clk new_AGEMA_reg_buffer_4484 ( .C (clk), .D (new_AGEMA_signal_5985), .Q (new_AGEMA_signal_10336) ) ;
    buf_clk new_AGEMA_reg_buffer_4485 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_M27), .Q (new_AGEMA_signal_10337) ) ;
    buf_clk new_AGEMA_reg_buffer_4486 ( .C (clk), .D (new_AGEMA_signal_5987), .Q (new_AGEMA_signal_10338) ) ;
    buf_clk new_AGEMA_reg_buffer_4487 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_M24), .Q (new_AGEMA_signal_10339) ) ;
    buf_clk new_AGEMA_reg_buffer_4488 ( .C (clk), .D (new_AGEMA_signal_6083), .Q (new_AGEMA_signal_10340) ) ;
    buf_clk new_AGEMA_reg_buffer_4489 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_M21), .Q (new_AGEMA_signal_10341) ) ;
    buf_clk new_AGEMA_reg_buffer_4490 ( .C (clk), .D (new_AGEMA_signal_5911), .Q (new_AGEMA_signal_10342) ) ;
    buf_clk new_AGEMA_reg_buffer_4491 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_M23), .Q (new_AGEMA_signal_10343) ) ;
    buf_clk new_AGEMA_reg_buffer_4492 ( .C (clk), .D (new_AGEMA_signal_5989), .Q (new_AGEMA_signal_10344) ) ;
    buf_clk new_AGEMA_reg_buffer_4493 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_M27), .Q (new_AGEMA_signal_10345) ) ;
    buf_clk new_AGEMA_reg_buffer_4494 ( .C (clk), .D (new_AGEMA_signal_5991), .Q (new_AGEMA_signal_10346) ) ;
    buf_clk new_AGEMA_reg_buffer_4495 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_M24), .Q (new_AGEMA_signal_10347) ) ;
    buf_clk new_AGEMA_reg_buffer_4496 ( .C (clk), .D (new_AGEMA_signal_6088), .Q (new_AGEMA_signal_10348) ) ;
    buf_clk new_AGEMA_reg_buffer_4497 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21), .Q (new_AGEMA_signal_10349) ) ;
    buf_clk new_AGEMA_reg_buffer_4498 ( .C (clk), .D (new_AGEMA_signal_5835), .Q (new_AGEMA_signal_10350) ) ;
    buf_clk new_AGEMA_reg_buffer_4499 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23), .Q (new_AGEMA_signal_10351) ) ;
    buf_clk new_AGEMA_reg_buffer_4500 ( .C (clk), .D (new_AGEMA_signal_5913), .Q (new_AGEMA_signal_10352) ) ;
    buf_clk new_AGEMA_reg_buffer_4501 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27), .Q (new_AGEMA_signal_10353) ) ;
    buf_clk new_AGEMA_reg_buffer_4502 ( .C (clk), .D (new_AGEMA_signal_5915), .Q (new_AGEMA_signal_10354) ) ;
    buf_clk new_AGEMA_reg_buffer_4503 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24), .Q (new_AGEMA_signal_10355) ) ;
    buf_clk new_AGEMA_reg_buffer_4504 ( .C (clk), .D (new_AGEMA_signal_5993), .Q (new_AGEMA_signal_10356) ) ;
    buf_clk new_AGEMA_reg_buffer_4505 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21), .Q (new_AGEMA_signal_10357) ) ;
    buf_clk new_AGEMA_reg_buffer_4506 ( .C (clk), .D (new_AGEMA_signal_5839), .Q (new_AGEMA_signal_10358) ) ;
    buf_clk new_AGEMA_reg_buffer_4507 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23), .Q (new_AGEMA_signal_10359) ) ;
    buf_clk new_AGEMA_reg_buffer_4508 ( .C (clk), .D (new_AGEMA_signal_5917), .Q (new_AGEMA_signal_10360) ) ;
    buf_clk new_AGEMA_reg_buffer_4509 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27), .Q (new_AGEMA_signal_10361) ) ;
    buf_clk new_AGEMA_reg_buffer_4510 ( .C (clk), .D (new_AGEMA_signal_5919), .Q (new_AGEMA_signal_10362) ) ;
    buf_clk new_AGEMA_reg_buffer_4511 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24), .Q (new_AGEMA_signal_10363) ) ;
    buf_clk new_AGEMA_reg_buffer_4512 ( .C (clk), .D (new_AGEMA_signal_5998), .Q (new_AGEMA_signal_10364) ) ;
    buf_clk new_AGEMA_reg_buffer_4513 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21), .Q (new_AGEMA_signal_10365) ) ;
    buf_clk new_AGEMA_reg_buffer_4514 ( .C (clk), .D (new_AGEMA_signal_5843), .Q (new_AGEMA_signal_10366) ) ;
    buf_clk new_AGEMA_reg_buffer_4515 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23), .Q (new_AGEMA_signal_10367) ) ;
    buf_clk new_AGEMA_reg_buffer_4516 ( .C (clk), .D (new_AGEMA_signal_5921), .Q (new_AGEMA_signal_10368) ) ;
    buf_clk new_AGEMA_reg_buffer_4517 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27), .Q (new_AGEMA_signal_10369) ) ;
    buf_clk new_AGEMA_reg_buffer_4518 ( .C (clk), .D (new_AGEMA_signal_5923), .Q (new_AGEMA_signal_10370) ) ;
    buf_clk new_AGEMA_reg_buffer_4519 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24), .Q (new_AGEMA_signal_10371) ) ;
    buf_clk new_AGEMA_reg_buffer_4520 ( .C (clk), .D (new_AGEMA_signal_6003), .Q (new_AGEMA_signal_10372) ) ;
    buf_clk new_AGEMA_reg_buffer_4521 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21), .Q (new_AGEMA_signal_10373) ) ;
    buf_clk new_AGEMA_reg_buffer_4522 ( .C (clk), .D (new_AGEMA_signal_5847), .Q (new_AGEMA_signal_10374) ) ;
    buf_clk new_AGEMA_reg_buffer_4523 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23), .Q (new_AGEMA_signal_10375) ) ;
    buf_clk new_AGEMA_reg_buffer_4524 ( .C (clk), .D (new_AGEMA_signal_5925), .Q (new_AGEMA_signal_10376) ) ;
    buf_clk new_AGEMA_reg_buffer_4525 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27), .Q (new_AGEMA_signal_10377) ) ;
    buf_clk new_AGEMA_reg_buffer_4526 ( .C (clk), .D (new_AGEMA_signal_5927), .Q (new_AGEMA_signal_10378) ) ;
    buf_clk new_AGEMA_reg_buffer_4527 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24), .Q (new_AGEMA_signal_10379) ) ;
    buf_clk new_AGEMA_reg_buffer_4528 ( .C (clk), .D (new_AGEMA_signal_6008), .Q (new_AGEMA_signal_10380) ) ;
    buf_clk new_AGEMA_reg_buffer_4690 ( .C (clk), .D (new_AGEMA_signal_10541), .Q (new_AGEMA_signal_10542) ) ;
    buf_clk new_AGEMA_reg_buffer_4694 ( .C (clk), .D (new_AGEMA_signal_10545), .Q (new_AGEMA_signal_10546) ) ;
    buf_clk new_AGEMA_reg_buffer_4698 ( .C (clk), .D (new_AGEMA_signal_10549), .Q (new_AGEMA_signal_10550) ) ;
    buf_clk new_AGEMA_reg_buffer_4702 ( .C (clk), .D (new_AGEMA_signal_10553), .Q (new_AGEMA_signal_10554) ) ;
    buf_clk new_AGEMA_reg_buffer_4706 ( .C (clk), .D (new_AGEMA_signal_10557), .Q (new_AGEMA_signal_10558) ) ;
    buf_clk new_AGEMA_reg_buffer_4710 ( .C (clk), .D (new_AGEMA_signal_10561), .Q (new_AGEMA_signal_10562) ) ;
    buf_clk new_AGEMA_reg_buffer_4714 ( .C (clk), .D (new_AGEMA_signal_10565), .Q (new_AGEMA_signal_10566) ) ;
    buf_clk new_AGEMA_reg_buffer_4718 ( .C (clk), .D (new_AGEMA_signal_10569), .Q (new_AGEMA_signal_10570) ) ;
    buf_clk new_AGEMA_reg_buffer_4722 ( .C (clk), .D (new_AGEMA_signal_10573), .Q (new_AGEMA_signal_10574) ) ;
    buf_clk new_AGEMA_reg_buffer_4726 ( .C (clk), .D (new_AGEMA_signal_10577), .Q (new_AGEMA_signal_10578) ) ;
    buf_clk new_AGEMA_reg_buffer_4730 ( .C (clk), .D (new_AGEMA_signal_10581), .Q (new_AGEMA_signal_10582) ) ;
    buf_clk new_AGEMA_reg_buffer_4734 ( .C (clk), .D (new_AGEMA_signal_10585), .Q (new_AGEMA_signal_10586) ) ;
    buf_clk new_AGEMA_reg_buffer_4738 ( .C (clk), .D (new_AGEMA_signal_10589), .Q (new_AGEMA_signal_10590) ) ;
    buf_clk new_AGEMA_reg_buffer_4742 ( .C (clk), .D (new_AGEMA_signal_10593), .Q (new_AGEMA_signal_10594) ) ;
    buf_clk new_AGEMA_reg_buffer_4746 ( .C (clk), .D (new_AGEMA_signal_10597), .Q (new_AGEMA_signal_10598) ) ;
    buf_clk new_AGEMA_reg_buffer_4750 ( .C (clk), .D (new_AGEMA_signal_10601), .Q (new_AGEMA_signal_10602) ) ;
    buf_clk new_AGEMA_reg_buffer_4754 ( .C (clk), .D (new_AGEMA_signal_10605), .Q (new_AGEMA_signal_10606) ) ;
    buf_clk new_AGEMA_reg_buffer_4758 ( .C (clk), .D (new_AGEMA_signal_10609), .Q (new_AGEMA_signal_10610) ) ;
    buf_clk new_AGEMA_reg_buffer_4762 ( .C (clk), .D (new_AGEMA_signal_10613), .Q (new_AGEMA_signal_10614) ) ;
    buf_clk new_AGEMA_reg_buffer_4766 ( .C (clk), .D (new_AGEMA_signal_10617), .Q (new_AGEMA_signal_10618) ) ;
    buf_clk new_AGEMA_reg_buffer_4770 ( .C (clk), .D (new_AGEMA_signal_10621), .Q (new_AGEMA_signal_10622) ) ;
    buf_clk new_AGEMA_reg_buffer_4774 ( .C (clk), .D (new_AGEMA_signal_10625), .Q (new_AGEMA_signal_10626) ) ;
    buf_clk new_AGEMA_reg_buffer_4778 ( .C (clk), .D (new_AGEMA_signal_10629), .Q (new_AGEMA_signal_10630) ) ;
    buf_clk new_AGEMA_reg_buffer_4782 ( .C (clk), .D (new_AGEMA_signal_10633), .Q (new_AGEMA_signal_10634) ) ;
    buf_clk new_AGEMA_reg_buffer_4786 ( .C (clk), .D (new_AGEMA_signal_10637), .Q (new_AGEMA_signal_10638) ) ;
    buf_clk new_AGEMA_reg_buffer_4790 ( .C (clk), .D (new_AGEMA_signal_10641), .Q (new_AGEMA_signal_10642) ) ;
    buf_clk new_AGEMA_reg_buffer_4794 ( .C (clk), .D (new_AGEMA_signal_10645), .Q (new_AGEMA_signal_10646) ) ;
    buf_clk new_AGEMA_reg_buffer_4798 ( .C (clk), .D (new_AGEMA_signal_10649), .Q (new_AGEMA_signal_10650) ) ;
    buf_clk new_AGEMA_reg_buffer_4802 ( .C (clk), .D (new_AGEMA_signal_10653), .Q (new_AGEMA_signal_10654) ) ;
    buf_clk new_AGEMA_reg_buffer_4806 ( .C (clk), .D (new_AGEMA_signal_10657), .Q (new_AGEMA_signal_10658) ) ;
    buf_clk new_AGEMA_reg_buffer_4810 ( .C (clk), .D (new_AGEMA_signal_10661), .Q (new_AGEMA_signal_10662) ) ;
    buf_clk new_AGEMA_reg_buffer_4814 ( .C (clk), .D (new_AGEMA_signal_10665), .Q (new_AGEMA_signal_10666) ) ;
    buf_clk new_AGEMA_reg_buffer_4818 ( .C (clk), .D (new_AGEMA_signal_10669), .Q (new_AGEMA_signal_10670) ) ;
    buf_clk new_AGEMA_reg_buffer_4822 ( .C (clk), .D (new_AGEMA_signal_10673), .Q (new_AGEMA_signal_10674) ) ;
    buf_clk new_AGEMA_reg_buffer_4826 ( .C (clk), .D (new_AGEMA_signal_10677), .Q (new_AGEMA_signal_10678) ) ;
    buf_clk new_AGEMA_reg_buffer_4830 ( .C (clk), .D (new_AGEMA_signal_10681), .Q (new_AGEMA_signal_10682) ) ;
    buf_clk new_AGEMA_reg_buffer_4834 ( .C (clk), .D (new_AGEMA_signal_10685), .Q (new_AGEMA_signal_10686) ) ;
    buf_clk new_AGEMA_reg_buffer_4838 ( .C (clk), .D (new_AGEMA_signal_10689), .Q (new_AGEMA_signal_10690) ) ;
    buf_clk new_AGEMA_reg_buffer_4842 ( .C (clk), .D (new_AGEMA_signal_10693), .Q (new_AGEMA_signal_10694) ) ;
    buf_clk new_AGEMA_reg_buffer_4846 ( .C (clk), .D (new_AGEMA_signal_10697), .Q (new_AGEMA_signal_10698) ) ;
    buf_clk new_AGEMA_reg_buffer_4850 ( .C (clk), .D (new_AGEMA_signal_10701), .Q (new_AGEMA_signal_10702) ) ;
    buf_clk new_AGEMA_reg_buffer_4854 ( .C (clk), .D (new_AGEMA_signal_10705), .Q (new_AGEMA_signal_10706) ) ;
    buf_clk new_AGEMA_reg_buffer_4858 ( .C (clk), .D (new_AGEMA_signal_10709), .Q (new_AGEMA_signal_10710) ) ;
    buf_clk new_AGEMA_reg_buffer_4862 ( .C (clk), .D (new_AGEMA_signal_10713), .Q (new_AGEMA_signal_10714) ) ;
    buf_clk new_AGEMA_reg_buffer_4866 ( .C (clk), .D (new_AGEMA_signal_10717), .Q (new_AGEMA_signal_10718) ) ;
    buf_clk new_AGEMA_reg_buffer_4870 ( .C (clk), .D (new_AGEMA_signal_10721), .Q (new_AGEMA_signal_10722) ) ;
    buf_clk new_AGEMA_reg_buffer_4874 ( .C (clk), .D (new_AGEMA_signal_10725), .Q (new_AGEMA_signal_10726) ) ;
    buf_clk new_AGEMA_reg_buffer_4878 ( .C (clk), .D (new_AGEMA_signal_10729), .Q (new_AGEMA_signal_10730) ) ;
    buf_clk new_AGEMA_reg_buffer_4882 ( .C (clk), .D (new_AGEMA_signal_10733), .Q (new_AGEMA_signal_10734) ) ;
    buf_clk new_AGEMA_reg_buffer_4886 ( .C (clk), .D (new_AGEMA_signal_10737), .Q (new_AGEMA_signal_10738) ) ;
    buf_clk new_AGEMA_reg_buffer_4890 ( .C (clk), .D (new_AGEMA_signal_10741), .Q (new_AGEMA_signal_10742) ) ;
    buf_clk new_AGEMA_reg_buffer_4894 ( .C (clk), .D (new_AGEMA_signal_10745), .Q (new_AGEMA_signal_10746) ) ;
    buf_clk new_AGEMA_reg_buffer_4898 ( .C (clk), .D (new_AGEMA_signal_10749), .Q (new_AGEMA_signal_10750) ) ;
    buf_clk new_AGEMA_reg_buffer_4902 ( .C (clk), .D (new_AGEMA_signal_10753), .Q (new_AGEMA_signal_10754) ) ;
    buf_clk new_AGEMA_reg_buffer_4906 ( .C (clk), .D (new_AGEMA_signal_10757), .Q (new_AGEMA_signal_10758) ) ;
    buf_clk new_AGEMA_reg_buffer_4910 ( .C (clk), .D (new_AGEMA_signal_10761), .Q (new_AGEMA_signal_10762) ) ;
    buf_clk new_AGEMA_reg_buffer_4914 ( .C (clk), .D (new_AGEMA_signal_10765), .Q (new_AGEMA_signal_10766) ) ;
    buf_clk new_AGEMA_reg_buffer_4918 ( .C (clk), .D (new_AGEMA_signal_10769), .Q (new_AGEMA_signal_10770) ) ;
    buf_clk new_AGEMA_reg_buffer_4922 ( .C (clk), .D (new_AGEMA_signal_10773), .Q (new_AGEMA_signal_10774) ) ;
    buf_clk new_AGEMA_reg_buffer_4926 ( .C (clk), .D (new_AGEMA_signal_10777), .Q (new_AGEMA_signal_10778) ) ;
    buf_clk new_AGEMA_reg_buffer_4930 ( .C (clk), .D (new_AGEMA_signal_10781), .Q (new_AGEMA_signal_10782) ) ;
    buf_clk new_AGEMA_reg_buffer_4934 ( .C (clk), .D (new_AGEMA_signal_10785), .Q (new_AGEMA_signal_10786) ) ;
    buf_clk new_AGEMA_reg_buffer_4938 ( .C (clk), .D (new_AGEMA_signal_10789), .Q (new_AGEMA_signal_10790) ) ;
    buf_clk new_AGEMA_reg_buffer_4942 ( .C (clk), .D (new_AGEMA_signal_10793), .Q (new_AGEMA_signal_10794) ) ;
    buf_clk new_AGEMA_reg_buffer_4946 ( .C (clk), .D (new_AGEMA_signal_10797), .Q (new_AGEMA_signal_10798) ) ;
    buf_clk new_AGEMA_reg_buffer_4950 ( .C (clk), .D (new_AGEMA_signal_10801), .Q (new_AGEMA_signal_10802) ) ;
    buf_clk new_AGEMA_reg_buffer_4954 ( .C (clk), .D (new_AGEMA_signal_10805), .Q (new_AGEMA_signal_10806) ) ;
    buf_clk new_AGEMA_reg_buffer_4958 ( .C (clk), .D (new_AGEMA_signal_10809), .Q (new_AGEMA_signal_10810) ) ;
    buf_clk new_AGEMA_reg_buffer_4962 ( .C (clk), .D (new_AGEMA_signal_10813), .Q (new_AGEMA_signal_10814) ) ;
    buf_clk new_AGEMA_reg_buffer_4966 ( .C (clk), .D (new_AGEMA_signal_10817), .Q (new_AGEMA_signal_10818) ) ;
    buf_clk new_AGEMA_reg_buffer_4970 ( .C (clk), .D (new_AGEMA_signal_10821), .Q (new_AGEMA_signal_10822) ) ;
    buf_clk new_AGEMA_reg_buffer_4974 ( .C (clk), .D (new_AGEMA_signal_10825), .Q (new_AGEMA_signal_10826) ) ;
    buf_clk new_AGEMA_reg_buffer_4978 ( .C (clk), .D (new_AGEMA_signal_10829), .Q (new_AGEMA_signal_10830) ) ;
    buf_clk new_AGEMA_reg_buffer_4982 ( .C (clk), .D (new_AGEMA_signal_10833), .Q (new_AGEMA_signal_10834) ) ;
    buf_clk new_AGEMA_reg_buffer_4986 ( .C (clk), .D (new_AGEMA_signal_10837), .Q (new_AGEMA_signal_10838) ) ;
    buf_clk new_AGEMA_reg_buffer_4990 ( .C (clk), .D (new_AGEMA_signal_10841), .Q (new_AGEMA_signal_10842) ) ;
    buf_clk new_AGEMA_reg_buffer_4994 ( .C (clk), .D (new_AGEMA_signal_10845), .Q (new_AGEMA_signal_10846) ) ;
    buf_clk new_AGEMA_reg_buffer_4998 ( .C (clk), .D (new_AGEMA_signal_10849), .Q (new_AGEMA_signal_10850) ) ;
    buf_clk new_AGEMA_reg_buffer_5002 ( .C (clk), .D (new_AGEMA_signal_10853), .Q (new_AGEMA_signal_10854) ) ;
    buf_clk new_AGEMA_reg_buffer_5006 ( .C (clk), .D (new_AGEMA_signal_10857), .Q (new_AGEMA_signal_10858) ) ;
    buf_clk new_AGEMA_reg_buffer_5010 ( .C (clk), .D (new_AGEMA_signal_10861), .Q (new_AGEMA_signal_10862) ) ;
    buf_clk new_AGEMA_reg_buffer_5014 ( .C (clk), .D (new_AGEMA_signal_10865), .Q (new_AGEMA_signal_10866) ) ;
    buf_clk new_AGEMA_reg_buffer_5018 ( .C (clk), .D (new_AGEMA_signal_10869), .Q (new_AGEMA_signal_10870) ) ;
    buf_clk new_AGEMA_reg_buffer_5022 ( .C (clk), .D (new_AGEMA_signal_10873), .Q (new_AGEMA_signal_10874) ) ;
    buf_clk new_AGEMA_reg_buffer_5026 ( .C (clk), .D (new_AGEMA_signal_10877), .Q (new_AGEMA_signal_10878) ) ;
    buf_clk new_AGEMA_reg_buffer_5030 ( .C (clk), .D (new_AGEMA_signal_10881), .Q (new_AGEMA_signal_10882) ) ;
    buf_clk new_AGEMA_reg_buffer_5034 ( .C (clk), .D (new_AGEMA_signal_10885), .Q (new_AGEMA_signal_10886) ) ;
    buf_clk new_AGEMA_reg_buffer_5038 ( .C (clk), .D (new_AGEMA_signal_10889), .Q (new_AGEMA_signal_10890) ) ;
    buf_clk new_AGEMA_reg_buffer_5042 ( .C (clk), .D (new_AGEMA_signal_10893), .Q (new_AGEMA_signal_10894) ) ;
    buf_clk new_AGEMA_reg_buffer_5046 ( .C (clk), .D (new_AGEMA_signal_10897), .Q (new_AGEMA_signal_10898) ) ;
    buf_clk new_AGEMA_reg_buffer_5050 ( .C (clk), .D (new_AGEMA_signal_10901), .Q (new_AGEMA_signal_10902) ) ;
    buf_clk new_AGEMA_reg_buffer_5054 ( .C (clk), .D (new_AGEMA_signal_10905), .Q (new_AGEMA_signal_10906) ) ;
    buf_clk new_AGEMA_reg_buffer_5058 ( .C (clk), .D (new_AGEMA_signal_10909), .Q (new_AGEMA_signal_10910) ) ;
    buf_clk new_AGEMA_reg_buffer_5062 ( .C (clk), .D (new_AGEMA_signal_10913), .Q (new_AGEMA_signal_10914) ) ;
    buf_clk new_AGEMA_reg_buffer_5066 ( .C (clk), .D (new_AGEMA_signal_10917), .Q (new_AGEMA_signal_10918) ) ;
    buf_clk new_AGEMA_reg_buffer_5070 ( .C (clk), .D (new_AGEMA_signal_10921), .Q (new_AGEMA_signal_10922) ) ;
    buf_clk new_AGEMA_reg_buffer_5074 ( .C (clk), .D (new_AGEMA_signal_10925), .Q (new_AGEMA_signal_10926) ) ;
    buf_clk new_AGEMA_reg_buffer_5078 ( .C (clk), .D (new_AGEMA_signal_10929), .Q (new_AGEMA_signal_10930) ) ;
    buf_clk new_AGEMA_reg_buffer_5082 ( .C (clk), .D (new_AGEMA_signal_10933), .Q (new_AGEMA_signal_10934) ) ;
    buf_clk new_AGEMA_reg_buffer_5086 ( .C (clk), .D (new_AGEMA_signal_10937), .Q (new_AGEMA_signal_10938) ) ;
    buf_clk new_AGEMA_reg_buffer_5090 ( .C (clk), .D (new_AGEMA_signal_10941), .Q (new_AGEMA_signal_10942) ) ;
    buf_clk new_AGEMA_reg_buffer_5094 ( .C (clk), .D (new_AGEMA_signal_10945), .Q (new_AGEMA_signal_10946) ) ;
    buf_clk new_AGEMA_reg_buffer_5098 ( .C (clk), .D (new_AGEMA_signal_10949), .Q (new_AGEMA_signal_10950) ) ;
    buf_clk new_AGEMA_reg_buffer_5102 ( .C (clk), .D (new_AGEMA_signal_10953), .Q (new_AGEMA_signal_10954) ) ;
    buf_clk new_AGEMA_reg_buffer_5106 ( .C (clk), .D (new_AGEMA_signal_10957), .Q (new_AGEMA_signal_10958) ) ;
    buf_clk new_AGEMA_reg_buffer_5110 ( .C (clk), .D (new_AGEMA_signal_10961), .Q (new_AGEMA_signal_10962) ) ;
    buf_clk new_AGEMA_reg_buffer_5114 ( .C (clk), .D (new_AGEMA_signal_10965), .Q (new_AGEMA_signal_10966) ) ;
    buf_clk new_AGEMA_reg_buffer_5118 ( .C (clk), .D (new_AGEMA_signal_10969), .Q (new_AGEMA_signal_10970) ) ;
    buf_clk new_AGEMA_reg_buffer_5122 ( .C (clk), .D (new_AGEMA_signal_10973), .Q (new_AGEMA_signal_10974) ) ;
    buf_clk new_AGEMA_reg_buffer_5126 ( .C (clk), .D (new_AGEMA_signal_10977), .Q (new_AGEMA_signal_10978) ) ;
    buf_clk new_AGEMA_reg_buffer_5130 ( .C (clk), .D (new_AGEMA_signal_10981), .Q (new_AGEMA_signal_10982) ) ;
    buf_clk new_AGEMA_reg_buffer_5134 ( .C (clk), .D (new_AGEMA_signal_10985), .Q (new_AGEMA_signal_10986) ) ;
    buf_clk new_AGEMA_reg_buffer_5138 ( .C (clk), .D (new_AGEMA_signal_10989), .Q (new_AGEMA_signal_10990) ) ;
    buf_clk new_AGEMA_reg_buffer_5142 ( .C (clk), .D (new_AGEMA_signal_10993), .Q (new_AGEMA_signal_10994) ) ;
    buf_clk new_AGEMA_reg_buffer_5146 ( .C (clk), .D (new_AGEMA_signal_10997), .Q (new_AGEMA_signal_10998) ) ;
    buf_clk new_AGEMA_reg_buffer_5150 ( .C (clk), .D (new_AGEMA_signal_11001), .Q (new_AGEMA_signal_11002) ) ;
    buf_clk new_AGEMA_reg_buffer_5154 ( .C (clk), .D (new_AGEMA_signal_11005), .Q (new_AGEMA_signal_11006) ) ;
    buf_clk new_AGEMA_reg_buffer_5158 ( .C (clk), .D (new_AGEMA_signal_11009), .Q (new_AGEMA_signal_11010) ) ;
    buf_clk new_AGEMA_reg_buffer_5162 ( .C (clk), .D (new_AGEMA_signal_11013), .Q (new_AGEMA_signal_11014) ) ;
    buf_clk new_AGEMA_reg_buffer_5166 ( .C (clk), .D (new_AGEMA_signal_11017), .Q (new_AGEMA_signal_11018) ) ;
    buf_clk new_AGEMA_reg_buffer_5170 ( .C (clk), .D (new_AGEMA_signal_11021), .Q (new_AGEMA_signal_11022) ) ;
    buf_clk new_AGEMA_reg_buffer_5174 ( .C (clk), .D (new_AGEMA_signal_11025), .Q (new_AGEMA_signal_11026) ) ;
    buf_clk new_AGEMA_reg_buffer_5178 ( .C (clk), .D (new_AGEMA_signal_11029), .Q (new_AGEMA_signal_11030) ) ;
    buf_clk new_AGEMA_reg_buffer_5182 ( .C (clk), .D (new_AGEMA_signal_11033), .Q (new_AGEMA_signal_11034) ) ;
    buf_clk new_AGEMA_reg_buffer_5186 ( .C (clk), .D (new_AGEMA_signal_11037), .Q (new_AGEMA_signal_11038) ) ;
    buf_clk new_AGEMA_reg_buffer_5190 ( .C (clk), .D (new_AGEMA_signal_11041), .Q (new_AGEMA_signal_11042) ) ;
    buf_clk new_AGEMA_reg_buffer_5194 ( .C (clk), .D (new_AGEMA_signal_11045), .Q (new_AGEMA_signal_11046) ) ;
    buf_clk new_AGEMA_reg_buffer_5198 ( .C (clk), .D (new_AGEMA_signal_11049), .Q (new_AGEMA_signal_11050) ) ;
    buf_clk new_AGEMA_reg_buffer_5202 ( .C (clk), .D (new_AGEMA_signal_11053), .Q (new_AGEMA_signal_11054) ) ;
    buf_clk new_AGEMA_reg_buffer_5206 ( .C (clk), .D (new_AGEMA_signal_11057), .Q (new_AGEMA_signal_11058) ) ;
    buf_clk new_AGEMA_reg_buffer_5210 ( .C (clk), .D (new_AGEMA_signal_11061), .Q (new_AGEMA_signal_11062) ) ;
    buf_clk new_AGEMA_reg_buffer_5214 ( .C (clk), .D (new_AGEMA_signal_11065), .Q (new_AGEMA_signal_11066) ) ;
    buf_clk new_AGEMA_reg_buffer_5218 ( .C (clk), .D (new_AGEMA_signal_11069), .Q (new_AGEMA_signal_11070) ) ;
    buf_clk new_AGEMA_reg_buffer_5222 ( .C (clk), .D (new_AGEMA_signal_11073), .Q (new_AGEMA_signal_11074) ) ;
    buf_clk new_AGEMA_reg_buffer_5226 ( .C (clk), .D (new_AGEMA_signal_11077), .Q (new_AGEMA_signal_11078) ) ;
    buf_clk new_AGEMA_reg_buffer_5230 ( .C (clk), .D (new_AGEMA_signal_11081), .Q (new_AGEMA_signal_11082) ) ;
    buf_clk new_AGEMA_reg_buffer_5234 ( .C (clk), .D (new_AGEMA_signal_11085), .Q (new_AGEMA_signal_11086) ) ;
    buf_clk new_AGEMA_reg_buffer_5238 ( .C (clk), .D (new_AGEMA_signal_11089), .Q (new_AGEMA_signal_11090) ) ;
    buf_clk new_AGEMA_reg_buffer_5242 ( .C (clk), .D (new_AGEMA_signal_11093), .Q (new_AGEMA_signal_11094) ) ;
    buf_clk new_AGEMA_reg_buffer_5246 ( .C (clk), .D (new_AGEMA_signal_11097), .Q (new_AGEMA_signal_11098) ) ;
    buf_clk new_AGEMA_reg_buffer_5250 ( .C (clk), .D (new_AGEMA_signal_11101), .Q (new_AGEMA_signal_11102) ) ;
    buf_clk new_AGEMA_reg_buffer_5254 ( .C (clk), .D (new_AGEMA_signal_11105), .Q (new_AGEMA_signal_11106) ) ;
    buf_clk new_AGEMA_reg_buffer_5258 ( .C (clk), .D (new_AGEMA_signal_11109), .Q (new_AGEMA_signal_11110) ) ;
    buf_clk new_AGEMA_reg_buffer_5262 ( .C (clk), .D (new_AGEMA_signal_11113), .Q (new_AGEMA_signal_11114) ) ;
    buf_clk new_AGEMA_reg_buffer_5266 ( .C (clk), .D (new_AGEMA_signal_11117), .Q (new_AGEMA_signal_11118) ) ;
    buf_clk new_AGEMA_reg_buffer_5270 ( .C (clk), .D (new_AGEMA_signal_11121), .Q (new_AGEMA_signal_11122) ) ;
    buf_clk new_AGEMA_reg_buffer_5274 ( .C (clk), .D (new_AGEMA_signal_11125), .Q (new_AGEMA_signal_11126) ) ;
    buf_clk new_AGEMA_reg_buffer_5278 ( .C (clk), .D (new_AGEMA_signal_11129), .Q (new_AGEMA_signal_11130) ) ;
    buf_clk new_AGEMA_reg_buffer_5282 ( .C (clk), .D (new_AGEMA_signal_11133), .Q (new_AGEMA_signal_11134) ) ;
    buf_clk new_AGEMA_reg_buffer_5286 ( .C (clk), .D (new_AGEMA_signal_11137), .Q (new_AGEMA_signal_11138) ) ;
    buf_clk new_AGEMA_reg_buffer_5290 ( .C (clk), .D (new_AGEMA_signal_11141), .Q (new_AGEMA_signal_11142) ) ;
    buf_clk new_AGEMA_reg_buffer_5294 ( .C (clk), .D (new_AGEMA_signal_11145), .Q (new_AGEMA_signal_11146) ) ;
    buf_clk new_AGEMA_reg_buffer_5298 ( .C (clk), .D (new_AGEMA_signal_11149), .Q (new_AGEMA_signal_11150) ) ;
    buf_clk new_AGEMA_reg_buffer_5302 ( .C (clk), .D (new_AGEMA_signal_11153), .Q (new_AGEMA_signal_11154) ) ;
    buf_clk new_AGEMA_reg_buffer_5306 ( .C (clk), .D (new_AGEMA_signal_11157), .Q (new_AGEMA_signal_11158) ) ;
    buf_clk new_AGEMA_reg_buffer_5310 ( .C (clk), .D (new_AGEMA_signal_11161), .Q (new_AGEMA_signal_11162) ) ;
    buf_clk new_AGEMA_reg_buffer_5314 ( .C (clk), .D (new_AGEMA_signal_11165), .Q (new_AGEMA_signal_11166) ) ;
    buf_clk new_AGEMA_reg_buffer_5318 ( .C (clk), .D (new_AGEMA_signal_11169), .Q (new_AGEMA_signal_11170) ) ;
    buf_clk new_AGEMA_reg_buffer_5322 ( .C (clk), .D (new_AGEMA_signal_11173), .Q (new_AGEMA_signal_11174) ) ;
    buf_clk new_AGEMA_reg_buffer_5326 ( .C (clk), .D (new_AGEMA_signal_11177), .Q (new_AGEMA_signal_11178) ) ;
    buf_clk new_AGEMA_reg_buffer_5330 ( .C (clk), .D (new_AGEMA_signal_11181), .Q (new_AGEMA_signal_11182) ) ;
    buf_clk new_AGEMA_reg_buffer_5334 ( .C (clk), .D (new_AGEMA_signal_11185), .Q (new_AGEMA_signal_11186) ) ;
    buf_clk new_AGEMA_reg_buffer_5338 ( .C (clk), .D (new_AGEMA_signal_11189), .Q (new_AGEMA_signal_11190) ) ;
    buf_clk new_AGEMA_reg_buffer_5342 ( .C (clk), .D (new_AGEMA_signal_11193), .Q (new_AGEMA_signal_11194) ) ;
    buf_clk new_AGEMA_reg_buffer_5346 ( .C (clk), .D (new_AGEMA_signal_11197), .Q (new_AGEMA_signal_11198) ) ;
    buf_clk new_AGEMA_reg_buffer_5350 ( .C (clk), .D (new_AGEMA_signal_11201), .Q (new_AGEMA_signal_11202) ) ;
    buf_clk new_AGEMA_reg_buffer_5354 ( .C (clk), .D (new_AGEMA_signal_11205), .Q (new_AGEMA_signal_11206) ) ;
    buf_clk new_AGEMA_reg_buffer_5358 ( .C (clk), .D (new_AGEMA_signal_11209), .Q (new_AGEMA_signal_11210) ) ;
    buf_clk new_AGEMA_reg_buffer_5362 ( .C (clk), .D (new_AGEMA_signal_11213), .Q (new_AGEMA_signal_11214) ) ;
    buf_clk new_AGEMA_reg_buffer_5366 ( .C (clk), .D (new_AGEMA_signal_11217), .Q (new_AGEMA_signal_11218) ) ;
    buf_clk new_AGEMA_reg_buffer_5370 ( .C (clk), .D (new_AGEMA_signal_11221), .Q (new_AGEMA_signal_11222) ) ;
    buf_clk new_AGEMA_reg_buffer_5374 ( .C (clk), .D (new_AGEMA_signal_11225), .Q (new_AGEMA_signal_11226) ) ;
    buf_clk new_AGEMA_reg_buffer_5378 ( .C (clk), .D (new_AGEMA_signal_11229), .Q (new_AGEMA_signal_11230) ) ;
    buf_clk new_AGEMA_reg_buffer_5382 ( .C (clk), .D (new_AGEMA_signal_11233), .Q (new_AGEMA_signal_11234) ) ;
    buf_clk new_AGEMA_reg_buffer_5386 ( .C (clk), .D (new_AGEMA_signal_11237), .Q (new_AGEMA_signal_11238) ) ;
    buf_clk new_AGEMA_reg_buffer_5390 ( .C (clk), .D (new_AGEMA_signal_11241), .Q (new_AGEMA_signal_11242) ) ;
    buf_clk new_AGEMA_reg_buffer_5394 ( .C (clk), .D (new_AGEMA_signal_11245), .Q (new_AGEMA_signal_11246) ) ;
    buf_clk new_AGEMA_reg_buffer_5398 ( .C (clk), .D (new_AGEMA_signal_11249), .Q (new_AGEMA_signal_11250) ) ;
    buf_clk new_AGEMA_reg_buffer_5402 ( .C (clk), .D (new_AGEMA_signal_11253), .Q (new_AGEMA_signal_11254) ) ;
    buf_clk new_AGEMA_reg_buffer_5406 ( .C (clk), .D (new_AGEMA_signal_11257), .Q (new_AGEMA_signal_11258) ) ;
    buf_clk new_AGEMA_reg_buffer_5410 ( .C (clk), .D (new_AGEMA_signal_11261), .Q (new_AGEMA_signal_11262) ) ;
    buf_clk new_AGEMA_reg_buffer_5414 ( .C (clk), .D (new_AGEMA_signal_11265), .Q (new_AGEMA_signal_11266) ) ;
    buf_clk new_AGEMA_reg_buffer_5418 ( .C (clk), .D (new_AGEMA_signal_11269), .Q (new_AGEMA_signal_11270) ) ;
    buf_clk new_AGEMA_reg_buffer_5422 ( .C (clk), .D (new_AGEMA_signal_11273), .Q (new_AGEMA_signal_11274) ) ;
    buf_clk new_AGEMA_reg_buffer_5426 ( .C (clk), .D (new_AGEMA_signal_11277), .Q (new_AGEMA_signal_11278) ) ;
    buf_clk new_AGEMA_reg_buffer_5430 ( .C (clk), .D (new_AGEMA_signal_11281), .Q (new_AGEMA_signal_11282) ) ;
    buf_clk new_AGEMA_reg_buffer_5434 ( .C (clk), .D (new_AGEMA_signal_11285), .Q (new_AGEMA_signal_11286) ) ;
    buf_clk new_AGEMA_reg_buffer_5438 ( .C (clk), .D (new_AGEMA_signal_11289), .Q (new_AGEMA_signal_11290) ) ;
    buf_clk new_AGEMA_reg_buffer_5442 ( .C (clk), .D (new_AGEMA_signal_11293), .Q (new_AGEMA_signal_11294) ) ;
    buf_clk new_AGEMA_reg_buffer_5446 ( .C (clk), .D (new_AGEMA_signal_11297), .Q (new_AGEMA_signal_11298) ) ;
    buf_clk new_AGEMA_reg_buffer_5450 ( .C (clk), .D (new_AGEMA_signal_11301), .Q (new_AGEMA_signal_11302) ) ;
    buf_clk new_AGEMA_reg_buffer_5454 ( .C (clk), .D (new_AGEMA_signal_11305), .Q (new_AGEMA_signal_11306) ) ;
    buf_clk new_AGEMA_reg_buffer_5458 ( .C (clk), .D (new_AGEMA_signal_11309), .Q (new_AGEMA_signal_11310) ) ;
    buf_clk new_AGEMA_reg_buffer_5462 ( .C (clk), .D (new_AGEMA_signal_11313), .Q (new_AGEMA_signal_11314) ) ;
    buf_clk new_AGEMA_reg_buffer_5466 ( .C (clk), .D (new_AGEMA_signal_11317), .Q (new_AGEMA_signal_11318) ) ;
    buf_clk new_AGEMA_reg_buffer_5470 ( .C (clk), .D (new_AGEMA_signal_11321), .Q (new_AGEMA_signal_11322) ) ;
    buf_clk new_AGEMA_reg_buffer_5474 ( .C (clk), .D (new_AGEMA_signal_11325), .Q (new_AGEMA_signal_11326) ) ;
    buf_clk new_AGEMA_reg_buffer_5478 ( .C (clk), .D (new_AGEMA_signal_11329), .Q (new_AGEMA_signal_11330) ) ;
    buf_clk new_AGEMA_reg_buffer_5482 ( .C (clk), .D (new_AGEMA_signal_11333), .Q (new_AGEMA_signal_11334) ) ;
    buf_clk new_AGEMA_reg_buffer_5486 ( .C (clk), .D (new_AGEMA_signal_11337), .Q (new_AGEMA_signal_11338) ) ;
    buf_clk new_AGEMA_reg_buffer_5490 ( .C (clk), .D (new_AGEMA_signal_11341), .Q (new_AGEMA_signal_11342) ) ;
    buf_clk new_AGEMA_reg_buffer_5494 ( .C (clk), .D (new_AGEMA_signal_11345), .Q (new_AGEMA_signal_11346) ) ;
    buf_clk new_AGEMA_reg_buffer_5498 ( .C (clk), .D (new_AGEMA_signal_11349), .Q (new_AGEMA_signal_11350) ) ;
    buf_clk new_AGEMA_reg_buffer_5502 ( .C (clk), .D (new_AGEMA_signal_11353), .Q (new_AGEMA_signal_11354) ) ;
    buf_clk new_AGEMA_reg_buffer_5506 ( .C (clk), .D (new_AGEMA_signal_11357), .Q (new_AGEMA_signal_11358) ) ;
    buf_clk new_AGEMA_reg_buffer_5510 ( .C (clk), .D (new_AGEMA_signal_11361), .Q (new_AGEMA_signal_11362) ) ;
    buf_clk new_AGEMA_reg_buffer_5514 ( .C (clk), .D (new_AGEMA_signal_11365), .Q (new_AGEMA_signal_11366) ) ;
    buf_clk new_AGEMA_reg_buffer_5518 ( .C (clk), .D (new_AGEMA_signal_11369), .Q (new_AGEMA_signal_11370) ) ;
    buf_clk new_AGEMA_reg_buffer_5522 ( .C (clk), .D (new_AGEMA_signal_11373), .Q (new_AGEMA_signal_11374) ) ;
    buf_clk new_AGEMA_reg_buffer_5526 ( .C (clk), .D (new_AGEMA_signal_11377), .Q (new_AGEMA_signal_11378) ) ;
    buf_clk new_AGEMA_reg_buffer_5530 ( .C (clk), .D (new_AGEMA_signal_11381), .Q (new_AGEMA_signal_11382) ) ;
    buf_clk new_AGEMA_reg_buffer_5534 ( .C (clk), .D (new_AGEMA_signal_11385), .Q (new_AGEMA_signal_11386) ) ;
    buf_clk new_AGEMA_reg_buffer_5538 ( .C (clk), .D (new_AGEMA_signal_11389), .Q (new_AGEMA_signal_11390) ) ;
    buf_clk new_AGEMA_reg_buffer_5542 ( .C (clk), .D (new_AGEMA_signal_11393), .Q (new_AGEMA_signal_11394) ) ;
    buf_clk new_AGEMA_reg_buffer_5546 ( .C (clk), .D (new_AGEMA_signal_11397), .Q (new_AGEMA_signal_11398) ) ;
    buf_clk new_AGEMA_reg_buffer_5550 ( .C (clk), .D (new_AGEMA_signal_11401), .Q (new_AGEMA_signal_11402) ) ;
    buf_clk new_AGEMA_reg_buffer_5554 ( .C (clk), .D (new_AGEMA_signal_11405), .Q (new_AGEMA_signal_11406) ) ;
    buf_clk new_AGEMA_reg_buffer_5558 ( .C (clk), .D (new_AGEMA_signal_11409), .Q (new_AGEMA_signal_11410) ) ;
    buf_clk new_AGEMA_reg_buffer_5562 ( .C (clk), .D (new_AGEMA_signal_11413), .Q (new_AGEMA_signal_11414) ) ;
    buf_clk new_AGEMA_reg_buffer_5566 ( .C (clk), .D (new_AGEMA_signal_11417), .Q (new_AGEMA_signal_11418) ) ;
    buf_clk new_AGEMA_reg_buffer_5570 ( .C (clk), .D (new_AGEMA_signal_11421), .Q (new_AGEMA_signal_11422) ) ;
    buf_clk new_AGEMA_reg_buffer_5574 ( .C (clk), .D (new_AGEMA_signal_11425), .Q (new_AGEMA_signal_11426) ) ;
    buf_clk new_AGEMA_reg_buffer_5578 ( .C (clk), .D (new_AGEMA_signal_11429), .Q (new_AGEMA_signal_11430) ) ;
    buf_clk new_AGEMA_reg_buffer_5582 ( .C (clk), .D (new_AGEMA_signal_11433), .Q (new_AGEMA_signal_11434) ) ;
    buf_clk new_AGEMA_reg_buffer_5586 ( .C (clk), .D (new_AGEMA_signal_11437), .Q (new_AGEMA_signal_11438) ) ;
    buf_clk new_AGEMA_reg_buffer_5590 ( .C (clk), .D (new_AGEMA_signal_11441), .Q (new_AGEMA_signal_11442) ) ;
    buf_clk new_AGEMA_reg_buffer_5594 ( .C (clk), .D (new_AGEMA_signal_11445), .Q (new_AGEMA_signal_11446) ) ;
    buf_clk new_AGEMA_reg_buffer_5598 ( .C (clk), .D (new_AGEMA_signal_11449), .Q (new_AGEMA_signal_11450) ) ;
    buf_clk new_AGEMA_reg_buffer_5602 ( .C (clk), .D (new_AGEMA_signal_11453), .Q (new_AGEMA_signal_11454) ) ;
    buf_clk new_AGEMA_reg_buffer_5606 ( .C (clk), .D (new_AGEMA_signal_11457), .Q (new_AGEMA_signal_11458) ) ;
    buf_clk new_AGEMA_reg_buffer_5610 ( .C (clk), .D (new_AGEMA_signal_11461), .Q (new_AGEMA_signal_11462) ) ;
    buf_clk new_AGEMA_reg_buffer_5614 ( .C (clk), .D (new_AGEMA_signal_11465), .Q (new_AGEMA_signal_11466) ) ;
    buf_clk new_AGEMA_reg_buffer_5618 ( .C (clk), .D (new_AGEMA_signal_11469), .Q (new_AGEMA_signal_11470) ) ;
    buf_clk new_AGEMA_reg_buffer_5622 ( .C (clk), .D (new_AGEMA_signal_11473), .Q (new_AGEMA_signal_11474) ) ;
    buf_clk new_AGEMA_reg_buffer_5626 ( .C (clk), .D (new_AGEMA_signal_11477), .Q (new_AGEMA_signal_11478) ) ;
    buf_clk new_AGEMA_reg_buffer_5630 ( .C (clk), .D (new_AGEMA_signal_11481), .Q (new_AGEMA_signal_11482) ) ;
    buf_clk new_AGEMA_reg_buffer_5634 ( .C (clk), .D (new_AGEMA_signal_11485), .Q (new_AGEMA_signal_11486) ) ;
    buf_clk new_AGEMA_reg_buffer_5638 ( .C (clk), .D (new_AGEMA_signal_11489), .Q (new_AGEMA_signal_11490) ) ;
    buf_clk new_AGEMA_reg_buffer_5642 ( .C (clk), .D (new_AGEMA_signal_11493), .Q (new_AGEMA_signal_11494) ) ;
    buf_clk new_AGEMA_reg_buffer_5646 ( .C (clk), .D (new_AGEMA_signal_11497), .Q (new_AGEMA_signal_11498) ) ;
    buf_clk new_AGEMA_reg_buffer_5650 ( .C (clk), .D (new_AGEMA_signal_11501), .Q (new_AGEMA_signal_11502) ) ;
    buf_clk new_AGEMA_reg_buffer_5654 ( .C (clk), .D (new_AGEMA_signal_11505), .Q (new_AGEMA_signal_11506) ) ;
    buf_clk new_AGEMA_reg_buffer_5658 ( .C (clk), .D (new_AGEMA_signal_11509), .Q (new_AGEMA_signal_11510) ) ;
    buf_clk new_AGEMA_reg_buffer_5662 ( .C (clk), .D (new_AGEMA_signal_11513), .Q (new_AGEMA_signal_11514) ) ;
    buf_clk new_AGEMA_reg_buffer_5666 ( .C (clk), .D (new_AGEMA_signal_11517), .Q (new_AGEMA_signal_11518) ) ;
    buf_clk new_AGEMA_reg_buffer_5670 ( .C (clk), .D (new_AGEMA_signal_11521), .Q (new_AGEMA_signal_11522) ) ;
    buf_clk new_AGEMA_reg_buffer_5674 ( .C (clk), .D (new_AGEMA_signal_11525), .Q (new_AGEMA_signal_11526) ) ;
    buf_clk new_AGEMA_reg_buffer_5678 ( .C (clk), .D (new_AGEMA_signal_11529), .Q (new_AGEMA_signal_11530) ) ;
    buf_clk new_AGEMA_reg_buffer_5682 ( .C (clk), .D (new_AGEMA_signal_11533), .Q (new_AGEMA_signal_11534) ) ;
    buf_clk new_AGEMA_reg_buffer_5686 ( .C (clk), .D (new_AGEMA_signal_11537), .Q (new_AGEMA_signal_11538) ) ;
    buf_clk new_AGEMA_reg_buffer_5690 ( .C (clk), .D (new_AGEMA_signal_11541), .Q (new_AGEMA_signal_11542) ) ;
    buf_clk new_AGEMA_reg_buffer_5694 ( .C (clk), .D (new_AGEMA_signal_11545), .Q (new_AGEMA_signal_11546) ) ;
    buf_clk new_AGEMA_reg_buffer_5698 ( .C (clk), .D (new_AGEMA_signal_11549), .Q (new_AGEMA_signal_11550) ) ;
    buf_clk new_AGEMA_reg_buffer_5702 ( .C (clk), .D (new_AGEMA_signal_11553), .Q (new_AGEMA_signal_11554) ) ;
    buf_clk new_AGEMA_reg_buffer_5706 ( .C (clk), .D (new_AGEMA_signal_11557), .Q (new_AGEMA_signal_11558) ) ;
    buf_clk new_AGEMA_reg_buffer_5710 ( .C (clk), .D (new_AGEMA_signal_11561), .Q (new_AGEMA_signal_11562) ) ;
    buf_clk new_AGEMA_reg_buffer_5714 ( .C (clk), .D (new_AGEMA_signal_11565), .Q (new_AGEMA_signal_11566) ) ;
    buf_clk new_AGEMA_reg_buffer_5718 ( .C (clk), .D (new_AGEMA_signal_11569), .Q (new_AGEMA_signal_11570) ) ;
    buf_clk new_AGEMA_reg_buffer_5722 ( .C (clk), .D (new_AGEMA_signal_11573), .Q (new_AGEMA_signal_11574) ) ;
    buf_clk new_AGEMA_reg_buffer_5726 ( .C (clk), .D (new_AGEMA_signal_11577), .Q (new_AGEMA_signal_11578) ) ;
    buf_clk new_AGEMA_reg_buffer_5730 ( .C (clk), .D (new_AGEMA_signal_11581), .Q (new_AGEMA_signal_11582) ) ;
    buf_clk new_AGEMA_reg_buffer_5734 ( .C (clk), .D (new_AGEMA_signal_11585), .Q (new_AGEMA_signal_11586) ) ;
    buf_clk new_AGEMA_reg_buffer_5738 ( .C (clk), .D (new_AGEMA_signal_11589), .Q (new_AGEMA_signal_11590) ) ;
    buf_clk new_AGEMA_reg_buffer_5742 ( .C (clk), .D (new_AGEMA_signal_11593), .Q (new_AGEMA_signal_11594) ) ;
    buf_clk new_AGEMA_reg_buffer_5746 ( .C (clk), .D (new_AGEMA_signal_11597), .Q (new_AGEMA_signal_11598) ) ;
    buf_clk new_AGEMA_reg_buffer_5749 ( .C (clk), .D (new_AGEMA_signal_11600), .Q (new_AGEMA_signal_11601) ) ;
    buf_clk new_AGEMA_reg_buffer_5752 ( .C (clk), .D (new_AGEMA_signal_11603), .Q (new_AGEMA_signal_11604) ) ;
    buf_clk new_AGEMA_reg_buffer_5755 ( .C (clk), .D (new_AGEMA_signal_11606), .Q (new_AGEMA_signal_11607) ) ;
    buf_clk new_AGEMA_reg_buffer_5758 ( .C (clk), .D (new_AGEMA_signal_11609), .Q (new_AGEMA_signal_11610) ) ;
    buf_clk new_AGEMA_reg_buffer_5761 ( .C (clk), .D (new_AGEMA_signal_11612), .Q (new_AGEMA_signal_11613) ) ;
    buf_clk new_AGEMA_reg_buffer_5764 ( .C (clk), .D (new_AGEMA_signal_11615), .Q (new_AGEMA_signal_11616) ) ;
    buf_clk new_AGEMA_reg_buffer_5767 ( .C (clk), .D (new_AGEMA_signal_11618), .Q (new_AGEMA_signal_11619) ) ;
    buf_clk new_AGEMA_reg_buffer_5770 ( .C (clk), .D (new_AGEMA_signal_11621), .Q (new_AGEMA_signal_11622) ) ;
    buf_clk new_AGEMA_reg_buffer_5773 ( .C (clk), .D (new_AGEMA_signal_11624), .Q (new_AGEMA_signal_11625) ) ;
    buf_clk new_AGEMA_reg_buffer_5776 ( .C (clk), .D (new_AGEMA_signal_11627), .Q (new_AGEMA_signal_11628) ) ;
    buf_clk new_AGEMA_reg_buffer_5779 ( .C (clk), .D (new_AGEMA_signal_11630), .Q (new_AGEMA_signal_11631) ) ;
    buf_clk new_AGEMA_reg_buffer_5782 ( .C (clk), .D (new_AGEMA_signal_11633), .Q (new_AGEMA_signal_11634) ) ;
    buf_clk new_AGEMA_reg_buffer_5785 ( .C (clk), .D (new_AGEMA_signal_11636), .Q (new_AGEMA_signal_11637) ) ;
    buf_clk new_AGEMA_reg_buffer_5788 ( .C (clk), .D (new_AGEMA_signal_11639), .Q (new_AGEMA_signal_11640) ) ;
    buf_clk new_AGEMA_reg_buffer_5791 ( .C (clk), .D (new_AGEMA_signal_11642), .Q (new_AGEMA_signal_11643) ) ;
    buf_clk new_AGEMA_reg_buffer_5794 ( .C (clk), .D (new_AGEMA_signal_11645), .Q (new_AGEMA_signal_11646) ) ;
    buf_clk new_AGEMA_reg_buffer_5797 ( .C (clk), .D (new_AGEMA_signal_11648), .Q (new_AGEMA_signal_11649) ) ;
    buf_clk new_AGEMA_reg_buffer_5800 ( .C (clk), .D (new_AGEMA_signal_11651), .Q (new_AGEMA_signal_11652) ) ;
    buf_clk new_AGEMA_reg_buffer_5803 ( .C (clk), .D (new_AGEMA_signal_11654), .Q (new_AGEMA_signal_11655) ) ;
    buf_clk new_AGEMA_reg_buffer_5806 ( .C (clk), .D (new_AGEMA_signal_11657), .Q (new_AGEMA_signal_11658) ) ;
    buf_clk new_AGEMA_reg_buffer_5809 ( .C (clk), .D (new_AGEMA_signal_11660), .Q (new_AGEMA_signal_11661) ) ;
    buf_clk new_AGEMA_reg_buffer_5812 ( .C (clk), .D (new_AGEMA_signal_11663), .Q (new_AGEMA_signal_11664) ) ;
    buf_clk new_AGEMA_reg_buffer_5815 ( .C (clk), .D (new_AGEMA_signal_11666), .Q (new_AGEMA_signal_11667) ) ;
    buf_clk new_AGEMA_reg_buffer_5818 ( .C (clk), .D (new_AGEMA_signal_11669), .Q (new_AGEMA_signal_11670) ) ;
    buf_clk new_AGEMA_reg_buffer_5821 ( .C (clk), .D (new_AGEMA_signal_11672), .Q (new_AGEMA_signal_11673) ) ;
    buf_clk new_AGEMA_reg_buffer_5824 ( .C (clk), .D (new_AGEMA_signal_11675), .Q (new_AGEMA_signal_11676) ) ;
    buf_clk new_AGEMA_reg_buffer_5827 ( .C (clk), .D (new_AGEMA_signal_11678), .Q (new_AGEMA_signal_11679) ) ;
    buf_clk new_AGEMA_reg_buffer_5830 ( .C (clk), .D (new_AGEMA_signal_11681), .Q (new_AGEMA_signal_11682) ) ;
    buf_clk new_AGEMA_reg_buffer_5833 ( .C (clk), .D (new_AGEMA_signal_11684), .Q (new_AGEMA_signal_11685) ) ;
    buf_clk new_AGEMA_reg_buffer_5836 ( .C (clk), .D (new_AGEMA_signal_11687), .Q (new_AGEMA_signal_11688) ) ;
    buf_clk new_AGEMA_reg_buffer_5839 ( .C (clk), .D (new_AGEMA_signal_11690), .Q (new_AGEMA_signal_11691) ) ;
    buf_clk new_AGEMA_reg_buffer_5842 ( .C (clk), .D (new_AGEMA_signal_11693), .Q (new_AGEMA_signal_11694) ) ;
    buf_clk new_AGEMA_reg_buffer_5845 ( .C (clk), .D (new_AGEMA_signal_11696), .Q (new_AGEMA_signal_11697) ) ;
    buf_clk new_AGEMA_reg_buffer_5848 ( .C (clk), .D (new_AGEMA_signal_11699), .Q (new_AGEMA_signal_11700) ) ;
    buf_clk new_AGEMA_reg_buffer_5851 ( .C (clk), .D (new_AGEMA_signal_11702), .Q (new_AGEMA_signal_11703) ) ;
    buf_clk new_AGEMA_reg_buffer_5854 ( .C (clk), .D (new_AGEMA_signal_11705), .Q (new_AGEMA_signal_11706) ) ;
    buf_clk new_AGEMA_reg_buffer_5857 ( .C (clk), .D (new_AGEMA_signal_11708), .Q (new_AGEMA_signal_11709) ) ;
    buf_clk new_AGEMA_reg_buffer_5860 ( .C (clk), .D (new_AGEMA_signal_11711), .Q (new_AGEMA_signal_11712) ) ;
    buf_clk new_AGEMA_reg_buffer_5863 ( .C (clk), .D (new_AGEMA_signal_11714), .Q (new_AGEMA_signal_11715) ) ;
    buf_clk new_AGEMA_reg_buffer_5866 ( .C (clk), .D (new_AGEMA_signal_11717), .Q (new_AGEMA_signal_11718) ) ;
    buf_clk new_AGEMA_reg_buffer_5869 ( .C (clk), .D (new_AGEMA_signal_11720), .Q (new_AGEMA_signal_11721) ) ;
    buf_clk new_AGEMA_reg_buffer_5872 ( .C (clk), .D (new_AGEMA_signal_11723), .Q (new_AGEMA_signal_11724) ) ;
    buf_clk new_AGEMA_reg_buffer_5875 ( .C (clk), .D (new_AGEMA_signal_11726), .Q (new_AGEMA_signal_11727) ) ;
    buf_clk new_AGEMA_reg_buffer_5878 ( .C (clk), .D (new_AGEMA_signal_11729), .Q (new_AGEMA_signal_11730) ) ;
    buf_clk new_AGEMA_reg_buffer_5881 ( .C (clk), .D (new_AGEMA_signal_11732), .Q (new_AGEMA_signal_11733) ) ;
    buf_clk new_AGEMA_reg_buffer_5884 ( .C (clk), .D (new_AGEMA_signal_11735), .Q (new_AGEMA_signal_11736) ) ;
    buf_clk new_AGEMA_reg_buffer_5887 ( .C (clk), .D (new_AGEMA_signal_11738), .Q (new_AGEMA_signal_11739) ) ;
    buf_clk new_AGEMA_reg_buffer_5890 ( .C (clk), .D (new_AGEMA_signal_11741), .Q (new_AGEMA_signal_11742) ) ;
    buf_clk new_AGEMA_reg_buffer_5893 ( .C (clk), .D (new_AGEMA_signal_11744), .Q (new_AGEMA_signal_11745) ) ;
    buf_clk new_AGEMA_reg_buffer_5896 ( .C (clk), .D (new_AGEMA_signal_11747), .Q (new_AGEMA_signal_11748) ) ;
    buf_clk new_AGEMA_reg_buffer_5899 ( .C (clk), .D (new_AGEMA_signal_11750), .Q (new_AGEMA_signal_11751) ) ;
    buf_clk new_AGEMA_reg_buffer_5902 ( .C (clk), .D (new_AGEMA_signal_11753), .Q (new_AGEMA_signal_11754) ) ;
    buf_clk new_AGEMA_reg_buffer_5905 ( .C (clk), .D (new_AGEMA_signal_11756), .Q (new_AGEMA_signal_11757) ) ;
    buf_clk new_AGEMA_reg_buffer_5908 ( .C (clk), .D (new_AGEMA_signal_11759), .Q (new_AGEMA_signal_11760) ) ;
    buf_clk new_AGEMA_reg_buffer_5911 ( .C (clk), .D (new_AGEMA_signal_11762), .Q (new_AGEMA_signal_11763) ) ;
    buf_clk new_AGEMA_reg_buffer_5914 ( .C (clk), .D (new_AGEMA_signal_11765), .Q (new_AGEMA_signal_11766) ) ;
    buf_clk new_AGEMA_reg_buffer_5917 ( .C (clk), .D (new_AGEMA_signal_11768), .Q (new_AGEMA_signal_11769) ) ;
    buf_clk new_AGEMA_reg_buffer_5920 ( .C (clk), .D (new_AGEMA_signal_11771), .Q (new_AGEMA_signal_11772) ) ;
    buf_clk new_AGEMA_reg_buffer_5923 ( .C (clk), .D (new_AGEMA_signal_11774), .Q (new_AGEMA_signal_11775) ) ;
    buf_clk new_AGEMA_reg_buffer_5926 ( .C (clk), .D (new_AGEMA_signal_11777), .Q (new_AGEMA_signal_11778) ) ;
    buf_clk new_AGEMA_reg_buffer_5929 ( .C (clk), .D (new_AGEMA_signal_11780), .Q (new_AGEMA_signal_11781) ) ;
    buf_clk new_AGEMA_reg_buffer_5932 ( .C (clk), .D (new_AGEMA_signal_11783), .Q (new_AGEMA_signal_11784) ) ;
    buf_clk new_AGEMA_reg_buffer_5935 ( .C (clk), .D (new_AGEMA_signal_11786), .Q (new_AGEMA_signal_11787) ) ;
    buf_clk new_AGEMA_reg_buffer_5938 ( .C (clk), .D (new_AGEMA_signal_11789), .Q (new_AGEMA_signal_11790) ) ;
    buf_clk new_AGEMA_reg_buffer_5941 ( .C (clk), .D (new_AGEMA_signal_11792), .Q (new_AGEMA_signal_11793) ) ;
    buf_clk new_AGEMA_reg_buffer_5944 ( .C (clk), .D (new_AGEMA_signal_11795), .Q (new_AGEMA_signal_11796) ) ;
    buf_clk new_AGEMA_reg_buffer_5947 ( .C (clk), .D (new_AGEMA_signal_11798), .Q (new_AGEMA_signal_11799) ) ;
    buf_clk new_AGEMA_reg_buffer_5950 ( .C (clk), .D (new_AGEMA_signal_11801), .Q (new_AGEMA_signal_11802) ) ;
    buf_clk new_AGEMA_reg_buffer_5953 ( .C (clk), .D (new_AGEMA_signal_11804), .Q (new_AGEMA_signal_11805) ) ;
    buf_clk new_AGEMA_reg_buffer_5956 ( .C (clk), .D (new_AGEMA_signal_11807), .Q (new_AGEMA_signal_11808) ) ;
    buf_clk new_AGEMA_reg_buffer_5959 ( .C (clk), .D (new_AGEMA_signal_11810), .Q (new_AGEMA_signal_11811) ) ;
    buf_clk new_AGEMA_reg_buffer_5962 ( .C (clk), .D (new_AGEMA_signal_11813), .Q (new_AGEMA_signal_11814) ) ;
    buf_clk new_AGEMA_reg_buffer_5965 ( .C (clk), .D (new_AGEMA_signal_11816), .Q (new_AGEMA_signal_11817) ) ;
    buf_clk new_AGEMA_reg_buffer_5968 ( .C (clk), .D (new_AGEMA_signal_11819), .Q (new_AGEMA_signal_11820) ) ;
    buf_clk new_AGEMA_reg_buffer_5971 ( .C (clk), .D (new_AGEMA_signal_11822), .Q (new_AGEMA_signal_11823) ) ;
    buf_clk new_AGEMA_reg_buffer_5974 ( .C (clk), .D (new_AGEMA_signal_11825), .Q (new_AGEMA_signal_11826) ) ;
    buf_clk new_AGEMA_reg_buffer_5977 ( .C (clk), .D (new_AGEMA_signal_11828), .Q (new_AGEMA_signal_11829) ) ;
    buf_clk new_AGEMA_reg_buffer_5980 ( .C (clk), .D (new_AGEMA_signal_11831), .Q (new_AGEMA_signal_11832) ) ;
    buf_clk new_AGEMA_reg_buffer_5983 ( .C (clk), .D (new_AGEMA_signal_11834), .Q (new_AGEMA_signal_11835) ) ;
    buf_clk new_AGEMA_reg_buffer_5986 ( .C (clk), .D (new_AGEMA_signal_11837), .Q (new_AGEMA_signal_11838) ) ;
    buf_clk new_AGEMA_reg_buffer_5989 ( .C (clk), .D (new_AGEMA_signal_11840), .Q (new_AGEMA_signal_11841) ) ;
    buf_clk new_AGEMA_reg_buffer_5992 ( .C (clk), .D (new_AGEMA_signal_11843), .Q (new_AGEMA_signal_11844) ) ;
    buf_clk new_AGEMA_reg_buffer_5995 ( .C (clk), .D (new_AGEMA_signal_11846), .Q (new_AGEMA_signal_11847) ) ;
    buf_clk new_AGEMA_reg_buffer_5998 ( .C (clk), .D (new_AGEMA_signal_11849), .Q (new_AGEMA_signal_11850) ) ;
    buf_clk new_AGEMA_reg_buffer_6001 ( .C (clk), .D (new_AGEMA_signal_11852), .Q (new_AGEMA_signal_11853) ) ;
    buf_clk new_AGEMA_reg_buffer_6004 ( .C (clk), .D (new_AGEMA_signal_11855), .Q (new_AGEMA_signal_11856) ) ;
    buf_clk new_AGEMA_reg_buffer_6007 ( .C (clk), .D (new_AGEMA_signal_11858), .Q (new_AGEMA_signal_11859) ) ;
    buf_clk new_AGEMA_reg_buffer_6010 ( .C (clk), .D (new_AGEMA_signal_11861), .Q (new_AGEMA_signal_11862) ) ;
    buf_clk new_AGEMA_reg_buffer_6013 ( .C (clk), .D (new_AGEMA_signal_11864), .Q (new_AGEMA_signal_11865) ) ;
    buf_clk new_AGEMA_reg_buffer_6016 ( .C (clk), .D (new_AGEMA_signal_11867), .Q (new_AGEMA_signal_11868) ) ;
    buf_clk new_AGEMA_reg_buffer_6019 ( .C (clk), .D (new_AGEMA_signal_11870), .Q (new_AGEMA_signal_11871) ) ;
    buf_clk new_AGEMA_reg_buffer_6022 ( .C (clk), .D (new_AGEMA_signal_11873), .Q (new_AGEMA_signal_11874) ) ;
    buf_clk new_AGEMA_reg_buffer_6025 ( .C (clk), .D (new_AGEMA_signal_11876), .Q (new_AGEMA_signal_11877) ) ;
    buf_clk new_AGEMA_reg_buffer_6028 ( .C (clk), .D (new_AGEMA_signal_11879), .Q (new_AGEMA_signal_11880) ) ;
    buf_clk new_AGEMA_reg_buffer_6031 ( .C (clk), .D (new_AGEMA_signal_11882), .Q (new_AGEMA_signal_11883) ) ;
    buf_clk new_AGEMA_reg_buffer_6034 ( .C (clk), .D (new_AGEMA_signal_11885), .Q (new_AGEMA_signal_11886) ) ;
    buf_clk new_AGEMA_reg_buffer_6037 ( .C (clk), .D (new_AGEMA_signal_11888), .Q (new_AGEMA_signal_11889) ) ;
    buf_clk new_AGEMA_reg_buffer_6040 ( .C (clk), .D (new_AGEMA_signal_11891), .Q (new_AGEMA_signal_11892) ) ;
    buf_clk new_AGEMA_reg_buffer_6043 ( .C (clk), .D (new_AGEMA_signal_11894), .Q (new_AGEMA_signal_11895) ) ;
    buf_clk new_AGEMA_reg_buffer_6046 ( .C (clk), .D (new_AGEMA_signal_11897), .Q (new_AGEMA_signal_11898) ) ;
    buf_clk new_AGEMA_reg_buffer_6049 ( .C (clk), .D (new_AGEMA_signal_11900), .Q (new_AGEMA_signal_11901) ) ;
    buf_clk new_AGEMA_reg_buffer_6052 ( .C (clk), .D (new_AGEMA_signal_11903), .Q (new_AGEMA_signal_11904) ) ;
    buf_clk new_AGEMA_reg_buffer_6055 ( .C (clk), .D (new_AGEMA_signal_11906), .Q (new_AGEMA_signal_11907) ) ;
    buf_clk new_AGEMA_reg_buffer_6058 ( .C (clk), .D (new_AGEMA_signal_11909), .Q (new_AGEMA_signal_11910) ) ;
    buf_clk new_AGEMA_reg_buffer_6061 ( .C (clk), .D (new_AGEMA_signal_11912), .Q (new_AGEMA_signal_11913) ) ;
    buf_clk new_AGEMA_reg_buffer_6064 ( .C (clk), .D (new_AGEMA_signal_11915), .Q (new_AGEMA_signal_11916) ) ;
    buf_clk new_AGEMA_reg_buffer_6067 ( .C (clk), .D (new_AGEMA_signal_11918), .Q (new_AGEMA_signal_11919) ) ;
    buf_clk new_AGEMA_reg_buffer_6070 ( .C (clk), .D (new_AGEMA_signal_11921), .Q (new_AGEMA_signal_11922) ) ;
    buf_clk new_AGEMA_reg_buffer_6073 ( .C (clk), .D (new_AGEMA_signal_11924), .Q (new_AGEMA_signal_11925) ) ;
    buf_clk new_AGEMA_reg_buffer_6076 ( .C (clk), .D (new_AGEMA_signal_11927), .Q (new_AGEMA_signal_11928) ) ;
    buf_clk new_AGEMA_reg_buffer_6079 ( .C (clk), .D (new_AGEMA_signal_11930), .Q (new_AGEMA_signal_11931) ) ;
    buf_clk new_AGEMA_reg_buffer_6082 ( .C (clk), .D (new_AGEMA_signal_11933), .Q (new_AGEMA_signal_11934) ) ;
    buf_clk new_AGEMA_reg_buffer_6085 ( .C (clk), .D (new_AGEMA_signal_11936), .Q (new_AGEMA_signal_11937) ) ;
    buf_clk new_AGEMA_reg_buffer_6088 ( .C (clk), .D (new_AGEMA_signal_11939), .Q (new_AGEMA_signal_11940) ) ;
    buf_clk new_AGEMA_reg_buffer_6091 ( .C (clk), .D (new_AGEMA_signal_11942), .Q (new_AGEMA_signal_11943) ) ;
    buf_clk new_AGEMA_reg_buffer_6094 ( .C (clk), .D (new_AGEMA_signal_11945), .Q (new_AGEMA_signal_11946) ) ;
    buf_clk new_AGEMA_reg_buffer_6097 ( .C (clk), .D (new_AGEMA_signal_11948), .Q (new_AGEMA_signal_11949) ) ;
    buf_clk new_AGEMA_reg_buffer_6100 ( .C (clk), .D (new_AGEMA_signal_11951), .Q (new_AGEMA_signal_11952) ) ;
    buf_clk new_AGEMA_reg_buffer_6103 ( .C (clk), .D (new_AGEMA_signal_11954), .Q (new_AGEMA_signal_11955) ) ;
    buf_clk new_AGEMA_reg_buffer_6106 ( .C (clk), .D (new_AGEMA_signal_11957), .Q (new_AGEMA_signal_11958) ) ;
    buf_clk new_AGEMA_reg_buffer_6109 ( .C (clk), .D (new_AGEMA_signal_11960), .Q (new_AGEMA_signal_11961) ) ;
    buf_clk new_AGEMA_reg_buffer_6112 ( .C (clk), .D (new_AGEMA_signal_11963), .Q (new_AGEMA_signal_11964) ) ;
    buf_clk new_AGEMA_reg_buffer_6115 ( .C (clk), .D (new_AGEMA_signal_11966), .Q (new_AGEMA_signal_11967) ) ;
    buf_clk new_AGEMA_reg_buffer_6118 ( .C (clk), .D (new_AGEMA_signal_11969), .Q (new_AGEMA_signal_11970) ) ;
    buf_clk new_AGEMA_reg_buffer_6121 ( .C (clk), .D (new_AGEMA_signal_11972), .Q (new_AGEMA_signal_11973) ) ;
    buf_clk new_AGEMA_reg_buffer_6124 ( .C (clk), .D (new_AGEMA_signal_11975), .Q (new_AGEMA_signal_11976) ) ;
    buf_clk new_AGEMA_reg_buffer_6127 ( .C (clk), .D (new_AGEMA_signal_11978), .Q (new_AGEMA_signal_11979) ) ;
    buf_clk new_AGEMA_reg_buffer_6130 ( .C (clk), .D (new_AGEMA_signal_11981), .Q (new_AGEMA_signal_11982) ) ;
    buf_clk new_AGEMA_reg_buffer_6133 ( .C (clk), .D (new_AGEMA_signal_11984), .Q (new_AGEMA_signal_11985) ) ;
    buf_clk new_AGEMA_reg_buffer_6136 ( .C (clk), .D (new_AGEMA_signal_11987), .Q (new_AGEMA_signal_11988) ) ;
    buf_clk new_AGEMA_reg_buffer_6139 ( .C (clk), .D (new_AGEMA_signal_11990), .Q (new_AGEMA_signal_11991) ) ;
    buf_clk new_AGEMA_reg_buffer_6142 ( .C (clk), .D (new_AGEMA_signal_11993), .Q (new_AGEMA_signal_11994) ) ;
    buf_clk new_AGEMA_reg_buffer_6145 ( .C (clk), .D (new_AGEMA_signal_11996), .Q (new_AGEMA_signal_11997) ) ;
    buf_clk new_AGEMA_reg_buffer_6148 ( .C (clk), .D (new_AGEMA_signal_11999), .Q (new_AGEMA_signal_12000) ) ;
    buf_clk new_AGEMA_reg_buffer_6151 ( .C (clk), .D (new_AGEMA_signal_12002), .Q (new_AGEMA_signal_12003) ) ;
    buf_clk new_AGEMA_reg_buffer_6154 ( .C (clk), .D (new_AGEMA_signal_12005), .Q (new_AGEMA_signal_12006) ) ;
    buf_clk new_AGEMA_reg_buffer_6157 ( .C (clk), .D (new_AGEMA_signal_12008), .Q (new_AGEMA_signal_12009) ) ;
    buf_clk new_AGEMA_reg_buffer_6160 ( .C (clk), .D (new_AGEMA_signal_12011), .Q (new_AGEMA_signal_12012) ) ;
    buf_clk new_AGEMA_reg_buffer_6163 ( .C (clk), .D (new_AGEMA_signal_12014), .Q (new_AGEMA_signal_12015) ) ;
    buf_clk new_AGEMA_reg_buffer_6166 ( .C (clk), .D (new_AGEMA_signal_12017), .Q (new_AGEMA_signal_12018) ) ;
    buf_clk new_AGEMA_reg_buffer_6169 ( .C (clk), .D (new_AGEMA_signal_12020), .Q (new_AGEMA_signal_12021) ) ;
    buf_clk new_AGEMA_reg_buffer_6172 ( .C (clk), .D (new_AGEMA_signal_12023), .Q (new_AGEMA_signal_12024) ) ;
    buf_clk new_AGEMA_reg_buffer_6175 ( .C (clk), .D (new_AGEMA_signal_12026), .Q (new_AGEMA_signal_12027) ) ;
    buf_clk new_AGEMA_reg_buffer_6178 ( .C (clk), .D (new_AGEMA_signal_12029), .Q (new_AGEMA_signal_12030) ) ;
    buf_clk new_AGEMA_reg_buffer_6181 ( .C (clk), .D (new_AGEMA_signal_12032), .Q (new_AGEMA_signal_12033) ) ;
    buf_clk new_AGEMA_reg_buffer_6184 ( .C (clk), .D (new_AGEMA_signal_12035), .Q (new_AGEMA_signal_12036) ) ;
    buf_clk new_AGEMA_reg_buffer_6187 ( .C (clk), .D (new_AGEMA_signal_12038), .Q (new_AGEMA_signal_12039) ) ;
    buf_clk new_AGEMA_reg_buffer_6190 ( .C (clk), .D (new_AGEMA_signal_12041), .Q (new_AGEMA_signal_12042) ) ;
    buf_clk new_AGEMA_reg_buffer_6193 ( .C (clk), .D (new_AGEMA_signal_12044), .Q (new_AGEMA_signal_12045) ) ;
    buf_clk new_AGEMA_reg_buffer_6196 ( .C (clk), .D (new_AGEMA_signal_12047), .Q (new_AGEMA_signal_12048) ) ;
    buf_clk new_AGEMA_reg_buffer_6199 ( .C (clk), .D (new_AGEMA_signal_12050), .Q (new_AGEMA_signal_12051) ) ;
    buf_clk new_AGEMA_reg_buffer_6202 ( .C (clk), .D (new_AGEMA_signal_12053), .Q (new_AGEMA_signal_12054) ) ;
    buf_clk new_AGEMA_reg_buffer_6205 ( .C (clk), .D (new_AGEMA_signal_12056), .Q (new_AGEMA_signal_12057) ) ;
    buf_clk new_AGEMA_reg_buffer_6208 ( .C (clk), .D (new_AGEMA_signal_12059), .Q (new_AGEMA_signal_12060) ) ;
    buf_clk new_AGEMA_reg_buffer_6211 ( .C (clk), .D (new_AGEMA_signal_12062), .Q (new_AGEMA_signal_12063) ) ;
    buf_clk new_AGEMA_reg_buffer_6214 ( .C (clk), .D (new_AGEMA_signal_12065), .Q (new_AGEMA_signal_12066) ) ;
    buf_clk new_AGEMA_reg_buffer_6217 ( .C (clk), .D (new_AGEMA_signal_12068), .Q (new_AGEMA_signal_12069) ) ;
    buf_clk new_AGEMA_reg_buffer_6220 ( .C (clk), .D (new_AGEMA_signal_12071), .Q (new_AGEMA_signal_12072) ) ;
    buf_clk new_AGEMA_reg_buffer_6223 ( .C (clk), .D (new_AGEMA_signal_12074), .Q (new_AGEMA_signal_12075) ) ;
    buf_clk new_AGEMA_reg_buffer_6226 ( .C (clk), .D (new_AGEMA_signal_12077), .Q (new_AGEMA_signal_12078) ) ;
    buf_clk new_AGEMA_reg_buffer_6229 ( .C (clk), .D (new_AGEMA_signal_12080), .Q (new_AGEMA_signal_12081) ) ;
    buf_clk new_AGEMA_reg_buffer_6232 ( .C (clk), .D (new_AGEMA_signal_12083), .Q (new_AGEMA_signal_12084) ) ;
    buf_clk new_AGEMA_reg_buffer_6235 ( .C (clk), .D (new_AGEMA_signal_12086), .Q (new_AGEMA_signal_12087) ) ;
    buf_clk new_AGEMA_reg_buffer_6238 ( .C (clk), .D (new_AGEMA_signal_12089), .Q (new_AGEMA_signal_12090) ) ;
    buf_clk new_AGEMA_reg_buffer_6241 ( .C (clk), .D (new_AGEMA_signal_12092), .Q (new_AGEMA_signal_12093) ) ;
    buf_clk new_AGEMA_reg_buffer_6244 ( .C (clk), .D (new_AGEMA_signal_12095), .Q (new_AGEMA_signal_12096) ) ;
    buf_clk new_AGEMA_reg_buffer_6247 ( .C (clk), .D (new_AGEMA_signal_12098), .Q (new_AGEMA_signal_12099) ) ;
    buf_clk new_AGEMA_reg_buffer_6250 ( .C (clk), .D (new_AGEMA_signal_12101), .Q (new_AGEMA_signal_12102) ) ;
    buf_clk new_AGEMA_reg_buffer_6253 ( .C (clk), .D (new_AGEMA_signal_12104), .Q (new_AGEMA_signal_12105) ) ;
    buf_clk new_AGEMA_reg_buffer_6256 ( .C (clk), .D (new_AGEMA_signal_12107), .Q (new_AGEMA_signal_12108) ) ;
    buf_clk new_AGEMA_reg_buffer_6259 ( .C (clk), .D (new_AGEMA_signal_12110), .Q (new_AGEMA_signal_12111) ) ;
    buf_clk new_AGEMA_reg_buffer_6262 ( .C (clk), .D (new_AGEMA_signal_12113), .Q (new_AGEMA_signal_12114) ) ;
    buf_clk new_AGEMA_reg_buffer_6265 ( .C (clk), .D (new_AGEMA_signal_12116), .Q (new_AGEMA_signal_12117) ) ;
    buf_clk new_AGEMA_reg_buffer_6268 ( .C (clk), .D (new_AGEMA_signal_12119), .Q (new_AGEMA_signal_12120) ) ;
    buf_clk new_AGEMA_reg_buffer_6271 ( .C (clk), .D (new_AGEMA_signal_12122), .Q (new_AGEMA_signal_12123) ) ;
    buf_clk new_AGEMA_reg_buffer_6274 ( .C (clk), .D (new_AGEMA_signal_12125), .Q (new_AGEMA_signal_12126) ) ;
    buf_clk new_AGEMA_reg_buffer_6277 ( .C (clk), .D (new_AGEMA_signal_12128), .Q (new_AGEMA_signal_12129) ) ;
    buf_clk new_AGEMA_reg_buffer_6280 ( .C (clk), .D (new_AGEMA_signal_12131), .Q (new_AGEMA_signal_12132) ) ;
    buf_clk new_AGEMA_reg_buffer_6283 ( .C (clk), .D (new_AGEMA_signal_12134), .Q (new_AGEMA_signal_12135) ) ;
    buf_clk new_AGEMA_reg_buffer_6286 ( .C (clk), .D (new_AGEMA_signal_12137), .Q (new_AGEMA_signal_12138) ) ;
    buf_clk new_AGEMA_reg_buffer_6289 ( .C (clk), .D (new_AGEMA_signal_12140), .Q (new_AGEMA_signal_12141) ) ;
    buf_clk new_AGEMA_reg_buffer_6292 ( .C (clk), .D (new_AGEMA_signal_12143), .Q (new_AGEMA_signal_12144) ) ;
    buf_clk new_AGEMA_reg_buffer_6295 ( .C (clk), .D (new_AGEMA_signal_12146), .Q (new_AGEMA_signal_12147) ) ;
    buf_clk new_AGEMA_reg_buffer_6298 ( .C (clk), .D (new_AGEMA_signal_12149), .Q (new_AGEMA_signal_12150) ) ;
    buf_clk new_AGEMA_reg_buffer_6301 ( .C (clk), .D (new_AGEMA_signal_12152), .Q (new_AGEMA_signal_12153) ) ;
    buf_clk new_AGEMA_reg_buffer_6304 ( .C (clk), .D (new_AGEMA_signal_12155), .Q (new_AGEMA_signal_12156) ) ;
    buf_clk new_AGEMA_reg_buffer_6307 ( .C (clk), .D (new_AGEMA_signal_12158), .Q (new_AGEMA_signal_12159) ) ;
    buf_clk new_AGEMA_reg_buffer_6310 ( .C (clk), .D (new_AGEMA_signal_12161), .Q (new_AGEMA_signal_12162) ) ;
    buf_clk new_AGEMA_reg_buffer_6313 ( .C (clk), .D (new_AGEMA_signal_12164), .Q (new_AGEMA_signal_12165) ) ;
    buf_clk new_AGEMA_reg_buffer_6316 ( .C (clk), .D (new_AGEMA_signal_12167), .Q (new_AGEMA_signal_12168) ) ;
    buf_clk new_AGEMA_reg_buffer_6319 ( .C (clk), .D (new_AGEMA_signal_12170), .Q (new_AGEMA_signal_12171) ) ;
    buf_clk new_AGEMA_reg_buffer_6322 ( .C (clk), .D (new_AGEMA_signal_12173), .Q (new_AGEMA_signal_12174) ) ;
    buf_clk new_AGEMA_reg_buffer_6325 ( .C (clk), .D (new_AGEMA_signal_12176), .Q (new_AGEMA_signal_12177) ) ;
    buf_clk new_AGEMA_reg_buffer_6328 ( .C (clk), .D (new_AGEMA_signal_12179), .Q (new_AGEMA_signal_12180) ) ;
    buf_clk new_AGEMA_reg_buffer_6331 ( .C (clk), .D (new_AGEMA_signal_12182), .Q (new_AGEMA_signal_12183) ) ;
    buf_clk new_AGEMA_reg_buffer_6334 ( .C (clk), .D (new_AGEMA_signal_12185), .Q (new_AGEMA_signal_12186) ) ;
    buf_clk new_AGEMA_reg_buffer_6337 ( .C (clk), .D (new_AGEMA_signal_12188), .Q (new_AGEMA_signal_12189) ) ;
    buf_clk new_AGEMA_reg_buffer_6340 ( .C (clk), .D (new_AGEMA_signal_12191), .Q (new_AGEMA_signal_12192) ) ;
    buf_clk new_AGEMA_reg_buffer_6343 ( .C (clk), .D (new_AGEMA_signal_12194), .Q (new_AGEMA_signal_12195) ) ;
    buf_clk new_AGEMA_reg_buffer_6346 ( .C (clk), .D (new_AGEMA_signal_12197), .Q (new_AGEMA_signal_12198) ) ;
    buf_clk new_AGEMA_reg_buffer_6349 ( .C (clk), .D (new_AGEMA_signal_12200), .Q (new_AGEMA_signal_12201) ) ;
    buf_clk new_AGEMA_reg_buffer_6352 ( .C (clk), .D (new_AGEMA_signal_12203), .Q (new_AGEMA_signal_12204) ) ;
    buf_clk new_AGEMA_reg_buffer_6355 ( .C (clk), .D (new_AGEMA_signal_12206), .Q (new_AGEMA_signal_12207) ) ;
    buf_clk new_AGEMA_reg_buffer_6358 ( .C (clk), .D (new_AGEMA_signal_12209), .Q (new_AGEMA_signal_12210) ) ;
    buf_clk new_AGEMA_reg_buffer_6361 ( .C (clk), .D (new_AGEMA_signal_12212), .Q (new_AGEMA_signal_12213) ) ;
    buf_clk new_AGEMA_reg_buffer_6364 ( .C (clk), .D (new_AGEMA_signal_12215), .Q (new_AGEMA_signal_12216) ) ;
    buf_clk new_AGEMA_reg_buffer_6367 ( .C (clk), .D (new_AGEMA_signal_12218), .Q (new_AGEMA_signal_12219) ) ;
    buf_clk new_AGEMA_reg_buffer_6370 ( .C (clk), .D (new_AGEMA_signal_12221), .Q (new_AGEMA_signal_12222) ) ;
    buf_clk new_AGEMA_reg_buffer_6373 ( .C (clk), .D (new_AGEMA_signal_12224), .Q (new_AGEMA_signal_12225) ) ;
    buf_clk new_AGEMA_reg_buffer_6376 ( .C (clk), .D (new_AGEMA_signal_12227), .Q (new_AGEMA_signal_12228) ) ;
    buf_clk new_AGEMA_reg_buffer_6379 ( .C (clk), .D (new_AGEMA_signal_12230), .Q (new_AGEMA_signal_12231) ) ;
    buf_clk new_AGEMA_reg_buffer_6382 ( .C (clk), .D (new_AGEMA_signal_12233), .Q (new_AGEMA_signal_12234) ) ;
    buf_clk new_AGEMA_reg_buffer_6385 ( .C (clk), .D (new_AGEMA_signal_12236), .Q (new_AGEMA_signal_12237) ) ;
    buf_clk new_AGEMA_reg_buffer_6388 ( .C (clk), .D (new_AGEMA_signal_12239), .Q (new_AGEMA_signal_12240) ) ;
    buf_clk new_AGEMA_reg_buffer_6391 ( .C (clk), .D (new_AGEMA_signal_12242), .Q (new_AGEMA_signal_12243) ) ;
    buf_clk new_AGEMA_reg_buffer_6394 ( .C (clk), .D (new_AGEMA_signal_12245), .Q (new_AGEMA_signal_12246) ) ;
    buf_clk new_AGEMA_reg_buffer_6397 ( .C (clk), .D (new_AGEMA_signal_12248), .Q (new_AGEMA_signal_12249) ) ;
    buf_clk new_AGEMA_reg_buffer_6400 ( .C (clk), .D (new_AGEMA_signal_12251), .Q (new_AGEMA_signal_12252) ) ;
    buf_clk new_AGEMA_reg_buffer_6403 ( .C (clk), .D (new_AGEMA_signal_12254), .Q (new_AGEMA_signal_12255) ) ;
    buf_clk new_AGEMA_reg_buffer_6406 ( .C (clk), .D (new_AGEMA_signal_12257), .Q (new_AGEMA_signal_12258) ) ;
    buf_clk new_AGEMA_reg_buffer_6409 ( .C (clk), .D (new_AGEMA_signal_12260), .Q (new_AGEMA_signal_12261) ) ;
    buf_clk new_AGEMA_reg_buffer_6412 ( .C (clk), .D (new_AGEMA_signal_12263), .Q (new_AGEMA_signal_12264) ) ;
    buf_clk new_AGEMA_reg_buffer_6415 ( .C (clk), .D (new_AGEMA_signal_12266), .Q (new_AGEMA_signal_12267) ) ;
    buf_clk new_AGEMA_reg_buffer_6418 ( .C (clk), .D (new_AGEMA_signal_12269), .Q (new_AGEMA_signal_12270) ) ;
    buf_clk new_AGEMA_reg_buffer_6421 ( .C (clk), .D (new_AGEMA_signal_12272), .Q (new_AGEMA_signal_12273) ) ;
    buf_clk new_AGEMA_reg_buffer_6424 ( .C (clk), .D (new_AGEMA_signal_12275), .Q (new_AGEMA_signal_12276) ) ;
    buf_clk new_AGEMA_reg_buffer_6427 ( .C (clk), .D (new_AGEMA_signal_12278), .Q (new_AGEMA_signal_12279) ) ;
    buf_clk new_AGEMA_reg_buffer_6430 ( .C (clk), .D (new_AGEMA_signal_12281), .Q (new_AGEMA_signal_12282) ) ;
    buf_clk new_AGEMA_reg_buffer_6433 ( .C (clk), .D (new_AGEMA_signal_12284), .Q (new_AGEMA_signal_12285) ) ;
    buf_clk new_AGEMA_reg_buffer_6436 ( .C (clk), .D (new_AGEMA_signal_12287), .Q (new_AGEMA_signal_12288) ) ;
    buf_clk new_AGEMA_reg_buffer_6439 ( .C (clk), .D (new_AGEMA_signal_12290), .Q (new_AGEMA_signal_12291) ) ;
    buf_clk new_AGEMA_reg_buffer_6442 ( .C (clk), .D (new_AGEMA_signal_12293), .Q (new_AGEMA_signal_12294) ) ;
    buf_clk new_AGEMA_reg_buffer_6445 ( .C (clk), .D (new_AGEMA_signal_12296), .Q (new_AGEMA_signal_12297) ) ;
    buf_clk new_AGEMA_reg_buffer_6448 ( .C (clk), .D (new_AGEMA_signal_12299), .Q (new_AGEMA_signal_12300) ) ;
    buf_clk new_AGEMA_reg_buffer_6451 ( .C (clk), .D (new_AGEMA_signal_12302), .Q (new_AGEMA_signal_12303) ) ;
    buf_clk new_AGEMA_reg_buffer_6454 ( .C (clk), .D (new_AGEMA_signal_12305), .Q (new_AGEMA_signal_12306) ) ;
    buf_clk new_AGEMA_reg_buffer_6457 ( .C (clk), .D (new_AGEMA_signal_12308), .Q (new_AGEMA_signal_12309) ) ;
    buf_clk new_AGEMA_reg_buffer_6460 ( .C (clk), .D (new_AGEMA_signal_12311), .Q (new_AGEMA_signal_12312) ) ;
    buf_clk new_AGEMA_reg_buffer_6463 ( .C (clk), .D (new_AGEMA_signal_12314), .Q (new_AGEMA_signal_12315) ) ;
    buf_clk new_AGEMA_reg_buffer_6466 ( .C (clk), .D (new_AGEMA_signal_12317), .Q (new_AGEMA_signal_12318) ) ;
    buf_clk new_AGEMA_reg_buffer_6469 ( .C (clk), .D (new_AGEMA_signal_12320), .Q (new_AGEMA_signal_12321) ) ;
    buf_clk new_AGEMA_reg_buffer_6472 ( .C (clk), .D (new_AGEMA_signal_12323), .Q (new_AGEMA_signal_12324) ) ;
    buf_clk new_AGEMA_reg_buffer_6475 ( .C (clk), .D (new_AGEMA_signal_12326), .Q (new_AGEMA_signal_12327) ) ;
    buf_clk new_AGEMA_reg_buffer_6478 ( .C (clk), .D (new_AGEMA_signal_12329), .Q (new_AGEMA_signal_12330) ) ;
    buf_clk new_AGEMA_reg_buffer_6481 ( .C (clk), .D (new_AGEMA_signal_12332), .Q (new_AGEMA_signal_12333) ) ;
    buf_clk new_AGEMA_reg_buffer_6484 ( .C (clk), .D (new_AGEMA_signal_12335), .Q (new_AGEMA_signal_12336) ) ;
    buf_clk new_AGEMA_reg_buffer_6487 ( .C (clk), .D (new_AGEMA_signal_12338), .Q (new_AGEMA_signal_12339) ) ;
    buf_clk new_AGEMA_reg_buffer_6490 ( .C (clk), .D (new_AGEMA_signal_12341), .Q (new_AGEMA_signal_12342) ) ;
    buf_clk new_AGEMA_reg_buffer_6493 ( .C (clk), .D (new_AGEMA_signal_12344), .Q (new_AGEMA_signal_12345) ) ;
    buf_clk new_AGEMA_reg_buffer_6496 ( .C (clk), .D (new_AGEMA_signal_12347), .Q (new_AGEMA_signal_12348) ) ;
    buf_clk new_AGEMA_reg_buffer_6499 ( .C (clk), .D (new_AGEMA_signal_12350), .Q (new_AGEMA_signal_12351) ) ;
    buf_clk new_AGEMA_reg_buffer_6502 ( .C (clk), .D (new_AGEMA_signal_12353), .Q (new_AGEMA_signal_12354) ) ;
    buf_clk new_AGEMA_reg_buffer_6505 ( .C (clk), .D (new_AGEMA_signal_12356), .Q (new_AGEMA_signal_12357) ) ;
    buf_clk new_AGEMA_reg_buffer_6508 ( .C (clk), .D (new_AGEMA_signal_12359), .Q (new_AGEMA_signal_12360) ) ;
    buf_clk new_AGEMA_reg_buffer_6511 ( .C (clk), .D (new_AGEMA_signal_12362), .Q (new_AGEMA_signal_12363) ) ;
    buf_clk new_AGEMA_reg_buffer_6514 ( .C (clk), .D (new_AGEMA_signal_12365), .Q (new_AGEMA_signal_12366) ) ;
    buf_clk new_AGEMA_reg_buffer_6517 ( .C (clk), .D (new_AGEMA_signal_12368), .Q (new_AGEMA_signal_12369) ) ;
    buf_clk new_AGEMA_reg_buffer_6520 ( .C (clk), .D (new_AGEMA_signal_12371), .Q (new_AGEMA_signal_12372) ) ;
    buf_clk new_AGEMA_reg_buffer_6523 ( .C (clk), .D (new_AGEMA_signal_12374), .Q (new_AGEMA_signal_12375) ) ;
    buf_clk new_AGEMA_reg_buffer_6526 ( .C (clk), .D (new_AGEMA_signal_12377), .Q (new_AGEMA_signal_12378) ) ;
    buf_clk new_AGEMA_reg_buffer_6529 ( .C (clk), .D (new_AGEMA_signal_12380), .Q (new_AGEMA_signal_12381) ) ;
    buf_clk new_AGEMA_reg_buffer_6532 ( .C (clk), .D (new_AGEMA_signal_12383), .Q (new_AGEMA_signal_12384) ) ;
    buf_clk new_AGEMA_reg_buffer_6535 ( .C (clk), .D (new_AGEMA_signal_12386), .Q (new_AGEMA_signal_12387) ) ;
    buf_clk new_AGEMA_reg_buffer_6538 ( .C (clk), .D (new_AGEMA_signal_12389), .Q (new_AGEMA_signal_12390) ) ;
    buf_clk new_AGEMA_reg_buffer_6541 ( .C (clk), .D (new_AGEMA_signal_12392), .Q (new_AGEMA_signal_12393) ) ;
    buf_clk new_AGEMA_reg_buffer_6544 ( .C (clk), .D (new_AGEMA_signal_12395), .Q (new_AGEMA_signal_12396) ) ;
    buf_clk new_AGEMA_reg_buffer_6547 ( .C (clk), .D (new_AGEMA_signal_12398), .Q (new_AGEMA_signal_12399) ) ;
    buf_clk new_AGEMA_reg_buffer_6550 ( .C (clk), .D (new_AGEMA_signal_12401), .Q (new_AGEMA_signal_12402) ) ;
    buf_clk new_AGEMA_reg_buffer_6553 ( .C (clk), .D (new_AGEMA_signal_12404), .Q (new_AGEMA_signal_12405) ) ;
    buf_clk new_AGEMA_reg_buffer_6556 ( .C (clk), .D (new_AGEMA_signal_12407), .Q (new_AGEMA_signal_12408) ) ;
    buf_clk new_AGEMA_reg_buffer_6559 ( .C (clk), .D (new_AGEMA_signal_12410), .Q (new_AGEMA_signal_12411) ) ;
    buf_clk new_AGEMA_reg_buffer_6562 ( .C (clk), .D (new_AGEMA_signal_12413), .Q (new_AGEMA_signal_12414) ) ;
    buf_clk new_AGEMA_reg_buffer_6565 ( .C (clk), .D (new_AGEMA_signal_12416), .Q (new_AGEMA_signal_12417) ) ;
    buf_clk new_AGEMA_reg_buffer_6568 ( .C (clk), .D (new_AGEMA_signal_12419), .Q (new_AGEMA_signal_12420) ) ;
    buf_clk new_AGEMA_reg_buffer_6571 ( .C (clk), .D (new_AGEMA_signal_12422), .Q (new_AGEMA_signal_12423) ) ;
    buf_clk new_AGEMA_reg_buffer_6574 ( .C (clk), .D (new_AGEMA_signal_12425), .Q (new_AGEMA_signal_12426) ) ;
    buf_clk new_AGEMA_reg_buffer_6577 ( .C (clk), .D (new_AGEMA_signal_12428), .Q (new_AGEMA_signal_12429) ) ;
    buf_clk new_AGEMA_reg_buffer_6580 ( .C (clk), .D (new_AGEMA_signal_12431), .Q (new_AGEMA_signal_12432) ) ;
    buf_clk new_AGEMA_reg_buffer_6583 ( .C (clk), .D (new_AGEMA_signal_12434), .Q (new_AGEMA_signal_12435) ) ;
    buf_clk new_AGEMA_reg_buffer_6586 ( .C (clk), .D (new_AGEMA_signal_12437), .Q (new_AGEMA_signal_12438) ) ;
    buf_clk new_AGEMA_reg_buffer_6589 ( .C (clk), .D (new_AGEMA_signal_12440), .Q (new_AGEMA_signal_12441) ) ;
    buf_clk new_AGEMA_reg_buffer_6592 ( .C (clk), .D (new_AGEMA_signal_12443), .Q (new_AGEMA_signal_12444) ) ;
    buf_clk new_AGEMA_reg_buffer_6595 ( .C (clk), .D (new_AGEMA_signal_12446), .Q (new_AGEMA_signal_12447) ) ;
    buf_clk new_AGEMA_reg_buffer_6598 ( .C (clk), .D (new_AGEMA_signal_12449), .Q (new_AGEMA_signal_12450) ) ;
    buf_clk new_AGEMA_reg_buffer_6601 ( .C (clk), .D (new_AGEMA_signal_12452), .Q (new_AGEMA_signal_12453) ) ;
    buf_clk new_AGEMA_reg_buffer_6604 ( .C (clk), .D (new_AGEMA_signal_12455), .Q (new_AGEMA_signal_12456) ) ;
    buf_clk new_AGEMA_reg_buffer_6607 ( .C (clk), .D (new_AGEMA_signal_12458), .Q (new_AGEMA_signal_12459) ) ;
    buf_clk new_AGEMA_reg_buffer_6610 ( .C (clk), .D (new_AGEMA_signal_12461), .Q (new_AGEMA_signal_12462) ) ;
    buf_clk new_AGEMA_reg_buffer_6613 ( .C (clk), .D (new_AGEMA_signal_12464), .Q (new_AGEMA_signal_12465) ) ;
    buf_clk new_AGEMA_reg_buffer_6616 ( .C (clk), .D (new_AGEMA_signal_12467), .Q (new_AGEMA_signal_12468) ) ;
    buf_clk new_AGEMA_reg_buffer_6619 ( .C (clk), .D (new_AGEMA_signal_12470), .Q (new_AGEMA_signal_12471) ) ;
    buf_clk new_AGEMA_reg_buffer_6622 ( .C (clk), .D (new_AGEMA_signal_12473), .Q (new_AGEMA_signal_12474) ) ;
    buf_clk new_AGEMA_reg_buffer_6625 ( .C (clk), .D (new_AGEMA_signal_12476), .Q (new_AGEMA_signal_12477) ) ;
    buf_clk new_AGEMA_reg_buffer_6628 ( .C (clk), .D (new_AGEMA_signal_12479), .Q (new_AGEMA_signal_12480) ) ;
    buf_clk new_AGEMA_reg_buffer_6631 ( .C (clk), .D (new_AGEMA_signal_12482), .Q (new_AGEMA_signal_12483) ) ;
    buf_clk new_AGEMA_reg_buffer_6634 ( .C (clk), .D (new_AGEMA_signal_12485), .Q (new_AGEMA_signal_12486) ) ;
    buf_clk new_AGEMA_reg_buffer_6637 ( .C (clk), .D (new_AGEMA_signal_12488), .Q (new_AGEMA_signal_12489) ) ;
    buf_clk new_AGEMA_reg_buffer_6640 ( .C (clk), .D (new_AGEMA_signal_12491), .Q (new_AGEMA_signal_12492) ) ;
    buf_clk new_AGEMA_reg_buffer_6643 ( .C (clk), .D (new_AGEMA_signal_12494), .Q (new_AGEMA_signal_12495) ) ;
    buf_clk new_AGEMA_reg_buffer_6646 ( .C (clk), .D (new_AGEMA_signal_12497), .Q (new_AGEMA_signal_12498) ) ;
    buf_clk new_AGEMA_reg_buffer_6649 ( .C (clk), .D (new_AGEMA_signal_12500), .Q (new_AGEMA_signal_12501) ) ;
    buf_clk new_AGEMA_reg_buffer_6652 ( .C (clk), .D (new_AGEMA_signal_12503), .Q (new_AGEMA_signal_12504) ) ;
    buf_clk new_AGEMA_reg_buffer_6655 ( .C (clk), .D (new_AGEMA_signal_12506), .Q (new_AGEMA_signal_12507) ) ;
    buf_clk new_AGEMA_reg_buffer_6658 ( .C (clk), .D (new_AGEMA_signal_12509), .Q (new_AGEMA_signal_12510) ) ;
    buf_clk new_AGEMA_reg_buffer_6661 ( .C (clk), .D (new_AGEMA_signal_12512), .Q (new_AGEMA_signal_12513) ) ;
    buf_clk new_AGEMA_reg_buffer_6664 ( .C (clk), .D (new_AGEMA_signal_12515), .Q (new_AGEMA_signal_12516) ) ;
    buf_clk new_AGEMA_reg_buffer_6667 ( .C (clk), .D (new_AGEMA_signal_12518), .Q (new_AGEMA_signal_12519) ) ;
    buf_clk new_AGEMA_reg_buffer_6670 ( .C (clk), .D (new_AGEMA_signal_12521), .Q (new_AGEMA_signal_12522) ) ;
    buf_clk new_AGEMA_reg_buffer_6673 ( .C (clk), .D (new_AGEMA_signal_12524), .Q (new_AGEMA_signal_12525) ) ;
    buf_clk new_AGEMA_reg_buffer_6676 ( .C (clk), .D (new_AGEMA_signal_12527), .Q (new_AGEMA_signal_12528) ) ;
    buf_clk new_AGEMA_reg_buffer_6679 ( .C (clk), .D (new_AGEMA_signal_12530), .Q (new_AGEMA_signal_12531) ) ;
    buf_clk new_AGEMA_reg_buffer_6682 ( .C (clk), .D (new_AGEMA_signal_12533), .Q (new_AGEMA_signal_12534) ) ;
    buf_clk new_AGEMA_reg_buffer_6685 ( .C (clk), .D (new_AGEMA_signal_12536), .Q (new_AGEMA_signal_12537) ) ;
    buf_clk new_AGEMA_reg_buffer_6688 ( .C (clk), .D (new_AGEMA_signal_12539), .Q (new_AGEMA_signal_12540) ) ;
    buf_clk new_AGEMA_reg_buffer_6691 ( .C (clk), .D (new_AGEMA_signal_12542), .Q (new_AGEMA_signal_12543) ) ;
    buf_clk new_AGEMA_reg_buffer_6694 ( .C (clk), .D (new_AGEMA_signal_12545), .Q (new_AGEMA_signal_12546) ) ;
    buf_clk new_AGEMA_reg_buffer_6697 ( .C (clk), .D (new_AGEMA_signal_12548), .Q (new_AGEMA_signal_12549) ) ;
    buf_clk new_AGEMA_reg_buffer_6700 ( .C (clk), .D (new_AGEMA_signal_12551), .Q (new_AGEMA_signal_12552) ) ;
    buf_clk new_AGEMA_reg_buffer_6703 ( .C (clk), .D (new_AGEMA_signal_12554), .Q (new_AGEMA_signal_12555) ) ;
    buf_clk new_AGEMA_reg_buffer_6706 ( .C (clk), .D (new_AGEMA_signal_12557), .Q (new_AGEMA_signal_12558) ) ;
    buf_clk new_AGEMA_reg_buffer_6709 ( .C (clk), .D (new_AGEMA_signal_12560), .Q (new_AGEMA_signal_12561) ) ;
    buf_clk new_AGEMA_reg_buffer_6712 ( .C (clk), .D (new_AGEMA_signal_12563), .Q (new_AGEMA_signal_12564) ) ;
    buf_clk new_AGEMA_reg_buffer_6715 ( .C (clk), .D (new_AGEMA_signal_12566), .Q (new_AGEMA_signal_12567) ) ;
    buf_clk new_AGEMA_reg_buffer_6718 ( .C (clk), .D (new_AGEMA_signal_12569), .Q (new_AGEMA_signal_12570) ) ;
    buf_clk new_AGEMA_reg_buffer_6721 ( .C (clk), .D (new_AGEMA_signal_12572), .Q (new_AGEMA_signal_12573) ) ;
    buf_clk new_AGEMA_reg_buffer_6724 ( .C (clk), .D (new_AGEMA_signal_12575), .Q (new_AGEMA_signal_12576) ) ;
    buf_clk new_AGEMA_reg_buffer_6727 ( .C (clk), .D (new_AGEMA_signal_12578), .Q (new_AGEMA_signal_12579) ) ;
    buf_clk new_AGEMA_reg_buffer_6730 ( .C (clk), .D (new_AGEMA_signal_12581), .Q (new_AGEMA_signal_12582) ) ;
    buf_clk new_AGEMA_reg_buffer_6733 ( .C (clk), .D (new_AGEMA_signal_12584), .Q (new_AGEMA_signal_12585) ) ;
    buf_clk new_AGEMA_reg_buffer_6736 ( .C (clk), .D (new_AGEMA_signal_12587), .Q (new_AGEMA_signal_12588) ) ;
    buf_clk new_AGEMA_reg_buffer_6739 ( .C (clk), .D (new_AGEMA_signal_12590), .Q (new_AGEMA_signal_12591) ) ;
    buf_clk new_AGEMA_reg_buffer_6742 ( .C (clk), .D (new_AGEMA_signal_12593), .Q (new_AGEMA_signal_12594) ) ;
    buf_clk new_AGEMA_reg_buffer_6745 ( .C (clk), .D (new_AGEMA_signal_12596), .Q (new_AGEMA_signal_12597) ) ;
    buf_clk new_AGEMA_reg_buffer_6748 ( .C (clk), .D (new_AGEMA_signal_12599), .Q (new_AGEMA_signal_12600) ) ;
    buf_clk new_AGEMA_reg_buffer_6751 ( .C (clk), .D (new_AGEMA_signal_12602), .Q (new_AGEMA_signal_12603) ) ;
    buf_clk new_AGEMA_reg_buffer_6754 ( .C (clk), .D (new_AGEMA_signal_12605), .Q (new_AGEMA_signal_12606) ) ;
    buf_clk new_AGEMA_reg_buffer_6757 ( .C (clk), .D (new_AGEMA_signal_12608), .Q (new_AGEMA_signal_12609) ) ;
    buf_clk new_AGEMA_reg_buffer_6760 ( .C (clk), .D (new_AGEMA_signal_12611), .Q (new_AGEMA_signal_12612) ) ;
    buf_clk new_AGEMA_reg_buffer_6763 ( .C (clk), .D (new_AGEMA_signal_12614), .Q (new_AGEMA_signal_12615) ) ;
    buf_clk new_AGEMA_reg_buffer_6766 ( .C (clk), .D (new_AGEMA_signal_12617), .Q (new_AGEMA_signal_12618) ) ;
    buf_clk new_AGEMA_reg_buffer_6769 ( .C (clk), .D (new_AGEMA_signal_12620), .Q (new_AGEMA_signal_12621) ) ;
    buf_clk new_AGEMA_reg_buffer_6772 ( .C (clk), .D (new_AGEMA_signal_12623), .Q (new_AGEMA_signal_12624) ) ;
    buf_clk new_AGEMA_reg_buffer_6775 ( .C (clk), .D (new_AGEMA_signal_12626), .Q (new_AGEMA_signal_12627) ) ;
    buf_clk new_AGEMA_reg_buffer_6778 ( .C (clk), .D (new_AGEMA_signal_12629), .Q (new_AGEMA_signal_12630) ) ;
    buf_clk new_AGEMA_reg_buffer_6781 ( .C (clk), .D (new_AGEMA_signal_12632), .Q (new_AGEMA_signal_12633) ) ;
    buf_clk new_AGEMA_reg_buffer_6784 ( .C (clk), .D (new_AGEMA_signal_12635), .Q (new_AGEMA_signal_12636) ) ;
    buf_clk new_AGEMA_reg_buffer_6787 ( .C (clk), .D (new_AGEMA_signal_12638), .Q (new_AGEMA_signal_12639) ) ;
    buf_clk new_AGEMA_reg_buffer_6790 ( .C (clk), .D (new_AGEMA_signal_12641), .Q (new_AGEMA_signal_12642) ) ;
    buf_clk new_AGEMA_reg_buffer_6793 ( .C (clk), .D (new_AGEMA_signal_12644), .Q (new_AGEMA_signal_12645) ) ;
    buf_clk new_AGEMA_reg_buffer_6796 ( .C (clk), .D (new_AGEMA_signal_12647), .Q (new_AGEMA_signal_12648) ) ;
    buf_clk new_AGEMA_reg_buffer_6799 ( .C (clk), .D (new_AGEMA_signal_12650), .Q (new_AGEMA_signal_12651) ) ;
    buf_clk new_AGEMA_reg_buffer_6802 ( .C (clk), .D (new_AGEMA_signal_12653), .Q (new_AGEMA_signal_12654) ) ;
    buf_clk new_AGEMA_reg_buffer_6805 ( .C (clk), .D (new_AGEMA_signal_12656), .Q (new_AGEMA_signal_12657) ) ;
    buf_clk new_AGEMA_reg_buffer_6808 ( .C (clk), .D (new_AGEMA_signal_12659), .Q (new_AGEMA_signal_12660) ) ;
    buf_clk new_AGEMA_reg_buffer_6811 ( .C (clk), .D (new_AGEMA_signal_12662), .Q (new_AGEMA_signal_12663) ) ;
    buf_clk new_AGEMA_reg_buffer_6814 ( .C (clk), .D (new_AGEMA_signal_12665), .Q (new_AGEMA_signal_12666) ) ;
    buf_clk new_AGEMA_reg_buffer_6817 ( .C (clk), .D (new_AGEMA_signal_12668), .Q (new_AGEMA_signal_12669) ) ;
    buf_clk new_AGEMA_reg_buffer_6820 ( .C (clk), .D (new_AGEMA_signal_12671), .Q (new_AGEMA_signal_12672) ) ;
    buf_clk new_AGEMA_reg_buffer_6823 ( .C (clk), .D (new_AGEMA_signal_12674), .Q (new_AGEMA_signal_12675) ) ;
    buf_clk new_AGEMA_reg_buffer_6826 ( .C (clk), .D (new_AGEMA_signal_12677), .Q (new_AGEMA_signal_12678) ) ;
    buf_clk new_AGEMA_reg_buffer_6829 ( .C (clk), .D (new_AGEMA_signal_12680), .Q (new_AGEMA_signal_12681) ) ;
    buf_clk new_AGEMA_reg_buffer_6832 ( .C (clk), .D (new_AGEMA_signal_12683), .Q (new_AGEMA_signal_12684) ) ;
    buf_clk new_AGEMA_reg_buffer_6835 ( .C (clk), .D (new_AGEMA_signal_12686), .Q (new_AGEMA_signal_12687) ) ;
    buf_clk new_AGEMA_reg_buffer_6838 ( .C (clk), .D (new_AGEMA_signal_12689), .Q (new_AGEMA_signal_12690) ) ;
    buf_clk new_AGEMA_reg_buffer_6841 ( .C (clk), .D (new_AGEMA_signal_12692), .Q (new_AGEMA_signal_12693) ) ;
    buf_clk new_AGEMA_reg_buffer_6844 ( .C (clk), .D (new_AGEMA_signal_12695), .Q (new_AGEMA_signal_12696) ) ;
    buf_clk new_AGEMA_reg_buffer_6847 ( .C (clk), .D (new_AGEMA_signal_12698), .Q (new_AGEMA_signal_12699) ) ;
    buf_clk new_AGEMA_reg_buffer_6850 ( .C (clk), .D (new_AGEMA_signal_12701), .Q (new_AGEMA_signal_12702) ) ;
    buf_clk new_AGEMA_reg_buffer_6853 ( .C (clk), .D (new_AGEMA_signal_12704), .Q (new_AGEMA_signal_12705) ) ;
    buf_clk new_AGEMA_reg_buffer_6856 ( .C (clk), .D (new_AGEMA_signal_12707), .Q (new_AGEMA_signal_12708) ) ;
    buf_clk new_AGEMA_reg_buffer_6859 ( .C (clk), .D (new_AGEMA_signal_12710), .Q (new_AGEMA_signal_12711) ) ;
    buf_clk new_AGEMA_reg_buffer_6862 ( .C (clk), .D (new_AGEMA_signal_12713), .Q (new_AGEMA_signal_12714) ) ;
    buf_clk new_AGEMA_reg_buffer_6865 ( .C (clk), .D (new_AGEMA_signal_12716), .Q (new_AGEMA_signal_12717) ) ;
    buf_clk new_AGEMA_reg_buffer_6868 ( .C (clk), .D (new_AGEMA_signal_12719), .Q (new_AGEMA_signal_12720) ) ;
    buf_clk new_AGEMA_reg_buffer_6871 ( .C (clk), .D (new_AGEMA_signal_12722), .Q (new_AGEMA_signal_12723) ) ;
    buf_clk new_AGEMA_reg_buffer_6874 ( .C (clk), .D (new_AGEMA_signal_12725), .Q (new_AGEMA_signal_12726) ) ;
    buf_clk new_AGEMA_reg_buffer_6877 ( .C (clk), .D (new_AGEMA_signal_12728), .Q (new_AGEMA_signal_12729) ) ;
    buf_clk new_AGEMA_reg_buffer_6880 ( .C (clk), .D (new_AGEMA_signal_12731), .Q (new_AGEMA_signal_12732) ) ;
    buf_clk new_AGEMA_reg_buffer_6883 ( .C (clk), .D (new_AGEMA_signal_12734), .Q (new_AGEMA_signal_12735) ) ;
    buf_clk new_AGEMA_reg_buffer_6886 ( .C (clk), .D (new_AGEMA_signal_12737), .Q (new_AGEMA_signal_12738) ) ;
    buf_clk new_AGEMA_reg_buffer_6889 ( .C (clk), .D (new_AGEMA_signal_12740), .Q (new_AGEMA_signal_12741) ) ;
    buf_clk new_AGEMA_reg_buffer_6892 ( .C (clk), .D (new_AGEMA_signal_12743), .Q (new_AGEMA_signal_12744) ) ;
    buf_clk new_AGEMA_reg_buffer_6895 ( .C (clk), .D (new_AGEMA_signal_12746), .Q (new_AGEMA_signal_12747) ) ;
    buf_clk new_AGEMA_reg_buffer_6898 ( .C (clk), .D (new_AGEMA_signal_12749), .Q (new_AGEMA_signal_12750) ) ;
    buf_clk new_AGEMA_reg_buffer_6901 ( .C (clk), .D (new_AGEMA_signal_12752), .Q (new_AGEMA_signal_12753) ) ;
    buf_clk new_AGEMA_reg_buffer_6904 ( .C (clk), .D (new_AGEMA_signal_12755), .Q (new_AGEMA_signal_12756) ) ;
    buf_clk new_AGEMA_reg_buffer_6907 ( .C (clk), .D (new_AGEMA_signal_12758), .Q (new_AGEMA_signal_12759) ) ;
    buf_clk new_AGEMA_reg_buffer_6910 ( .C (clk), .D (new_AGEMA_signal_12761), .Q (new_AGEMA_signal_12762) ) ;
    buf_clk new_AGEMA_reg_buffer_6913 ( .C (clk), .D (new_AGEMA_signal_12764), .Q (new_AGEMA_signal_12765) ) ;
    buf_clk new_AGEMA_reg_buffer_6916 ( .C (clk), .D (new_AGEMA_signal_12767), .Q (new_AGEMA_signal_12768) ) ;
    buf_clk new_AGEMA_reg_buffer_6919 ( .C (clk), .D (new_AGEMA_signal_12770), .Q (new_AGEMA_signal_12771) ) ;
    buf_clk new_AGEMA_reg_buffer_6922 ( .C (clk), .D (new_AGEMA_signal_12773), .Q (new_AGEMA_signal_12774) ) ;
    buf_clk new_AGEMA_reg_buffer_6925 ( .C (clk), .D (new_AGEMA_signal_12776), .Q (new_AGEMA_signal_12777) ) ;
    buf_clk new_AGEMA_reg_buffer_6928 ( .C (clk), .D (new_AGEMA_signal_12779), .Q (new_AGEMA_signal_12780) ) ;
    buf_clk new_AGEMA_reg_buffer_6931 ( .C (clk), .D (new_AGEMA_signal_12782), .Q (new_AGEMA_signal_12783) ) ;
    buf_clk new_AGEMA_reg_buffer_6934 ( .C (clk), .D (new_AGEMA_signal_12785), .Q (new_AGEMA_signal_12786) ) ;
    buf_clk new_AGEMA_reg_buffer_6937 ( .C (clk), .D (new_AGEMA_signal_12788), .Q (new_AGEMA_signal_12789) ) ;
    buf_clk new_AGEMA_reg_buffer_6940 ( .C (clk), .D (new_AGEMA_signal_12791), .Q (new_AGEMA_signal_12792) ) ;
    buf_clk new_AGEMA_reg_buffer_6943 ( .C (clk), .D (new_AGEMA_signal_12794), .Q (new_AGEMA_signal_12795) ) ;
    buf_clk new_AGEMA_reg_buffer_6946 ( .C (clk), .D (new_AGEMA_signal_12797), .Q (new_AGEMA_signal_12798) ) ;
    buf_clk new_AGEMA_reg_buffer_6949 ( .C (clk), .D (new_AGEMA_signal_12800), .Q (new_AGEMA_signal_12801) ) ;
    buf_clk new_AGEMA_reg_buffer_6952 ( .C (clk), .D (new_AGEMA_signal_12803), .Q (new_AGEMA_signal_12804) ) ;
    buf_clk new_AGEMA_reg_buffer_6955 ( .C (clk), .D (new_AGEMA_signal_12806), .Q (new_AGEMA_signal_12807) ) ;
    buf_clk new_AGEMA_reg_buffer_6958 ( .C (clk), .D (new_AGEMA_signal_12809), .Q (new_AGEMA_signal_12810) ) ;
    buf_clk new_AGEMA_reg_buffer_6961 ( .C (clk), .D (new_AGEMA_signal_12812), .Q (new_AGEMA_signal_12813) ) ;
    buf_clk new_AGEMA_reg_buffer_6964 ( .C (clk), .D (new_AGEMA_signal_12815), .Q (new_AGEMA_signal_12816) ) ;
    buf_clk new_AGEMA_reg_buffer_6967 ( .C (clk), .D (new_AGEMA_signal_12818), .Q (new_AGEMA_signal_12819) ) ;
    buf_clk new_AGEMA_reg_buffer_6970 ( .C (clk), .D (new_AGEMA_signal_12821), .Q (new_AGEMA_signal_12822) ) ;
    buf_clk new_AGEMA_reg_buffer_6973 ( .C (clk), .D (new_AGEMA_signal_12824), .Q (new_AGEMA_signal_12825) ) ;
    buf_clk new_AGEMA_reg_buffer_6976 ( .C (clk), .D (new_AGEMA_signal_12827), .Q (new_AGEMA_signal_12828) ) ;
    buf_clk new_AGEMA_reg_buffer_6979 ( .C (clk), .D (new_AGEMA_signal_12830), .Q (new_AGEMA_signal_12831) ) ;
    buf_clk new_AGEMA_reg_buffer_6982 ( .C (clk), .D (new_AGEMA_signal_12833), .Q (new_AGEMA_signal_12834) ) ;
    buf_clk new_AGEMA_reg_buffer_6985 ( .C (clk), .D (new_AGEMA_signal_12836), .Q (new_AGEMA_signal_12837) ) ;
    buf_clk new_AGEMA_reg_buffer_6988 ( .C (clk), .D (new_AGEMA_signal_12839), .Q (new_AGEMA_signal_12840) ) ;
    buf_clk new_AGEMA_reg_buffer_6991 ( .C (clk), .D (new_AGEMA_signal_12842), .Q (new_AGEMA_signal_12843) ) ;
    buf_clk new_AGEMA_reg_buffer_6994 ( .C (clk), .D (new_AGEMA_signal_12845), .Q (new_AGEMA_signal_12846) ) ;
    buf_clk new_AGEMA_reg_buffer_6997 ( .C (clk), .D (new_AGEMA_signal_12848), .Q (new_AGEMA_signal_12849) ) ;
    buf_clk new_AGEMA_reg_buffer_7000 ( .C (clk), .D (new_AGEMA_signal_12851), .Q (new_AGEMA_signal_12852) ) ;
    buf_clk new_AGEMA_reg_buffer_7003 ( .C (clk), .D (new_AGEMA_signal_12854), .Q (new_AGEMA_signal_12855) ) ;
    buf_clk new_AGEMA_reg_buffer_7006 ( .C (clk), .D (new_AGEMA_signal_12857), .Q (new_AGEMA_signal_12858) ) ;
    buf_clk new_AGEMA_reg_buffer_7009 ( .C (clk), .D (new_AGEMA_signal_12860), .Q (new_AGEMA_signal_12861) ) ;
    buf_clk new_AGEMA_reg_buffer_7012 ( .C (clk), .D (new_AGEMA_signal_12863), .Q (new_AGEMA_signal_12864) ) ;
    buf_clk new_AGEMA_reg_buffer_7015 ( .C (clk), .D (new_AGEMA_signal_12866), .Q (new_AGEMA_signal_12867) ) ;
    buf_clk new_AGEMA_reg_buffer_7018 ( .C (clk), .D (new_AGEMA_signal_12869), .Q (new_AGEMA_signal_12870) ) ;
    buf_clk new_AGEMA_reg_buffer_7021 ( .C (clk), .D (new_AGEMA_signal_12872), .Q (new_AGEMA_signal_12873) ) ;
    buf_clk new_AGEMA_reg_buffer_7024 ( .C (clk), .D (new_AGEMA_signal_12875), .Q (new_AGEMA_signal_12876) ) ;
    buf_clk new_AGEMA_reg_buffer_7027 ( .C (clk), .D (new_AGEMA_signal_12878), .Q (new_AGEMA_signal_12879) ) ;
    buf_clk new_AGEMA_reg_buffer_7030 ( .C (clk), .D (new_AGEMA_signal_12881), .Q (new_AGEMA_signal_12882) ) ;
    buf_clk new_AGEMA_reg_buffer_7033 ( .C (clk), .D (new_AGEMA_signal_12884), .Q (new_AGEMA_signal_12885) ) ;
    buf_clk new_AGEMA_reg_buffer_7036 ( .C (clk), .D (new_AGEMA_signal_12887), .Q (new_AGEMA_signal_12888) ) ;
    buf_clk new_AGEMA_reg_buffer_7039 ( .C (clk), .D (new_AGEMA_signal_12890), .Q (new_AGEMA_signal_12891) ) ;
    buf_clk new_AGEMA_reg_buffer_7042 ( .C (clk), .D (new_AGEMA_signal_12893), .Q (new_AGEMA_signal_12894) ) ;
    buf_clk new_AGEMA_reg_buffer_7045 ( .C (clk), .D (new_AGEMA_signal_12896), .Q (new_AGEMA_signal_12897) ) ;
    buf_clk new_AGEMA_reg_buffer_7048 ( .C (clk), .D (new_AGEMA_signal_12899), .Q (new_AGEMA_signal_12900) ) ;
    buf_clk new_AGEMA_reg_buffer_7051 ( .C (clk), .D (new_AGEMA_signal_12902), .Q (new_AGEMA_signal_12903) ) ;
    buf_clk new_AGEMA_reg_buffer_7054 ( .C (clk), .D (new_AGEMA_signal_12905), .Q (new_AGEMA_signal_12906) ) ;
    buf_clk new_AGEMA_reg_buffer_7057 ( .C (clk), .D (new_AGEMA_signal_12908), .Q (new_AGEMA_signal_12909) ) ;
    buf_clk new_AGEMA_reg_buffer_7060 ( .C (clk), .D (new_AGEMA_signal_12911), .Q (new_AGEMA_signal_12912) ) ;
    buf_clk new_AGEMA_reg_buffer_7063 ( .C (clk), .D (new_AGEMA_signal_12914), .Q (new_AGEMA_signal_12915) ) ;
    buf_clk new_AGEMA_reg_buffer_7066 ( .C (clk), .D (new_AGEMA_signal_12917), .Q (new_AGEMA_signal_12918) ) ;
    buf_clk new_AGEMA_reg_buffer_7069 ( .C (clk), .D (new_AGEMA_signal_12920), .Q (new_AGEMA_signal_12921) ) ;
    buf_clk new_AGEMA_reg_buffer_7072 ( .C (clk), .D (new_AGEMA_signal_12923), .Q (new_AGEMA_signal_12924) ) ;
    buf_clk new_AGEMA_reg_buffer_7075 ( .C (clk), .D (new_AGEMA_signal_12926), .Q (new_AGEMA_signal_12927) ) ;
    buf_clk new_AGEMA_reg_buffer_7078 ( .C (clk), .D (new_AGEMA_signal_12929), .Q (new_AGEMA_signal_12930) ) ;
    buf_clk new_AGEMA_reg_buffer_7081 ( .C (clk), .D (new_AGEMA_signal_12932), .Q (new_AGEMA_signal_12933) ) ;
    buf_clk new_AGEMA_reg_buffer_7084 ( .C (clk), .D (new_AGEMA_signal_12935), .Q (new_AGEMA_signal_12936) ) ;
    buf_clk new_AGEMA_reg_buffer_7087 ( .C (clk), .D (new_AGEMA_signal_12938), .Q (new_AGEMA_signal_12939) ) ;
    buf_clk new_AGEMA_reg_buffer_7090 ( .C (clk), .D (new_AGEMA_signal_12941), .Q (new_AGEMA_signal_12942) ) ;
    buf_clk new_AGEMA_reg_buffer_7093 ( .C (clk), .D (new_AGEMA_signal_12944), .Q (new_AGEMA_signal_12945) ) ;
    buf_clk new_AGEMA_reg_buffer_7096 ( .C (clk), .D (new_AGEMA_signal_12947), .Q (new_AGEMA_signal_12948) ) ;
    buf_clk new_AGEMA_reg_buffer_7099 ( .C (clk), .D (new_AGEMA_signal_12950), .Q (new_AGEMA_signal_12951) ) ;
    buf_clk new_AGEMA_reg_buffer_7102 ( .C (clk), .D (new_AGEMA_signal_12953), .Q (new_AGEMA_signal_12954) ) ;
    buf_clk new_AGEMA_reg_buffer_7105 ( .C (clk), .D (new_AGEMA_signal_12956), .Q (new_AGEMA_signal_12957) ) ;
    buf_clk new_AGEMA_reg_buffer_7108 ( .C (clk), .D (new_AGEMA_signal_12959), .Q (new_AGEMA_signal_12960) ) ;
    buf_clk new_AGEMA_reg_buffer_7111 ( .C (clk), .D (new_AGEMA_signal_12962), .Q (new_AGEMA_signal_12963) ) ;
    buf_clk new_AGEMA_reg_buffer_7114 ( .C (clk), .D (new_AGEMA_signal_12965), .Q (new_AGEMA_signal_12966) ) ;
    buf_clk new_AGEMA_reg_buffer_7117 ( .C (clk), .D (new_AGEMA_signal_12968), .Q (new_AGEMA_signal_12969) ) ;
    buf_clk new_AGEMA_reg_buffer_7120 ( .C (clk), .D (new_AGEMA_signal_12971), .Q (new_AGEMA_signal_12972) ) ;
    buf_clk new_AGEMA_reg_buffer_7123 ( .C (clk), .D (new_AGEMA_signal_12974), .Q (new_AGEMA_signal_12975) ) ;
    buf_clk new_AGEMA_reg_buffer_7126 ( .C (clk), .D (new_AGEMA_signal_12977), .Q (new_AGEMA_signal_12978) ) ;
    buf_clk new_AGEMA_reg_buffer_7129 ( .C (clk), .D (new_AGEMA_signal_12980), .Q (new_AGEMA_signal_12981) ) ;
    buf_clk new_AGEMA_reg_buffer_7132 ( .C (clk), .D (new_AGEMA_signal_12983), .Q (new_AGEMA_signal_12984) ) ;
    buf_clk new_AGEMA_reg_buffer_7135 ( .C (clk), .D (new_AGEMA_signal_12986), .Q (new_AGEMA_signal_12987) ) ;
    buf_clk new_AGEMA_reg_buffer_7138 ( .C (clk), .D (new_AGEMA_signal_12989), .Q (new_AGEMA_signal_12990) ) ;
    buf_clk new_AGEMA_reg_buffer_7141 ( .C (clk), .D (new_AGEMA_signal_12992), .Q (new_AGEMA_signal_12993) ) ;
    buf_clk new_AGEMA_reg_buffer_7144 ( .C (clk), .D (new_AGEMA_signal_12995), .Q (new_AGEMA_signal_12996) ) ;
    buf_clk new_AGEMA_reg_buffer_7147 ( .C (clk), .D (new_AGEMA_signal_12998), .Q (new_AGEMA_signal_12999) ) ;
    buf_clk new_AGEMA_reg_buffer_7150 ( .C (clk), .D (new_AGEMA_signal_13001), .Q (new_AGEMA_signal_13002) ) ;
    buf_clk new_AGEMA_reg_buffer_7153 ( .C (clk), .D (new_AGEMA_signal_13004), .Q (new_AGEMA_signal_13005) ) ;
    buf_clk new_AGEMA_reg_buffer_7156 ( .C (clk), .D (new_AGEMA_signal_13007), .Q (new_AGEMA_signal_13008) ) ;
    buf_clk new_AGEMA_reg_buffer_7159 ( .C (clk), .D (new_AGEMA_signal_13010), .Q (new_AGEMA_signal_13011) ) ;
    buf_clk new_AGEMA_reg_buffer_7162 ( .C (clk), .D (new_AGEMA_signal_13013), .Q (new_AGEMA_signal_13014) ) ;
    buf_clk new_AGEMA_reg_buffer_7165 ( .C (clk), .D (new_AGEMA_signal_13016), .Q (new_AGEMA_signal_13017) ) ;
    buf_clk new_AGEMA_reg_buffer_7168 ( .C (clk), .D (new_AGEMA_signal_13019), .Q (new_AGEMA_signal_13020) ) ;
    buf_clk new_AGEMA_reg_buffer_7171 ( .C (clk), .D (new_AGEMA_signal_13022), .Q (new_AGEMA_signal_13023) ) ;
    buf_clk new_AGEMA_reg_buffer_7174 ( .C (clk), .D (new_AGEMA_signal_13025), .Q (new_AGEMA_signal_13026) ) ;
    buf_clk new_AGEMA_reg_buffer_7177 ( .C (clk), .D (new_AGEMA_signal_13028), .Q (new_AGEMA_signal_13029) ) ;
    buf_clk new_AGEMA_reg_buffer_7180 ( .C (clk), .D (new_AGEMA_signal_13031), .Q (new_AGEMA_signal_13032) ) ;
    buf_clk new_AGEMA_reg_buffer_7183 ( .C (clk), .D (new_AGEMA_signal_13034), .Q (new_AGEMA_signal_13035) ) ;
    buf_clk new_AGEMA_reg_buffer_7186 ( .C (clk), .D (new_AGEMA_signal_13037), .Q (new_AGEMA_signal_13038) ) ;
    buf_clk new_AGEMA_reg_buffer_7189 ( .C (clk), .D (new_AGEMA_signal_13040), .Q (new_AGEMA_signal_13041) ) ;
    buf_clk new_AGEMA_reg_buffer_7192 ( .C (clk), .D (new_AGEMA_signal_13043), .Q (new_AGEMA_signal_13044) ) ;
    buf_clk new_AGEMA_reg_buffer_7195 ( .C (clk), .D (new_AGEMA_signal_13046), .Q (new_AGEMA_signal_13047) ) ;
    buf_clk new_AGEMA_reg_buffer_7198 ( .C (clk), .D (new_AGEMA_signal_13049), .Q (new_AGEMA_signal_13050) ) ;
    buf_clk new_AGEMA_reg_buffer_7201 ( .C (clk), .D (new_AGEMA_signal_13052), .Q (new_AGEMA_signal_13053) ) ;
    buf_clk new_AGEMA_reg_buffer_7204 ( .C (clk), .D (new_AGEMA_signal_13055), .Q (new_AGEMA_signal_13056) ) ;
    buf_clk new_AGEMA_reg_buffer_7207 ( .C (clk), .D (new_AGEMA_signal_13058), .Q (new_AGEMA_signal_13059) ) ;
    buf_clk new_AGEMA_reg_buffer_7210 ( .C (clk), .D (new_AGEMA_signal_13061), .Q (new_AGEMA_signal_13062) ) ;
    buf_clk new_AGEMA_reg_buffer_7213 ( .C (clk), .D (new_AGEMA_signal_13064), .Q (new_AGEMA_signal_13065) ) ;
    buf_clk new_AGEMA_reg_buffer_7216 ( .C (clk), .D (new_AGEMA_signal_13067), .Q (new_AGEMA_signal_13068) ) ;
    buf_clk new_AGEMA_reg_buffer_7219 ( .C (clk), .D (new_AGEMA_signal_13070), .Q (new_AGEMA_signal_13071) ) ;
    buf_clk new_AGEMA_reg_buffer_7222 ( .C (clk), .D (new_AGEMA_signal_13073), .Q (new_AGEMA_signal_13074) ) ;
    buf_clk new_AGEMA_reg_buffer_7225 ( .C (clk), .D (new_AGEMA_signal_13076), .Q (new_AGEMA_signal_13077) ) ;
    buf_clk new_AGEMA_reg_buffer_7228 ( .C (clk), .D (new_AGEMA_signal_13079), .Q (new_AGEMA_signal_13080) ) ;
    buf_clk new_AGEMA_reg_buffer_7231 ( .C (clk), .D (new_AGEMA_signal_13082), .Q (new_AGEMA_signal_13083) ) ;
    buf_clk new_AGEMA_reg_buffer_7234 ( .C (clk), .D (new_AGEMA_signal_13085), .Q (new_AGEMA_signal_13086) ) ;
    buf_clk new_AGEMA_reg_buffer_7237 ( .C (clk), .D (new_AGEMA_signal_13088), .Q (new_AGEMA_signal_13089) ) ;
    buf_clk new_AGEMA_reg_buffer_7240 ( .C (clk), .D (new_AGEMA_signal_13091), .Q (new_AGEMA_signal_13092) ) ;
    buf_clk new_AGEMA_reg_buffer_7243 ( .C (clk), .D (new_AGEMA_signal_13094), .Q (new_AGEMA_signal_13095) ) ;
    buf_clk new_AGEMA_reg_buffer_7246 ( .C (clk), .D (new_AGEMA_signal_13097), .Q (new_AGEMA_signal_13098) ) ;
    buf_clk new_AGEMA_reg_buffer_7249 ( .C (clk), .D (new_AGEMA_signal_13100), .Q (new_AGEMA_signal_13101) ) ;
    buf_clk new_AGEMA_reg_buffer_7252 ( .C (clk), .D (new_AGEMA_signal_13103), .Q (new_AGEMA_signal_13104) ) ;
    buf_clk new_AGEMA_reg_buffer_7255 ( .C (clk), .D (new_AGEMA_signal_13106), .Q (new_AGEMA_signal_13107) ) ;
    buf_clk new_AGEMA_reg_buffer_7258 ( .C (clk), .D (new_AGEMA_signal_13109), .Q (new_AGEMA_signal_13110) ) ;
    buf_clk new_AGEMA_reg_buffer_7261 ( .C (clk), .D (new_AGEMA_signal_13112), .Q (new_AGEMA_signal_13113) ) ;
    buf_clk new_AGEMA_reg_buffer_7264 ( .C (clk), .D (new_AGEMA_signal_13115), .Q (new_AGEMA_signal_13116) ) ;
    buf_clk new_AGEMA_reg_buffer_7267 ( .C (clk), .D (new_AGEMA_signal_13118), .Q (new_AGEMA_signal_13119) ) ;
    buf_clk new_AGEMA_reg_buffer_7270 ( .C (clk), .D (new_AGEMA_signal_13121), .Q (new_AGEMA_signal_13122) ) ;
    buf_clk new_AGEMA_reg_buffer_7273 ( .C (clk), .D (new_AGEMA_signal_13124), .Q (new_AGEMA_signal_13125) ) ;
    buf_clk new_AGEMA_reg_buffer_7276 ( .C (clk), .D (new_AGEMA_signal_13127), .Q (new_AGEMA_signal_13128) ) ;
    buf_clk new_AGEMA_reg_buffer_7279 ( .C (clk), .D (new_AGEMA_signal_13130), .Q (new_AGEMA_signal_13131) ) ;
    buf_clk new_AGEMA_reg_buffer_7282 ( .C (clk), .D (new_AGEMA_signal_13133), .Q (new_AGEMA_signal_13134) ) ;
    buf_clk new_AGEMA_reg_buffer_7285 ( .C (clk), .D (new_AGEMA_signal_13136), .Q (new_AGEMA_signal_13137) ) ;
    buf_clk new_AGEMA_reg_buffer_7288 ( .C (clk), .D (new_AGEMA_signal_13139), .Q (new_AGEMA_signal_13140) ) ;
    buf_clk new_AGEMA_reg_buffer_7291 ( .C (clk), .D (new_AGEMA_signal_13142), .Q (new_AGEMA_signal_13143) ) ;
    buf_clk new_AGEMA_reg_buffer_7294 ( .C (clk), .D (new_AGEMA_signal_13145), .Q (new_AGEMA_signal_13146) ) ;
    buf_clk new_AGEMA_reg_buffer_7297 ( .C (clk), .D (new_AGEMA_signal_13148), .Q (new_AGEMA_signal_13149) ) ;
    buf_clk new_AGEMA_reg_buffer_7300 ( .C (clk), .D (new_AGEMA_signal_13151), .Q (new_AGEMA_signal_13152) ) ;
    buf_clk new_AGEMA_reg_buffer_7303 ( .C (clk), .D (new_AGEMA_signal_13154), .Q (new_AGEMA_signal_13155) ) ;
    buf_clk new_AGEMA_reg_buffer_7306 ( .C (clk), .D (new_AGEMA_signal_13157), .Q (new_AGEMA_signal_13158) ) ;
    buf_clk new_AGEMA_reg_buffer_7309 ( .C (clk), .D (new_AGEMA_signal_13160), .Q (new_AGEMA_signal_13161) ) ;
    buf_clk new_AGEMA_reg_buffer_7312 ( .C (clk), .D (new_AGEMA_signal_13163), .Q (new_AGEMA_signal_13164) ) ;
    buf_clk new_AGEMA_reg_buffer_7315 ( .C (clk), .D (new_AGEMA_signal_13166), .Q (new_AGEMA_signal_13167) ) ;
    buf_clk new_AGEMA_reg_buffer_7318 ( .C (clk), .D (new_AGEMA_signal_13169), .Q (new_AGEMA_signal_13170) ) ;
    buf_clk new_AGEMA_reg_buffer_7321 ( .C (clk), .D (new_AGEMA_signal_13172), .Q (new_AGEMA_signal_13173) ) ;
    buf_clk new_AGEMA_reg_buffer_7324 ( .C (clk), .D (new_AGEMA_signal_13175), .Q (new_AGEMA_signal_13176) ) ;
    buf_clk new_AGEMA_reg_buffer_7327 ( .C (clk), .D (new_AGEMA_signal_13178), .Q (new_AGEMA_signal_13179) ) ;
    buf_clk new_AGEMA_reg_buffer_7330 ( .C (clk), .D (new_AGEMA_signal_13181), .Q (new_AGEMA_signal_13182) ) ;
    buf_clk new_AGEMA_reg_buffer_7333 ( .C (clk), .D (new_AGEMA_signal_13184), .Q (new_AGEMA_signal_13185) ) ;
    buf_clk new_AGEMA_reg_buffer_7336 ( .C (clk), .D (new_AGEMA_signal_13187), .Q (new_AGEMA_signal_13188) ) ;
    buf_clk new_AGEMA_reg_buffer_7339 ( .C (clk), .D (new_AGEMA_signal_13190), .Q (new_AGEMA_signal_13191) ) ;
    buf_clk new_AGEMA_reg_buffer_7342 ( .C (clk), .D (new_AGEMA_signal_13193), .Q (new_AGEMA_signal_13194) ) ;
    buf_clk new_AGEMA_reg_buffer_7345 ( .C (clk), .D (new_AGEMA_signal_13196), .Q (new_AGEMA_signal_13197) ) ;
    buf_clk new_AGEMA_reg_buffer_7348 ( .C (clk), .D (new_AGEMA_signal_13199), .Q (new_AGEMA_signal_13200) ) ;
    buf_clk new_AGEMA_reg_buffer_7351 ( .C (clk), .D (new_AGEMA_signal_13202), .Q (new_AGEMA_signal_13203) ) ;
    buf_clk new_AGEMA_reg_buffer_7354 ( .C (clk), .D (new_AGEMA_signal_13205), .Q (new_AGEMA_signal_13206) ) ;
    buf_clk new_AGEMA_reg_buffer_7357 ( .C (clk), .D (new_AGEMA_signal_13208), .Q (new_AGEMA_signal_13209) ) ;
    buf_clk new_AGEMA_reg_buffer_7360 ( .C (clk), .D (new_AGEMA_signal_13211), .Q (new_AGEMA_signal_13212) ) ;
    buf_clk new_AGEMA_reg_buffer_7363 ( .C (clk), .D (new_AGEMA_signal_13214), .Q (new_AGEMA_signal_13215) ) ;
    buf_clk new_AGEMA_reg_buffer_7366 ( .C (clk), .D (new_AGEMA_signal_13217), .Q (new_AGEMA_signal_13218) ) ;
    buf_clk new_AGEMA_reg_buffer_7369 ( .C (clk), .D (new_AGEMA_signal_13220), .Q (new_AGEMA_signal_13221) ) ;
    buf_clk new_AGEMA_reg_buffer_7372 ( .C (clk), .D (new_AGEMA_signal_13223), .Q (new_AGEMA_signal_13224) ) ;
    buf_clk new_AGEMA_reg_buffer_7375 ( .C (clk), .D (new_AGEMA_signal_13226), .Q (new_AGEMA_signal_13227) ) ;
    buf_clk new_AGEMA_reg_buffer_7378 ( .C (clk), .D (new_AGEMA_signal_13229), .Q (new_AGEMA_signal_13230) ) ;
    buf_clk new_AGEMA_reg_buffer_7381 ( .C (clk), .D (new_AGEMA_signal_13232), .Q (new_AGEMA_signal_13233) ) ;
    buf_clk new_AGEMA_reg_buffer_7384 ( .C (clk), .D (new_AGEMA_signal_13235), .Q (new_AGEMA_signal_13236) ) ;
    buf_clk new_AGEMA_reg_buffer_7387 ( .C (clk), .D (new_AGEMA_signal_13238), .Q (new_AGEMA_signal_13239) ) ;
    buf_clk new_AGEMA_reg_buffer_7390 ( .C (clk), .D (new_AGEMA_signal_13241), .Q (new_AGEMA_signal_13242) ) ;
    buf_clk new_AGEMA_reg_buffer_7393 ( .C (clk), .D (new_AGEMA_signal_13244), .Q (new_AGEMA_signal_13245) ) ;
    buf_clk new_AGEMA_reg_buffer_7396 ( .C (clk), .D (new_AGEMA_signal_13247), .Q (new_AGEMA_signal_13248) ) ;
    buf_clk new_AGEMA_reg_buffer_7399 ( .C (clk), .D (new_AGEMA_signal_13250), .Q (new_AGEMA_signal_13251) ) ;
    buf_clk new_AGEMA_reg_buffer_7402 ( .C (clk), .D (new_AGEMA_signal_13253), .Q (new_AGEMA_signal_13254) ) ;
    buf_clk new_AGEMA_reg_buffer_7405 ( .C (clk), .D (new_AGEMA_signal_13256), .Q (new_AGEMA_signal_13257) ) ;
    buf_clk new_AGEMA_reg_buffer_7408 ( .C (clk), .D (new_AGEMA_signal_13259), .Q (new_AGEMA_signal_13260) ) ;
    buf_clk new_AGEMA_reg_buffer_7411 ( .C (clk), .D (new_AGEMA_signal_13262), .Q (new_AGEMA_signal_13263) ) ;
    buf_clk new_AGEMA_reg_buffer_7414 ( .C (clk), .D (new_AGEMA_signal_13265), .Q (new_AGEMA_signal_13266) ) ;
    buf_clk new_AGEMA_reg_buffer_7417 ( .C (clk), .D (new_AGEMA_signal_13268), .Q (new_AGEMA_signal_13269) ) ;
    buf_clk new_AGEMA_reg_buffer_7420 ( .C (clk), .D (new_AGEMA_signal_13271), .Q (new_AGEMA_signal_13272) ) ;
    buf_clk new_AGEMA_reg_buffer_7423 ( .C (clk), .D (new_AGEMA_signal_13274), .Q (new_AGEMA_signal_13275) ) ;
    buf_clk new_AGEMA_reg_buffer_7426 ( .C (clk), .D (new_AGEMA_signal_13277), .Q (new_AGEMA_signal_13278) ) ;
    buf_clk new_AGEMA_reg_buffer_7429 ( .C (clk), .D (new_AGEMA_signal_13280), .Q (new_AGEMA_signal_13281) ) ;
    buf_clk new_AGEMA_reg_buffer_7432 ( .C (clk), .D (new_AGEMA_signal_13283), .Q (new_AGEMA_signal_13284) ) ;
    buf_clk new_AGEMA_reg_buffer_7435 ( .C (clk), .D (new_AGEMA_signal_13286), .Q (new_AGEMA_signal_13287) ) ;
    buf_clk new_AGEMA_reg_buffer_7438 ( .C (clk), .D (new_AGEMA_signal_13289), .Q (new_AGEMA_signal_13290) ) ;
    buf_clk new_AGEMA_reg_buffer_7441 ( .C (clk), .D (new_AGEMA_signal_13292), .Q (new_AGEMA_signal_13293) ) ;
    buf_clk new_AGEMA_reg_buffer_7444 ( .C (clk), .D (new_AGEMA_signal_13295), .Q (new_AGEMA_signal_13296) ) ;
    buf_clk new_AGEMA_reg_buffer_7447 ( .C (clk), .D (new_AGEMA_signal_13298), .Q (new_AGEMA_signal_13299) ) ;
    buf_clk new_AGEMA_reg_buffer_7450 ( .C (clk), .D (new_AGEMA_signal_13301), .Q (new_AGEMA_signal_13302) ) ;
    buf_clk new_AGEMA_reg_buffer_7453 ( .C (clk), .D (new_AGEMA_signal_13304), .Q (new_AGEMA_signal_13305) ) ;
    buf_clk new_AGEMA_reg_buffer_7456 ( .C (clk), .D (new_AGEMA_signal_13307), .Q (new_AGEMA_signal_13308) ) ;
    buf_clk new_AGEMA_reg_buffer_7459 ( .C (clk), .D (new_AGEMA_signal_13310), .Q (new_AGEMA_signal_13311) ) ;
    buf_clk new_AGEMA_reg_buffer_7462 ( .C (clk), .D (new_AGEMA_signal_13313), .Q (new_AGEMA_signal_13314) ) ;
    buf_clk new_AGEMA_reg_buffer_7465 ( .C (clk), .D (new_AGEMA_signal_13316), .Q (new_AGEMA_signal_13317) ) ;
    buf_clk new_AGEMA_reg_buffer_7468 ( .C (clk), .D (new_AGEMA_signal_13319), .Q (new_AGEMA_signal_13320) ) ;
    buf_clk new_AGEMA_reg_buffer_7471 ( .C (clk), .D (new_AGEMA_signal_13322), .Q (new_AGEMA_signal_13323) ) ;
    buf_clk new_AGEMA_reg_buffer_7474 ( .C (clk), .D (new_AGEMA_signal_13325), .Q (new_AGEMA_signal_13326) ) ;
    buf_clk new_AGEMA_reg_buffer_7478 ( .C (clk), .D (new_AGEMA_signal_13329), .Q (new_AGEMA_signal_13330) ) ;
    buf_clk new_AGEMA_reg_buffer_7482 ( .C (clk), .D (new_AGEMA_signal_13333), .Q (new_AGEMA_signal_13334) ) ;
    buf_clk new_AGEMA_reg_buffer_7486 ( .C (clk), .D (new_AGEMA_signal_13337), .Q (new_AGEMA_signal_13338) ) ;
    buf_clk new_AGEMA_reg_buffer_7490 ( .C (clk), .D (new_AGEMA_signal_13341), .Q (new_AGEMA_signal_13342) ) ;
    buf_clk new_AGEMA_reg_buffer_7494 ( .C (clk), .D (new_AGEMA_signal_13345), .Q (new_AGEMA_signal_13346) ) ;
    buf_clk new_AGEMA_reg_buffer_7498 ( .C (clk), .D (new_AGEMA_signal_13349), .Q (new_AGEMA_signal_13350) ) ;
    buf_clk new_AGEMA_reg_buffer_7502 ( .C (clk), .D (new_AGEMA_signal_13353), .Q (new_AGEMA_signal_13354) ) ;
    buf_clk new_AGEMA_reg_buffer_7506 ( .C (clk), .D (new_AGEMA_signal_13357), .Q (new_AGEMA_signal_13358) ) ;
    buf_clk new_AGEMA_reg_buffer_7510 ( .C (clk), .D (new_AGEMA_signal_13361), .Q (new_AGEMA_signal_13362) ) ;
    buf_clk new_AGEMA_reg_buffer_7514 ( .C (clk), .D (new_AGEMA_signal_13365), .Q (new_AGEMA_signal_13366) ) ;
    buf_clk new_AGEMA_reg_buffer_7518 ( .C (clk), .D (new_AGEMA_signal_13369), .Q (new_AGEMA_signal_13370) ) ;
    buf_clk new_AGEMA_reg_buffer_7522 ( .C (clk), .D (new_AGEMA_signal_13373), .Q (new_AGEMA_signal_13374) ) ;
    buf_clk new_AGEMA_reg_buffer_7526 ( .C (clk), .D (new_AGEMA_signal_13377), .Q (new_AGEMA_signal_13378) ) ;
    buf_clk new_AGEMA_reg_buffer_7530 ( .C (clk), .D (new_AGEMA_signal_13381), .Q (new_AGEMA_signal_13382) ) ;
    buf_clk new_AGEMA_reg_buffer_7534 ( .C (clk), .D (new_AGEMA_signal_13385), .Q (new_AGEMA_signal_13386) ) ;
    buf_clk new_AGEMA_reg_buffer_7538 ( .C (clk), .D (new_AGEMA_signal_13389), .Q (new_AGEMA_signal_13390) ) ;
    buf_clk new_AGEMA_reg_buffer_7542 ( .C (clk), .D (new_AGEMA_signal_13393), .Q (new_AGEMA_signal_13394) ) ;
    buf_clk new_AGEMA_reg_buffer_7546 ( .C (clk), .D (new_AGEMA_signal_13397), .Q (new_AGEMA_signal_13398) ) ;
    buf_clk new_AGEMA_reg_buffer_7550 ( .C (clk), .D (new_AGEMA_signal_13401), .Q (new_AGEMA_signal_13402) ) ;
    buf_clk new_AGEMA_reg_buffer_7554 ( .C (clk), .D (new_AGEMA_signal_13405), .Q (new_AGEMA_signal_13406) ) ;
    buf_clk new_AGEMA_reg_buffer_7558 ( .C (clk), .D (new_AGEMA_signal_13409), .Q (new_AGEMA_signal_13410) ) ;
    buf_clk new_AGEMA_reg_buffer_7562 ( .C (clk), .D (new_AGEMA_signal_13413), .Q (new_AGEMA_signal_13414) ) ;
    buf_clk new_AGEMA_reg_buffer_7566 ( .C (clk), .D (new_AGEMA_signal_13417), .Q (new_AGEMA_signal_13418) ) ;
    buf_clk new_AGEMA_reg_buffer_7570 ( .C (clk), .D (new_AGEMA_signal_13421), .Q (new_AGEMA_signal_13422) ) ;
    buf_clk new_AGEMA_reg_buffer_7574 ( .C (clk), .D (new_AGEMA_signal_13425), .Q (new_AGEMA_signal_13426) ) ;
    buf_clk new_AGEMA_reg_buffer_7578 ( .C (clk), .D (new_AGEMA_signal_13429), .Q (new_AGEMA_signal_13430) ) ;
    buf_clk new_AGEMA_reg_buffer_7582 ( .C (clk), .D (new_AGEMA_signal_13433), .Q (new_AGEMA_signal_13434) ) ;
    buf_clk new_AGEMA_reg_buffer_7586 ( .C (clk), .D (new_AGEMA_signal_13437), .Q (new_AGEMA_signal_13438) ) ;
    buf_clk new_AGEMA_reg_buffer_7590 ( .C (clk), .D (new_AGEMA_signal_13441), .Q (new_AGEMA_signal_13442) ) ;
    buf_clk new_AGEMA_reg_buffer_7594 ( .C (clk), .D (new_AGEMA_signal_13445), .Q (new_AGEMA_signal_13446) ) ;
    buf_clk new_AGEMA_reg_buffer_7598 ( .C (clk), .D (new_AGEMA_signal_13449), .Q (new_AGEMA_signal_13450) ) ;
    buf_clk new_AGEMA_reg_buffer_7602 ( .C (clk), .D (new_AGEMA_signal_13453), .Q (new_AGEMA_signal_13454) ) ;
    buf_clk new_AGEMA_reg_buffer_7606 ( .C (clk), .D (new_AGEMA_signal_13457), .Q (new_AGEMA_signal_13458) ) ;
    buf_clk new_AGEMA_reg_buffer_7610 ( .C (clk), .D (new_AGEMA_signal_13461), .Q (new_AGEMA_signal_13462) ) ;
    buf_clk new_AGEMA_reg_buffer_7614 ( .C (clk), .D (new_AGEMA_signal_13465), .Q (new_AGEMA_signal_13466) ) ;
    buf_clk new_AGEMA_reg_buffer_7618 ( .C (clk), .D (new_AGEMA_signal_13469), .Q (new_AGEMA_signal_13470) ) ;
    buf_clk new_AGEMA_reg_buffer_7622 ( .C (clk), .D (new_AGEMA_signal_13473), .Q (new_AGEMA_signal_13474) ) ;
    buf_clk new_AGEMA_reg_buffer_7626 ( .C (clk), .D (new_AGEMA_signal_13477), .Q (new_AGEMA_signal_13478) ) ;
    buf_clk new_AGEMA_reg_buffer_7630 ( .C (clk), .D (new_AGEMA_signal_13481), .Q (new_AGEMA_signal_13482) ) ;
    buf_clk new_AGEMA_reg_buffer_7634 ( .C (clk), .D (new_AGEMA_signal_13485), .Q (new_AGEMA_signal_13486) ) ;
    buf_clk new_AGEMA_reg_buffer_7638 ( .C (clk), .D (new_AGEMA_signal_13489), .Q (new_AGEMA_signal_13490) ) ;
    buf_clk new_AGEMA_reg_buffer_7642 ( .C (clk), .D (new_AGEMA_signal_13493), .Q (new_AGEMA_signal_13494) ) ;
    buf_clk new_AGEMA_reg_buffer_7646 ( .C (clk), .D (new_AGEMA_signal_13497), .Q (new_AGEMA_signal_13498) ) ;
    buf_clk new_AGEMA_reg_buffer_7650 ( .C (clk), .D (new_AGEMA_signal_13501), .Q (new_AGEMA_signal_13502) ) ;
    buf_clk new_AGEMA_reg_buffer_7654 ( .C (clk), .D (new_AGEMA_signal_13505), .Q (new_AGEMA_signal_13506) ) ;
    buf_clk new_AGEMA_reg_buffer_7658 ( .C (clk), .D (new_AGEMA_signal_13509), .Q (new_AGEMA_signal_13510) ) ;
    buf_clk new_AGEMA_reg_buffer_7662 ( .C (clk), .D (new_AGEMA_signal_13513), .Q (new_AGEMA_signal_13514) ) ;
    buf_clk new_AGEMA_reg_buffer_7666 ( .C (clk), .D (new_AGEMA_signal_13517), .Q (new_AGEMA_signal_13518) ) ;
    buf_clk new_AGEMA_reg_buffer_7670 ( .C (clk), .D (new_AGEMA_signal_13521), .Q (new_AGEMA_signal_13522) ) ;
    buf_clk new_AGEMA_reg_buffer_7674 ( .C (clk), .D (new_AGEMA_signal_13525), .Q (new_AGEMA_signal_13526) ) ;
    buf_clk new_AGEMA_reg_buffer_7678 ( .C (clk), .D (new_AGEMA_signal_13529), .Q (new_AGEMA_signal_13530) ) ;
    buf_clk new_AGEMA_reg_buffer_7682 ( .C (clk), .D (new_AGEMA_signal_13533), .Q (new_AGEMA_signal_13534) ) ;
    buf_clk new_AGEMA_reg_buffer_7686 ( .C (clk), .D (new_AGEMA_signal_13537), .Q (new_AGEMA_signal_13538) ) ;
    buf_clk new_AGEMA_reg_buffer_7690 ( .C (clk), .D (new_AGEMA_signal_13541), .Q (new_AGEMA_signal_13542) ) ;
    buf_clk new_AGEMA_reg_buffer_7694 ( .C (clk), .D (new_AGEMA_signal_13545), .Q (new_AGEMA_signal_13546) ) ;
    buf_clk new_AGEMA_reg_buffer_7698 ( .C (clk), .D (new_AGEMA_signal_13549), .Q (new_AGEMA_signal_13550) ) ;
    buf_clk new_AGEMA_reg_buffer_7702 ( .C (clk), .D (new_AGEMA_signal_13553), .Q (new_AGEMA_signal_13554) ) ;
    buf_clk new_AGEMA_reg_buffer_7706 ( .C (clk), .D (new_AGEMA_signal_13557), .Q (new_AGEMA_signal_13558) ) ;
    buf_clk new_AGEMA_reg_buffer_7710 ( .C (clk), .D (new_AGEMA_signal_13561), .Q (new_AGEMA_signal_13562) ) ;
    buf_clk new_AGEMA_reg_buffer_7714 ( .C (clk), .D (new_AGEMA_signal_13565), .Q (new_AGEMA_signal_13566) ) ;
    buf_clk new_AGEMA_reg_buffer_7718 ( .C (clk), .D (new_AGEMA_signal_13569), .Q (new_AGEMA_signal_13570) ) ;
    buf_clk new_AGEMA_reg_buffer_7722 ( .C (clk), .D (new_AGEMA_signal_13573), .Q (new_AGEMA_signal_13574) ) ;
    buf_clk new_AGEMA_reg_buffer_7726 ( .C (clk), .D (new_AGEMA_signal_13577), .Q (new_AGEMA_signal_13578) ) ;
    buf_clk new_AGEMA_reg_buffer_7730 ( .C (clk), .D (new_AGEMA_signal_13581), .Q (new_AGEMA_signal_13582) ) ;
    buf_clk new_AGEMA_reg_buffer_7734 ( .C (clk), .D (new_AGEMA_signal_13585), .Q (new_AGEMA_signal_13586) ) ;
    buf_clk new_AGEMA_reg_buffer_7738 ( .C (clk), .D (new_AGEMA_signal_13589), .Q (new_AGEMA_signal_13590) ) ;
    buf_clk new_AGEMA_reg_buffer_7742 ( .C (clk), .D (new_AGEMA_signal_13593), .Q (new_AGEMA_signal_13594) ) ;
    buf_clk new_AGEMA_reg_buffer_7746 ( .C (clk), .D (new_AGEMA_signal_13597), .Q (new_AGEMA_signal_13598) ) ;
    buf_clk new_AGEMA_reg_buffer_7750 ( .C (clk), .D (new_AGEMA_signal_13601), .Q (new_AGEMA_signal_13602) ) ;
    buf_clk new_AGEMA_reg_buffer_7754 ( .C (clk), .D (new_AGEMA_signal_13605), .Q (new_AGEMA_signal_13606) ) ;
    buf_clk new_AGEMA_reg_buffer_7758 ( .C (clk), .D (new_AGEMA_signal_13609), .Q (new_AGEMA_signal_13610) ) ;
    buf_clk new_AGEMA_reg_buffer_7762 ( .C (clk), .D (new_AGEMA_signal_13613), .Q (new_AGEMA_signal_13614) ) ;
    buf_clk new_AGEMA_reg_buffer_7766 ( .C (clk), .D (new_AGEMA_signal_13617), .Q (new_AGEMA_signal_13618) ) ;
    buf_clk new_AGEMA_reg_buffer_7770 ( .C (clk), .D (new_AGEMA_signal_13621), .Q (new_AGEMA_signal_13622) ) ;
    buf_clk new_AGEMA_reg_buffer_7774 ( .C (clk), .D (new_AGEMA_signal_13625), .Q (new_AGEMA_signal_13626) ) ;
    buf_clk new_AGEMA_reg_buffer_7778 ( .C (clk), .D (new_AGEMA_signal_13629), .Q (new_AGEMA_signal_13630) ) ;
    buf_clk new_AGEMA_reg_buffer_7782 ( .C (clk), .D (new_AGEMA_signal_13633), .Q (new_AGEMA_signal_13634) ) ;
    buf_clk new_AGEMA_reg_buffer_7786 ( .C (clk), .D (new_AGEMA_signal_13637), .Q (new_AGEMA_signal_13638) ) ;
    buf_clk new_AGEMA_reg_buffer_7790 ( .C (clk), .D (new_AGEMA_signal_13641), .Q (new_AGEMA_signal_13642) ) ;
    buf_clk new_AGEMA_reg_buffer_7794 ( .C (clk), .D (new_AGEMA_signal_13645), .Q (new_AGEMA_signal_13646) ) ;
    buf_clk new_AGEMA_reg_buffer_7798 ( .C (clk), .D (new_AGEMA_signal_13649), .Q (new_AGEMA_signal_13650) ) ;
    buf_clk new_AGEMA_reg_buffer_7802 ( .C (clk), .D (new_AGEMA_signal_13653), .Q (new_AGEMA_signal_13654) ) ;
    buf_clk new_AGEMA_reg_buffer_7806 ( .C (clk), .D (new_AGEMA_signal_13657), .Q (new_AGEMA_signal_13658) ) ;
    buf_clk new_AGEMA_reg_buffer_7810 ( .C (clk), .D (new_AGEMA_signal_13661), .Q (new_AGEMA_signal_13662) ) ;
    buf_clk new_AGEMA_reg_buffer_7814 ( .C (clk), .D (new_AGEMA_signal_13665), .Q (new_AGEMA_signal_13666) ) ;
    buf_clk new_AGEMA_reg_buffer_7818 ( .C (clk), .D (new_AGEMA_signal_13669), .Q (new_AGEMA_signal_13670) ) ;
    buf_clk new_AGEMA_reg_buffer_7822 ( .C (clk), .D (new_AGEMA_signal_13673), .Q (new_AGEMA_signal_13674) ) ;
    buf_clk new_AGEMA_reg_buffer_7826 ( .C (clk), .D (new_AGEMA_signal_13677), .Q (new_AGEMA_signal_13678) ) ;
    buf_clk new_AGEMA_reg_buffer_7830 ( .C (clk), .D (new_AGEMA_signal_13681), .Q (new_AGEMA_signal_13682) ) ;
    buf_clk new_AGEMA_reg_buffer_7834 ( .C (clk), .D (new_AGEMA_signal_13685), .Q (new_AGEMA_signal_13686) ) ;
    buf_clk new_AGEMA_reg_buffer_7838 ( .C (clk), .D (new_AGEMA_signal_13689), .Q (new_AGEMA_signal_13690) ) ;
    buf_clk new_AGEMA_reg_buffer_7842 ( .C (clk), .D (new_AGEMA_signal_13693), .Q (new_AGEMA_signal_13694) ) ;
    buf_clk new_AGEMA_reg_buffer_7846 ( .C (clk), .D (new_AGEMA_signal_13697), .Q (new_AGEMA_signal_13698) ) ;
    buf_clk new_AGEMA_reg_buffer_7850 ( .C (clk), .D (new_AGEMA_signal_13701), .Q (new_AGEMA_signal_13702) ) ;
    buf_clk new_AGEMA_reg_buffer_7854 ( .C (clk), .D (new_AGEMA_signal_13705), .Q (new_AGEMA_signal_13706) ) ;
    buf_clk new_AGEMA_reg_buffer_7858 ( .C (clk), .D (new_AGEMA_signal_13709), .Q (new_AGEMA_signal_13710) ) ;
    buf_clk new_AGEMA_reg_buffer_7862 ( .C (clk), .D (new_AGEMA_signal_13713), .Q (new_AGEMA_signal_13714) ) ;
    buf_clk new_AGEMA_reg_buffer_7866 ( .C (clk), .D (new_AGEMA_signal_13717), .Q (new_AGEMA_signal_13718) ) ;
    buf_clk new_AGEMA_reg_buffer_7870 ( .C (clk), .D (new_AGEMA_signal_13721), .Q (new_AGEMA_signal_13722) ) ;
    buf_clk new_AGEMA_reg_buffer_7874 ( .C (clk), .D (new_AGEMA_signal_13725), .Q (new_AGEMA_signal_13726) ) ;
    buf_clk new_AGEMA_reg_buffer_7878 ( .C (clk), .D (new_AGEMA_signal_13729), .Q (new_AGEMA_signal_13730) ) ;
    buf_clk new_AGEMA_reg_buffer_7882 ( .C (clk), .D (new_AGEMA_signal_13733), .Q (new_AGEMA_signal_13734) ) ;
    buf_clk new_AGEMA_reg_buffer_7886 ( .C (clk), .D (new_AGEMA_signal_13737), .Q (new_AGEMA_signal_13738) ) ;
    buf_clk new_AGEMA_reg_buffer_7890 ( .C (clk), .D (new_AGEMA_signal_13741), .Q (new_AGEMA_signal_13742) ) ;
    buf_clk new_AGEMA_reg_buffer_7894 ( .C (clk), .D (new_AGEMA_signal_13745), .Q (new_AGEMA_signal_13746) ) ;
    buf_clk new_AGEMA_reg_buffer_7898 ( .C (clk), .D (new_AGEMA_signal_13749), .Q (new_AGEMA_signal_13750) ) ;
    buf_clk new_AGEMA_reg_buffer_7902 ( .C (clk), .D (new_AGEMA_signal_13753), .Q (new_AGEMA_signal_13754) ) ;
    buf_clk new_AGEMA_reg_buffer_7906 ( .C (clk), .D (new_AGEMA_signal_13757), .Q (new_AGEMA_signal_13758) ) ;
    buf_clk new_AGEMA_reg_buffer_7910 ( .C (clk), .D (new_AGEMA_signal_13761), .Q (new_AGEMA_signal_13762) ) ;
    buf_clk new_AGEMA_reg_buffer_7914 ( .C (clk), .D (new_AGEMA_signal_13765), .Q (new_AGEMA_signal_13766) ) ;
    buf_clk new_AGEMA_reg_buffer_7918 ( .C (clk), .D (new_AGEMA_signal_13769), .Q (new_AGEMA_signal_13770) ) ;
    buf_clk new_AGEMA_reg_buffer_7922 ( .C (clk), .D (new_AGEMA_signal_13773), .Q (new_AGEMA_signal_13774) ) ;
    buf_clk new_AGEMA_reg_buffer_7926 ( .C (clk), .D (new_AGEMA_signal_13777), .Q (new_AGEMA_signal_13778) ) ;
    buf_clk new_AGEMA_reg_buffer_7930 ( .C (clk), .D (new_AGEMA_signal_13781), .Q (new_AGEMA_signal_13782) ) ;
    buf_clk new_AGEMA_reg_buffer_7934 ( .C (clk), .D (new_AGEMA_signal_13785), .Q (new_AGEMA_signal_13786) ) ;
    buf_clk new_AGEMA_reg_buffer_7938 ( .C (clk), .D (new_AGEMA_signal_13789), .Q (new_AGEMA_signal_13790) ) ;
    buf_clk new_AGEMA_reg_buffer_7942 ( .C (clk), .D (new_AGEMA_signal_13793), .Q (new_AGEMA_signal_13794) ) ;
    buf_clk new_AGEMA_reg_buffer_7946 ( .C (clk), .D (new_AGEMA_signal_13797), .Q (new_AGEMA_signal_13798) ) ;
    buf_clk new_AGEMA_reg_buffer_7950 ( .C (clk), .D (new_AGEMA_signal_13801), .Q (new_AGEMA_signal_13802) ) ;
    buf_clk new_AGEMA_reg_buffer_7954 ( .C (clk), .D (new_AGEMA_signal_13805), .Q (new_AGEMA_signal_13806) ) ;
    buf_clk new_AGEMA_reg_buffer_7958 ( .C (clk), .D (new_AGEMA_signal_13809), .Q (new_AGEMA_signal_13810) ) ;
    buf_clk new_AGEMA_reg_buffer_7962 ( .C (clk), .D (new_AGEMA_signal_13813), .Q (new_AGEMA_signal_13814) ) ;
    buf_clk new_AGEMA_reg_buffer_7966 ( .C (clk), .D (new_AGEMA_signal_13817), .Q (new_AGEMA_signal_13818) ) ;
    buf_clk new_AGEMA_reg_buffer_7970 ( .C (clk), .D (new_AGEMA_signal_13821), .Q (new_AGEMA_signal_13822) ) ;
    buf_clk new_AGEMA_reg_buffer_7974 ( .C (clk), .D (new_AGEMA_signal_13825), .Q (new_AGEMA_signal_13826) ) ;
    buf_clk new_AGEMA_reg_buffer_7978 ( .C (clk), .D (new_AGEMA_signal_13829), .Q (new_AGEMA_signal_13830) ) ;
    buf_clk new_AGEMA_reg_buffer_7982 ( .C (clk), .D (new_AGEMA_signal_13833), .Q (new_AGEMA_signal_13834) ) ;
    buf_clk new_AGEMA_reg_buffer_7986 ( .C (clk), .D (new_AGEMA_signal_13837), .Q (new_AGEMA_signal_13838) ) ;
    buf_clk new_AGEMA_reg_buffer_7990 ( .C (clk), .D (new_AGEMA_signal_13841), .Q (new_AGEMA_signal_13842) ) ;
    buf_clk new_AGEMA_reg_buffer_7994 ( .C (clk), .D (new_AGEMA_signal_13845), .Q (new_AGEMA_signal_13846) ) ;
    buf_clk new_AGEMA_reg_buffer_7998 ( .C (clk), .D (new_AGEMA_signal_13849), .Q (new_AGEMA_signal_13850) ) ;
    buf_clk new_AGEMA_reg_buffer_8002 ( .C (clk), .D (new_AGEMA_signal_13853), .Q (new_AGEMA_signal_13854) ) ;
    buf_clk new_AGEMA_reg_buffer_8006 ( .C (clk), .D (new_AGEMA_signal_13857), .Q (new_AGEMA_signal_13858) ) ;
    buf_clk new_AGEMA_reg_buffer_8010 ( .C (clk), .D (new_AGEMA_signal_13861), .Q (new_AGEMA_signal_13862) ) ;
    buf_clk new_AGEMA_reg_buffer_8014 ( .C (clk), .D (new_AGEMA_signal_13865), .Q (new_AGEMA_signal_13866) ) ;
    buf_clk new_AGEMA_reg_buffer_8018 ( .C (clk), .D (new_AGEMA_signal_13869), .Q (new_AGEMA_signal_13870) ) ;
    buf_clk new_AGEMA_reg_buffer_8022 ( .C (clk), .D (new_AGEMA_signal_13873), .Q (new_AGEMA_signal_13874) ) ;
    buf_clk new_AGEMA_reg_buffer_8026 ( .C (clk), .D (new_AGEMA_signal_13877), .Q (new_AGEMA_signal_13878) ) ;
    buf_clk new_AGEMA_reg_buffer_8030 ( .C (clk), .D (new_AGEMA_signal_13881), .Q (new_AGEMA_signal_13882) ) ;
    buf_clk new_AGEMA_reg_buffer_8034 ( .C (clk), .D (new_AGEMA_signal_13885), .Q (new_AGEMA_signal_13886) ) ;
    buf_clk new_AGEMA_reg_buffer_8038 ( .C (clk), .D (new_AGEMA_signal_13889), .Q (new_AGEMA_signal_13890) ) ;
    buf_clk new_AGEMA_reg_buffer_8042 ( .C (clk), .D (new_AGEMA_signal_13893), .Q (new_AGEMA_signal_13894) ) ;
    buf_clk new_AGEMA_reg_buffer_8046 ( .C (clk), .D (new_AGEMA_signal_13897), .Q (new_AGEMA_signal_13898) ) ;
    buf_clk new_AGEMA_reg_buffer_8050 ( .C (clk), .D (new_AGEMA_signal_13901), .Q (new_AGEMA_signal_13902) ) ;
    buf_clk new_AGEMA_reg_buffer_8054 ( .C (clk), .D (new_AGEMA_signal_13905), .Q (new_AGEMA_signal_13906) ) ;
    buf_clk new_AGEMA_reg_buffer_8058 ( .C (clk), .D (new_AGEMA_signal_13909), .Q (new_AGEMA_signal_13910) ) ;
    buf_clk new_AGEMA_reg_buffer_8062 ( .C (clk), .D (new_AGEMA_signal_13913), .Q (new_AGEMA_signal_13914) ) ;
    buf_clk new_AGEMA_reg_buffer_8066 ( .C (clk), .D (new_AGEMA_signal_13917), .Q (new_AGEMA_signal_13918) ) ;
    buf_clk new_AGEMA_reg_buffer_8070 ( .C (clk), .D (new_AGEMA_signal_13921), .Q (new_AGEMA_signal_13922) ) ;
    buf_clk new_AGEMA_reg_buffer_8074 ( .C (clk), .D (new_AGEMA_signal_13925), .Q (new_AGEMA_signal_13926) ) ;
    buf_clk new_AGEMA_reg_buffer_8078 ( .C (clk), .D (new_AGEMA_signal_13929), .Q (new_AGEMA_signal_13930) ) ;
    buf_clk new_AGEMA_reg_buffer_8082 ( .C (clk), .D (new_AGEMA_signal_13933), .Q (new_AGEMA_signal_13934) ) ;
    buf_clk new_AGEMA_reg_buffer_8086 ( .C (clk), .D (new_AGEMA_signal_13937), .Q (new_AGEMA_signal_13938) ) ;
    buf_clk new_AGEMA_reg_buffer_8090 ( .C (clk), .D (new_AGEMA_signal_13941), .Q (new_AGEMA_signal_13942) ) ;
    buf_clk new_AGEMA_reg_buffer_8094 ( .C (clk), .D (new_AGEMA_signal_13945), .Q (new_AGEMA_signal_13946) ) ;
    buf_clk new_AGEMA_reg_buffer_8098 ( .C (clk), .D (new_AGEMA_signal_13949), .Q (new_AGEMA_signal_13950) ) ;
    buf_clk new_AGEMA_reg_buffer_8102 ( .C (clk), .D (new_AGEMA_signal_13953), .Q (new_AGEMA_signal_13954) ) ;
    buf_clk new_AGEMA_reg_buffer_8106 ( .C (clk), .D (new_AGEMA_signal_13957), .Q (new_AGEMA_signal_13958) ) ;
    buf_clk new_AGEMA_reg_buffer_8110 ( .C (clk), .D (new_AGEMA_signal_13961), .Q (new_AGEMA_signal_13962) ) ;
    buf_clk new_AGEMA_reg_buffer_8114 ( .C (clk), .D (new_AGEMA_signal_13965), .Q (new_AGEMA_signal_13966) ) ;
    buf_clk new_AGEMA_reg_buffer_8118 ( .C (clk), .D (new_AGEMA_signal_13969), .Q (new_AGEMA_signal_13970) ) ;
    buf_clk new_AGEMA_reg_buffer_8122 ( .C (clk), .D (new_AGEMA_signal_13973), .Q (new_AGEMA_signal_13974) ) ;
    buf_clk new_AGEMA_reg_buffer_8126 ( .C (clk), .D (new_AGEMA_signal_13977), .Q (new_AGEMA_signal_13978) ) ;
    buf_clk new_AGEMA_reg_buffer_8130 ( .C (clk), .D (new_AGEMA_signal_13981), .Q (new_AGEMA_signal_13982) ) ;
    buf_clk new_AGEMA_reg_buffer_8134 ( .C (clk), .D (new_AGEMA_signal_13985), .Q (new_AGEMA_signal_13986) ) ;
    buf_clk new_AGEMA_reg_buffer_8138 ( .C (clk), .D (new_AGEMA_signal_13989), .Q (new_AGEMA_signal_13990) ) ;
    buf_clk new_AGEMA_reg_buffer_8142 ( .C (clk), .D (new_AGEMA_signal_13993), .Q (new_AGEMA_signal_13994) ) ;
    buf_clk new_AGEMA_reg_buffer_8146 ( .C (clk), .D (new_AGEMA_signal_13997), .Q (new_AGEMA_signal_13998) ) ;
    buf_clk new_AGEMA_reg_buffer_8150 ( .C (clk), .D (new_AGEMA_signal_14001), .Q (new_AGEMA_signal_14002) ) ;
    buf_clk new_AGEMA_reg_buffer_8154 ( .C (clk), .D (new_AGEMA_signal_14005), .Q (new_AGEMA_signal_14006) ) ;
    buf_clk new_AGEMA_reg_buffer_8158 ( .C (clk), .D (new_AGEMA_signal_14009), .Q (new_AGEMA_signal_14010) ) ;
    buf_clk new_AGEMA_reg_buffer_8162 ( .C (clk), .D (new_AGEMA_signal_14013), .Q (new_AGEMA_signal_14014) ) ;
    buf_clk new_AGEMA_reg_buffer_8166 ( .C (clk), .D (new_AGEMA_signal_14017), .Q (new_AGEMA_signal_14018) ) ;
    buf_clk new_AGEMA_reg_buffer_8170 ( .C (clk), .D (new_AGEMA_signal_14021), .Q (new_AGEMA_signal_14022) ) ;
    buf_clk new_AGEMA_reg_buffer_8174 ( .C (clk), .D (new_AGEMA_signal_14025), .Q (new_AGEMA_signal_14026) ) ;
    buf_clk new_AGEMA_reg_buffer_8178 ( .C (clk), .D (new_AGEMA_signal_14029), .Q (new_AGEMA_signal_14030) ) ;
    buf_clk new_AGEMA_reg_buffer_8182 ( .C (clk), .D (new_AGEMA_signal_14033), .Q (new_AGEMA_signal_14034) ) ;
    buf_clk new_AGEMA_reg_buffer_8186 ( .C (clk), .D (new_AGEMA_signal_14037), .Q (new_AGEMA_signal_14038) ) ;
    buf_clk new_AGEMA_reg_buffer_8190 ( .C (clk), .D (new_AGEMA_signal_14041), .Q (new_AGEMA_signal_14042) ) ;
    buf_clk new_AGEMA_reg_buffer_8194 ( .C (clk), .D (new_AGEMA_signal_14045), .Q (new_AGEMA_signal_14046) ) ;
    buf_clk new_AGEMA_reg_buffer_8198 ( .C (clk), .D (new_AGEMA_signal_14049), .Q (new_AGEMA_signal_14050) ) ;
    buf_clk new_AGEMA_reg_buffer_8202 ( .C (clk), .D (new_AGEMA_signal_14053), .Q (new_AGEMA_signal_14054) ) ;
    buf_clk new_AGEMA_reg_buffer_8206 ( .C (clk), .D (new_AGEMA_signal_14057), .Q (new_AGEMA_signal_14058) ) ;
    buf_clk new_AGEMA_reg_buffer_8210 ( .C (clk), .D (new_AGEMA_signal_14061), .Q (new_AGEMA_signal_14062) ) ;
    buf_clk new_AGEMA_reg_buffer_8214 ( .C (clk), .D (new_AGEMA_signal_14065), .Q (new_AGEMA_signal_14066) ) ;
    buf_clk new_AGEMA_reg_buffer_8218 ( .C (clk), .D (new_AGEMA_signal_14069), .Q (new_AGEMA_signal_14070) ) ;
    buf_clk new_AGEMA_reg_buffer_8222 ( .C (clk), .D (new_AGEMA_signal_14073), .Q (new_AGEMA_signal_14074) ) ;
    buf_clk new_AGEMA_reg_buffer_8226 ( .C (clk), .D (new_AGEMA_signal_14077), .Q (new_AGEMA_signal_14078) ) ;
    buf_clk new_AGEMA_reg_buffer_8230 ( .C (clk), .D (new_AGEMA_signal_14081), .Q (new_AGEMA_signal_14082) ) ;
    buf_clk new_AGEMA_reg_buffer_8234 ( .C (clk), .D (new_AGEMA_signal_14085), .Q (new_AGEMA_signal_14086) ) ;
    buf_clk new_AGEMA_reg_buffer_8238 ( .C (clk), .D (new_AGEMA_signal_14089), .Q (new_AGEMA_signal_14090) ) ;
    buf_clk new_AGEMA_reg_buffer_8242 ( .C (clk), .D (new_AGEMA_signal_14093), .Q (new_AGEMA_signal_14094) ) ;
    buf_clk new_AGEMA_reg_buffer_8246 ( .C (clk), .D (new_AGEMA_signal_14097), .Q (new_AGEMA_signal_14098) ) ;
    buf_clk new_AGEMA_reg_buffer_8250 ( .C (clk), .D (new_AGEMA_signal_14101), .Q (new_AGEMA_signal_14102) ) ;
    buf_clk new_AGEMA_reg_buffer_8254 ( .C (clk), .D (new_AGEMA_signal_14105), .Q (new_AGEMA_signal_14106) ) ;
    buf_clk new_AGEMA_reg_buffer_8258 ( .C (clk), .D (new_AGEMA_signal_14109), .Q (new_AGEMA_signal_14110) ) ;
    buf_clk new_AGEMA_reg_buffer_8262 ( .C (clk), .D (new_AGEMA_signal_14113), .Q (new_AGEMA_signal_14114) ) ;
    buf_clk new_AGEMA_reg_buffer_8266 ( .C (clk), .D (new_AGEMA_signal_14117), .Q (new_AGEMA_signal_14118) ) ;
    buf_clk new_AGEMA_reg_buffer_8270 ( .C (clk), .D (new_AGEMA_signal_14121), .Q (new_AGEMA_signal_14122) ) ;
    buf_clk new_AGEMA_reg_buffer_8274 ( .C (clk), .D (new_AGEMA_signal_14125), .Q (new_AGEMA_signal_14126) ) ;
    buf_clk new_AGEMA_reg_buffer_8278 ( .C (clk), .D (new_AGEMA_signal_14129), .Q (new_AGEMA_signal_14130) ) ;
    buf_clk new_AGEMA_reg_buffer_8282 ( .C (clk), .D (new_AGEMA_signal_14133), .Q (new_AGEMA_signal_14134) ) ;
    buf_clk new_AGEMA_reg_buffer_8286 ( .C (clk), .D (new_AGEMA_signal_14137), .Q (new_AGEMA_signal_14138) ) ;
    buf_clk new_AGEMA_reg_buffer_8290 ( .C (clk), .D (new_AGEMA_signal_14141), .Q (new_AGEMA_signal_14142) ) ;
    buf_clk new_AGEMA_reg_buffer_8294 ( .C (clk), .D (new_AGEMA_signal_14145), .Q (new_AGEMA_signal_14146) ) ;
    buf_clk new_AGEMA_reg_buffer_8298 ( .C (clk), .D (new_AGEMA_signal_14149), .Q (new_AGEMA_signal_14150) ) ;
    buf_clk new_AGEMA_reg_buffer_8302 ( .C (clk), .D (new_AGEMA_signal_14153), .Q (new_AGEMA_signal_14154) ) ;
    buf_clk new_AGEMA_reg_buffer_8306 ( .C (clk), .D (new_AGEMA_signal_14157), .Q (new_AGEMA_signal_14158) ) ;
    buf_clk new_AGEMA_reg_buffer_8310 ( .C (clk), .D (new_AGEMA_signal_14161), .Q (new_AGEMA_signal_14162) ) ;
    buf_clk new_AGEMA_reg_buffer_8314 ( .C (clk), .D (new_AGEMA_signal_14165), .Q (new_AGEMA_signal_14166) ) ;
    buf_clk new_AGEMA_reg_buffer_8318 ( .C (clk), .D (new_AGEMA_signal_14169), .Q (new_AGEMA_signal_14170) ) ;
    buf_clk new_AGEMA_reg_buffer_8322 ( .C (clk), .D (new_AGEMA_signal_14173), .Q (new_AGEMA_signal_14174) ) ;
    buf_clk new_AGEMA_reg_buffer_8326 ( .C (clk), .D (new_AGEMA_signal_14177), .Q (new_AGEMA_signal_14178) ) ;
    buf_clk new_AGEMA_reg_buffer_8330 ( .C (clk), .D (new_AGEMA_signal_14181), .Q (new_AGEMA_signal_14182) ) ;
    buf_clk new_AGEMA_reg_buffer_8334 ( .C (clk), .D (new_AGEMA_signal_14185), .Q (new_AGEMA_signal_14186) ) ;
    buf_clk new_AGEMA_reg_buffer_8338 ( .C (clk), .D (new_AGEMA_signal_14189), .Q (new_AGEMA_signal_14190) ) ;
    buf_clk new_AGEMA_reg_buffer_8342 ( .C (clk), .D (new_AGEMA_signal_14193), .Q (new_AGEMA_signal_14194) ) ;
    buf_clk new_AGEMA_reg_buffer_8346 ( .C (clk), .D (new_AGEMA_signal_14197), .Q (new_AGEMA_signal_14198) ) ;
    buf_clk new_AGEMA_reg_buffer_8350 ( .C (clk), .D (new_AGEMA_signal_14201), .Q (new_AGEMA_signal_14202) ) ;
    buf_clk new_AGEMA_reg_buffer_8354 ( .C (clk), .D (new_AGEMA_signal_14205), .Q (new_AGEMA_signal_14206) ) ;
    buf_clk new_AGEMA_reg_buffer_8358 ( .C (clk), .D (new_AGEMA_signal_14209), .Q (new_AGEMA_signal_14210) ) ;
    buf_clk new_AGEMA_reg_buffer_8362 ( .C (clk), .D (new_AGEMA_signal_14213), .Q (new_AGEMA_signal_14214) ) ;
    buf_clk new_AGEMA_reg_buffer_8366 ( .C (clk), .D (new_AGEMA_signal_14217), .Q (new_AGEMA_signal_14218) ) ;
    buf_clk new_AGEMA_reg_buffer_8370 ( .C (clk), .D (new_AGEMA_signal_14221), .Q (new_AGEMA_signal_14222) ) ;
    buf_clk new_AGEMA_reg_buffer_8374 ( .C (clk), .D (new_AGEMA_signal_14225), .Q (new_AGEMA_signal_14226) ) ;
    buf_clk new_AGEMA_reg_buffer_8378 ( .C (clk), .D (new_AGEMA_signal_14229), .Q (new_AGEMA_signal_14230) ) ;
    buf_clk new_AGEMA_reg_buffer_8382 ( .C (clk), .D (new_AGEMA_signal_14233), .Q (new_AGEMA_signal_14234) ) ;
    buf_clk new_AGEMA_reg_buffer_8386 ( .C (clk), .D (new_AGEMA_signal_14237), .Q (new_AGEMA_signal_14238) ) ;
    buf_clk new_AGEMA_reg_buffer_8390 ( .C (clk), .D (new_AGEMA_signal_14241), .Q (new_AGEMA_signal_14242) ) ;
    buf_clk new_AGEMA_reg_buffer_8394 ( .C (clk), .D (new_AGEMA_signal_14245), .Q (new_AGEMA_signal_14246) ) ;
    buf_clk new_AGEMA_reg_buffer_8398 ( .C (clk), .D (new_AGEMA_signal_14249), .Q (new_AGEMA_signal_14250) ) ;
    buf_clk new_AGEMA_reg_buffer_8402 ( .C (clk), .D (new_AGEMA_signal_14253), .Q (new_AGEMA_signal_14254) ) ;
    buf_clk new_AGEMA_reg_buffer_8406 ( .C (clk), .D (new_AGEMA_signal_14257), .Q (new_AGEMA_signal_14258) ) ;
    buf_clk new_AGEMA_reg_buffer_8410 ( .C (clk), .D (new_AGEMA_signal_14261), .Q (new_AGEMA_signal_14262) ) ;
    buf_clk new_AGEMA_reg_buffer_8414 ( .C (clk), .D (new_AGEMA_signal_14265), .Q (new_AGEMA_signal_14266) ) ;
    buf_clk new_AGEMA_reg_buffer_8418 ( .C (clk), .D (new_AGEMA_signal_14269), .Q (new_AGEMA_signal_14270) ) ;
    buf_clk new_AGEMA_reg_buffer_8422 ( .C (clk), .D (new_AGEMA_signal_14273), .Q (new_AGEMA_signal_14274) ) ;
    buf_clk new_AGEMA_reg_buffer_8426 ( .C (clk), .D (new_AGEMA_signal_14277), .Q (new_AGEMA_signal_14278) ) ;
    buf_clk new_AGEMA_reg_buffer_8430 ( .C (clk), .D (new_AGEMA_signal_14281), .Q (new_AGEMA_signal_14282) ) ;
    buf_clk new_AGEMA_reg_buffer_8434 ( .C (clk), .D (new_AGEMA_signal_14285), .Q (new_AGEMA_signal_14286) ) ;
    buf_clk new_AGEMA_reg_buffer_8438 ( .C (clk), .D (new_AGEMA_signal_14289), .Q (new_AGEMA_signal_14290) ) ;
    buf_clk new_AGEMA_reg_buffer_8442 ( .C (clk), .D (new_AGEMA_signal_14293), .Q (new_AGEMA_signal_14294) ) ;
    buf_clk new_AGEMA_reg_buffer_8446 ( .C (clk), .D (new_AGEMA_signal_14297), .Q (new_AGEMA_signal_14298) ) ;
    buf_clk new_AGEMA_reg_buffer_8450 ( .C (clk), .D (new_AGEMA_signal_14301), .Q (new_AGEMA_signal_14302) ) ;
    buf_clk new_AGEMA_reg_buffer_8454 ( .C (clk), .D (new_AGEMA_signal_14305), .Q (new_AGEMA_signal_14306) ) ;
    buf_clk new_AGEMA_reg_buffer_8458 ( .C (clk), .D (new_AGEMA_signal_14309), .Q (new_AGEMA_signal_14310) ) ;
    buf_clk new_AGEMA_reg_buffer_8462 ( .C (clk), .D (new_AGEMA_signal_14313), .Q (new_AGEMA_signal_14314) ) ;
    buf_clk new_AGEMA_reg_buffer_8466 ( .C (clk), .D (new_AGEMA_signal_14317), .Q (new_AGEMA_signal_14318) ) ;
    buf_clk new_AGEMA_reg_buffer_8470 ( .C (clk), .D (new_AGEMA_signal_14321), .Q (new_AGEMA_signal_14322) ) ;
    buf_clk new_AGEMA_reg_buffer_8474 ( .C (clk), .D (new_AGEMA_signal_14325), .Q (new_AGEMA_signal_14326) ) ;
    buf_clk new_AGEMA_reg_buffer_8478 ( .C (clk), .D (new_AGEMA_signal_14329), .Q (new_AGEMA_signal_14330) ) ;
    buf_clk new_AGEMA_reg_buffer_8482 ( .C (clk), .D (new_AGEMA_signal_14333), .Q (new_AGEMA_signal_14334) ) ;
    buf_clk new_AGEMA_reg_buffer_8486 ( .C (clk), .D (new_AGEMA_signal_14337), .Q (new_AGEMA_signal_14338) ) ;
    buf_clk new_AGEMA_reg_buffer_8490 ( .C (clk), .D (new_AGEMA_signal_14341), .Q (new_AGEMA_signal_14342) ) ;
    buf_clk new_AGEMA_reg_buffer_8494 ( .C (clk), .D (new_AGEMA_signal_14345), .Q (new_AGEMA_signal_14346) ) ;
    buf_clk new_AGEMA_reg_buffer_8498 ( .C (clk), .D (new_AGEMA_signal_14349), .Q (new_AGEMA_signal_14350) ) ;
    buf_clk new_AGEMA_reg_buffer_8502 ( .C (clk), .D (new_AGEMA_signal_14353), .Q (new_AGEMA_signal_14354) ) ;
    buf_clk new_AGEMA_reg_buffer_8506 ( .C (clk), .D (new_AGEMA_signal_14357), .Q (new_AGEMA_signal_14358) ) ;
    buf_clk new_AGEMA_reg_buffer_8510 ( .C (clk), .D (new_AGEMA_signal_14361), .Q (new_AGEMA_signal_14362) ) ;
    buf_clk new_AGEMA_reg_buffer_8514 ( .C (clk), .D (new_AGEMA_signal_14365), .Q (new_AGEMA_signal_14366) ) ;
    buf_clk new_AGEMA_reg_buffer_8518 ( .C (clk), .D (new_AGEMA_signal_14369), .Q (new_AGEMA_signal_14370) ) ;
    buf_clk new_AGEMA_reg_buffer_8522 ( .C (clk), .D (new_AGEMA_signal_14373), .Q (new_AGEMA_signal_14374) ) ;
    buf_clk new_AGEMA_reg_buffer_8526 ( .C (clk), .D (new_AGEMA_signal_14377), .Q (new_AGEMA_signal_14378) ) ;
    buf_clk new_AGEMA_reg_buffer_8530 ( .C (clk), .D (new_AGEMA_signal_14381), .Q (new_AGEMA_signal_14382) ) ;
    buf_clk new_AGEMA_reg_buffer_8534 ( .C (clk), .D (new_AGEMA_signal_14385), .Q (new_AGEMA_signal_14386) ) ;
    buf_clk new_AGEMA_reg_buffer_8538 ( .C (clk), .D (new_AGEMA_signal_14389), .Q (new_AGEMA_signal_14390) ) ;
    buf_clk new_AGEMA_reg_buffer_8542 ( .C (clk), .D (new_AGEMA_signal_14393), .Q (new_AGEMA_signal_14394) ) ;
    buf_clk new_AGEMA_reg_buffer_8546 ( .C (clk), .D (new_AGEMA_signal_14397), .Q (new_AGEMA_signal_14398) ) ;
    buf_clk new_AGEMA_reg_buffer_8550 ( .C (clk), .D (new_AGEMA_signal_14401), .Q (new_AGEMA_signal_14402) ) ;
    buf_clk new_AGEMA_reg_buffer_8554 ( .C (clk), .D (new_AGEMA_signal_14405), .Q (new_AGEMA_signal_14406) ) ;
    buf_clk new_AGEMA_reg_buffer_8558 ( .C (clk), .D (new_AGEMA_signal_14409), .Q (new_AGEMA_signal_14410) ) ;
    buf_clk new_AGEMA_reg_buffer_8562 ( .C (clk), .D (new_AGEMA_signal_14413), .Q (new_AGEMA_signal_14414) ) ;
    buf_clk new_AGEMA_reg_buffer_8566 ( .C (clk), .D (new_AGEMA_signal_14417), .Q (new_AGEMA_signal_14418) ) ;
    buf_clk new_AGEMA_reg_buffer_8570 ( .C (clk), .D (new_AGEMA_signal_14421), .Q (new_AGEMA_signal_14422) ) ;
    buf_clk new_AGEMA_reg_buffer_8574 ( .C (clk), .D (new_AGEMA_signal_14425), .Q (new_AGEMA_signal_14426) ) ;
    buf_clk new_AGEMA_reg_buffer_8578 ( .C (clk), .D (new_AGEMA_signal_14429), .Q (new_AGEMA_signal_14430) ) ;
    buf_clk new_AGEMA_reg_buffer_8582 ( .C (clk), .D (new_AGEMA_signal_14433), .Q (new_AGEMA_signal_14434) ) ;
    buf_clk new_AGEMA_reg_buffer_8586 ( .C (clk), .D (new_AGEMA_signal_14437), .Q (new_AGEMA_signal_14438) ) ;
    buf_clk new_AGEMA_reg_buffer_8590 ( .C (clk), .D (new_AGEMA_signal_14441), .Q (new_AGEMA_signal_14442) ) ;
    buf_clk new_AGEMA_reg_buffer_8594 ( .C (clk), .D (new_AGEMA_signal_14445), .Q (new_AGEMA_signal_14446) ) ;
    buf_clk new_AGEMA_reg_buffer_8598 ( .C (clk), .D (new_AGEMA_signal_14449), .Q (new_AGEMA_signal_14450) ) ;
    buf_clk new_AGEMA_reg_buffer_8602 ( .C (clk), .D (new_AGEMA_signal_14453), .Q (new_AGEMA_signal_14454) ) ;
    buf_clk new_AGEMA_reg_buffer_8606 ( .C (clk), .D (new_AGEMA_signal_14457), .Q (new_AGEMA_signal_14458) ) ;
    buf_clk new_AGEMA_reg_buffer_8610 ( .C (clk), .D (new_AGEMA_signal_14461), .Q (new_AGEMA_signal_14462) ) ;
    buf_clk new_AGEMA_reg_buffer_8614 ( .C (clk), .D (new_AGEMA_signal_14465), .Q (new_AGEMA_signal_14466) ) ;
    buf_clk new_AGEMA_reg_buffer_8618 ( .C (clk), .D (new_AGEMA_signal_14469), .Q (new_AGEMA_signal_14470) ) ;
    buf_clk new_AGEMA_reg_buffer_8622 ( .C (clk), .D (new_AGEMA_signal_14473), .Q (new_AGEMA_signal_14474) ) ;
    buf_clk new_AGEMA_reg_buffer_8626 ( .C (clk), .D (new_AGEMA_signal_14477), .Q (new_AGEMA_signal_14478) ) ;
    buf_clk new_AGEMA_reg_buffer_8630 ( .C (clk), .D (new_AGEMA_signal_14481), .Q (new_AGEMA_signal_14482) ) ;
    buf_clk new_AGEMA_reg_buffer_8634 ( .C (clk), .D (new_AGEMA_signal_14485), .Q (new_AGEMA_signal_14486) ) ;
    buf_clk new_AGEMA_reg_buffer_8638 ( .C (clk), .D (new_AGEMA_signal_14489), .Q (new_AGEMA_signal_14490) ) ;
    buf_clk new_AGEMA_reg_buffer_8642 ( .C (clk), .D (new_AGEMA_signal_14493), .Q (new_AGEMA_signal_14494) ) ;
    buf_clk new_AGEMA_reg_buffer_8646 ( .C (clk), .D (new_AGEMA_signal_14497), .Q (new_AGEMA_signal_14498) ) ;
    buf_clk new_AGEMA_reg_buffer_8650 ( .C (clk), .D (new_AGEMA_signal_14501), .Q (new_AGEMA_signal_14502) ) ;
    buf_clk new_AGEMA_reg_buffer_8654 ( .C (clk), .D (new_AGEMA_signal_14505), .Q (new_AGEMA_signal_14506) ) ;
    buf_clk new_AGEMA_reg_buffer_8658 ( .C (clk), .D (new_AGEMA_signal_14509), .Q (new_AGEMA_signal_14510) ) ;
    buf_clk new_AGEMA_reg_buffer_8662 ( .C (clk), .D (new_AGEMA_signal_14513), .Q (new_AGEMA_signal_14514) ) ;
    buf_clk new_AGEMA_reg_buffer_8666 ( .C (clk), .D (new_AGEMA_signal_14517), .Q (new_AGEMA_signal_14518) ) ;
    buf_clk new_AGEMA_reg_buffer_8670 ( .C (clk), .D (new_AGEMA_signal_14521), .Q (new_AGEMA_signal_14522) ) ;
    buf_clk new_AGEMA_reg_buffer_8674 ( .C (clk), .D (new_AGEMA_signal_14525), .Q (new_AGEMA_signal_14526) ) ;
    buf_clk new_AGEMA_reg_buffer_8678 ( .C (clk), .D (new_AGEMA_signal_14529), .Q (new_AGEMA_signal_14530) ) ;
    buf_clk new_AGEMA_reg_buffer_8682 ( .C (clk), .D (new_AGEMA_signal_14533), .Q (new_AGEMA_signal_14534) ) ;
    buf_clk new_AGEMA_reg_buffer_8686 ( .C (clk), .D (new_AGEMA_signal_14537), .Q (new_AGEMA_signal_14538) ) ;
    buf_clk new_AGEMA_reg_buffer_8690 ( .C (clk), .D (new_AGEMA_signal_14541), .Q (new_AGEMA_signal_14542) ) ;
    buf_clk new_AGEMA_reg_buffer_8694 ( .C (clk), .D (new_AGEMA_signal_14545), .Q (new_AGEMA_signal_14546) ) ;
    buf_clk new_AGEMA_reg_buffer_8698 ( .C (clk), .D (new_AGEMA_signal_14549), .Q (new_AGEMA_signal_14550) ) ;
    buf_clk new_AGEMA_reg_buffer_8702 ( .C (clk), .D (new_AGEMA_signal_14553), .Q (new_AGEMA_signal_14554) ) ;
    buf_clk new_AGEMA_reg_buffer_8706 ( .C (clk), .D (new_AGEMA_signal_14557), .Q (new_AGEMA_signal_14558) ) ;
    buf_clk new_AGEMA_reg_buffer_8710 ( .C (clk), .D (new_AGEMA_signal_14561), .Q (new_AGEMA_signal_14562) ) ;
    buf_clk new_AGEMA_reg_buffer_8714 ( .C (clk), .D (new_AGEMA_signal_14565), .Q (new_AGEMA_signal_14566) ) ;
    buf_clk new_AGEMA_reg_buffer_8718 ( .C (clk), .D (new_AGEMA_signal_14569), .Q (new_AGEMA_signal_14570) ) ;
    buf_clk new_AGEMA_reg_buffer_8722 ( .C (clk), .D (new_AGEMA_signal_14573), .Q (new_AGEMA_signal_14574) ) ;
    buf_clk new_AGEMA_reg_buffer_8726 ( .C (clk), .D (new_AGEMA_signal_14577), .Q (new_AGEMA_signal_14578) ) ;
    buf_clk new_AGEMA_reg_buffer_8730 ( .C (clk), .D (new_AGEMA_signal_14581), .Q (new_AGEMA_signal_14582) ) ;
    buf_clk new_AGEMA_reg_buffer_8734 ( .C (clk), .D (new_AGEMA_signal_14585), .Q (new_AGEMA_signal_14586) ) ;
    buf_clk new_AGEMA_reg_buffer_8738 ( .C (clk), .D (new_AGEMA_signal_14589), .Q (new_AGEMA_signal_14590) ) ;
    buf_clk new_AGEMA_reg_buffer_8742 ( .C (clk), .D (new_AGEMA_signal_14593), .Q (new_AGEMA_signal_14594) ) ;
    buf_clk new_AGEMA_reg_buffer_8746 ( .C (clk), .D (new_AGEMA_signal_14597), .Q (new_AGEMA_signal_14598) ) ;
    buf_clk new_AGEMA_reg_buffer_8750 ( .C (clk), .D (new_AGEMA_signal_14601), .Q (new_AGEMA_signal_14602) ) ;
    buf_clk new_AGEMA_reg_buffer_8754 ( .C (clk), .D (new_AGEMA_signal_14605), .Q (new_AGEMA_signal_14606) ) ;
    buf_clk new_AGEMA_reg_buffer_8758 ( .C (clk), .D (new_AGEMA_signal_14609), .Q (new_AGEMA_signal_14610) ) ;
    buf_clk new_AGEMA_reg_buffer_8762 ( .C (clk), .D (new_AGEMA_signal_14613), .Q (new_AGEMA_signal_14614) ) ;
    buf_clk new_AGEMA_reg_buffer_8766 ( .C (clk), .D (new_AGEMA_signal_14617), .Q (new_AGEMA_signal_14618) ) ;
    buf_clk new_AGEMA_reg_buffer_8770 ( .C (clk), .D (new_AGEMA_signal_14621), .Q (new_AGEMA_signal_14622) ) ;
    buf_clk new_AGEMA_reg_buffer_8774 ( .C (clk), .D (new_AGEMA_signal_14625), .Q (new_AGEMA_signal_14626) ) ;
    buf_clk new_AGEMA_reg_buffer_8778 ( .C (clk), .D (new_AGEMA_signal_14629), .Q (new_AGEMA_signal_14630) ) ;
    buf_clk new_AGEMA_reg_buffer_8782 ( .C (clk), .D (new_AGEMA_signal_14633), .Q (new_AGEMA_signal_14634) ) ;
    buf_clk new_AGEMA_reg_buffer_8786 ( .C (clk), .D (new_AGEMA_signal_14637), .Q (new_AGEMA_signal_14638) ) ;
    buf_clk new_AGEMA_reg_buffer_8790 ( .C (clk), .D (new_AGEMA_signal_14641), .Q (new_AGEMA_signal_14642) ) ;
    buf_clk new_AGEMA_reg_buffer_8794 ( .C (clk), .D (new_AGEMA_signal_14645), .Q (new_AGEMA_signal_14646) ) ;
    buf_clk new_AGEMA_reg_buffer_8798 ( .C (clk), .D (new_AGEMA_signal_14649), .Q (new_AGEMA_signal_14650) ) ;
    buf_clk new_AGEMA_reg_buffer_8802 ( .C (clk), .D (new_AGEMA_signal_14653), .Q (new_AGEMA_signal_14654) ) ;
    buf_clk new_AGEMA_reg_buffer_8806 ( .C (clk), .D (new_AGEMA_signal_14657), .Q (new_AGEMA_signal_14658) ) ;
    buf_clk new_AGEMA_reg_buffer_8810 ( .C (clk), .D (new_AGEMA_signal_14661), .Q (new_AGEMA_signal_14662) ) ;
    buf_clk new_AGEMA_reg_buffer_8814 ( .C (clk), .D (new_AGEMA_signal_14665), .Q (new_AGEMA_signal_14666) ) ;
    buf_clk new_AGEMA_reg_buffer_8818 ( .C (clk), .D (new_AGEMA_signal_14669), .Q (new_AGEMA_signal_14670) ) ;
    buf_clk new_AGEMA_reg_buffer_8822 ( .C (clk), .D (new_AGEMA_signal_14673), .Q (new_AGEMA_signal_14674) ) ;
    buf_clk new_AGEMA_reg_buffer_8826 ( .C (clk), .D (new_AGEMA_signal_14677), .Q (new_AGEMA_signal_14678) ) ;
    buf_clk new_AGEMA_reg_buffer_8830 ( .C (clk), .D (new_AGEMA_signal_14681), .Q (new_AGEMA_signal_14682) ) ;
    buf_clk new_AGEMA_reg_buffer_8834 ( .C (clk), .D (new_AGEMA_signal_14685), .Q (new_AGEMA_signal_14686) ) ;
    buf_clk new_AGEMA_reg_buffer_8838 ( .C (clk), .D (new_AGEMA_signal_14689), .Q (new_AGEMA_signal_14690) ) ;
    buf_clk new_AGEMA_reg_buffer_8842 ( .C (clk), .D (new_AGEMA_signal_14693), .Q (new_AGEMA_signal_14694) ) ;
    buf_clk new_AGEMA_reg_buffer_8846 ( .C (clk), .D (new_AGEMA_signal_14697), .Q (new_AGEMA_signal_14698) ) ;
    buf_clk new_AGEMA_reg_buffer_8850 ( .C (clk), .D (new_AGEMA_signal_14701), .Q (new_AGEMA_signal_14702) ) ;
    buf_clk new_AGEMA_reg_buffer_8854 ( .C (clk), .D (new_AGEMA_signal_14705), .Q (new_AGEMA_signal_14706) ) ;
    buf_clk new_AGEMA_reg_buffer_8858 ( .C (clk), .D (new_AGEMA_signal_14709), .Q (new_AGEMA_signal_14710) ) ;
    buf_clk new_AGEMA_reg_buffer_8862 ( .C (clk), .D (new_AGEMA_signal_14713), .Q (new_AGEMA_signal_14714) ) ;
    buf_clk new_AGEMA_reg_buffer_8866 ( .C (clk), .D (new_AGEMA_signal_14717), .Q (new_AGEMA_signal_14718) ) ;
    buf_clk new_AGEMA_reg_buffer_8870 ( .C (clk), .D (new_AGEMA_signal_14721), .Q (new_AGEMA_signal_14722) ) ;
    buf_clk new_AGEMA_reg_buffer_8874 ( .C (clk), .D (new_AGEMA_signal_14725), .Q (new_AGEMA_signal_14726) ) ;
    buf_clk new_AGEMA_reg_buffer_8878 ( .C (clk), .D (new_AGEMA_signal_14729), .Q (new_AGEMA_signal_14730) ) ;
    buf_clk new_AGEMA_reg_buffer_8882 ( .C (clk), .D (new_AGEMA_signal_14733), .Q (new_AGEMA_signal_14734) ) ;
    buf_clk new_AGEMA_reg_buffer_8886 ( .C (clk), .D (new_AGEMA_signal_14737), .Q (new_AGEMA_signal_14738) ) ;
    buf_clk new_AGEMA_reg_buffer_8890 ( .C (clk), .D (new_AGEMA_signal_14741), .Q (new_AGEMA_signal_14742) ) ;
    buf_clk new_AGEMA_reg_buffer_8894 ( .C (clk), .D (new_AGEMA_signal_14745), .Q (new_AGEMA_signal_14746) ) ;
    buf_clk new_AGEMA_reg_buffer_8898 ( .C (clk), .D (new_AGEMA_signal_14749), .Q (new_AGEMA_signal_14750) ) ;
    buf_clk new_AGEMA_reg_buffer_8902 ( .C (clk), .D (new_AGEMA_signal_14753), .Q (new_AGEMA_signal_14754) ) ;
    buf_clk new_AGEMA_reg_buffer_8906 ( .C (clk), .D (new_AGEMA_signal_14757), .Q (new_AGEMA_signal_14758) ) ;
    buf_clk new_AGEMA_reg_buffer_8910 ( .C (clk), .D (new_AGEMA_signal_14761), .Q (new_AGEMA_signal_14762) ) ;
    buf_clk new_AGEMA_reg_buffer_8914 ( .C (clk), .D (new_AGEMA_signal_14765), .Q (new_AGEMA_signal_14766) ) ;
    buf_clk new_AGEMA_reg_buffer_8918 ( .C (clk), .D (new_AGEMA_signal_14769), .Q (new_AGEMA_signal_14770) ) ;
    buf_clk new_AGEMA_reg_buffer_8922 ( .C (clk), .D (new_AGEMA_signal_14773), .Q (new_AGEMA_signal_14774) ) ;
    buf_clk new_AGEMA_reg_buffer_8926 ( .C (clk), .D (new_AGEMA_signal_14777), .Q (new_AGEMA_signal_14778) ) ;
    buf_clk new_AGEMA_reg_buffer_8930 ( .C (clk), .D (new_AGEMA_signal_14781), .Q (new_AGEMA_signal_14782) ) ;
    buf_clk new_AGEMA_reg_buffer_8934 ( .C (clk), .D (new_AGEMA_signal_14785), .Q (new_AGEMA_signal_14786) ) ;
    buf_clk new_AGEMA_reg_buffer_8938 ( .C (clk), .D (new_AGEMA_signal_14789), .Q (new_AGEMA_signal_14790) ) ;
    buf_clk new_AGEMA_reg_buffer_8942 ( .C (clk), .D (new_AGEMA_signal_14793), .Q (new_AGEMA_signal_14794) ) ;
    buf_clk new_AGEMA_reg_buffer_8946 ( .C (clk), .D (new_AGEMA_signal_14797), .Q (new_AGEMA_signal_14798) ) ;
    buf_clk new_AGEMA_reg_buffer_8950 ( .C (clk), .D (new_AGEMA_signal_14801), .Q (new_AGEMA_signal_14802) ) ;
    buf_clk new_AGEMA_reg_buffer_8954 ( .C (clk), .D (new_AGEMA_signal_14805), .Q (new_AGEMA_signal_14806) ) ;
    buf_clk new_AGEMA_reg_buffer_8958 ( .C (clk), .D (new_AGEMA_signal_14809), .Q (new_AGEMA_signal_14810) ) ;
    buf_clk new_AGEMA_reg_buffer_8962 ( .C (clk), .D (new_AGEMA_signal_14813), .Q (new_AGEMA_signal_14814) ) ;
    buf_clk new_AGEMA_reg_buffer_8966 ( .C (clk), .D (new_AGEMA_signal_14817), .Q (new_AGEMA_signal_14818) ) ;
    buf_clk new_AGEMA_reg_buffer_8970 ( .C (clk), .D (new_AGEMA_signal_14821), .Q (new_AGEMA_signal_14822) ) ;
    buf_clk new_AGEMA_reg_buffer_8974 ( .C (clk), .D (new_AGEMA_signal_14825), .Q (new_AGEMA_signal_14826) ) ;
    buf_clk new_AGEMA_reg_buffer_8978 ( .C (clk), .D (new_AGEMA_signal_14829), .Q (new_AGEMA_signal_14830) ) ;
    buf_clk new_AGEMA_reg_buffer_8982 ( .C (clk), .D (new_AGEMA_signal_14833), .Q (new_AGEMA_signal_14834) ) ;
    buf_clk new_AGEMA_reg_buffer_8986 ( .C (clk), .D (new_AGEMA_signal_14837), .Q (new_AGEMA_signal_14838) ) ;
    buf_clk new_AGEMA_reg_buffer_8990 ( .C (clk), .D (new_AGEMA_signal_14841), .Q (new_AGEMA_signal_14842) ) ;
    buf_clk new_AGEMA_reg_buffer_8994 ( .C (clk), .D (new_AGEMA_signal_14845), .Q (new_AGEMA_signal_14846) ) ;
    buf_clk new_AGEMA_reg_buffer_8998 ( .C (clk), .D (new_AGEMA_signal_14849), .Q (new_AGEMA_signal_14850) ) ;
    buf_clk new_AGEMA_reg_buffer_9002 ( .C (clk), .D (new_AGEMA_signal_14853), .Q (new_AGEMA_signal_14854) ) ;
    buf_clk new_AGEMA_reg_buffer_9006 ( .C (clk), .D (new_AGEMA_signal_14857), .Q (new_AGEMA_signal_14858) ) ;
    buf_clk new_AGEMA_reg_buffer_9010 ( .C (clk), .D (new_AGEMA_signal_14861), .Q (new_AGEMA_signal_14862) ) ;
    buf_clk new_AGEMA_reg_buffer_9014 ( .C (clk), .D (new_AGEMA_signal_14865), .Q (new_AGEMA_signal_14866) ) ;
    buf_clk new_AGEMA_reg_buffer_9018 ( .C (clk), .D (new_AGEMA_signal_14869), .Q (new_AGEMA_signal_14870) ) ;
    buf_clk new_AGEMA_reg_buffer_9022 ( .C (clk), .D (new_AGEMA_signal_14873), .Q (new_AGEMA_signal_14874) ) ;
    buf_clk new_AGEMA_reg_buffer_9026 ( .C (clk), .D (new_AGEMA_signal_14877), .Q (new_AGEMA_signal_14878) ) ;
    buf_clk new_AGEMA_reg_buffer_9030 ( .C (clk), .D (new_AGEMA_signal_14881), .Q (new_AGEMA_signal_14882) ) ;
    buf_clk new_AGEMA_reg_buffer_9034 ( .C (clk), .D (new_AGEMA_signal_14885), .Q (new_AGEMA_signal_14886) ) ;
    buf_clk new_AGEMA_reg_buffer_9038 ( .C (clk), .D (new_AGEMA_signal_14889), .Q (new_AGEMA_signal_14890) ) ;
    buf_clk new_AGEMA_reg_buffer_9042 ( .C (clk), .D (new_AGEMA_signal_14893), .Q (new_AGEMA_signal_14894) ) ;
    buf_clk new_AGEMA_reg_buffer_9046 ( .C (clk), .D (new_AGEMA_signal_14897), .Q (new_AGEMA_signal_14898) ) ;
    buf_clk new_AGEMA_reg_buffer_9050 ( .C (clk), .D (new_AGEMA_signal_14901), .Q (new_AGEMA_signal_14902) ) ;
    buf_clk new_AGEMA_reg_buffer_9054 ( .C (clk), .D (new_AGEMA_signal_14905), .Q (new_AGEMA_signal_14906) ) ;
    buf_clk new_AGEMA_reg_buffer_9058 ( .C (clk), .D (new_AGEMA_signal_14909), .Q (new_AGEMA_signal_14910) ) ;
    buf_clk new_AGEMA_reg_buffer_9062 ( .C (clk), .D (new_AGEMA_signal_14913), .Q (new_AGEMA_signal_14914) ) ;
    buf_clk new_AGEMA_reg_buffer_9066 ( .C (clk), .D (new_AGEMA_signal_14917), .Q (new_AGEMA_signal_14918) ) ;
    buf_clk new_AGEMA_reg_buffer_9070 ( .C (clk), .D (new_AGEMA_signal_14921), .Q (new_AGEMA_signal_14922) ) ;
    buf_clk new_AGEMA_reg_buffer_9074 ( .C (clk), .D (new_AGEMA_signal_14925), .Q (new_AGEMA_signal_14926) ) ;
    buf_clk new_AGEMA_reg_buffer_9078 ( .C (clk), .D (new_AGEMA_signal_14929), .Q (new_AGEMA_signal_14930) ) ;
    buf_clk new_AGEMA_reg_buffer_9082 ( .C (clk), .D (new_AGEMA_signal_14933), .Q (new_AGEMA_signal_14934) ) ;
    buf_clk new_AGEMA_reg_buffer_9086 ( .C (clk), .D (new_AGEMA_signal_14937), .Q (new_AGEMA_signal_14938) ) ;
    buf_clk new_AGEMA_reg_buffer_9090 ( .C (clk), .D (new_AGEMA_signal_14941), .Q (new_AGEMA_signal_14942) ) ;
    buf_clk new_AGEMA_reg_buffer_9094 ( .C (clk), .D (new_AGEMA_signal_14945), .Q (new_AGEMA_signal_14946) ) ;
    buf_clk new_AGEMA_reg_buffer_9098 ( .C (clk), .D (new_AGEMA_signal_14949), .Q (new_AGEMA_signal_14950) ) ;
    buf_clk new_AGEMA_reg_buffer_9102 ( .C (clk), .D (new_AGEMA_signal_14953), .Q (new_AGEMA_signal_14954) ) ;
    buf_clk new_AGEMA_reg_buffer_9106 ( .C (clk), .D (new_AGEMA_signal_14957), .Q (new_AGEMA_signal_14958) ) ;
    buf_clk new_AGEMA_reg_buffer_9110 ( .C (clk), .D (new_AGEMA_signal_14961), .Q (new_AGEMA_signal_14962) ) ;
    buf_clk new_AGEMA_reg_buffer_9114 ( .C (clk), .D (new_AGEMA_signal_14965), .Q (new_AGEMA_signal_14966) ) ;
    buf_clk new_AGEMA_reg_buffer_9118 ( .C (clk), .D (new_AGEMA_signal_14969), .Q (new_AGEMA_signal_14970) ) ;
    buf_clk new_AGEMA_reg_buffer_9122 ( .C (clk), .D (new_AGEMA_signal_14973), .Q (new_AGEMA_signal_14974) ) ;
    buf_clk new_AGEMA_reg_buffer_9126 ( .C (clk), .D (new_AGEMA_signal_14977), .Q (new_AGEMA_signal_14978) ) ;
    buf_clk new_AGEMA_reg_buffer_9130 ( .C (clk), .D (new_AGEMA_signal_14981), .Q (new_AGEMA_signal_14982) ) ;
    buf_clk new_AGEMA_reg_buffer_9134 ( .C (clk), .D (new_AGEMA_signal_14985), .Q (new_AGEMA_signal_14986) ) ;
    buf_clk new_AGEMA_reg_buffer_9138 ( .C (clk), .D (new_AGEMA_signal_14989), .Q (new_AGEMA_signal_14990) ) ;
    buf_clk new_AGEMA_reg_buffer_9142 ( .C (clk), .D (new_AGEMA_signal_14993), .Q (new_AGEMA_signal_14994) ) ;
    buf_clk new_AGEMA_reg_buffer_9146 ( .C (clk), .D (new_AGEMA_signal_14997), .Q (new_AGEMA_signal_14998) ) ;
    buf_clk new_AGEMA_reg_buffer_9150 ( .C (clk), .D (new_AGEMA_signal_15001), .Q (new_AGEMA_signal_15002) ) ;
    buf_clk new_AGEMA_reg_buffer_9154 ( .C (clk), .D (new_AGEMA_signal_15005), .Q (new_AGEMA_signal_15006) ) ;
    buf_clk new_AGEMA_reg_buffer_9158 ( .C (clk), .D (new_AGEMA_signal_15009), .Q (new_AGEMA_signal_15010) ) ;
    buf_clk new_AGEMA_reg_buffer_9162 ( .C (clk), .D (new_AGEMA_signal_15013), .Q (new_AGEMA_signal_15014) ) ;
    buf_clk new_AGEMA_reg_buffer_9166 ( .C (clk), .D (new_AGEMA_signal_15017), .Q (new_AGEMA_signal_15018) ) ;
    buf_clk new_AGEMA_reg_buffer_9170 ( .C (clk), .D (new_AGEMA_signal_15021), .Q (new_AGEMA_signal_15022) ) ;
    buf_clk new_AGEMA_reg_buffer_9174 ( .C (clk), .D (new_AGEMA_signal_15025), .Q (new_AGEMA_signal_15026) ) ;
    buf_clk new_AGEMA_reg_buffer_9178 ( .C (clk), .D (new_AGEMA_signal_15029), .Q (new_AGEMA_signal_15030) ) ;
    buf_clk new_AGEMA_reg_buffer_9182 ( .C (clk), .D (new_AGEMA_signal_15033), .Q (new_AGEMA_signal_15034) ) ;
    buf_clk new_AGEMA_reg_buffer_9186 ( .C (clk), .D (new_AGEMA_signal_15037), .Q (new_AGEMA_signal_15038) ) ;
    buf_clk new_AGEMA_reg_buffer_9190 ( .C (clk), .D (new_AGEMA_signal_15041), .Q (new_AGEMA_signal_15042) ) ;
    buf_clk new_AGEMA_reg_buffer_9194 ( .C (clk), .D (new_AGEMA_signal_15045), .Q (new_AGEMA_signal_15046) ) ;
    buf_clk new_AGEMA_reg_buffer_9198 ( .C (clk), .D (new_AGEMA_signal_15049), .Q (new_AGEMA_signal_15050) ) ;
    buf_clk new_AGEMA_reg_buffer_9202 ( .C (clk), .D (new_AGEMA_signal_15053), .Q (new_AGEMA_signal_15054) ) ;
    buf_clk new_AGEMA_reg_buffer_9206 ( .C (clk), .D (new_AGEMA_signal_15057), .Q (new_AGEMA_signal_15058) ) ;
    buf_clk new_AGEMA_reg_buffer_9210 ( .C (clk), .D (new_AGEMA_signal_15061), .Q (new_AGEMA_signal_15062) ) ;
    buf_clk new_AGEMA_reg_buffer_9214 ( .C (clk), .D (new_AGEMA_signal_15065), .Q (new_AGEMA_signal_15066) ) ;
    buf_clk new_AGEMA_reg_buffer_9218 ( .C (clk), .D (new_AGEMA_signal_15069), .Q (new_AGEMA_signal_15070) ) ;
    buf_clk new_AGEMA_reg_buffer_9222 ( .C (clk), .D (new_AGEMA_signal_15073), .Q (new_AGEMA_signal_15074) ) ;
    buf_clk new_AGEMA_reg_buffer_9226 ( .C (clk), .D (new_AGEMA_signal_15077), .Q (new_AGEMA_signal_15078) ) ;
    buf_clk new_AGEMA_reg_buffer_9230 ( .C (clk), .D (new_AGEMA_signal_15081), .Q (new_AGEMA_signal_15082) ) ;
    buf_clk new_AGEMA_reg_buffer_9234 ( .C (clk), .D (new_AGEMA_signal_15085), .Q (new_AGEMA_signal_15086) ) ;
    buf_clk new_AGEMA_reg_buffer_9238 ( .C (clk), .D (new_AGEMA_signal_15089), .Q (new_AGEMA_signal_15090) ) ;
    buf_clk new_AGEMA_reg_buffer_9242 ( .C (clk), .D (new_AGEMA_signal_15093), .Q (new_AGEMA_signal_15094) ) ;
    buf_clk new_AGEMA_reg_buffer_9246 ( .C (clk), .D (new_AGEMA_signal_15097), .Q (new_AGEMA_signal_15098) ) ;
    buf_clk new_AGEMA_reg_buffer_9250 ( .C (clk), .D (new_AGEMA_signal_15101), .Q (new_AGEMA_signal_15102) ) ;
    buf_clk new_AGEMA_reg_buffer_9254 ( .C (clk), .D (new_AGEMA_signal_15105), .Q (new_AGEMA_signal_15106) ) ;
    buf_clk new_AGEMA_reg_buffer_9258 ( .C (clk), .D (new_AGEMA_signal_15109), .Q (new_AGEMA_signal_15110) ) ;
    buf_clk new_AGEMA_reg_buffer_9262 ( .C (clk), .D (new_AGEMA_signal_15113), .Q (new_AGEMA_signal_15114) ) ;
    buf_clk new_AGEMA_reg_buffer_9266 ( .C (clk), .D (new_AGEMA_signal_15117), .Q (new_AGEMA_signal_15118) ) ;
    buf_clk new_AGEMA_reg_buffer_9270 ( .C (clk), .D (new_AGEMA_signal_15121), .Q (new_AGEMA_signal_15122) ) ;
    buf_clk new_AGEMA_reg_buffer_9274 ( .C (clk), .D (new_AGEMA_signal_15125), .Q (new_AGEMA_signal_15126) ) ;
    buf_clk new_AGEMA_reg_buffer_9278 ( .C (clk), .D (new_AGEMA_signal_15129), .Q (new_AGEMA_signal_15130) ) ;
    buf_clk new_AGEMA_reg_buffer_9282 ( .C (clk), .D (new_AGEMA_signal_15133), .Q (new_AGEMA_signal_15134) ) ;
    buf_clk new_AGEMA_reg_buffer_9286 ( .C (clk), .D (new_AGEMA_signal_15137), .Q (new_AGEMA_signal_15138) ) ;
    buf_clk new_AGEMA_reg_buffer_9290 ( .C (clk), .D (new_AGEMA_signal_15141), .Q (new_AGEMA_signal_15142) ) ;
    buf_clk new_AGEMA_reg_buffer_9294 ( .C (clk), .D (new_AGEMA_signal_15145), .Q (new_AGEMA_signal_15146) ) ;
    buf_clk new_AGEMA_reg_buffer_9298 ( .C (clk), .D (new_AGEMA_signal_15149), .Q (new_AGEMA_signal_15150) ) ;
    buf_clk new_AGEMA_reg_buffer_9302 ( .C (clk), .D (new_AGEMA_signal_15153), .Q (new_AGEMA_signal_15154) ) ;
    buf_clk new_AGEMA_reg_buffer_9306 ( .C (clk), .D (new_AGEMA_signal_15157), .Q (new_AGEMA_signal_15158) ) ;
    buf_clk new_AGEMA_reg_buffer_9310 ( .C (clk), .D (new_AGEMA_signal_15161), .Q (new_AGEMA_signal_15162) ) ;
    buf_clk new_AGEMA_reg_buffer_9314 ( .C (clk), .D (new_AGEMA_signal_15165), .Q (new_AGEMA_signal_15166) ) ;
    buf_clk new_AGEMA_reg_buffer_9318 ( .C (clk), .D (new_AGEMA_signal_15169), .Q (new_AGEMA_signal_15170) ) ;
    buf_clk new_AGEMA_reg_buffer_9322 ( .C (clk), .D (new_AGEMA_signal_15173), .Q (new_AGEMA_signal_15174) ) ;
    buf_clk new_AGEMA_reg_buffer_9326 ( .C (clk), .D (new_AGEMA_signal_15177), .Q (new_AGEMA_signal_15178) ) ;
    buf_clk new_AGEMA_reg_buffer_9330 ( .C (clk), .D (new_AGEMA_signal_15181), .Q (new_AGEMA_signal_15182) ) ;
    buf_clk new_AGEMA_reg_buffer_9334 ( .C (clk), .D (new_AGEMA_signal_15185), .Q (new_AGEMA_signal_15186) ) ;
    buf_clk new_AGEMA_reg_buffer_9338 ( .C (clk), .D (new_AGEMA_signal_15189), .Q (new_AGEMA_signal_15190) ) ;
    buf_clk new_AGEMA_reg_buffer_9342 ( .C (clk), .D (new_AGEMA_signal_15193), .Q (new_AGEMA_signal_15194) ) ;
    buf_clk new_AGEMA_reg_buffer_9346 ( .C (clk), .D (new_AGEMA_signal_15197), .Q (new_AGEMA_signal_15198) ) ;
    buf_clk new_AGEMA_reg_buffer_9350 ( .C (clk), .D (new_AGEMA_signal_15201), .Q (new_AGEMA_signal_15202) ) ;
    buf_clk new_AGEMA_reg_buffer_9354 ( .C (clk), .D (new_AGEMA_signal_15205), .Q (new_AGEMA_signal_15206) ) ;
    buf_clk new_AGEMA_reg_buffer_9358 ( .C (clk), .D (new_AGEMA_signal_15209), .Q (new_AGEMA_signal_15210) ) ;
    buf_clk new_AGEMA_reg_buffer_9362 ( .C (clk), .D (new_AGEMA_signal_15213), .Q (new_AGEMA_signal_15214) ) ;
    buf_clk new_AGEMA_reg_buffer_9366 ( .C (clk), .D (new_AGEMA_signal_15217), .Q (new_AGEMA_signal_15218) ) ;
    buf_clk new_AGEMA_reg_buffer_9370 ( .C (clk), .D (new_AGEMA_signal_15221), .Q (new_AGEMA_signal_15222) ) ;
    buf_clk new_AGEMA_reg_buffer_9374 ( .C (clk), .D (new_AGEMA_signal_15225), .Q (new_AGEMA_signal_15226) ) ;
    buf_clk new_AGEMA_reg_buffer_9378 ( .C (clk), .D (new_AGEMA_signal_15229), .Q (new_AGEMA_signal_15230) ) ;
    buf_clk new_AGEMA_reg_buffer_9382 ( .C (clk), .D (new_AGEMA_signal_15233), .Q (new_AGEMA_signal_15234) ) ;
    buf_clk new_AGEMA_reg_buffer_9386 ( .C (clk), .D (new_AGEMA_signal_15237), .Q (new_AGEMA_signal_15238) ) ;
    buf_clk new_AGEMA_reg_buffer_9390 ( .C (clk), .D (new_AGEMA_signal_15241), .Q (new_AGEMA_signal_15242) ) ;
    buf_clk new_AGEMA_reg_buffer_9394 ( .C (clk), .D (new_AGEMA_signal_15245), .Q (new_AGEMA_signal_15246) ) ;
    buf_clk new_AGEMA_reg_buffer_9398 ( .C (clk), .D (new_AGEMA_signal_15249), .Q (new_AGEMA_signal_15250) ) ;
    buf_clk new_AGEMA_reg_buffer_9402 ( .C (clk), .D (new_AGEMA_signal_15253), .Q (new_AGEMA_signal_15254) ) ;
    buf_clk new_AGEMA_reg_buffer_9406 ( .C (clk), .D (new_AGEMA_signal_15257), .Q (new_AGEMA_signal_15258) ) ;
    buf_clk new_AGEMA_reg_buffer_9410 ( .C (clk), .D (new_AGEMA_signal_15261), .Q (new_AGEMA_signal_15262) ) ;
    buf_clk new_AGEMA_reg_buffer_9414 ( .C (clk), .D (new_AGEMA_signal_15265), .Q (new_AGEMA_signal_15266) ) ;
    buf_clk new_AGEMA_reg_buffer_9418 ( .C (clk), .D (new_AGEMA_signal_15269), .Q (new_AGEMA_signal_15270) ) ;
    buf_clk new_AGEMA_reg_buffer_9422 ( .C (clk), .D (new_AGEMA_signal_15273), .Q (new_AGEMA_signal_15274) ) ;
    buf_clk new_AGEMA_reg_buffer_9426 ( .C (clk), .D (new_AGEMA_signal_15277), .Q (new_AGEMA_signal_15278) ) ;
    buf_clk new_AGEMA_reg_buffer_9430 ( .C (clk), .D (new_AGEMA_signal_15281), .Q (new_AGEMA_signal_15282) ) ;
    buf_clk new_AGEMA_reg_buffer_9434 ( .C (clk), .D (new_AGEMA_signal_15285), .Q (new_AGEMA_signal_15286) ) ;
    buf_clk new_AGEMA_reg_buffer_9438 ( .C (clk), .D (new_AGEMA_signal_15289), .Q (new_AGEMA_signal_15290) ) ;
    buf_clk new_AGEMA_reg_buffer_9442 ( .C (clk), .D (new_AGEMA_signal_15293), .Q (new_AGEMA_signal_15294) ) ;
    buf_clk new_AGEMA_reg_buffer_9446 ( .C (clk), .D (new_AGEMA_signal_15297), .Q (new_AGEMA_signal_15298) ) ;
    buf_clk new_AGEMA_reg_buffer_9450 ( .C (clk), .D (new_AGEMA_signal_15301), .Q (new_AGEMA_signal_15302) ) ;
    buf_clk new_AGEMA_reg_buffer_9454 ( .C (clk), .D (new_AGEMA_signal_15305), .Q (new_AGEMA_signal_15306) ) ;
    buf_clk new_AGEMA_reg_buffer_9458 ( .C (clk), .D (new_AGEMA_signal_15309), .Q (new_AGEMA_signal_15310) ) ;
    buf_clk new_AGEMA_reg_buffer_9462 ( .C (clk), .D (new_AGEMA_signal_15313), .Q (new_AGEMA_signal_15314) ) ;
    buf_clk new_AGEMA_reg_buffer_9466 ( .C (clk), .D (new_AGEMA_signal_15317), .Q (new_AGEMA_signal_15318) ) ;
    buf_clk new_AGEMA_reg_buffer_9470 ( .C (clk), .D (new_AGEMA_signal_15321), .Q (new_AGEMA_signal_15322) ) ;
    buf_clk new_AGEMA_reg_buffer_9474 ( .C (clk), .D (new_AGEMA_signal_15325), .Q (new_AGEMA_signal_15326) ) ;
    buf_clk new_AGEMA_reg_buffer_9478 ( .C (clk), .D (new_AGEMA_signal_15329), .Q (new_AGEMA_signal_15330) ) ;
    buf_clk new_AGEMA_reg_buffer_9482 ( .C (clk), .D (new_AGEMA_signal_15333), .Q (new_AGEMA_signal_15334) ) ;
    buf_clk new_AGEMA_reg_buffer_9486 ( .C (clk), .D (new_AGEMA_signal_15337), .Q (new_AGEMA_signal_15338) ) ;
    buf_clk new_AGEMA_reg_buffer_9490 ( .C (clk), .D (new_AGEMA_signal_15341), .Q (new_AGEMA_signal_15342) ) ;
    buf_clk new_AGEMA_reg_buffer_9494 ( .C (clk), .D (new_AGEMA_signal_15345), .Q (new_AGEMA_signal_15346) ) ;
    buf_clk new_AGEMA_reg_buffer_9498 ( .C (clk), .D (new_AGEMA_signal_15349), .Q (new_AGEMA_signal_15350) ) ;
    buf_clk new_AGEMA_reg_buffer_9502 ( .C (clk), .D (new_AGEMA_signal_15353), .Q (new_AGEMA_signal_15354) ) ;
    buf_clk new_AGEMA_reg_buffer_9506 ( .C (clk), .D (new_AGEMA_signal_15357), .Q (new_AGEMA_signal_15358) ) ;
    buf_clk new_AGEMA_reg_buffer_9510 ( .C (clk), .D (new_AGEMA_signal_15361), .Q (new_AGEMA_signal_15362) ) ;
    buf_clk new_AGEMA_reg_buffer_9514 ( .C (clk), .D (new_AGEMA_signal_15365), .Q (new_AGEMA_signal_15366) ) ;
    buf_clk new_AGEMA_reg_buffer_9518 ( .C (clk), .D (new_AGEMA_signal_15369), .Q (new_AGEMA_signal_15370) ) ;
    buf_clk new_AGEMA_reg_buffer_9522 ( .C (clk), .D (new_AGEMA_signal_15373), .Q (new_AGEMA_signal_15374) ) ;
    buf_clk new_AGEMA_reg_buffer_9526 ( .C (clk), .D (new_AGEMA_signal_15377), .Q (new_AGEMA_signal_15378) ) ;
    buf_clk new_AGEMA_reg_buffer_9530 ( .C (clk), .D (new_AGEMA_signal_15381), .Q (new_AGEMA_signal_15382) ) ;
    buf_clk new_AGEMA_reg_buffer_9534 ( .C (clk), .D (new_AGEMA_signal_15385), .Q (new_AGEMA_signal_15386) ) ;
    buf_clk new_AGEMA_reg_buffer_9538 ( .C (clk), .D (new_AGEMA_signal_15389), .Q (new_AGEMA_signal_15390) ) ;
    buf_clk new_AGEMA_reg_buffer_9542 ( .C (clk), .D (new_AGEMA_signal_15393), .Q (new_AGEMA_signal_15394) ) ;
    buf_clk new_AGEMA_reg_buffer_9546 ( .C (clk), .D (new_AGEMA_signal_15397), .Q (new_AGEMA_signal_15398) ) ;
    buf_clk new_AGEMA_reg_buffer_9550 ( .C (clk), .D (new_AGEMA_signal_15401), .Q (new_AGEMA_signal_15402) ) ;
    buf_clk new_AGEMA_reg_buffer_9554 ( .C (clk), .D (new_AGEMA_signal_15405), .Q (new_AGEMA_signal_15406) ) ;
    buf_clk new_AGEMA_reg_buffer_9557 ( .C (clk), .D (new_AGEMA_signal_15408), .Q (new_AGEMA_signal_15409) ) ;
    buf_clk new_AGEMA_reg_buffer_9560 ( .C (clk), .D (new_AGEMA_signal_15411), .Q (new_AGEMA_signal_15412) ) ;
    buf_clk new_AGEMA_reg_buffer_9563 ( .C (clk), .D (new_AGEMA_signal_15414), .Q (new_AGEMA_signal_15415) ) ;
    buf_clk new_AGEMA_reg_buffer_9566 ( .C (clk), .D (new_AGEMA_signal_15417), .Q (new_AGEMA_signal_15418) ) ;
    buf_clk new_AGEMA_reg_buffer_9569 ( .C (clk), .D (new_AGEMA_signal_15420), .Q (new_AGEMA_signal_15421) ) ;
    buf_clk new_AGEMA_reg_buffer_9572 ( .C (clk), .D (new_AGEMA_signal_15423), .Q (new_AGEMA_signal_15424) ) ;
    buf_clk new_AGEMA_reg_buffer_9575 ( .C (clk), .D (new_AGEMA_signal_15426), .Q (new_AGEMA_signal_15427) ) ;
    buf_clk new_AGEMA_reg_buffer_9578 ( .C (clk), .D (new_AGEMA_signal_15429), .Q (new_AGEMA_signal_15430) ) ;
    buf_clk new_AGEMA_reg_buffer_9581 ( .C (clk), .D (new_AGEMA_signal_15432), .Q (new_AGEMA_signal_15433) ) ;
    buf_clk new_AGEMA_reg_buffer_9584 ( .C (clk), .D (new_AGEMA_signal_15435), .Q (new_AGEMA_signal_15436) ) ;
    buf_clk new_AGEMA_reg_buffer_9587 ( .C (clk), .D (new_AGEMA_signal_15438), .Q (new_AGEMA_signal_15439) ) ;
    buf_clk new_AGEMA_reg_buffer_9590 ( .C (clk), .D (new_AGEMA_signal_15441), .Q (new_AGEMA_signal_15442) ) ;
    buf_clk new_AGEMA_reg_buffer_9593 ( .C (clk), .D (new_AGEMA_signal_15444), .Q (new_AGEMA_signal_15445) ) ;
    buf_clk new_AGEMA_reg_buffer_9596 ( .C (clk), .D (new_AGEMA_signal_15447), .Q (new_AGEMA_signal_15448) ) ;
    buf_clk new_AGEMA_reg_buffer_9599 ( .C (clk), .D (new_AGEMA_signal_15450), .Q (new_AGEMA_signal_15451) ) ;
    buf_clk new_AGEMA_reg_buffer_9602 ( .C (clk), .D (new_AGEMA_signal_15453), .Q (new_AGEMA_signal_15454) ) ;
    buf_clk new_AGEMA_reg_buffer_9605 ( .C (clk), .D (new_AGEMA_signal_15456), .Q (new_AGEMA_signal_15457) ) ;
    buf_clk new_AGEMA_reg_buffer_9608 ( .C (clk), .D (new_AGEMA_signal_15459), .Q (new_AGEMA_signal_15460) ) ;
    buf_clk new_AGEMA_reg_buffer_9611 ( .C (clk), .D (new_AGEMA_signal_15462), .Q (new_AGEMA_signal_15463) ) ;
    buf_clk new_AGEMA_reg_buffer_9614 ( .C (clk), .D (new_AGEMA_signal_15465), .Q (new_AGEMA_signal_15466) ) ;
    buf_clk new_AGEMA_reg_buffer_9617 ( .C (clk), .D (new_AGEMA_signal_15468), .Q (new_AGEMA_signal_15469) ) ;
    buf_clk new_AGEMA_reg_buffer_9620 ( .C (clk), .D (new_AGEMA_signal_15471), .Q (new_AGEMA_signal_15472) ) ;
    buf_clk new_AGEMA_reg_buffer_9623 ( .C (clk), .D (new_AGEMA_signal_15474), .Q (new_AGEMA_signal_15475) ) ;
    buf_clk new_AGEMA_reg_buffer_9626 ( .C (clk), .D (new_AGEMA_signal_15477), .Q (new_AGEMA_signal_15478) ) ;
    buf_clk new_AGEMA_reg_buffer_9629 ( .C (clk), .D (new_AGEMA_signal_15480), .Q (new_AGEMA_signal_15481) ) ;
    buf_clk new_AGEMA_reg_buffer_9632 ( .C (clk), .D (new_AGEMA_signal_15483), .Q (new_AGEMA_signal_15484) ) ;
    buf_clk new_AGEMA_reg_buffer_9635 ( .C (clk), .D (new_AGEMA_signal_15486), .Q (new_AGEMA_signal_15487) ) ;
    buf_clk new_AGEMA_reg_buffer_9638 ( .C (clk), .D (new_AGEMA_signal_15489), .Q (new_AGEMA_signal_15490) ) ;
    buf_clk new_AGEMA_reg_buffer_9641 ( .C (clk), .D (new_AGEMA_signal_15492), .Q (new_AGEMA_signal_15493) ) ;
    buf_clk new_AGEMA_reg_buffer_9644 ( .C (clk), .D (new_AGEMA_signal_15495), .Q (new_AGEMA_signal_15496) ) ;
    buf_clk new_AGEMA_reg_buffer_9647 ( .C (clk), .D (new_AGEMA_signal_15498), .Q (new_AGEMA_signal_15499) ) ;
    buf_clk new_AGEMA_reg_buffer_9650 ( .C (clk), .D (new_AGEMA_signal_15501), .Q (new_AGEMA_signal_15502) ) ;
    buf_clk new_AGEMA_reg_buffer_9653 ( .C (clk), .D (new_AGEMA_signal_15504), .Q (new_AGEMA_signal_15505) ) ;
    buf_clk new_AGEMA_reg_buffer_9656 ( .C (clk), .D (new_AGEMA_signal_15507), .Q (new_AGEMA_signal_15508) ) ;
    buf_clk new_AGEMA_reg_buffer_9659 ( .C (clk), .D (new_AGEMA_signal_15510), .Q (new_AGEMA_signal_15511) ) ;
    buf_clk new_AGEMA_reg_buffer_9662 ( .C (clk), .D (new_AGEMA_signal_15513), .Q (new_AGEMA_signal_15514) ) ;
    buf_clk new_AGEMA_reg_buffer_9665 ( .C (clk), .D (new_AGEMA_signal_15516), .Q (new_AGEMA_signal_15517) ) ;
    buf_clk new_AGEMA_reg_buffer_9668 ( .C (clk), .D (new_AGEMA_signal_15519), .Q (new_AGEMA_signal_15520) ) ;
    buf_clk new_AGEMA_reg_buffer_9671 ( .C (clk), .D (new_AGEMA_signal_15522), .Q (new_AGEMA_signal_15523) ) ;
    buf_clk new_AGEMA_reg_buffer_9674 ( .C (clk), .D (new_AGEMA_signal_15525), .Q (new_AGEMA_signal_15526) ) ;
    buf_clk new_AGEMA_reg_buffer_9677 ( .C (clk), .D (new_AGEMA_signal_15528), .Q (new_AGEMA_signal_15529) ) ;
    buf_clk new_AGEMA_reg_buffer_9680 ( .C (clk), .D (new_AGEMA_signal_15531), .Q (new_AGEMA_signal_15532) ) ;
    buf_clk new_AGEMA_reg_buffer_9683 ( .C (clk), .D (new_AGEMA_signal_15534), .Q (new_AGEMA_signal_15535) ) ;
    buf_clk new_AGEMA_reg_buffer_9686 ( .C (clk), .D (new_AGEMA_signal_15537), .Q (new_AGEMA_signal_15538) ) ;
    buf_clk new_AGEMA_reg_buffer_9689 ( .C (clk), .D (new_AGEMA_signal_15540), .Q (new_AGEMA_signal_15541) ) ;
    buf_clk new_AGEMA_reg_buffer_9692 ( .C (clk), .D (new_AGEMA_signal_15543), .Q (new_AGEMA_signal_15544) ) ;
    buf_clk new_AGEMA_reg_buffer_9695 ( .C (clk), .D (new_AGEMA_signal_15546), .Q (new_AGEMA_signal_15547) ) ;
    buf_clk new_AGEMA_reg_buffer_9698 ( .C (clk), .D (new_AGEMA_signal_15549), .Q (new_AGEMA_signal_15550) ) ;
    buf_clk new_AGEMA_reg_buffer_9701 ( .C (clk), .D (new_AGEMA_signal_15552), .Q (new_AGEMA_signal_15553) ) ;
    buf_clk new_AGEMA_reg_buffer_9704 ( .C (clk), .D (new_AGEMA_signal_15555), .Q (new_AGEMA_signal_15556) ) ;
    buf_clk new_AGEMA_reg_buffer_9707 ( .C (clk), .D (new_AGEMA_signal_15558), .Q (new_AGEMA_signal_15559) ) ;
    buf_clk new_AGEMA_reg_buffer_9710 ( .C (clk), .D (new_AGEMA_signal_15561), .Q (new_AGEMA_signal_15562) ) ;
    buf_clk new_AGEMA_reg_buffer_9713 ( .C (clk), .D (new_AGEMA_signal_15564), .Q (new_AGEMA_signal_15565) ) ;
    buf_clk new_AGEMA_reg_buffer_9716 ( .C (clk), .D (new_AGEMA_signal_15567), .Q (new_AGEMA_signal_15568) ) ;
    buf_clk new_AGEMA_reg_buffer_9719 ( .C (clk), .D (new_AGEMA_signal_15570), .Q (new_AGEMA_signal_15571) ) ;
    buf_clk new_AGEMA_reg_buffer_9722 ( .C (clk), .D (new_AGEMA_signal_15573), .Q (new_AGEMA_signal_15574) ) ;
    buf_clk new_AGEMA_reg_buffer_9725 ( .C (clk), .D (new_AGEMA_signal_15576), .Q (new_AGEMA_signal_15577) ) ;
    buf_clk new_AGEMA_reg_buffer_9728 ( .C (clk), .D (new_AGEMA_signal_15579), .Q (new_AGEMA_signal_15580) ) ;
    buf_clk new_AGEMA_reg_buffer_9731 ( .C (clk), .D (new_AGEMA_signal_15582), .Q (new_AGEMA_signal_15583) ) ;
    buf_clk new_AGEMA_reg_buffer_9734 ( .C (clk), .D (new_AGEMA_signal_15585), .Q (new_AGEMA_signal_15586) ) ;
    buf_clk new_AGEMA_reg_buffer_9737 ( .C (clk), .D (new_AGEMA_signal_15588), .Q (new_AGEMA_signal_15589) ) ;
    buf_clk new_AGEMA_reg_buffer_9740 ( .C (clk), .D (new_AGEMA_signal_15591), .Q (new_AGEMA_signal_15592) ) ;
    buf_clk new_AGEMA_reg_buffer_9743 ( .C (clk), .D (new_AGEMA_signal_15594), .Q (new_AGEMA_signal_15595) ) ;
    buf_clk new_AGEMA_reg_buffer_9746 ( .C (clk), .D (new_AGEMA_signal_15597), .Q (new_AGEMA_signal_15598) ) ;
    buf_clk new_AGEMA_reg_buffer_9749 ( .C (clk), .D (new_AGEMA_signal_15600), .Q (new_AGEMA_signal_15601) ) ;
    buf_clk new_AGEMA_reg_buffer_9752 ( .C (clk), .D (new_AGEMA_signal_15603), .Q (new_AGEMA_signal_15604) ) ;
    buf_clk new_AGEMA_reg_buffer_9755 ( .C (clk), .D (new_AGEMA_signal_15606), .Q (new_AGEMA_signal_15607) ) ;
    buf_clk new_AGEMA_reg_buffer_9758 ( .C (clk), .D (new_AGEMA_signal_15609), .Q (new_AGEMA_signal_15610) ) ;
    buf_clk new_AGEMA_reg_buffer_9761 ( .C (clk), .D (new_AGEMA_signal_15612), .Q (new_AGEMA_signal_15613) ) ;
    buf_clk new_AGEMA_reg_buffer_9764 ( .C (clk), .D (new_AGEMA_signal_15615), .Q (new_AGEMA_signal_15616) ) ;
    buf_clk new_AGEMA_reg_buffer_9767 ( .C (clk), .D (new_AGEMA_signal_15618), .Q (new_AGEMA_signal_15619) ) ;
    buf_clk new_AGEMA_reg_buffer_9770 ( .C (clk), .D (new_AGEMA_signal_15621), .Q (new_AGEMA_signal_15622) ) ;
    buf_clk new_AGEMA_reg_buffer_9773 ( .C (clk), .D (new_AGEMA_signal_15624), .Q (new_AGEMA_signal_15625) ) ;
    buf_clk new_AGEMA_reg_buffer_9776 ( .C (clk), .D (new_AGEMA_signal_15627), .Q (new_AGEMA_signal_15628) ) ;
    buf_clk new_AGEMA_reg_buffer_9779 ( .C (clk), .D (new_AGEMA_signal_15630), .Q (new_AGEMA_signal_15631) ) ;
    buf_clk new_AGEMA_reg_buffer_9782 ( .C (clk), .D (new_AGEMA_signal_15633), .Q (new_AGEMA_signal_15634) ) ;
    buf_clk new_AGEMA_reg_buffer_9785 ( .C (clk), .D (new_AGEMA_signal_15636), .Q (new_AGEMA_signal_15637) ) ;
    buf_clk new_AGEMA_reg_buffer_9788 ( .C (clk), .D (new_AGEMA_signal_15639), .Q (new_AGEMA_signal_15640) ) ;
    buf_clk new_AGEMA_reg_buffer_9791 ( .C (clk), .D (new_AGEMA_signal_15642), .Q (new_AGEMA_signal_15643) ) ;
    buf_clk new_AGEMA_reg_buffer_9794 ( .C (clk), .D (new_AGEMA_signal_15645), .Q (new_AGEMA_signal_15646) ) ;
    buf_clk new_AGEMA_reg_buffer_9797 ( .C (clk), .D (new_AGEMA_signal_15648), .Q (new_AGEMA_signal_15649) ) ;
    buf_clk new_AGEMA_reg_buffer_9800 ( .C (clk), .D (new_AGEMA_signal_15651), .Q (new_AGEMA_signal_15652) ) ;
    buf_clk new_AGEMA_reg_buffer_9803 ( .C (clk), .D (new_AGEMA_signal_15654), .Q (new_AGEMA_signal_15655) ) ;
    buf_clk new_AGEMA_reg_buffer_9806 ( .C (clk), .D (new_AGEMA_signal_15657), .Q (new_AGEMA_signal_15658) ) ;
    buf_clk new_AGEMA_reg_buffer_9809 ( .C (clk), .D (new_AGEMA_signal_15660), .Q (new_AGEMA_signal_15661) ) ;
    buf_clk new_AGEMA_reg_buffer_9812 ( .C (clk), .D (new_AGEMA_signal_15663), .Q (new_AGEMA_signal_15664) ) ;
    buf_clk new_AGEMA_reg_buffer_9815 ( .C (clk), .D (new_AGEMA_signal_15666), .Q (new_AGEMA_signal_15667) ) ;
    buf_clk new_AGEMA_reg_buffer_9818 ( .C (clk), .D (new_AGEMA_signal_15669), .Q (new_AGEMA_signal_15670) ) ;
    buf_clk new_AGEMA_reg_buffer_9821 ( .C (clk), .D (new_AGEMA_signal_15672), .Q (new_AGEMA_signal_15673) ) ;
    buf_clk new_AGEMA_reg_buffer_9824 ( .C (clk), .D (new_AGEMA_signal_15675), .Q (new_AGEMA_signal_15676) ) ;
    buf_clk new_AGEMA_reg_buffer_9827 ( .C (clk), .D (new_AGEMA_signal_15678), .Q (new_AGEMA_signal_15679) ) ;
    buf_clk new_AGEMA_reg_buffer_9830 ( .C (clk), .D (new_AGEMA_signal_15681), .Q (new_AGEMA_signal_15682) ) ;
    buf_clk new_AGEMA_reg_buffer_9833 ( .C (clk), .D (new_AGEMA_signal_15684), .Q (new_AGEMA_signal_15685) ) ;
    buf_clk new_AGEMA_reg_buffer_9836 ( .C (clk), .D (new_AGEMA_signal_15687), .Q (new_AGEMA_signal_15688) ) ;
    buf_clk new_AGEMA_reg_buffer_9839 ( .C (clk), .D (new_AGEMA_signal_15690), .Q (new_AGEMA_signal_15691) ) ;
    buf_clk new_AGEMA_reg_buffer_9842 ( .C (clk), .D (new_AGEMA_signal_15693), .Q (new_AGEMA_signal_15694) ) ;
    buf_clk new_AGEMA_reg_buffer_9845 ( .C (clk), .D (new_AGEMA_signal_15696), .Q (new_AGEMA_signal_15697) ) ;
    buf_clk new_AGEMA_reg_buffer_9848 ( .C (clk), .D (new_AGEMA_signal_15699), .Q (new_AGEMA_signal_15700) ) ;
    buf_clk new_AGEMA_reg_buffer_9851 ( .C (clk), .D (new_AGEMA_signal_15702), .Q (new_AGEMA_signal_15703) ) ;
    buf_clk new_AGEMA_reg_buffer_9854 ( .C (clk), .D (new_AGEMA_signal_15705), .Q (new_AGEMA_signal_15706) ) ;
    buf_clk new_AGEMA_reg_buffer_9857 ( .C (clk), .D (new_AGEMA_signal_15708), .Q (new_AGEMA_signal_15709) ) ;
    buf_clk new_AGEMA_reg_buffer_9860 ( .C (clk), .D (new_AGEMA_signal_15711), .Q (new_AGEMA_signal_15712) ) ;
    buf_clk new_AGEMA_reg_buffer_9863 ( .C (clk), .D (new_AGEMA_signal_15714), .Q (new_AGEMA_signal_15715) ) ;
    buf_clk new_AGEMA_reg_buffer_9866 ( .C (clk), .D (new_AGEMA_signal_15717), .Q (new_AGEMA_signal_15718) ) ;
    buf_clk new_AGEMA_reg_buffer_9869 ( .C (clk), .D (new_AGEMA_signal_15720), .Q (new_AGEMA_signal_15721) ) ;
    buf_clk new_AGEMA_reg_buffer_9872 ( .C (clk), .D (new_AGEMA_signal_15723), .Q (new_AGEMA_signal_15724) ) ;
    buf_clk new_AGEMA_reg_buffer_9875 ( .C (clk), .D (new_AGEMA_signal_15726), .Q (new_AGEMA_signal_15727) ) ;
    buf_clk new_AGEMA_reg_buffer_9878 ( .C (clk), .D (new_AGEMA_signal_15729), .Q (new_AGEMA_signal_15730) ) ;
    buf_clk new_AGEMA_reg_buffer_9881 ( .C (clk), .D (new_AGEMA_signal_15732), .Q (new_AGEMA_signal_15733) ) ;
    buf_clk new_AGEMA_reg_buffer_9884 ( .C (clk), .D (new_AGEMA_signal_15735), .Q (new_AGEMA_signal_15736) ) ;
    buf_clk new_AGEMA_reg_buffer_9887 ( .C (clk), .D (new_AGEMA_signal_15738), .Q (new_AGEMA_signal_15739) ) ;
    buf_clk new_AGEMA_reg_buffer_9890 ( .C (clk), .D (new_AGEMA_signal_15741), .Q (new_AGEMA_signal_15742) ) ;
    buf_clk new_AGEMA_reg_buffer_9893 ( .C (clk), .D (new_AGEMA_signal_15744), .Q (new_AGEMA_signal_15745) ) ;
    buf_clk new_AGEMA_reg_buffer_9896 ( .C (clk), .D (new_AGEMA_signal_15747), .Q (new_AGEMA_signal_15748) ) ;
    buf_clk new_AGEMA_reg_buffer_9899 ( .C (clk), .D (new_AGEMA_signal_15750), .Q (new_AGEMA_signal_15751) ) ;
    buf_clk new_AGEMA_reg_buffer_9902 ( .C (clk), .D (new_AGEMA_signal_15753), .Q (new_AGEMA_signal_15754) ) ;
    buf_clk new_AGEMA_reg_buffer_9905 ( .C (clk), .D (new_AGEMA_signal_15756), .Q (new_AGEMA_signal_15757) ) ;
    buf_clk new_AGEMA_reg_buffer_9908 ( .C (clk), .D (new_AGEMA_signal_15759), .Q (new_AGEMA_signal_15760) ) ;
    buf_clk new_AGEMA_reg_buffer_9911 ( .C (clk), .D (new_AGEMA_signal_15762), .Q (new_AGEMA_signal_15763) ) ;
    buf_clk new_AGEMA_reg_buffer_9914 ( .C (clk), .D (new_AGEMA_signal_15765), .Q (new_AGEMA_signal_15766) ) ;
    buf_clk new_AGEMA_reg_buffer_9917 ( .C (clk), .D (new_AGEMA_signal_15768), .Q (new_AGEMA_signal_15769) ) ;
    buf_clk new_AGEMA_reg_buffer_9920 ( .C (clk), .D (new_AGEMA_signal_15771), .Q (new_AGEMA_signal_15772) ) ;
    buf_clk new_AGEMA_reg_buffer_9923 ( .C (clk), .D (new_AGEMA_signal_15774), .Q (new_AGEMA_signal_15775) ) ;
    buf_clk new_AGEMA_reg_buffer_9926 ( .C (clk), .D (new_AGEMA_signal_15777), .Q (new_AGEMA_signal_15778) ) ;
    buf_clk new_AGEMA_reg_buffer_9929 ( .C (clk), .D (new_AGEMA_signal_15780), .Q (new_AGEMA_signal_15781) ) ;
    buf_clk new_AGEMA_reg_buffer_9932 ( .C (clk), .D (new_AGEMA_signal_15783), .Q (new_AGEMA_signal_15784) ) ;
    buf_clk new_AGEMA_reg_buffer_9935 ( .C (clk), .D (new_AGEMA_signal_15786), .Q (new_AGEMA_signal_15787) ) ;
    buf_clk new_AGEMA_reg_buffer_9938 ( .C (clk), .D (new_AGEMA_signal_15789), .Q (new_AGEMA_signal_15790) ) ;
    buf_clk new_AGEMA_reg_buffer_9941 ( .C (clk), .D (new_AGEMA_signal_15792), .Q (new_AGEMA_signal_15793) ) ;
    buf_clk new_AGEMA_reg_buffer_9944 ( .C (clk), .D (new_AGEMA_signal_15795), .Q (new_AGEMA_signal_15796) ) ;
    buf_clk new_AGEMA_reg_buffer_9947 ( .C (clk), .D (new_AGEMA_signal_15798), .Q (new_AGEMA_signal_15799) ) ;
    buf_clk new_AGEMA_reg_buffer_9950 ( .C (clk), .D (new_AGEMA_signal_15801), .Q (new_AGEMA_signal_15802) ) ;
    buf_clk new_AGEMA_reg_buffer_9953 ( .C (clk), .D (new_AGEMA_signal_15804), .Q (new_AGEMA_signal_15805) ) ;
    buf_clk new_AGEMA_reg_buffer_9956 ( .C (clk), .D (new_AGEMA_signal_15807), .Q (new_AGEMA_signal_15808) ) ;
    buf_clk new_AGEMA_reg_buffer_9959 ( .C (clk), .D (new_AGEMA_signal_15810), .Q (new_AGEMA_signal_15811) ) ;
    buf_clk new_AGEMA_reg_buffer_9962 ( .C (clk), .D (new_AGEMA_signal_15813), .Q (new_AGEMA_signal_15814) ) ;
    buf_clk new_AGEMA_reg_buffer_9966 ( .C (clk), .D (new_AGEMA_signal_15817), .Q (new_AGEMA_signal_15818) ) ;
    buf_clk new_AGEMA_reg_buffer_9970 ( .C (clk), .D (new_AGEMA_signal_15821), .Q (new_AGEMA_signal_15822) ) ;
    buf_clk new_AGEMA_reg_buffer_9974 ( .C (clk), .D (new_AGEMA_signal_15825), .Q (new_AGEMA_signal_15826) ) ;

    /* cells in depth 3 */
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M29_U1 ( .a ({new_AGEMA_signal_6015, SubBytesIns_Inst_Sbox_0_M28}), .b ({new_AGEMA_signal_10226, new_AGEMA_signal_10225}), .clk (clk), .r ({Fresh[481], Fresh[480]}), .c ({new_AGEMA_signal_6113, SubBytesIns_Inst_Sbox_0_M29}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M30_U1 ( .a ({new_AGEMA_signal_6014, SubBytesIns_Inst_Sbox_0_M26}), .b ({new_AGEMA_signal_10228, new_AGEMA_signal_10227}), .clk (clk), .r ({Fresh[483], Fresh[482]}), .c ({new_AGEMA_signal_6114, SubBytesIns_Inst_Sbox_0_M30}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M32_U1 ( .a ({new_AGEMA_signal_10226, new_AGEMA_signal_10225}), .b ({new_AGEMA_signal_6016, SubBytesIns_Inst_Sbox_0_M31}), .clk (clk), .r ({Fresh[485], Fresh[484]}), .c ({new_AGEMA_signal_6115, SubBytesIns_Inst_Sbox_0_M32}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M35_U1 ( .a ({new_AGEMA_signal_10228, new_AGEMA_signal_10227}), .b ({new_AGEMA_signal_5932, SubBytesIns_Inst_Sbox_0_M34}), .clk (clk), .r ({Fresh[487], Fresh[486]}), .c ({new_AGEMA_signal_6116, SubBytesIns_Inst_Sbox_0_M35}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M37_U1 ( .a ({new_AGEMA_signal_10382, new_AGEMA_signal_10381}), .b ({new_AGEMA_signal_6113, SubBytesIns_Inst_Sbox_0_M29}), .c ({new_AGEMA_signal_6209, SubBytesIns_Inst_Sbox_0_M37}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M38_U1 ( .a ({new_AGEMA_signal_6115, SubBytesIns_Inst_Sbox_0_M32}), .b ({new_AGEMA_signal_10384, new_AGEMA_signal_10383}), .c ({new_AGEMA_signal_6210, SubBytesIns_Inst_Sbox_0_M38}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M39_U1 ( .a ({new_AGEMA_signal_10386, new_AGEMA_signal_10385}), .b ({new_AGEMA_signal_6114, SubBytesIns_Inst_Sbox_0_M30}), .c ({new_AGEMA_signal_6211, SubBytesIns_Inst_Sbox_0_M39}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M40_U1 ( .a ({new_AGEMA_signal_6116, SubBytesIns_Inst_Sbox_0_M35}), .b ({new_AGEMA_signal_10388, new_AGEMA_signal_10387}), .c ({new_AGEMA_signal_6212, SubBytesIns_Inst_Sbox_0_M40}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M41_U1 ( .a ({new_AGEMA_signal_6210, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_6212, SubBytesIns_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_6321, SubBytesIns_Inst_Sbox_0_M41}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M42_U1 ( .a ({new_AGEMA_signal_6209, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_6211, SubBytesIns_Inst_Sbox_0_M39}), .c ({new_AGEMA_signal_6322, SubBytesIns_Inst_Sbox_0_M42}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M43_U1 ( .a ({new_AGEMA_signal_6209, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_6210, SubBytesIns_Inst_Sbox_0_M38}), .c ({new_AGEMA_signal_6323, SubBytesIns_Inst_Sbox_0_M43}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M44_U1 ( .a ({new_AGEMA_signal_6211, SubBytesIns_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_6212, SubBytesIns_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_6324, SubBytesIns_Inst_Sbox_0_M44}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M45_U1 ( .a ({new_AGEMA_signal_6322, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_6321, SubBytesIns_Inst_Sbox_0_M41}), .c ({new_AGEMA_signal_6561, SubBytesIns_Inst_Sbox_0_M45}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M29_U1 ( .a ({new_AGEMA_signal_6020, SubBytesIns_Inst_Sbox_1_M28}), .b ({new_AGEMA_signal_10234, new_AGEMA_signal_10233}), .clk (clk), .r ({Fresh[489], Fresh[488]}), .c ({new_AGEMA_signal_6118, SubBytesIns_Inst_Sbox_1_M29}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M30_U1 ( .a ({new_AGEMA_signal_6019, SubBytesIns_Inst_Sbox_1_M26}), .b ({new_AGEMA_signal_10236, new_AGEMA_signal_10235}), .clk (clk), .r ({Fresh[491], Fresh[490]}), .c ({new_AGEMA_signal_6119, SubBytesIns_Inst_Sbox_1_M30}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M32_U1 ( .a ({new_AGEMA_signal_10234, new_AGEMA_signal_10233}), .b ({new_AGEMA_signal_6021, SubBytesIns_Inst_Sbox_1_M31}), .clk (clk), .r ({Fresh[493], Fresh[492]}), .c ({new_AGEMA_signal_6120, SubBytesIns_Inst_Sbox_1_M32}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M35_U1 ( .a ({new_AGEMA_signal_10236, new_AGEMA_signal_10235}), .b ({new_AGEMA_signal_5936, SubBytesIns_Inst_Sbox_1_M34}), .clk (clk), .r ({Fresh[495], Fresh[494]}), .c ({new_AGEMA_signal_6121, SubBytesIns_Inst_Sbox_1_M35}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M37_U1 ( .a ({new_AGEMA_signal_10390, new_AGEMA_signal_10389}), .b ({new_AGEMA_signal_6118, SubBytesIns_Inst_Sbox_1_M29}), .c ({new_AGEMA_signal_6213, SubBytesIns_Inst_Sbox_1_M37}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M38_U1 ( .a ({new_AGEMA_signal_6120, SubBytesIns_Inst_Sbox_1_M32}), .b ({new_AGEMA_signal_10392, new_AGEMA_signal_10391}), .c ({new_AGEMA_signal_6214, SubBytesIns_Inst_Sbox_1_M38}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M39_U1 ( .a ({new_AGEMA_signal_10394, new_AGEMA_signal_10393}), .b ({new_AGEMA_signal_6119, SubBytesIns_Inst_Sbox_1_M30}), .c ({new_AGEMA_signal_6215, SubBytesIns_Inst_Sbox_1_M39}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M40_U1 ( .a ({new_AGEMA_signal_6121, SubBytesIns_Inst_Sbox_1_M35}), .b ({new_AGEMA_signal_10396, new_AGEMA_signal_10395}), .c ({new_AGEMA_signal_6216, SubBytesIns_Inst_Sbox_1_M40}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M41_U1 ( .a ({new_AGEMA_signal_6214, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_6216, SubBytesIns_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_6333, SubBytesIns_Inst_Sbox_1_M41}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M42_U1 ( .a ({new_AGEMA_signal_6213, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_6215, SubBytesIns_Inst_Sbox_1_M39}), .c ({new_AGEMA_signal_6334, SubBytesIns_Inst_Sbox_1_M42}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M43_U1 ( .a ({new_AGEMA_signal_6213, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_6214, SubBytesIns_Inst_Sbox_1_M38}), .c ({new_AGEMA_signal_6335, SubBytesIns_Inst_Sbox_1_M43}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M44_U1 ( .a ({new_AGEMA_signal_6215, SubBytesIns_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_6216, SubBytesIns_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_6336, SubBytesIns_Inst_Sbox_1_M44}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M45_U1 ( .a ({new_AGEMA_signal_6334, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_6333, SubBytesIns_Inst_Sbox_1_M41}), .c ({new_AGEMA_signal_6573, SubBytesIns_Inst_Sbox_1_M45}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M29_U1 ( .a ({new_AGEMA_signal_6025, SubBytesIns_Inst_Sbox_2_M28}), .b ({new_AGEMA_signal_10242, new_AGEMA_signal_10241}), .clk (clk), .r ({Fresh[497], Fresh[496]}), .c ({new_AGEMA_signal_6123, SubBytesIns_Inst_Sbox_2_M29}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M30_U1 ( .a ({new_AGEMA_signal_6024, SubBytesIns_Inst_Sbox_2_M26}), .b ({new_AGEMA_signal_10244, new_AGEMA_signal_10243}), .clk (clk), .r ({Fresh[499], Fresh[498]}), .c ({new_AGEMA_signal_6124, SubBytesIns_Inst_Sbox_2_M30}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M32_U1 ( .a ({new_AGEMA_signal_10242, new_AGEMA_signal_10241}), .b ({new_AGEMA_signal_6026, SubBytesIns_Inst_Sbox_2_M31}), .clk (clk), .r ({Fresh[501], Fresh[500]}), .c ({new_AGEMA_signal_6125, SubBytesIns_Inst_Sbox_2_M32}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M35_U1 ( .a ({new_AGEMA_signal_10244, new_AGEMA_signal_10243}), .b ({new_AGEMA_signal_5940, SubBytesIns_Inst_Sbox_2_M34}), .clk (clk), .r ({Fresh[503], Fresh[502]}), .c ({new_AGEMA_signal_6126, SubBytesIns_Inst_Sbox_2_M35}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M37_U1 ( .a ({new_AGEMA_signal_10398, new_AGEMA_signal_10397}), .b ({new_AGEMA_signal_6123, SubBytesIns_Inst_Sbox_2_M29}), .c ({new_AGEMA_signal_6217, SubBytesIns_Inst_Sbox_2_M37}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M38_U1 ( .a ({new_AGEMA_signal_6125, SubBytesIns_Inst_Sbox_2_M32}), .b ({new_AGEMA_signal_10400, new_AGEMA_signal_10399}), .c ({new_AGEMA_signal_6218, SubBytesIns_Inst_Sbox_2_M38}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M39_U1 ( .a ({new_AGEMA_signal_10402, new_AGEMA_signal_10401}), .b ({new_AGEMA_signal_6124, SubBytesIns_Inst_Sbox_2_M30}), .c ({new_AGEMA_signal_6219, SubBytesIns_Inst_Sbox_2_M39}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M40_U1 ( .a ({new_AGEMA_signal_6126, SubBytesIns_Inst_Sbox_2_M35}), .b ({new_AGEMA_signal_10404, new_AGEMA_signal_10403}), .c ({new_AGEMA_signal_6220, SubBytesIns_Inst_Sbox_2_M40}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M41_U1 ( .a ({new_AGEMA_signal_6218, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_6220, SubBytesIns_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_6345, SubBytesIns_Inst_Sbox_2_M41}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M42_U1 ( .a ({new_AGEMA_signal_6217, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_6219, SubBytesIns_Inst_Sbox_2_M39}), .c ({new_AGEMA_signal_6346, SubBytesIns_Inst_Sbox_2_M42}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M43_U1 ( .a ({new_AGEMA_signal_6217, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_6218, SubBytesIns_Inst_Sbox_2_M38}), .c ({new_AGEMA_signal_6347, SubBytesIns_Inst_Sbox_2_M43}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M44_U1 ( .a ({new_AGEMA_signal_6219, SubBytesIns_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_6220, SubBytesIns_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_6348, SubBytesIns_Inst_Sbox_2_M44}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M45_U1 ( .a ({new_AGEMA_signal_6346, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_6345, SubBytesIns_Inst_Sbox_2_M41}), .c ({new_AGEMA_signal_6585, SubBytesIns_Inst_Sbox_2_M45}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M29_U1 ( .a ({new_AGEMA_signal_6030, SubBytesIns_Inst_Sbox_3_M28}), .b ({new_AGEMA_signal_10250, new_AGEMA_signal_10249}), .clk (clk), .r ({Fresh[505], Fresh[504]}), .c ({new_AGEMA_signal_6128, SubBytesIns_Inst_Sbox_3_M29}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M30_U1 ( .a ({new_AGEMA_signal_6029, SubBytesIns_Inst_Sbox_3_M26}), .b ({new_AGEMA_signal_10252, new_AGEMA_signal_10251}), .clk (clk), .r ({Fresh[507], Fresh[506]}), .c ({new_AGEMA_signal_6129, SubBytesIns_Inst_Sbox_3_M30}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M32_U1 ( .a ({new_AGEMA_signal_10250, new_AGEMA_signal_10249}), .b ({new_AGEMA_signal_6031, SubBytesIns_Inst_Sbox_3_M31}), .clk (clk), .r ({Fresh[509], Fresh[508]}), .c ({new_AGEMA_signal_6130, SubBytesIns_Inst_Sbox_3_M32}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M35_U1 ( .a ({new_AGEMA_signal_10252, new_AGEMA_signal_10251}), .b ({new_AGEMA_signal_5944, SubBytesIns_Inst_Sbox_3_M34}), .clk (clk), .r ({Fresh[511], Fresh[510]}), .c ({new_AGEMA_signal_6131, SubBytesIns_Inst_Sbox_3_M35}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M37_U1 ( .a ({new_AGEMA_signal_10406, new_AGEMA_signal_10405}), .b ({new_AGEMA_signal_6128, SubBytesIns_Inst_Sbox_3_M29}), .c ({new_AGEMA_signal_6221, SubBytesIns_Inst_Sbox_3_M37}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M38_U1 ( .a ({new_AGEMA_signal_6130, SubBytesIns_Inst_Sbox_3_M32}), .b ({new_AGEMA_signal_10408, new_AGEMA_signal_10407}), .c ({new_AGEMA_signal_6222, SubBytesIns_Inst_Sbox_3_M38}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M39_U1 ( .a ({new_AGEMA_signal_10410, new_AGEMA_signal_10409}), .b ({new_AGEMA_signal_6129, SubBytesIns_Inst_Sbox_3_M30}), .c ({new_AGEMA_signal_6223, SubBytesIns_Inst_Sbox_3_M39}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M40_U1 ( .a ({new_AGEMA_signal_6131, SubBytesIns_Inst_Sbox_3_M35}), .b ({new_AGEMA_signal_10412, new_AGEMA_signal_10411}), .c ({new_AGEMA_signal_6224, SubBytesIns_Inst_Sbox_3_M40}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M41_U1 ( .a ({new_AGEMA_signal_6222, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_6224, SubBytesIns_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_6357, SubBytesIns_Inst_Sbox_3_M41}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M42_U1 ( .a ({new_AGEMA_signal_6221, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_6223, SubBytesIns_Inst_Sbox_3_M39}), .c ({new_AGEMA_signal_6358, SubBytesIns_Inst_Sbox_3_M42}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M43_U1 ( .a ({new_AGEMA_signal_6221, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_6222, SubBytesIns_Inst_Sbox_3_M38}), .c ({new_AGEMA_signal_6359, SubBytesIns_Inst_Sbox_3_M43}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M44_U1 ( .a ({new_AGEMA_signal_6223, SubBytesIns_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_6224, SubBytesIns_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_6360, SubBytesIns_Inst_Sbox_3_M44}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M45_U1 ( .a ({new_AGEMA_signal_6358, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_6357, SubBytesIns_Inst_Sbox_3_M41}), .c ({new_AGEMA_signal_6597, SubBytesIns_Inst_Sbox_3_M45}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M29_U1 ( .a ({new_AGEMA_signal_6035, SubBytesIns_Inst_Sbox_4_M28}), .b ({new_AGEMA_signal_10258, new_AGEMA_signal_10257}), .clk (clk), .r ({Fresh[513], Fresh[512]}), .c ({new_AGEMA_signal_6133, SubBytesIns_Inst_Sbox_4_M29}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M30_U1 ( .a ({new_AGEMA_signal_6034, SubBytesIns_Inst_Sbox_4_M26}), .b ({new_AGEMA_signal_10260, new_AGEMA_signal_10259}), .clk (clk), .r ({Fresh[515], Fresh[514]}), .c ({new_AGEMA_signal_6134, SubBytesIns_Inst_Sbox_4_M30}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M32_U1 ( .a ({new_AGEMA_signal_10258, new_AGEMA_signal_10257}), .b ({new_AGEMA_signal_6036, SubBytesIns_Inst_Sbox_4_M31}), .clk (clk), .r ({Fresh[517], Fresh[516]}), .c ({new_AGEMA_signal_6135, SubBytesIns_Inst_Sbox_4_M32}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M35_U1 ( .a ({new_AGEMA_signal_10260, new_AGEMA_signal_10259}), .b ({new_AGEMA_signal_5948, SubBytesIns_Inst_Sbox_4_M34}), .clk (clk), .r ({Fresh[519], Fresh[518]}), .c ({new_AGEMA_signal_6136, SubBytesIns_Inst_Sbox_4_M35}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M37_U1 ( .a ({new_AGEMA_signal_10414, new_AGEMA_signal_10413}), .b ({new_AGEMA_signal_6133, SubBytesIns_Inst_Sbox_4_M29}), .c ({new_AGEMA_signal_6225, SubBytesIns_Inst_Sbox_4_M37}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M38_U1 ( .a ({new_AGEMA_signal_6135, SubBytesIns_Inst_Sbox_4_M32}), .b ({new_AGEMA_signal_10416, new_AGEMA_signal_10415}), .c ({new_AGEMA_signal_6226, SubBytesIns_Inst_Sbox_4_M38}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M39_U1 ( .a ({new_AGEMA_signal_10418, new_AGEMA_signal_10417}), .b ({new_AGEMA_signal_6134, SubBytesIns_Inst_Sbox_4_M30}), .c ({new_AGEMA_signal_6227, SubBytesIns_Inst_Sbox_4_M39}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M40_U1 ( .a ({new_AGEMA_signal_6136, SubBytesIns_Inst_Sbox_4_M35}), .b ({new_AGEMA_signal_10420, new_AGEMA_signal_10419}), .c ({new_AGEMA_signal_6228, SubBytesIns_Inst_Sbox_4_M40}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M41_U1 ( .a ({new_AGEMA_signal_6226, SubBytesIns_Inst_Sbox_4_M38}), .b ({new_AGEMA_signal_6228, SubBytesIns_Inst_Sbox_4_M40}), .c ({new_AGEMA_signal_6369, SubBytesIns_Inst_Sbox_4_M41}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M42_U1 ( .a ({new_AGEMA_signal_6225, SubBytesIns_Inst_Sbox_4_M37}), .b ({new_AGEMA_signal_6227, SubBytesIns_Inst_Sbox_4_M39}), .c ({new_AGEMA_signal_6370, SubBytesIns_Inst_Sbox_4_M42}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M43_U1 ( .a ({new_AGEMA_signal_6225, SubBytesIns_Inst_Sbox_4_M37}), .b ({new_AGEMA_signal_6226, SubBytesIns_Inst_Sbox_4_M38}), .c ({new_AGEMA_signal_6371, SubBytesIns_Inst_Sbox_4_M43}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M44_U1 ( .a ({new_AGEMA_signal_6227, SubBytesIns_Inst_Sbox_4_M39}), .b ({new_AGEMA_signal_6228, SubBytesIns_Inst_Sbox_4_M40}), .c ({new_AGEMA_signal_6372, SubBytesIns_Inst_Sbox_4_M44}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M45_U1 ( .a ({new_AGEMA_signal_6370, SubBytesIns_Inst_Sbox_4_M42}), .b ({new_AGEMA_signal_6369, SubBytesIns_Inst_Sbox_4_M41}), .c ({new_AGEMA_signal_6609, SubBytesIns_Inst_Sbox_4_M45}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M29_U1 ( .a ({new_AGEMA_signal_6040, SubBytesIns_Inst_Sbox_5_M28}), .b ({new_AGEMA_signal_10266, new_AGEMA_signal_10265}), .clk (clk), .r ({Fresh[521], Fresh[520]}), .c ({new_AGEMA_signal_6138, SubBytesIns_Inst_Sbox_5_M29}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M30_U1 ( .a ({new_AGEMA_signal_6039, SubBytesIns_Inst_Sbox_5_M26}), .b ({new_AGEMA_signal_10268, new_AGEMA_signal_10267}), .clk (clk), .r ({Fresh[523], Fresh[522]}), .c ({new_AGEMA_signal_6139, SubBytesIns_Inst_Sbox_5_M30}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M32_U1 ( .a ({new_AGEMA_signal_10266, new_AGEMA_signal_10265}), .b ({new_AGEMA_signal_6041, SubBytesIns_Inst_Sbox_5_M31}), .clk (clk), .r ({Fresh[525], Fresh[524]}), .c ({new_AGEMA_signal_6140, SubBytesIns_Inst_Sbox_5_M32}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M35_U1 ( .a ({new_AGEMA_signal_10268, new_AGEMA_signal_10267}), .b ({new_AGEMA_signal_5952, SubBytesIns_Inst_Sbox_5_M34}), .clk (clk), .r ({Fresh[527], Fresh[526]}), .c ({new_AGEMA_signal_6141, SubBytesIns_Inst_Sbox_5_M35}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M37_U1 ( .a ({new_AGEMA_signal_10422, new_AGEMA_signal_10421}), .b ({new_AGEMA_signal_6138, SubBytesIns_Inst_Sbox_5_M29}), .c ({new_AGEMA_signal_6229, SubBytesIns_Inst_Sbox_5_M37}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M38_U1 ( .a ({new_AGEMA_signal_6140, SubBytesIns_Inst_Sbox_5_M32}), .b ({new_AGEMA_signal_10424, new_AGEMA_signal_10423}), .c ({new_AGEMA_signal_6230, SubBytesIns_Inst_Sbox_5_M38}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M39_U1 ( .a ({new_AGEMA_signal_10426, new_AGEMA_signal_10425}), .b ({new_AGEMA_signal_6139, SubBytesIns_Inst_Sbox_5_M30}), .c ({new_AGEMA_signal_6231, SubBytesIns_Inst_Sbox_5_M39}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M40_U1 ( .a ({new_AGEMA_signal_6141, SubBytesIns_Inst_Sbox_5_M35}), .b ({new_AGEMA_signal_10428, new_AGEMA_signal_10427}), .c ({new_AGEMA_signal_6232, SubBytesIns_Inst_Sbox_5_M40}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M41_U1 ( .a ({new_AGEMA_signal_6230, SubBytesIns_Inst_Sbox_5_M38}), .b ({new_AGEMA_signal_6232, SubBytesIns_Inst_Sbox_5_M40}), .c ({new_AGEMA_signal_6381, SubBytesIns_Inst_Sbox_5_M41}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M42_U1 ( .a ({new_AGEMA_signal_6229, SubBytesIns_Inst_Sbox_5_M37}), .b ({new_AGEMA_signal_6231, SubBytesIns_Inst_Sbox_5_M39}), .c ({new_AGEMA_signal_6382, SubBytesIns_Inst_Sbox_5_M42}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M43_U1 ( .a ({new_AGEMA_signal_6229, SubBytesIns_Inst_Sbox_5_M37}), .b ({new_AGEMA_signal_6230, SubBytesIns_Inst_Sbox_5_M38}), .c ({new_AGEMA_signal_6383, SubBytesIns_Inst_Sbox_5_M43}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M44_U1 ( .a ({new_AGEMA_signal_6231, SubBytesIns_Inst_Sbox_5_M39}), .b ({new_AGEMA_signal_6232, SubBytesIns_Inst_Sbox_5_M40}), .c ({new_AGEMA_signal_6384, SubBytesIns_Inst_Sbox_5_M44}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M45_U1 ( .a ({new_AGEMA_signal_6382, SubBytesIns_Inst_Sbox_5_M42}), .b ({new_AGEMA_signal_6381, SubBytesIns_Inst_Sbox_5_M41}), .c ({new_AGEMA_signal_6621, SubBytesIns_Inst_Sbox_5_M45}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M29_U1 ( .a ({new_AGEMA_signal_6045, SubBytesIns_Inst_Sbox_6_M28}), .b ({new_AGEMA_signal_10274, new_AGEMA_signal_10273}), .clk (clk), .r ({Fresh[529], Fresh[528]}), .c ({new_AGEMA_signal_6143, SubBytesIns_Inst_Sbox_6_M29}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M30_U1 ( .a ({new_AGEMA_signal_6044, SubBytesIns_Inst_Sbox_6_M26}), .b ({new_AGEMA_signal_10276, new_AGEMA_signal_10275}), .clk (clk), .r ({Fresh[531], Fresh[530]}), .c ({new_AGEMA_signal_6144, SubBytesIns_Inst_Sbox_6_M30}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M32_U1 ( .a ({new_AGEMA_signal_10274, new_AGEMA_signal_10273}), .b ({new_AGEMA_signal_6046, SubBytesIns_Inst_Sbox_6_M31}), .clk (clk), .r ({Fresh[533], Fresh[532]}), .c ({new_AGEMA_signal_6145, SubBytesIns_Inst_Sbox_6_M32}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M35_U1 ( .a ({new_AGEMA_signal_10276, new_AGEMA_signal_10275}), .b ({new_AGEMA_signal_5956, SubBytesIns_Inst_Sbox_6_M34}), .clk (clk), .r ({Fresh[535], Fresh[534]}), .c ({new_AGEMA_signal_6146, SubBytesIns_Inst_Sbox_6_M35}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M37_U1 ( .a ({new_AGEMA_signal_10430, new_AGEMA_signal_10429}), .b ({new_AGEMA_signal_6143, SubBytesIns_Inst_Sbox_6_M29}), .c ({new_AGEMA_signal_6233, SubBytesIns_Inst_Sbox_6_M37}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M38_U1 ( .a ({new_AGEMA_signal_6145, SubBytesIns_Inst_Sbox_6_M32}), .b ({new_AGEMA_signal_10432, new_AGEMA_signal_10431}), .c ({new_AGEMA_signal_6234, SubBytesIns_Inst_Sbox_6_M38}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M39_U1 ( .a ({new_AGEMA_signal_10434, new_AGEMA_signal_10433}), .b ({new_AGEMA_signal_6144, SubBytesIns_Inst_Sbox_6_M30}), .c ({new_AGEMA_signal_6235, SubBytesIns_Inst_Sbox_6_M39}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M40_U1 ( .a ({new_AGEMA_signal_6146, SubBytesIns_Inst_Sbox_6_M35}), .b ({new_AGEMA_signal_10436, new_AGEMA_signal_10435}), .c ({new_AGEMA_signal_6236, SubBytesIns_Inst_Sbox_6_M40}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M41_U1 ( .a ({new_AGEMA_signal_6234, SubBytesIns_Inst_Sbox_6_M38}), .b ({new_AGEMA_signal_6236, SubBytesIns_Inst_Sbox_6_M40}), .c ({new_AGEMA_signal_6393, SubBytesIns_Inst_Sbox_6_M41}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M42_U1 ( .a ({new_AGEMA_signal_6233, SubBytesIns_Inst_Sbox_6_M37}), .b ({new_AGEMA_signal_6235, SubBytesIns_Inst_Sbox_6_M39}), .c ({new_AGEMA_signal_6394, SubBytesIns_Inst_Sbox_6_M42}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M43_U1 ( .a ({new_AGEMA_signal_6233, SubBytesIns_Inst_Sbox_6_M37}), .b ({new_AGEMA_signal_6234, SubBytesIns_Inst_Sbox_6_M38}), .c ({new_AGEMA_signal_6395, SubBytesIns_Inst_Sbox_6_M43}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M44_U1 ( .a ({new_AGEMA_signal_6235, SubBytesIns_Inst_Sbox_6_M39}), .b ({new_AGEMA_signal_6236, SubBytesIns_Inst_Sbox_6_M40}), .c ({new_AGEMA_signal_6396, SubBytesIns_Inst_Sbox_6_M44}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M45_U1 ( .a ({new_AGEMA_signal_6394, SubBytesIns_Inst_Sbox_6_M42}), .b ({new_AGEMA_signal_6393, SubBytesIns_Inst_Sbox_6_M41}), .c ({new_AGEMA_signal_6633, SubBytesIns_Inst_Sbox_6_M45}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M29_U1 ( .a ({new_AGEMA_signal_6050, SubBytesIns_Inst_Sbox_7_M28}), .b ({new_AGEMA_signal_10282, new_AGEMA_signal_10281}), .clk (clk), .r ({Fresh[537], Fresh[536]}), .c ({new_AGEMA_signal_6148, SubBytesIns_Inst_Sbox_7_M29}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M30_U1 ( .a ({new_AGEMA_signal_6049, SubBytesIns_Inst_Sbox_7_M26}), .b ({new_AGEMA_signal_10284, new_AGEMA_signal_10283}), .clk (clk), .r ({Fresh[539], Fresh[538]}), .c ({new_AGEMA_signal_6149, SubBytesIns_Inst_Sbox_7_M30}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M32_U1 ( .a ({new_AGEMA_signal_10282, new_AGEMA_signal_10281}), .b ({new_AGEMA_signal_6051, SubBytesIns_Inst_Sbox_7_M31}), .clk (clk), .r ({Fresh[541], Fresh[540]}), .c ({new_AGEMA_signal_6150, SubBytesIns_Inst_Sbox_7_M32}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M35_U1 ( .a ({new_AGEMA_signal_10284, new_AGEMA_signal_10283}), .b ({new_AGEMA_signal_5960, SubBytesIns_Inst_Sbox_7_M34}), .clk (clk), .r ({Fresh[543], Fresh[542]}), .c ({new_AGEMA_signal_6151, SubBytesIns_Inst_Sbox_7_M35}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M37_U1 ( .a ({new_AGEMA_signal_10438, new_AGEMA_signal_10437}), .b ({new_AGEMA_signal_6148, SubBytesIns_Inst_Sbox_7_M29}), .c ({new_AGEMA_signal_6237, SubBytesIns_Inst_Sbox_7_M37}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M38_U1 ( .a ({new_AGEMA_signal_6150, SubBytesIns_Inst_Sbox_7_M32}), .b ({new_AGEMA_signal_10440, new_AGEMA_signal_10439}), .c ({new_AGEMA_signal_6238, SubBytesIns_Inst_Sbox_7_M38}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M39_U1 ( .a ({new_AGEMA_signal_10442, new_AGEMA_signal_10441}), .b ({new_AGEMA_signal_6149, SubBytesIns_Inst_Sbox_7_M30}), .c ({new_AGEMA_signal_6239, SubBytesIns_Inst_Sbox_7_M39}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M40_U1 ( .a ({new_AGEMA_signal_6151, SubBytesIns_Inst_Sbox_7_M35}), .b ({new_AGEMA_signal_10444, new_AGEMA_signal_10443}), .c ({new_AGEMA_signal_6240, SubBytesIns_Inst_Sbox_7_M40}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M41_U1 ( .a ({new_AGEMA_signal_6238, SubBytesIns_Inst_Sbox_7_M38}), .b ({new_AGEMA_signal_6240, SubBytesIns_Inst_Sbox_7_M40}), .c ({new_AGEMA_signal_6405, SubBytesIns_Inst_Sbox_7_M41}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M42_U1 ( .a ({new_AGEMA_signal_6237, SubBytesIns_Inst_Sbox_7_M37}), .b ({new_AGEMA_signal_6239, SubBytesIns_Inst_Sbox_7_M39}), .c ({new_AGEMA_signal_6406, SubBytesIns_Inst_Sbox_7_M42}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M43_U1 ( .a ({new_AGEMA_signal_6237, SubBytesIns_Inst_Sbox_7_M37}), .b ({new_AGEMA_signal_6238, SubBytesIns_Inst_Sbox_7_M38}), .c ({new_AGEMA_signal_6407, SubBytesIns_Inst_Sbox_7_M43}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M44_U1 ( .a ({new_AGEMA_signal_6239, SubBytesIns_Inst_Sbox_7_M39}), .b ({new_AGEMA_signal_6240, SubBytesIns_Inst_Sbox_7_M40}), .c ({new_AGEMA_signal_6408, SubBytesIns_Inst_Sbox_7_M44}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M45_U1 ( .a ({new_AGEMA_signal_6406, SubBytesIns_Inst_Sbox_7_M42}), .b ({new_AGEMA_signal_6405, SubBytesIns_Inst_Sbox_7_M41}), .c ({new_AGEMA_signal_6645, SubBytesIns_Inst_Sbox_7_M45}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M29_U1 ( .a ({new_AGEMA_signal_6055, SubBytesIns_Inst_Sbox_8_M28}), .b ({new_AGEMA_signal_10290, new_AGEMA_signal_10289}), .clk (clk), .r ({Fresh[545], Fresh[544]}), .c ({new_AGEMA_signal_6153, SubBytesIns_Inst_Sbox_8_M29}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M30_U1 ( .a ({new_AGEMA_signal_6054, SubBytesIns_Inst_Sbox_8_M26}), .b ({new_AGEMA_signal_10292, new_AGEMA_signal_10291}), .clk (clk), .r ({Fresh[547], Fresh[546]}), .c ({new_AGEMA_signal_6154, SubBytesIns_Inst_Sbox_8_M30}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M32_U1 ( .a ({new_AGEMA_signal_10290, new_AGEMA_signal_10289}), .b ({new_AGEMA_signal_6056, SubBytesIns_Inst_Sbox_8_M31}), .clk (clk), .r ({Fresh[549], Fresh[548]}), .c ({new_AGEMA_signal_6155, SubBytesIns_Inst_Sbox_8_M32}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M35_U1 ( .a ({new_AGEMA_signal_10292, new_AGEMA_signal_10291}), .b ({new_AGEMA_signal_5964, SubBytesIns_Inst_Sbox_8_M34}), .clk (clk), .r ({Fresh[551], Fresh[550]}), .c ({new_AGEMA_signal_6156, SubBytesIns_Inst_Sbox_8_M35}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M37_U1 ( .a ({new_AGEMA_signal_10446, new_AGEMA_signal_10445}), .b ({new_AGEMA_signal_6153, SubBytesIns_Inst_Sbox_8_M29}), .c ({new_AGEMA_signal_6241, SubBytesIns_Inst_Sbox_8_M37}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M38_U1 ( .a ({new_AGEMA_signal_6155, SubBytesIns_Inst_Sbox_8_M32}), .b ({new_AGEMA_signal_10448, new_AGEMA_signal_10447}), .c ({new_AGEMA_signal_6242, SubBytesIns_Inst_Sbox_8_M38}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M39_U1 ( .a ({new_AGEMA_signal_10450, new_AGEMA_signal_10449}), .b ({new_AGEMA_signal_6154, SubBytesIns_Inst_Sbox_8_M30}), .c ({new_AGEMA_signal_6243, SubBytesIns_Inst_Sbox_8_M39}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M40_U1 ( .a ({new_AGEMA_signal_6156, SubBytesIns_Inst_Sbox_8_M35}), .b ({new_AGEMA_signal_10452, new_AGEMA_signal_10451}), .c ({new_AGEMA_signal_6244, SubBytesIns_Inst_Sbox_8_M40}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M41_U1 ( .a ({new_AGEMA_signal_6242, SubBytesIns_Inst_Sbox_8_M38}), .b ({new_AGEMA_signal_6244, SubBytesIns_Inst_Sbox_8_M40}), .c ({new_AGEMA_signal_6417, SubBytesIns_Inst_Sbox_8_M41}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M42_U1 ( .a ({new_AGEMA_signal_6241, SubBytesIns_Inst_Sbox_8_M37}), .b ({new_AGEMA_signal_6243, SubBytesIns_Inst_Sbox_8_M39}), .c ({new_AGEMA_signal_6418, SubBytesIns_Inst_Sbox_8_M42}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M43_U1 ( .a ({new_AGEMA_signal_6241, SubBytesIns_Inst_Sbox_8_M37}), .b ({new_AGEMA_signal_6242, SubBytesIns_Inst_Sbox_8_M38}), .c ({new_AGEMA_signal_6419, SubBytesIns_Inst_Sbox_8_M43}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M44_U1 ( .a ({new_AGEMA_signal_6243, SubBytesIns_Inst_Sbox_8_M39}), .b ({new_AGEMA_signal_6244, SubBytesIns_Inst_Sbox_8_M40}), .c ({new_AGEMA_signal_6420, SubBytesIns_Inst_Sbox_8_M44}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M45_U1 ( .a ({new_AGEMA_signal_6418, SubBytesIns_Inst_Sbox_8_M42}), .b ({new_AGEMA_signal_6417, SubBytesIns_Inst_Sbox_8_M41}), .c ({new_AGEMA_signal_6657, SubBytesIns_Inst_Sbox_8_M45}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M29_U1 ( .a ({new_AGEMA_signal_6060, SubBytesIns_Inst_Sbox_9_M28}), .b ({new_AGEMA_signal_10298, new_AGEMA_signal_10297}), .clk (clk), .r ({Fresh[553], Fresh[552]}), .c ({new_AGEMA_signal_6158, SubBytesIns_Inst_Sbox_9_M29}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M30_U1 ( .a ({new_AGEMA_signal_6059, SubBytesIns_Inst_Sbox_9_M26}), .b ({new_AGEMA_signal_10300, new_AGEMA_signal_10299}), .clk (clk), .r ({Fresh[555], Fresh[554]}), .c ({new_AGEMA_signal_6159, SubBytesIns_Inst_Sbox_9_M30}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M32_U1 ( .a ({new_AGEMA_signal_10298, new_AGEMA_signal_10297}), .b ({new_AGEMA_signal_6061, SubBytesIns_Inst_Sbox_9_M31}), .clk (clk), .r ({Fresh[557], Fresh[556]}), .c ({new_AGEMA_signal_6160, SubBytesIns_Inst_Sbox_9_M32}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M35_U1 ( .a ({new_AGEMA_signal_10300, new_AGEMA_signal_10299}), .b ({new_AGEMA_signal_5968, SubBytesIns_Inst_Sbox_9_M34}), .clk (clk), .r ({Fresh[559], Fresh[558]}), .c ({new_AGEMA_signal_6161, SubBytesIns_Inst_Sbox_9_M35}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M37_U1 ( .a ({new_AGEMA_signal_10454, new_AGEMA_signal_10453}), .b ({new_AGEMA_signal_6158, SubBytesIns_Inst_Sbox_9_M29}), .c ({new_AGEMA_signal_6245, SubBytesIns_Inst_Sbox_9_M37}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M38_U1 ( .a ({new_AGEMA_signal_6160, SubBytesIns_Inst_Sbox_9_M32}), .b ({new_AGEMA_signal_10456, new_AGEMA_signal_10455}), .c ({new_AGEMA_signal_6246, SubBytesIns_Inst_Sbox_9_M38}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M39_U1 ( .a ({new_AGEMA_signal_10458, new_AGEMA_signal_10457}), .b ({new_AGEMA_signal_6159, SubBytesIns_Inst_Sbox_9_M30}), .c ({new_AGEMA_signal_6247, SubBytesIns_Inst_Sbox_9_M39}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M40_U1 ( .a ({new_AGEMA_signal_6161, SubBytesIns_Inst_Sbox_9_M35}), .b ({new_AGEMA_signal_10460, new_AGEMA_signal_10459}), .c ({new_AGEMA_signal_6248, SubBytesIns_Inst_Sbox_9_M40}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M41_U1 ( .a ({new_AGEMA_signal_6246, SubBytesIns_Inst_Sbox_9_M38}), .b ({new_AGEMA_signal_6248, SubBytesIns_Inst_Sbox_9_M40}), .c ({new_AGEMA_signal_6429, SubBytesIns_Inst_Sbox_9_M41}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M42_U1 ( .a ({new_AGEMA_signal_6245, SubBytesIns_Inst_Sbox_9_M37}), .b ({new_AGEMA_signal_6247, SubBytesIns_Inst_Sbox_9_M39}), .c ({new_AGEMA_signal_6430, SubBytesIns_Inst_Sbox_9_M42}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M43_U1 ( .a ({new_AGEMA_signal_6245, SubBytesIns_Inst_Sbox_9_M37}), .b ({new_AGEMA_signal_6246, SubBytesIns_Inst_Sbox_9_M38}), .c ({new_AGEMA_signal_6431, SubBytesIns_Inst_Sbox_9_M43}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M44_U1 ( .a ({new_AGEMA_signal_6247, SubBytesIns_Inst_Sbox_9_M39}), .b ({new_AGEMA_signal_6248, SubBytesIns_Inst_Sbox_9_M40}), .c ({new_AGEMA_signal_6432, SubBytesIns_Inst_Sbox_9_M44}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M45_U1 ( .a ({new_AGEMA_signal_6430, SubBytesIns_Inst_Sbox_9_M42}), .b ({new_AGEMA_signal_6429, SubBytesIns_Inst_Sbox_9_M41}), .c ({new_AGEMA_signal_6669, SubBytesIns_Inst_Sbox_9_M45}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M29_U1 ( .a ({new_AGEMA_signal_6065, SubBytesIns_Inst_Sbox_10_M28}), .b ({new_AGEMA_signal_10306, new_AGEMA_signal_10305}), .clk (clk), .r ({Fresh[561], Fresh[560]}), .c ({new_AGEMA_signal_6163, SubBytesIns_Inst_Sbox_10_M29}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M30_U1 ( .a ({new_AGEMA_signal_6064, SubBytesIns_Inst_Sbox_10_M26}), .b ({new_AGEMA_signal_10308, new_AGEMA_signal_10307}), .clk (clk), .r ({Fresh[563], Fresh[562]}), .c ({new_AGEMA_signal_6164, SubBytesIns_Inst_Sbox_10_M30}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M32_U1 ( .a ({new_AGEMA_signal_10306, new_AGEMA_signal_10305}), .b ({new_AGEMA_signal_6066, SubBytesIns_Inst_Sbox_10_M31}), .clk (clk), .r ({Fresh[565], Fresh[564]}), .c ({new_AGEMA_signal_6165, SubBytesIns_Inst_Sbox_10_M32}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M35_U1 ( .a ({new_AGEMA_signal_10308, new_AGEMA_signal_10307}), .b ({new_AGEMA_signal_5972, SubBytesIns_Inst_Sbox_10_M34}), .clk (clk), .r ({Fresh[567], Fresh[566]}), .c ({new_AGEMA_signal_6166, SubBytesIns_Inst_Sbox_10_M35}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M37_U1 ( .a ({new_AGEMA_signal_10462, new_AGEMA_signal_10461}), .b ({new_AGEMA_signal_6163, SubBytesIns_Inst_Sbox_10_M29}), .c ({new_AGEMA_signal_6249, SubBytesIns_Inst_Sbox_10_M37}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M38_U1 ( .a ({new_AGEMA_signal_6165, SubBytesIns_Inst_Sbox_10_M32}), .b ({new_AGEMA_signal_10464, new_AGEMA_signal_10463}), .c ({new_AGEMA_signal_6250, SubBytesIns_Inst_Sbox_10_M38}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M39_U1 ( .a ({new_AGEMA_signal_10466, new_AGEMA_signal_10465}), .b ({new_AGEMA_signal_6164, SubBytesIns_Inst_Sbox_10_M30}), .c ({new_AGEMA_signal_6251, SubBytesIns_Inst_Sbox_10_M39}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M40_U1 ( .a ({new_AGEMA_signal_6166, SubBytesIns_Inst_Sbox_10_M35}), .b ({new_AGEMA_signal_10468, new_AGEMA_signal_10467}), .c ({new_AGEMA_signal_6252, SubBytesIns_Inst_Sbox_10_M40}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M41_U1 ( .a ({new_AGEMA_signal_6250, SubBytesIns_Inst_Sbox_10_M38}), .b ({new_AGEMA_signal_6252, SubBytesIns_Inst_Sbox_10_M40}), .c ({new_AGEMA_signal_6441, SubBytesIns_Inst_Sbox_10_M41}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M42_U1 ( .a ({new_AGEMA_signal_6249, SubBytesIns_Inst_Sbox_10_M37}), .b ({new_AGEMA_signal_6251, SubBytesIns_Inst_Sbox_10_M39}), .c ({new_AGEMA_signal_6442, SubBytesIns_Inst_Sbox_10_M42}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M43_U1 ( .a ({new_AGEMA_signal_6249, SubBytesIns_Inst_Sbox_10_M37}), .b ({new_AGEMA_signal_6250, SubBytesIns_Inst_Sbox_10_M38}), .c ({new_AGEMA_signal_6443, SubBytesIns_Inst_Sbox_10_M43}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M44_U1 ( .a ({new_AGEMA_signal_6251, SubBytesIns_Inst_Sbox_10_M39}), .b ({new_AGEMA_signal_6252, SubBytesIns_Inst_Sbox_10_M40}), .c ({new_AGEMA_signal_6444, SubBytesIns_Inst_Sbox_10_M44}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M45_U1 ( .a ({new_AGEMA_signal_6442, SubBytesIns_Inst_Sbox_10_M42}), .b ({new_AGEMA_signal_6441, SubBytesIns_Inst_Sbox_10_M41}), .c ({new_AGEMA_signal_6681, SubBytesIns_Inst_Sbox_10_M45}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M29_U1 ( .a ({new_AGEMA_signal_6070, SubBytesIns_Inst_Sbox_11_M28}), .b ({new_AGEMA_signal_10314, new_AGEMA_signal_10313}), .clk (clk), .r ({Fresh[569], Fresh[568]}), .c ({new_AGEMA_signal_6168, SubBytesIns_Inst_Sbox_11_M29}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M30_U1 ( .a ({new_AGEMA_signal_6069, SubBytesIns_Inst_Sbox_11_M26}), .b ({new_AGEMA_signal_10316, new_AGEMA_signal_10315}), .clk (clk), .r ({Fresh[571], Fresh[570]}), .c ({new_AGEMA_signal_6169, SubBytesIns_Inst_Sbox_11_M30}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M32_U1 ( .a ({new_AGEMA_signal_10314, new_AGEMA_signal_10313}), .b ({new_AGEMA_signal_6071, SubBytesIns_Inst_Sbox_11_M31}), .clk (clk), .r ({Fresh[573], Fresh[572]}), .c ({new_AGEMA_signal_6170, SubBytesIns_Inst_Sbox_11_M32}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M35_U1 ( .a ({new_AGEMA_signal_10316, new_AGEMA_signal_10315}), .b ({new_AGEMA_signal_5976, SubBytesIns_Inst_Sbox_11_M34}), .clk (clk), .r ({Fresh[575], Fresh[574]}), .c ({new_AGEMA_signal_6171, SubBytesIns_Inst_Sbox_11_M35}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M37_U1 ( .a ({new_AGEMA_signal_10470, new_AGEMA_signal_10469}), .b ({new_AGEMA_signal_6168, SubBytesIns_Inst_Sbox_11_M29}), .c ({new_AGEMA_signal_6253, SubBytesIns_Inst_Sbox_11_M37}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M38_U1 ( .a ({new_AGEMA_signal_6170, SubBytesIns_Inst_Sbox_11_M32}), .b ({new_AGEMA_signal_10472, new_AGEMA_signal_10471}), .c ({new_AGEMA_signal_6254, SubBytesIns_Inst_Sbox_11_M38}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M39_U1 ( .a ({new_AGEMA_signal_10474, new_AGEMA_signal_10473}), .b ({new_AGEMA_signal_6169, SubBytesIns_Inst_Sbox_11_M30}), .c ({new_AGEMA_signal_6255, SubBytesIns_Inst_Sbox_11_M39}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M40_U1 ( .a ({new_AGEMA_signal_6171, SubBytesIns_Inst_Sbox_11_M35}), .b ({new_AGEMA_signal_10476, new_AGEMA_signal_10475}), .c ({new_AGEMA_signal_6256, SubBytesIns_Inst_Sbox_11_M40}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M41_U1 ( .a ({new_AGEMA_signal_6254, SubBytesIns_Inst_Sbox_11_M38}), .b ({new_AGEMA_signal_6256, SubBytesIns_Inst_Sbox_11_M40}), .c ({new_AGEMA_signal_6453, SubBytesIns_Inst_Sbox_11_M41}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M42_U1 ( .a ({new_AGEMA_signal_6253, SubBytesIns_Inst_Sbox_11_M37}), .b ({new_AGEMA_signal_6255, SubBytesIns_Inst_Sbox_11_M39}), .c ({new_AGEMA_signal_6454, SubBytesIns_Inst_Sbox_11_M42}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M43_U1 ( .a ({new_AGEMA_signal_6253, SubBytesIns_Inst_Sbox_11_M37}), .b ({new_AGEMA_signal_6254, SubBytesIns_Inst_Sbox_11_M38}), .c ({new_AGEMA_signal_6455, SubBytesIns_Inst_Sbox_11_M43}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M44_U1 ( .a ({new_AGEMA_signal_6255, SubBytesIns_Inst_Sbox_11_M39}), .b ({new_AGEMA_signal_6256, SubBytesIns_Inst_Sbox_11_M40}), .c ({new_AGEMA_signal_6456, SubBytesIns_Inst_Sbox_11_M44}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M45_U1 ( .a ({new_AGEMA_signal_6454, SubBytesIns_Inst_Sbox_11_M42}), .b ({new_AGEMA_signal_6453, SubBytesIns_Inst_Sbox_11_M41}), .c ({new_AGEMA_signal_6693, SubBytesIns_Inst_Sbox_11_M45}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M29_U1 ( .a ({new_AGEMA_signal_6075, SubBytesIns_Inst_Sbox_12_M28}), .b ({new_AGEMA_signal_10322, new_AGEMA_signal_10321}), .clk (clk), .r ({Fresh[577], Fresh[576]}), .c ({new_AGEMA_signal_6173, SubBytesIns_Inst_Sbox_12_M29}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M30_U1 ( .a ({new_AGEMA_signal_6074, SubBytesIns_Inst_Sbox_12_M26}), .b ({new_AGEMA_signal_10324, new_AGEMA_signal_10323}), .clk (clk), .r ({Fresh[579], Fresh[578]}), .c ({new_AGEMA_signal_6174, SubBytesIns_Inst_Sbox_12_M30}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M32_U1 ( .a ({new_AGEMA_signal_10322, new_AGEMA_signal_10321}), .b ({new_AGEMA_signal_6076, SubBytesIns_Inst_Sbox_12_M31}), .clk (clk), .r ({Fresh[581], Fresh[580]}), .c ({new_AGEMA_signal_6175, SubBytesIns_Inst_Sbox_12_M32}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M35_U1 ( .a ({new_AGEMA_signal_10324, new_AGEMA_signal_10323}), .b ({new_AGEMA_signal_5980, SubBytesIns_Inst_Sbox_12_M34}), .clk (clk), .r ({Fresh[583], Fresh[582]}), .c ({new_AGEMA_signal_6176, SubBytesIns_Inst_Sbox_12_M35}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M37_U1 ( .a ({new_AGEMA_signal_10478, new_AGEMA_signal_10477}), .b ({new_AGEMA_signal_6173, SubBytesIns_Inst_Sbox_12_M29}), .c ({new_AGEMA_signal_6257, SubBytesIns_Inst_Sbox_12_M37}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M38_U1 ( .a ({new_AGEMA_signal_6175, SubBytesIns_Inst_Sbox_12_M32}), .b ({new_AGEMA_signal_10480, new_AGEMA_signal_10479}), .c ({new_AGEMA_signal_6258, SubBytesIns_Inst_Sbox_12_M38}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M39_U1 ( .a ({new_AGEMA_signal_10482, new_AGEMA_signal_10481}), .b ({new_AGEMA_signal_6174, SubBytesIns_Inst_Sbox_12_M30}), .c ({new_AGEMA_signal_6259, SubBytesIns_Inst_Sbox_12_M39}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M40_U1 ( .a ({new_AGEMA_signal_6176, SubBytesIns_Inst_Sbox_12_M35}), .b ({new_AGEMA_signal_10484, new_AGEMA_signal_10483}), .c ({new_AGEMA_signal_6260, SubBytesIns_Inst_Sbox_12_M40}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M41_U1 ( .a ({new_AGEMA_signal_6258, SubBytesIns_Inst_Sbox_12_M38}), .b ({new_AGEMA_signal_6260, SubBytesIns_Inst_Sbox_12_M40}), .c ({new_AGEMA_signal_6465, SubBytesIns_Inst_Sbox_12_M41}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M42_U1 ( .a ({new_AGEMA_signal_6257, SubBytesIns_Inst_Sbox_12_M37}), .b ({new_AGEMA_signal_6259, SubBytesIns_Inst_Sbox_12_M39}), .c ({new_AGEMA_signal_6466, SubBytesIns_Inst_Sbox_12_M42}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M43_U1 ( .a ({new_AGEMA_signal_6257, SubBytesIns_Inst_Sbox_12_M37}), .b ({new_AGEMA_signal_6258, SubBytesIns_Inst_Sbox_12_M38}), .c ({new_AGEMA_signal_6467, SubBytesIns_Inst_Sbox_12_M43}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M44_U1 ( .a ({new_AGEMA_signal_6259, SubBytesIns_Inst_Sbox_12_M39}), .b ({new_AGEMA_signal_6260, SubBytesIns_Inst_Sbox_12_M40}), .c ({new_AGEMA_signal_6468, SubBytesIns_Inst_Sbox_12_M44}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M45_U1 ( .a ({new_AGEMA_signal_6466, SubBytesIns_Inst_Sbox_12_M42}), .b ({new_AGEMA_signal_6465, SubBytesIns_Inst_Sbox_12_M41}), .c ({new_AGEMA_signal_6705, SubBytesIns_Inst_Sbox_12_M45}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M29_U1 ( .a ({new_AGEMA_signal_6080, SubBytesIns_Inst_Sbox_13_M28}), .b ({new_AGEMA_signal_10330, new_AGEMA_signal_10329}), .clk (clk), .r ({Fresh[585], Fresh[584]}), .c ({new_AGEMA_signal_6178, SubBytesIns_Inst_Sbox_13_M29}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M30_U1 ( .a ({new_AGEMA_signal_6079, SubBytesIns_Inst_Sbox_13_M26}), .b ({new_AGEMA_signal_10332, new_AGEMA_signal_10331}), .clk (clk), .r ({Fresh[587], Fresh[586]}), .c ({new_AGEMA_signal_6179, SubBytesIns_Inst_Sbox_13_M30}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M32_U1 ( .a ({new_AGEMA_signal_10330, new_AGEMA_signal_10329}), .b ({new_AGEMA_signal_6081, SubBytesIns_Inst_Sbox_13_M31}), .clk (clk), .r ({Fresh[589], Fresh[588]}), .c ({new_AGEMA_signal_6180, SubBytesIns_Inst_Sbox_13_M32}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M35_U1 ( .a ({new_AGEMA_signal_10332, new_AGEMA_signal_10331}), .b ({new_AGEMA_signal_5984, SubBytesIns_Inst_Sbox_13_M34}), .clk (clk), .r ({Fresh[591], Fresh[590]}), .c ({new_AGEMA_signal_6181, SubBytesIns_Inst_Sbox_13_M35}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M37_U1 ( .a ({new_AGEMA_signal_10486, new_AGEMA_signal_10485}), .b ({new_AGEMA_signal_6178, SubBytesIns_Inst_Sbox_13_M29}), .c ({new_AGEMA_signal_6261, SubBytesIns_Inst_Sbox_13_M37}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M38_U1 ( .a ({new_AGEMA_signal_6180, SubBytesIns_Inst_Sbox_13_M32}), .b ({new_AGEMA_signal_10488, new_AGEMA_signal_10487}), .c ({new_AGEMA_signal_6262, SubBytesIns_Inst_Sbox_13_M38}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M39_U1 ( .a ({new_AGEMA_signal_10490, new_AGEMA_signal_10489}), .b ({new_AGEMA_signal_6179, SubBytesIns_Inst_Sbox_13_M30}), .c ({new_AGEMA_signal_6263, SubBytesIns_Inst_Sbox_13_M39}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M40_U1 ( .a ({new_AGEMA_signal_6181, SubBytesIns_Inst_Sbox_13_M35}), .b ({new_AGEMA_signal_10492, new_AGEMA_signal_10491}), .c ({new_AGEMA_signal_6264, SubBytesIns_Inst_Sbox_13_M40}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M41_U1 ( .a ({new_AGEMA_signal_6262, SubBytesIns_Inst_Sbox_13_M38}), .b ({new_AGEMA_signal_6264, SubBytesIns_Inst_Sbox_13_M40}), .c ({new_AGEMA_signal_6477, SubBytesIns_Inst_Sbox_13_M41}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M42_U1 ( .a ({new_AGEMA_signal_6261, SubBytesIns_Inst_Sbox_13_M37}), .b ({new_AGEMA_signal_6263, SubBytesIns_Inst_Sbox_13_M39}), .c ({new_AGEMA_signal_6478, SubBytesIns_Inst_Sbox_13_M42}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M43_U1 ( .a ({new_AGEMA_signal_6261, SubBytesIns_Inst_Sbox_13_M37}), .b ({new_AGEMA_signal_6262, SubBytesIns_Inst_Sbox_13_M38}), .c ({new_AGEMA_signal_6479, SubBytesIns_Inst_Sbox_13_M43}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M44_U1 ( .a ({new_AGEMA_signal_6263, SubBytesIns_Inst_Sbox_13_M39}), .b ({new_AGEMA_signal_6264, SubBytesIns_Inst_Sbox_13_M40}), .c ({new_AGEMA_signal_6480, SubBytesIns_Inst_Sbox_13_M44}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M45_U1 ( .a ({new_AGEMA_signal_6478, SubBytesIns_Inst_Sbox_13_M42}), .b ({new_AGEMA_signal_6477, SubBytesIns_Inst_Sbox_13_M41}), .c ({new_AGEMA_signal_6717, SubBytesIns_Inst_Sbox_13_M45}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M29_U1 ( .a ({new_AGEMA_signal_6085, SubBytesIns_Inst_Sbox_14_M28}), .b ({new_AGEMA_signal_10338, new_AGEMA_signal_10337}), .clk (clk), .r ({Fresh[593], Fresh[592]}), .c ({new_AGEMA_signal_6183, SubBytesIns_Inst_Sbox_14_M29}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M30_U1 ( .a ({new_AGEMA_signal_6084, SubBytesIns_Inst_Sbox_14_M26}), .b ({new_AGEMA_signal_10340, new_AGEMA_signal_10339}), .clk (clk), .r ({Fresh[595], Fresh[594]}), .c ({new_AGEMA_signal_6184, SubBytesIns_Inst_Sbox_14_M30}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M32_U1 ( .a ({new_AGEMA_signal_10338, new_AGEMA_signal_10337}), .b ({new_AGEMA_signal_6086, SubBytesIns_Inst_Sbox_14_M31}), .clk (clk), .r ({Fresh[597], Fresh[596]}), .c ({new_AGEMA_signal_6185, SubBytesIns_Inst_Sbox_14_M32}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M35_U1 ( .a ({new_AGEMA_signal_10340, new_AGEMA_signal_10339}), .b ({new_AGEMA_signal_5988, SubBytesIns_Inst_Sbox_14_M34}), .clk (clk), .r ({Fresh[599], Fresh[598]}), .c ({new_AGEMA_signal_6186, SubBytesIns_Inst_Sbox_14_M35}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M37_U1 ( .a ({new_AGEMA_signal_10494, new_AGEMA_signal_10493}), .b ({new_AGEMA_signal_6183, SubBytesIns_Inst_Sbox_14_M29}), .c ({new_AGEMA_signal_6265, SubBytesIns_Inst_Sbox_14_M37}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M38_U1 ( .a ({new_AGEMA_signal_6185, SubBytesIns_Inst_Sbox_14_M32}), .b ({new_AGEMA_signal_10496, new_AGEMA_signal_10495}), .c ({new_AGEMA_signal_6266, SubBytesIns_Inst_Sbox_14_M38}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M39_U1 ( .a ({new_AGEMA_signal_10498, new_AGEMA_signal_10497}), .b ({new_AGEMA_signal_6184, SubBytesIns_Inst_Sbox_14_M30}), .c ({new_AGEMA_signal_6267, SubBytesIns_Inst_Sbox_14_M39}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M40_U1 ( .a ({new_AGEMA_signal_6186, SubBytesIns_Inst_Sbox_14_M35}), .b ({new_AGEMA_signal_10500, new_AGEMA_signal_10499}), .c ({new_AGEMA_signal_6268, SubBytesIns_Inst_Sbox_14_M40}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M41_U1 ( .a ({new_AGEMA_signal_6266, SubBytesIns_Inst_Sbox_14_M38}), .b ({new_AGEMA_signal_6268, SubBytesIns_Inst_Sbox_14_M40}), .c ({new_AGEMA_signal_6489, SubBytesIns_Inst_Sbox_14_M41}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M42_U1 ( .a ({new_AGEMA_signal_6265, SubBytesIns_Inst_Sbox_14_M37}), .b ({new_AGEMA_signal_6267, SubBytesIns_Inst_Sbox_14_M39}), .c ({new_AGEMA_signal_6490, SubBytesIns_Inst_Sbox_14_M42}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M43_U1 ( .a ({new_AGEMA_signal_6265, SubBytesIns_Inst_Sbox_14_M37}), .b ({new_AGEMA_signal_6266, SubBytesIns_Inst_Sbox_14_M38}), .c ({new_AGEMA_signal_6491, SubBytesIns_Inst_Sbox_14_M43}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M44_U1 ( .a ({new_AGEMA_signal_6267, SubBytesIns_Inst_Sbox_14_M39}), .b ({new_AGEMA_signal_6268, SubBytesIns_Inst_Sbox_14_M40}), .c ({new_AGEMA_signal_6492, SubBytesIns_Inst_Sbox_14_M44}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M45_U1 ( .a ({new_AGEMA_signal_6490, SubBytesIns_Inst_Sbox_14_M42}), .b ({new_AGEMA_signal_6489, SubBytesIns_Inst_Sbox_14_M41}), .c ({new_AGEMA_signal_6729, SubBytesIns_Inst_Sbox_14_M45}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M29_U1 ( .a ({new_AGEMA_signal_6090, SubBytesIns_Inst_Sbox_15_M28}), .b ({new_AGEMA_signal_10346, new_AGEMA_signal_10345}), .clk (clk), .r ({Fresh[601], Fresh[600]}), .c ({new_AGEMA_signal_6188, SubBytesIns_Inst_Sbox_15_M29}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M30_U1 ( .a ({new_AGEMA_signal_6089, SubBytesIns_Inst_Sbox_15_M26}), .b ({new_AGEMA_signal_10348, new_AGEMA_signal_10347}), .clk (clk), .r ({Fresh[603], Fresh[602]}), .c ({new_AGEMA_signal_6189, SubBytesIns_Inst_Sbox_15_M30}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M32_U1 ( .a ({new_AGEMA_signal_10346, new_AGEMA_signal_10345}), .b ({new_AGEMA_signal_6091, SubBytesIns_Inst_Sbox_15_M31}), .clk (clk), .r ({Fresh[605], Fresh[604]}), .c ({new_AGEMA_signal_6190, SubBytesIns_Inst_Sbox_15_M32}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M35_U1 ( .a ({new_AGEMA_signal_10348, new_AGEMA_signal_10347}), .b ({new_AGEMA_signal_5992, SubBytesIns_Inst_Sbox_15_M34}), .clk (clk), .r ({Fresh[607], Fresh[606]}), .c ({new_AGEMA_signal_6191, SubBytesIns_Inst_Sbox_15_M35}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M37_U1 ( .a ({new_AGEMA_signal_10502, new_AGEMA_signal_10501}), .b ({new_AGEMA_signal_6188, SubBytesIns_Inst_Sbox_15_M29}), .c ({new_AGEMA_signal_6269, SubBytesIns_Inst_Sbox_15_M37}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M38_U1 ( .a ({new_AGEMA_signal_6190, SubBytesIns_Inst_Sbox_15_M32}), .b ({new_AGEMA_signal_10504, new_AGEMA_signal_10503}), .c ({new_AGEMA_signal_6270, SubBytesIns_Inst_Sbox_15_M38}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M39_U1 ( .a ({new_AGEMA_signal_10506, new_AGEMA_signal_10505}), .b ({new_AGEMA_signal_6189, SubBytesIns_Inst_Sbox_15_M30}), .c ({new_AGEMA_signal_6271, SubBytesIns_Inst_Sbox_15_M39}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M40_U1 ( .a ({new_AGEMA_signal_6191, SubBytesIns_Inst_Sbox_15_M35}), .b ({new_AGEMA_signal_10508, new_AGEMA_signal_10507}), .c ({new_AGEMA_signal_6272, SubBytesIns_Inst_Sbox_15_M40}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M41_U1 ( .a ({new_AGEMA_signal_6270, SubBytesIns_Inst_Sbox_15_M38}), .b ({new_AGEMA_signal_6272, SubBytesIns_Inst_Sbox_15_M40}), .c ({new_AGEMA_signal_6501, SubBytesIns_Inst_Sbox_15_M41}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M42_U1 ( .a ({new_AGEMA_signal_6269, SubBytesIns_Inst_Sbox_15_M37}), .b ({new_AGEMA_signal_6271, SubBytesIns_Inst_Sbox_15_M39}), .c ({new_AGEMA_signal_6502, SubBytesIns_Inst_Sbox_15_M42}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M43_U1 ( .a ({new_AGEMA_signal_6269, SubBytesIns_Inst_Sbox_15_M37}), .b ({new_AGEMA_signal_6270, SubBytesIns_Inst_Sbox_15_M38}), .c ({new_AGEMA_signal_6503, SubBytesIns_Inst_Sbox_15_M43}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M44_U1 ( .a ({new_AGEMA_signal_6271, SubBytesIns_Inst_Sbox_15_M39}), .b ({new_AGEMA_signal_6272, SubBytesIns_Inst_Sbox_15_M40}), .c ({new_AGEMA_signal_6504, SubBytesIns_Inst_Sbox_15_M44}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M45_U1 ( .a ({new_AGEMA_signal_6502, SubBytesIns_Inst_Sbox_15_M42}), .b ({new_AGEMA_signal_6501, SubBytesIns_Inst_Sbox_15_M41}), .c ({new_AGEMA_signal_6741, SubBytesIns_Inst_Sbox_15_M45}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M29_U1 ( .a ({new_AGEMA_signal_5995, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M28}), .b ({new_AGEMA_signal_10354, new_AGEMA_signal_10353}), .clk (clk), .r ({Fresh[609], Fresh[608]}), .c ({new_AGEMA_signal_6093, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M29}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M30_U1 ( .a ({new_AGEMA_signal_5994, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M26}), .b ({new_AGEMA_signal_10356, new_AGEMA_signal_10355}), .clk (clk), .r ({Fresh[611], Fresh[610]}), .c ({new_AGEMA_signal_6094, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M30}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M32_U1 ( .a ({new_AGEMA_signal_10354, new_AGEMA_signal_10353}), .b ({new_AGEMA_signal_5996, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M31}), .clk (clk), .r ({Fresh[613], Fresh[612]}), .c ({new_AGEMA_signal_6095, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M32}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M35_U1 ( .a ({new_AGEMA_signal_10356, new_AGEMA_signal_10355}), .b ({new_AGEMA_signal_5916, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M34}), .clk (clk), .r ({Fresh[615], Fresh[614]}), .c ({new_AGEMA_signal_6096, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M35}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M37_U1 ( .a ({new_AGEMA_signal_10510, new_AGEMA_signal_10509}), .b ({new_AGEMA_signal_6093, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M29}), .c ({new_AGEMA_signal_6193, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M38_U1 ( .a ({new_AGEMA_signal_6095, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M32}), .b ({new_AGEMA_signal_10512, new_AGEMA_signal_10511}), .c ({new_AGEMA_signal_6194, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M39_U1 ( .a ({new_AGEMA_signal_10514, new_AGEMA_signal_10513}), .b ({new_AGEMA_signal_6094, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M30}), .c ({new_AGEMA_signal_6195, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M40_U1 ( .a ({new_AGEMA_signal_6096, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M35}), .b ({new_AGEMA_signal_10516, new_AGEMA_signal_10515}), .c ({new_AGEMA_signal_6196, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M41_U1 ( .a ({new_AGEMA_signal_6194, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_6196, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_6273, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M42_U1 ( .a ({new_AGEMA_signal_6193, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_6195, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39}), .c ({new_AGEMA_signal_6274, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M43_U1 ( .a ({new_AGEMA_signal_6193, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_6194, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38}), .c ({new_AGEMA_signal_6275, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M44_U1 ( .a ({new_AGEMA_signal_6195, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_6196, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_6276, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M45_U1 ( .a ({new_AGEMA_signal_6274, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_6273, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41}), .c ({new_AGEMA_signal_6513, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M29_U1 ( .a ({new_AGEMA_signal_6000, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M28}), .b ({new_AGEMA_signal_10362, new_AGEMA_signal_10361}), .clk (clk), .r ({Fresh[617], Fresh[616]}), .c ({new_AGEMA_signal_6098, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M29}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M30_U1 ( .a ({new_AGEMA_signal_5999, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M26}), .b ({new_AGEMA_signal_10364, new_AGEMA_signal_10363}), .clk (clk), .r ({Fresh[619], Fresh[618]}), .c ({new_AGEMA_signal_6099, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M30}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M32_U1 ( .a ({new_AGEMA_signal_10362, new_AGEMA_signal_10361}), .b ({new_AGEMA_signal_6001, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M31}), .clk (clk), .r ({Fresh[621], Fresh[620]}), .c ({new_AGEMA_signal_6100, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M32}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M35_U1 ( .a ({new_AGEMA_signal_10364, new_AGEMA_signal_10363}), .b ({new_AGEMA_signal_5920, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M34}), .clk (clk), .r ({Fresh[623], Fresh[622]}), .c ({new_AGEMA_signal_6101, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M35}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M37_U1 ( .a ({new_AGEMA_signal_10518, new_AGEMA_signal_10517}), .b ({new_AGEMA_signal_6098, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M29}), .c ({new_AGEMA_signal_6197, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M38_U1 ( .a ({new_AGEMA_signal_6100, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M32}), .b ({new_AGEMA_signal_10520, new_AGEMA_signal_10519}), .c ({new_AGEMA_signal_6198, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M39_U1 ( .a ({new_AGEMA_signal_10522, new_AGEMA_signal_10521}), .b ({new_AGEMA_signal_6099, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M30}), .c ({new_AGEMA_signal_6199, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M40_U1 ( .a ({new_AGEMA_signal_6101, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M35}), .b ({new_AGEMA_signal_10524, new_AGEMA_signal_10523}), .c ({new_AGEMA_signal_6200, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M41_U1 ( .a ({new_AGEMA_signal_6198, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_6200, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_6285, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M42_U1 ( .a ({new_AGEMA_signal_6197, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_6199, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39}), .c ({new_AGEMA_signal_6286, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M43_U1 ( .a ({new_AGEMA_signal_6197, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_6198, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38}), .c ({new_AGEMA_signal_6287, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M44_U1 ( .a ({new_AGEMA_signal_6199, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_6200, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_6288, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M45_U1 ( .a ({new_AGEMA_signal_6286, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_6285, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41}), .c ({new_AGEMA_signal_6525, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M29_U1 ( .a ({new_AGEMA_signal_6005, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M28}), .b ({new_AGEMA_signal_10370, new_AGEMA_signal_10369}), .clk (clk), .r ({Fresh[625], Fresh[624]}), .c ({new_AGEMA_signal_6103, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M29}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M30_U1 ( .a ({new_AGEMA_signal_6004, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M26}), .b ({new_AGEMA_signal_10372, new_AGEMA_signal_10371}), .clk (clk), .r ({Fresh[627], Fresh[626]}), .c ({new_AGEMA_signal_6104, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M30}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M32_U1 ( .a ({new_AGEMA_signal_10370, new_AGEMA_signal_10369}), .b ({new_AGEMA_signal_6006, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M31}), .clk (clk), .r ({Fresh[629], Fresh[628]}), .c ({new_AGEMA_signal_6105, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M32}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M35_U1 ( .a ({new_AGEMA_signal_10372, new_AGEMA_signal_10371}), .b ({new_AGEMA_signal_5924, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M34}), .clk (clk), .r ({Fresh[631], Fresh[630]}), .c ({new_AGEMA_signal_6106, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M35}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M37_U1 ( .a ({new_AGEMA_signal_10526, new_AGEMA_signal_10525}), .b ({new_AGEMA_signal_6103, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M29}), .c ({new_AGEMA_signal_6201, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M38_U1 ( .a ({new_AGEMA_signal_6105, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M32}), .b ({new_AGEMA_signal_10528, new_AGEMA_signal_10527}), .c ({new_AGEMA_signal_6202, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M39_U1 ( .a ({new_AGEMA_signal_10530, new_AGEMA_signal_10529}), .b ({new_AGEMA_signal_6104, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M30}), .c ({new_AGEMA_signal_6203, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M40_U1 ( .a ({new_AGEMA_signal_6106, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M35}), .b ({new_AGEMA_signal_10532, new_AGEMA_signal_10531}), .c ({new_AGEMA_signal_6204, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M41_U1 ( .a ({new_AGEMA_signal_6202, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_6204, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_6297, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M42_U1 ( .a ({new_AGEMA_signal_6201, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_6203, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39}), .c ({new_AGEMA_signal_6298, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M43_U1 ( .a ({new_AGEMA_signal_6201, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_6202, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38}), .c ({new_AGEMA_signal_6299, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M44_U1 ( .a ({new_AGEMA_signal_6203, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_6204, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_6300, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M45_U1 ( .a ({new_AGEMA_signal_6298, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_6297, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41}), .c ({new_AGEMA_signal_6537, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M29_U1 ( .a ({new_AGEMA_signal_6010, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M28}), .b ({new_AGEMA_signal_10378, new_AGEMA_signal_10377}), .clk (clk), .r ({Fresh[633], Fresh[632]}), .c ({new_AGEMA_signal_6108, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M29}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M30_U1 ( .a ({new_AGEMA_signal_6009, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M26}), .b ({new_AGEMA_signal_10380, new_AGEMA_signal_10379}), .clk (clk), .r ({Fresh[635], Fresh[634]}), .c ({new_AGEMA_signal_6109, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M30}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M32_U1 ( .a ({new_AGEMA_signal_10378, new_AGEMA_signal_10377}), .b ({new_AGEMA_signal_6011, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M31}), .clk (clk), .r ({Fresh[637], Fresh[636]}), .c ({new_AGEMA_signal_6110, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M32}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M35_U1 ( .a ({new_AGEMA_signal_10380, new_AGEMA_signal_10379}), .b ({new_AGEMA_signal_5928, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M34}), .clk (clk), .r ({Fresh[639], Fresh[638]}), .c ({new_AGEMA_signal_6111, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M35}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M37_U1 ( .a ({new_AGEMA_signal_10534, new_AGEMA_signal_10533}), .b ({new_AGEMA_signal_6108, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M29}), .c ({new_AGEMA_signal_6205, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M38_U1 ( .a ({new_AGEMA_signal_6110, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M32}), .b ({new_AGEMA_signal_10536, new_AGEMA_signal_10535}), .c ({new_AGEMA_signal_6206, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M39_U1 ( .a ({new_AGEMA_signal_10538, new_AGEMA_signal_10537}), .b ({new_AGEMA_signal_6109, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M30}), .c ({new_AGEMA_signal_6207, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M40_U1 ( .a ({new_AGEMA_signal_6111, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M35}), .b ({new_AGEMA_signal_10540, new_AGEMA_signal_10539}), .c ({new_AGEMA_signal_6208, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M41_U1 ( .a ({new_AGEMA_signal_6206, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_6208, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_6309, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M42_U1 ( .a ({new_AGEMA_signal_6205, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_6207, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39}), .c ({new_AGEMA_signal_6310, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M43_U1 ( .a ({new_AGEMA_signal_6205, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_6206, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38}), .c ({new_AGEMA_signal_6311, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M44_U1 ( .a ({new_AGEMA_signal_6207, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_6208, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_6312, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M45_U1 ( .a ({new_AGEMA_signal_6310, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_6309, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41}), .c ({new_AGEMA_signal_6549, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45}) ) ;
    buf_clk new_AGEMA_reg_buffer_4529 ( .C (clk), .D (new_AGEMA_signal_10221), .Q (new_AGEMA_signal_10381) ) ;
    buf_clk new_AGEMA_reg_buffer_4530 ( .C (clk), .D (new_AGEMA_signal_10222), .Q (new_AGEMA_signal_10382) ) ;
    buf_clk new_AGEMA_reg_buffer_4531 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M33), .Q (new_AGEMA_signal_10383) ) ;
    buf_clk new_AGEMA_reg_buffer_4532 ( .C (clk), .D (new_AGEMA_signal_6017), .Q (new_AGEMA_signal_10384) ) ;
    buf_clk new_AGEMA_reg_buffer_4533 ( .C (clk), .D (new_AGEMA_signal_10223), .Q (new_AGEMA_signal_10385) ) ;
    buf_clk new_AGEMA_reg_buffer_4534 ( .C (clk), .D (new_AGEMA_signal_10224), .Q (new_AGEMA_signal_10386) ) ;
    buf_clk new_AGEMA_reg_buffer_4535 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M36), .Q (new_AGEMA_signal_10387) ) ;
    buf_clk new_AGEMA_reg_buffer_4536 ( .C (clk), .D (new_AGEMA_signal_6117), .Q (new_AGEMA_signal_10388) ) ;
    buf_clk new_AGEMA_reg_buffer_4537 ( .C (clk), .D (new_AGEMA_signal_10229), .Q (new_AGEMA_signal_10389) ) ;
    buf_clk new_AGEMA_reg_buffer_4538 ( .C (clk), .D (new_AGEMA_signal_10230), .Q (new_AGEMA_signal_10390) ) ;
    buf_clk new_AGEMA_reg_buffer_4539 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M33), .Q (new_AGEMA_signal_10391) ) ;
    buf_clk new_AGEMA_reg_buffer_4540 ( .C (clk), .D (new_AGEMA_signal_6022), .Q (new_AGEMA_signal_10392) ) ;
    buf_clk new_AGEMA_reg_buffer_4541 ( .C (clk), .D (new_AGEMA_signal_10231), .Q (new_AGEMA_signal_10393) ) ;
    buf_clk new_AGEMA_reg_buffer_4542 ( .C (clk), .D (new_AGEMA_signal_10232), .Q (new_AGEMA_signal_10394) ) ;
    buf_clk new_AGEMA_reg_buffer_4543 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M36), .Q (new_AGEMA_signal_10395) ) ;
    buf_clk new_AGEMA_reg_buffer_4544 ( .C (clk), .D (new_AGEMA_signal_6122), .Q (new_AGEMA_signal_10396) ) ;
    buf_clk new_AGEMA_reg_buffer_4545 ( .C (clk), .D (new_AGEMA_signal_10237), .Q (new_AGEMA_signal_10397) ) ;
    buf_clk new_AGEMA_reg_buffer_4546 ( .C (clk), .D (new_AGEMA_signal_10238), .Q (new_AGEMA_signal_10398) ) ;
    buf_clk new_AGEMA_reg_buffer_4547 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M33), .Q (new_AGEMA_signal_10399) ) ;
    buf_clk new_AGEMA_reg_buffer_4548 ( .C (clk), .D (new_AGEMA_signal_6027), .Q (new_AGEMA_signal_10400) ) ;
    buf_clk new_AGEMA_reg_buffer_4549 ( .C (clk), .D (new_AGEMA_signal_10239), .Q (new_AGEMA_signal_10401) ) ;
    buf_clk new_AGEMA_reg_buffer_4550 ( .C (clk), .D (new_AGEMA_signal_10240), .Q (new_AGEMA_signal_10402) ) ;
    buf_clk new_AGEMA_reg_buffer_4551 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M36), .Q (new_AGEMA_signal_10403) ) ;
    buf_clk new_AGEMA_reg_buffer_4552 ( .C (clk), .D (new_AGEMA_signal_6127), .Q (new_AGEMA_signal_10404) ) ;
    buf_clk new_AGEMA_reg_buffer_4553 ( .C (clk), .D (new_AGEMA_signal_10245), .Q (new_AGEMA_signal_10405) ) ;
    buf_clk new_AGEMA_reg_buffer_4554 ( .C (clk), .D (new_AGEMA_signal_10246), .Q (new_AGEMA_signal_10406) ) ;
    buf_clk new_AGEMA_reg_buffer_4555 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M33), .Q (new_AGEMA_signal_10407) ) ;
    buf_clk new_AGEMA_reg_buffer_4556 ( .C (clk), .D (new_AGEMA_signal_6032), .Q (new_AGEMA_signal_10408) ) ;
    buf_clk new_AGEMA_reg_buffer_4557 ( .C (clk), .D (new_AGEMA_signal_10247), .Q (new_AGEMA_signal_10409) ) ;
    buf_clk new_AGEMA_reg_buffer_4558 ( .C (clk), .D (new_AGEMA_signal_10248), .Q (new_AGEMA_signal_10410) ) ;
    buf_clk new_AGEMA_reg_buffer_4559 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M36), .Q (new_AGEMA_signal_10411) ) ;
    buf_clk new_AGEMA_reg_buffer_4560 ( .C (clk), .D (new_AGEMA_signal_6132), .Q (new_AGEMA_signal_10412) ) ;
    buf_clk new_AGEMA_reg_buffer_4561 ( .C (clk), .D (new_AGEMA_signal_10253), .Q (new_AGEMA_signal_10413) ) ;
    buf_clk new_AGEMA_reg_buffer_4562 ( .C (clk), .D (new_AGEMA_signal_10254), .Q (new_AGEMA_signal_10414) ) ;
    buf_clk new_AGEMA_reg_buffer_4563 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_M33), .Q (new_AGEMA_signal_10415) ) ;
    buf_clk new_AGEMA_reg_buffer_4564 ( .C (clk), .D (new_AGEMA_signal_6037), .Q (new_AGEMA_signal_10416) ) ;
    buf_clk new_AGEMA_reg_buffer_4565 ( .C (clk), .D (new_AGEMA_signal_10255), .Q (new_AGEMA_signal_10417) ) ;
    buf_clk new_AGEMA_reg_buffer_4566 ( .C (clk), .D (new_AGEMA_signal_10256), .Q (new_AGEMA_signal_10418) ) ;
    buf_clk new_AGEMA_reg_buffer_4567 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_M36), .Q (new_AGEMA_signal_10419) ) ;
    buf_clk new_AGEMA_reg_buffer_4568 ( .C (clk), .D (new_AGEMA_signal_6137), .Q (new_AGEMA_signal_10420) ) ;
    buf_clk new_AGEMA_reg_buffer_4569 ( .C (clk), .D (new_AGEMA_signal_10261), .Q (new_AGEMA_signal_10421) ) ;
    buf_clk new_AGEMA_reg_buffer_4570 ( .C (clk), .D (new_AGEMA_signal_10262), .Q (new_AGEMA_signal_10422) ) ;
    buf_clk new_AGEMA_reg_buffer_4571 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_M33), .Q (new_AGEMA_signal_10423) ) ;
    buf_clk new_AGEMA_reg_buffer_4572 ( .C (clk), .D (new_AGEMA_signal_6042), .Q (new_AGEMA_signal_10424) ) ;
    buf_clk new_AGEMA_reg_buffer_4573 ( .C (clk), .D (new_AGEMA_signal_10263), .Q (new_AGEMA_signal_10425) ) ;
    buf_clk new_AGEMA_reg_buffer_4574 ( .C (clk), .D (new_AGEMA_signal_10264), .Q (new_AGEMA_signal_10426) ) ;
    buf_clk new_AGEMA_reg_buffer_4575 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_M36), .Q (new_AGEMA_signal_10427) ) ;
    buf_clk new_AGEMA_reg_buffer_4576 ( .C (clk), .D (new_AGEMA_signal_6142), .Q (new_AGEMA_signal_10428) ) ;
    buf_clk new_AGEMA_reg_buffer_4577 ( .C (clk), .D (new_AGEMA_signal_10269), .Q (new_AGEMA_signal_10429) ) ;
    buf_clk new_AGEMA_reg_buffer_4578 ( .C (clk), .D (new_AGEMA_signal_10270), .Q (new_AGEMA_signal_10430) ) ;
    buf_clk new_AGEMA_reg_buffer_4579 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_M33), .Q (new_AGEMA_signal_10431) ) ;
    buf_clk new_AGEMA_reg_buffer_4580 ( .C (clk), .D (new_AGEMA_signal_6047), .Q (new_AGEMA_signal_10432) ) ;
    buf_clk new_AGEMA_reg_buffer_4581 ( .C (clk), .D (new_AGEMA_signal_10271), .Q (new_AGEMA_signal_10433) ) ;
    buf_clk new_AGEMA_reg_buffer_4582 ( .C (clk), .D (new_AGEMA_signal_10272), .Q (new_AGEMA_signal_10434) ) ;
    buf_clk new_AGEMA_reg_buffer_4583 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_M36), .Q (new_AGEMA_signal_10435) ) ;
    buf_clk new_AGEMA_reg_buffer_4584 ( .C (clk), .D (new_AGEMA_signal_6147), .Q (new_AGEMA_signal_10436) ) ;
    buf_clk new_AGEMA_reg_buffer_4585 ( .C (clk), .D (new_AGEMA_signal_10277), .Q (new_AGEMA_signal_10437) ) ;
    buf_clk new_AGEMA_reg_buffer_4586 ( .C (clk), .D (new_AGEMA_signal_10278), .Q (new_AGEMA_signal_10438) ) ;
    buf_clk new_AGEMA_reg_buffer_4587 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_M33), .Q (new_AGEMA_signal_10439) ) ;
    buf_clk new_AGEMA_reg_buffer_4588 ( .C (clk), .D (new_AGEMA_signal_6052), .Q (new_AGEMA_signal_10440) ) ;
    buf_clk new_AGEMA_reg_buffer_4589 ( .C (clk), .D (new_AGEMA_signal_10279), .Q (new_AGEMA_signal_10441) ) ;
    buf_clk new_AGEMA_reg_buffer_4590 ( .C (clk), .D (new_AGEMA_signal_10280), .Q (new_AGEMA_signal_10442) ) ;
    buf_clk new_AGEMA_reg_buffer_4591 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_M36), .Q (new_AGEMA_signal_10443) ) ;
    buf_clk new_AGEMA_reg_buffer_4592 ( .C (clk), .D (new_AGEMA_signal_6152), .Q (new_AGEMA_signal_10444) ) ;
    buf_clk new_AGEMA_reg_buffer_4593 ( .C (clk), .D (new_AGEMA_signal_10285), .Q (new_AGEMA_signal_10445) ) ;
    buf_clk new_AGEMA_reg_buffer_4594 ( .C (clk), .D (new_AGEMA_signal_10286), .Q (new_AGEMA_signal_10446) ) ;
    buf_clk new_AGEMA_reg_buffer_4595 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_M33), .Q (new_AGEMA_signal_10447) ) ;
    buf_clk new_AGEMA_reg_buffer_4596 ( .C (clk), .D (new_AGEMA_signal_6057), .Q (new_AGEMA_signal_10448) ) ;
    buf_clk new_AGEMA_reg_buffer_4597 ( .C (clk), .D (new_AGEMA_signal_10287), .Q (new_AGEMA_signal_10449) ) ;
    buf_clk new_AGEMA_reg_buffer_4598 ( .C (clk), .D (new_AGEMA_signal_10288), .Q (new_AGEMA_signal_10450) ) ;
    buf_clk new_AGEMA_reg_buffer_4599 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_M36), .Q (new_AGEMA_signal_10451) ) ;
    buf_clk new_AGEMA_reg_buffer_4600 ( .C (clk), .D (new_AGEMA_signal_6157), .Q (new_AGEMA_signal_10452) ) ;
    buf_clk new_AGEMA_reg_buffer_4601 ( .C (clk), .D (new_AGEMA_signal_10293), .Q (new_AGEMA_signal_10453) ) ;
    buf_clk new_AGEMA_reg_buffer_4602 ( .C (clk), .D (new_AGEMA_signal_10294), .Q (new_AGEMA_signal_10454) ) ;
    buf_clk new_AGEMA_reg_buffer_4603 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_M33), .Q (new_AGEMA_signal_10455) ) ;
    buf_clk new_AGEMA_reg_buffer_4604 ( .C (clk), .D (new_AGEMA_signal_6062), .Q (new_AGEMA_signal_10456) ) ;
    buf_clk new_AGEMA_reg_buffer_4605 ( .C (clk), .D (new_AGEMA_signal_10295), .Q (new_AGEMA_signal_10457) ) ;
    buf_clk new_AGEMA_reg_buffer_4606 ( .C (clk), .D (new_AGEMA_signal_10296), .Q (new_AGEMA_signal_10458) ) ;
    buf_clk new_AGEMA_reg_buffer_4607 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_M36), .Q (new_AGEMA_signal_10459) ) ;
    buf_clk new_AGEMA_reg_buffer_4608 ( .C (clk), .D (new_AGEMA_signal_6162), .Q (new_AGEMA_signal_10460) ) ;
    buf_clk new_AGEMA_reg_buffer_4609 ( .C (clk), .D (new_AGEMA_signal_10301), .Q (new_AGEMA_signal_10461) ) ;
    buf_clk new_AGEMA_reg_buffer_4610 ( .C (clk), .D (new_AGEMA_signal_10302), .Q (new_AGEMA_signal_10462) ) ;
    buf_clk new_AGEMA_reg_buffer_4611 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_M33), .Q (new_AGEMA_signal_10463) ) ;
    buf_clk new_AGEMA_reg_buffer_4612 ( .C (clk), .D (new_AGEMA_signal_6067), .Q (new_AGEMA_signal_10464) ) ;
    buf_clk new_AGEMA_reg_buffer_4613 ( .C (clk), .D (new_AGEMA_signal_10303), .Q (new_AGEMA_signal_10465) ) ;
    buf_clk new_AGEMA_reg_buffer_4614 ( .C (clk), .D (new_AGEMA_signal_10304), .Q (new_AGEMA_signal_10466) ) ;
    buf_clk new_AGEMA_reg_buffer_4615 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_M36), .Q (new_AGEMA_signal_10467) ) ;
    buf_clk new_AGEMA_reg_buffer_4616 ( .C (clk), .D (new_AGEMA_signal_6167), .Q (new_AGEMA_signal_10468) ) ;
    buf_clk new_AGEMA_reg_buffer_4617 ( .C (clk), .D (new_AGEMA_signal_10309), .Q (new_AGEMA_signal_10469) ) ;
    buf_clk new_AGEMA_reg_buffer_4618 ( .C (clk), .D (new_AGEMA_signal_10310), .Q (new_AGEMA_signal_10470) ) ;
    buf_clk new_AGEMA_reg_buffer_4619 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_M33), .Q (new_AGEMA_signal_10471) ) ;
    buf_clk new_AGEMA_reg_buffer_4620 ( .C (clk), .D (new_AGEMA_signal_6072), .Q (new_AGEMA_signal_10472) ) ;
    buf_clk new_AGEMA_reg_buffer_4621 ( .C (clk), .D (new_AGEMA_signal_10311), .Q (new_AGEMA_signal_10473) ) ;
    buf_clk new_AGEMA_reg_buffer_4622 ( .C (clk), .D (new_AGEMA_signal_10312), .Q (new_AGEMA_signal_10474) ) ;
    buf_clk new_AGEMA_reg_buffer_4623 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_M36), .Q (new_AGEMA_signal_10475) ) ;
    buf_clk new_AGEMA_reg_buffer_4624 ( .C (clk), .D (new_AGEMA_signal_6172), .Q (new_AGEMA_signal_10476) ) ;
    buf_clk new_AGEMA_reg_buffer_4625 ( .C (clk), .D (new_AGEMA_signal_10317), .Q (new_AGEMA_signal_10477) ) ;
    buf_clk new_AGEMA_reg_buffer_4626 ( .C (clk), .D (new_AGEMA_signal_10318), .Q (new_AGEMA_signal_10478) ) ;
    buf_clk new_AGEMA_reg_buffer_4627 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_M33), .Q (new_AGEMA_signal_10479) ) ;
    buf_clk new_AGEMA_reg_buffer_4628 ( .C (clk), .D (new_AGEMA_signal_6077), .Q (new_AGEMA_signal_10480) ) ;
    buf_clk new_AGEMA_reg_buffer_4629 ( .C (clk), .D (new_AGEMA_signal_10319), .Q (new_AGEMA_signal_10481) ) ;
    buf_clk new_AGEMA_reg_buffer_4630 ( .C (clk), .D (new_AGEMA_signal_10320), .Q (new_AGEMA_signal_10482) ) ;
    buf_clk new_AGEMA_reg_buffer_4631 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_M36), .Q (new_AGEMA_signal_10483) ) ;
    buf_clk new_AGEMA_reg_buffer_4632 ( .C (clk), .D (new_AGEMA_signal_6177), .Q (new_AGEMA_signal_10484) ) ;
    buf_clk new_AGEMA_reg_buffer_4633 ( .C (clk), .D (new_AGEMA_signal_10325), .Q (new_AGEMA_signal_10485) ) ;
    buf_clk new_AGEMA_reg_buffer_4634 ( .C (clk), .D (new_AGEMA_signal_10326), .Q (new_AGEMA_signal_10486) ) ;
    buf_clk new_AGEMA_reg_buffer_4635 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_M33), .Q (new_AGEMA_signal_10487) ) ;
    buf_clk new_AGEMA_reg_buffer_4636 ( .C (clk), .D (new_AGEMA_signal_6082), .Q (new_AGEMA_signal_10488) ) ;
    buf_clk new_AGEMA_reg_buffer_4637 ( .C (clk), .D (new_AGEMA_signal_10327), .Q (new_AGEMA_signal_10489) ) ;
    buf_clk new_AGEMA_reg_buffer_4638 ( .C (clk), .D (new_AGEMA_signal_10328), .Q (new_AGEMA_signal_10490) ) ;
    buf_clk new_AGEMA_reg_buffer_4639 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_M36), .Q (new_AGEMA_signal_10491) ) ;
    buf_clk new_AGEMA_reg_buffer_4640 ( .C (clk), .D (new_AGEMA_signal_6182), .Q (new_AGEMA_signal_10492) ) ;
    buf_clk new_AGEMA_reg_buffer_4641 ( .C (clk), .D (new_AGEMA_signal_10333), .Q (new_AGEMA_signal_10493) ) ;
    buf_clk new_AGEMA_reg_buffer_4642 ( .C (clk), .D (new_AGEMA_signal_10334), .Q (new_AGEMA_signal_10494) ) ;
    buf_clk new_AGEMA_reg_buffer_4643 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_M33), .Q (new_AGEMA_signal_10495) ) ;
    buf_clk new_AGEMA_reg_buffer_4644 ( .C (clk), .D (new_AGEMA_signal_6087), .Q (new_AGEMA_signal_10496) ) ;
    buf_clk new_AGEMA_reg_buffer_4645 ( .C (clk), .D (new_AGEMA_signal_10335), .Q (new_AGEMA_signal_10497) ) ;
    buf_clk new_AGEMA_reg_buffer_4646 ( .C (clk), .D (new_AGEMA_signal_10336), .Q (new_AGEMA_signal_10498) ) ;
    buf_clk new_AGEMA_reg_buffer_4647 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_M36), .Q (new_AGEMA_signal_10499) ) ;
    buf_clk new_AGEMA_reg_buffer_4648 ( .C (clk), .D (new_AGEMA_signal_6187), .Q (new_AGEMA_signal_10500) ) ;
    buf_clk new_AGEMA_reg_buffer_4649 ( .C (clk), .D (new_AGEMA_signal_10341), .Q (new_AGEMA_signal_10501) ) ;
    buf_clk new_AGEMA_reg_buffer_4650 ( .C (clk), .D (new_AGEMA_signal_10342), .Q (new_AGEMA_signal_10502) ) ;
    buf_clk new_AGEMA_reg_buffer_4651 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_M33), .Q (new_AGEMA_signal_10503) ) ;
    buf_clk new_AGEMA_reg_buffer_4652 ( .C (clk), .D (new_AGEMA_signal_6092), .Q (new_AGEMA_signal_10504) ) ;
    buf_clk new_AGEMA_reg_buffer_4653 ( .C (clk), .D (new_AGEMA_signal_10343), .Q (new_AGEMA_signal_10505) ) ;
    buf_clk new_AGEMA_reg_buffer_4654 ( .C (clk), .D (new_AGEMA_signal_10344), .Q (new_AGEMA_signal_10506) ) ;
    buf_clk new_AGEMA_reg_buffer_4655 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_M36), .Q (new_AGEMA_signal_10507) ) ;
    buf_clk new_AGEMA_reg_buffer_4656 ( .C (clk), .D (new_AGEMA_signal_6192), .Q (new_AGEMA_signal_10508) ) ;
    buf_clk new_AGEMA_reg_buffer_4657 ( .C (clk), .D (new_AGEMA_signal_10349), .Q (new_AGEMA_signal_10509) ) ;
    buf_clk new_AGEMA_reg_buffer_4658 ( .C (clk), .D (new_AGEMA_signal_10350), .Q (new_AGEMA_signal_10510) ) ;
    buf_clk new_AGEMA_reg_buffer_4659 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M33), .Q (new_AGEMA_signal_10511) ) ;
    buf_clk new_AGEMA_reg_buffer_4660 ( .C (clk), .D (new_AGEMA_signal_5997), .Q (new_AGEMA_signal_10512) ) ;
    buf_clk new_AGEMA_reg_buffer_4661 ( .C (clk), .D (new_AGEMA_signal_10351), .Q (new_AGEMA_signal_10513) ) ;
    buf_clk new_AGEMA_reg_buffer_4662 ( .C (clk), .D (new_AGEMA_signal_10352), .Q (new_AGEMA_signal_10514) ) ;
    buf_clk new_AGEMA_reg_buffer_4663 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M36), .Q (new_AGEMA_signal_10515) ) ;
    buf_clk new_AGEMA_reg_buffer_4664 ( .C (clk), .D (new_AGEMA_signal_6097), .Q (new_AGEMA_signal_10516) ) ;
    buf_clk new_AGEMA_reg_buffer_4665 ( .C (clk), .D (new_AGEMA_signal_10357), .Q (new_AGEMA_signal_10517) ) ;
    buf_clk new_AGEMA_reg_buffer_4666 ( .C (clk), .D (new_AGEMA_signal_10358), .Q (new_AGEMA_signal_10518) ) ;
    buf_clk new_AGEMA_reg_buffer_4667 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M33), .Q (new_AGEMA_signal_10519) ) ;
    buf_clk new_AGEMA_reg_buffer_4668 ( .C (clk), .D (new_AGEMA_signal_6002), .Q (new_AGEMA_signal_10520) ) ;
    buf_clk new_AGEMA_reg_buffer_4669 ( .C (clk), .D (new_AGEMA_signal_10359), .Q (new_AGEMA_signal_10521) ) ;
    buf_clk new_AGEMA_reg_buffer_4670 ( .C (clk), .D (new_AGEMA_signal_10360), .Q (new_AGEMA_signal_10522) ) ;
    buf_clk new_AGEMA_reg_buffer_4671 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M36), .Q (new_AGEMA_signal_10523) ) ;
    buf_clk new_AGEMA_reg_buffer_4672 ( .C (clk), .D (new_AGEMA_signal_6102), .Q (new_AGEMA_signal_10524) ) ;
    buf_clk new_AGEMA_reg_buffer_4673 ( .C (clk), .D (new_AGEMA_signal_10365), .Q (new_AGEMA_signal_10525) ) ;
    buf_clk new_AGEMA_reg_buffer_4674 ( .C (clk), .D (new_AGEMA_signal_10366), .Q (new_AGEMA_signal_10526) ) ;
    buf_clk new_AGEMA_reg_buffer_4675 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M33), .Q (new_AGEMA_signal_10527) ) ;
    buf_clk new_AGEMA_reg_buffer_4676 ( .C (clk), .D (new_AGEMA_signal_6007), .Q (new_AGEMA_signal_10528) ) ;
    buf_clk new_AGEMA_reg_buffer_4677 ( .C (clk), .D (new_AGEMA_signal_10367), .Q (new_AGEMA_signal_10529) ) ;
    buf_clk new_AGEMA_reg_buffer_4678 ( .C (clk), .D (new_AGEMA_signal_10368), .Q (new_AGEMA_signal_10530) ) ;
    buf_clk new_AGEMA_reg_buffer_4679 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M36), .Q (new_AGEMA_signal_10531) ) ;
    buf_clk new_AGEMA_reg_buffer_4680 ( .C (clk), .D (new_AGEMA_signal_6107), .Q (new_AGEMA_signal_10532) ) ;
    buf_clk new_AGEMA_reg_buffer_4681 ( .C (clk), .D (new_AGEMA_signal_10373), .Q (new_AGEMA_signal_10533) ) ;
    buf_clk new_AGEMA_reg_buffer_4682 ( .C (clk), .D (new_AGEMA_signal_10374), .Q (new_AGEMA_signal_10534) ) ;
    buf_clk new_AGEMA_reg_buffer_4683 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M33), .Q (new_AGEMA_signal_10535) ) ;
    buf_clk new_AGEMA_reg_buffer_4684 ( .C (clk), .D (new_AGEMA_signal_6012), .Q (new_AGEMA_signal_10536) ) ;
    buf_clk new_AGEMA_reg_buffer_4685 ( .C (clk), .D (new_AGEMA_signal_10375), .Q (new_AGEMA_signal_10537) ) ;
    buf_clk new_AGEMA_reg_buffer_4686 ( .C (clk), .D (new_AGEMA_signal_10376), .Q (new_AGEMA_signal_10538) ) ;
    buf_clk new_AGEMA_reg_buffer_4687 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M36), .Q (new_AGEMA_signal_10539) ) ;
    buf_clk new_AGEMA_reg_buffer_4688 ( .C (clk), .D (new_AGEMA_signal_6112), .Q (new_AGEMA_signal_10540) ) ;
    buf_clk new_AGEMA_reg_buffer_4691 ( .C (clk), .D (new_AGEMA_signal_10542), .Q (new_AGEMA_signal_10543) ) ;
    buf_clk new_AGEMA_reg_buffer_4695 ( .C (clk), .D (new_AGEMA_signal_10546), .Q (new_AGEMA_signal_10547) ) ;
    buf_clk new_AGEMA_reg_buffer_4699 ( .C (clk), .D (new_AGEMA_signal_10550), .Q (new_AGEMA_signal_10551) ) ;
    buf_clk new_AGEMA_reg_buffer_4703 ( .C (clk), .D (new_AGEMA_signal_10554), .Q (new_AGEMA_signal_10555) ) ;
    buf_clk new_AGEMA_reg_buffer_4707 ( .C (clk), .D (new_AGEMA_signal_10558), .Q (new_AGEMA_signal_10559) ) ;
    buf_clk new_AGEMA_reg_buffer_4711 ( .C (clk), .D (new_AGEMA_signal_10562), .Q (new_AGEMA_signal_10563) ) ;
    buf_clk new_AGEMA_reg_buffer_4715 ( .C (clk), .D (new_AGEMA_signal_10566), .Q (new_AGEMA_signal_10567) ) ;
    buf_clk new_AGEMA_reg_buffer_4719 ( .C (clk), .D (new_AGEMA_signal_10570), .Q (new_AGEMA_signal_10571) ) ;
    buf_clk new_AGEMA_reg_buffer_4723 ( .C (clk), .D (new_AGEMA_signal_10574), .Q (new_AGEMA_signal_10575) ) ;
    buf_clk new_AGEMA_reg_buffer_4727 ( .C (clk), .D (new_AGEMA_signal_10578), .Q (new_AGEMA_signal_10579) ) ;
    buf_clk new_AGEMA_reg_buffer_4731 ( .C (clk), .D (new_AGEMA_signal_10582), .Q (new_AGEMA_signal_10583) ) ;
    buf_clk new_AGEMA_reg_buffer_4735 ( .C (clk), .D (new_AGEMA_signal_10586), .Q (new_AGEMA_signal_10587) ) ;
    buf_clk new_AGEMA_reg_buffer_4739 ( .C (clk), .D (new_AGEMA_signal_10590), .Q (new_AGEMA_signal_10591) ) ;
    buf_clk new_AGEMA_reg_buffer_4743 ( .C (clk), .D (new_AGEMA_signal_10594), .Q (new_AGEMA_signal_10595) ) ;
    buf_clk new_AGEMA_reg_buffer_4747 ( .C (clk), .D (new_AGEMA_signal_10598), .Q (new_AGEMA_signal_10599) ) ;
    buf_clk new_AGEMA_reg_buffer_4751 ( .C (clk), .D (new_AGEMA_signal_10602), .Q (new_AGEMA_signal_10603) ) ;
    buf_clk new_AGEMA_reg_buffer_4755 ( .C (clk), .D (new_AGEMA_signal_10606), .Q (new_AGEMA_signal_10607) ) ;
    buf_clk new_AGEMA_reg_buffer_4759 ( .C (clk), .D (new_AGEMA_signal_10610), .Q (new_AGEMA_signal_10611) ) ;
    buf_clk new_AGEMA_reg_buffer_4763 ( .C (clk), .D (new_AGEMA_signal_10614), .Q (new_AGEMA_signal_10615) ) ;
    buf_clk new_AGEMA_reg_buffer_4767 ( .C (clk), .D (new_AGEMA_signal_10618), .Q (new_AGEMA_signal_10619) ) ;
    buf_clk new_AGEMA_reg_buffer_4771 ( .C (clk), .D (new_AGEMA_signal_10622), .Q (new_AGEMA_signal_10623) ) ;
    buf_clk new_AGEMA_reg_buffer_4775 ( .C (clk), .D (new_AGEMA_signal_10626), .Q (new_AGEMA_signal_10627) ) ;
    buf_clk new_AGEMA_reg_buffer_4779 ( .C (clk), .D (new_AGEMA_signal_10630), .Q (new_AGEMA_signal_10631) ) ;
    buf_clk new_AGEMA_reg_buffer_4783 ( .C (clk), .D (new_AGEMA_signal_10634), .Q (new_AGEMA_signal_10635) ) ;
    buf_clk new_AGEMA_reg_buffer_4787 ( .C (clk), .D (new_AGEMA_signal_10638), .Q (new_AGEMA_signal_10639) ) ;
    buf_clk new_AGEMA_reg_buffer_4791 ( .C (clk), .D (new_AGEMA_signal_10642), .Q (new_AGEMA_signal_10643) ) ;
    buf_clk new_AGEMA_reg_buffer_4795 ( .C (clk), .D (new_AGEMA_signal_10646), .Q (new_AGEMA_signal_10647) ) ;
    buf_clk new_AGEMA_reg_buffer_4799 ( .C (clk), .D (new_AGEMA_signal_10650), .Q (new_AGEMA_signal_10651) ) ;
    buf_clk new_AGEMA_reg_buffer_4803 ( .C (clk), .D (new_AGEMA_signal_10654), .Q (new_AGEMA_signal_10655) ) ;
    buf_clk new_AGEMA_reg_buffer_4807 ( .C (clk), .D (new_AGEMA_signal_10658), .Q (new_AGEMA_signal_10659) ) ;
    buf_clk new_AGEMA_reg_buffer_4811 ( .C (clk), .D (new_AGEMA_signal_10662), .Q (new_AGEMA_signal_10663) ) ;
    buf_clk new_AGEMA_reg_buffer_4815 ( .C (clk), .D (new_AGEMA_signal_10666), .Q (new_AGEMA_signal_10667) ) ;
    buf_clk new_AGEMA_reg_buffer_4819 ( .C (clk), .D (new_AGEMA_signal_10670), .Q (new_AGEMA_signal_10671) ) ;
    buf_clk new_AGEMA_reg_buffer_4823 ( .C (clk), .D (new_AGEMA_signal_10674), .Q (new_AGEMA_signal_10675) ) ;
    buf_clk new_AGEMA_reg_buffer_4827 ( .C (clk), .D (new_AGEMA_signal_10678), .Q (new_AGEMA_signal_10679) ) ;
    buf_clk new_AGEMA_reg_buffer_4831 ( .C (clk), .D (new_AGEMA_signal_10682), .Q (new_AGEMA_signal_10683) ) ;
    buf_clk new_AGEMA_reg_buffer_4835 ( .C (clk), .D (new_AGEMA_signal_10686), .Q (new_AGEMA_signal_10687) ) ;
    buf_clk new_AGEMA_reg_buffer_4839 ( .C (clk), .D (new_AGEMA_signal_10690), .Q (new_AGEMA_signal_10691) ) ;
    buf_clk new_AGEMA_reg_buffer_4843 ( .C (clk), .D (new_AGEMA_signal_10694), .Q (new_AGEMA_signal_10695) ) ;
    buf_clk new_AGEMA_reg_buffer_4847 ( .C (clk), .D (new_AGEMA_signal_10698), .Q (new_AGEMA_signal_10699) ) ;
    buf_clk new_AGEMA_reg_buffer_4851 ( .C (clk), .D (new_AGEMA_signal_10702), .Q (new_AGEMA_signal_10703) ) ;
    buf_clk new_AGEMA_reg_buffer_4855 ( .C (clk), .D (new_AGEMA_signal_10706), .Q (new_AGEMA_signal_10707) ) ;
    buf_clk new_AGEMA_reg_buffer_4859 ( .C (clk), .D (new_AGEMA_signal_10710), .Q (new_AGEMA_signal_10711) ) ;
    buf_clk new_AGEMA_reg_buffer_4863 ( .C (clk), .D (new_AGEMA_signal_10714), .Q (new_AGEMA_signal_10715) ) ;
    buf_clk new_AGEMA_reg_buffer_4867 ( .C (clk), .D (new_AGEMA_signal_10718), .Q (new_AGEMA_signal_10719) ) ;
    buf_clk new_AGEMA_reg_buffer_4871 ( .C (clk), .D (new_AGEMA_signal_10722), .Q (new_AGEMA_signal_10723) ) ;
    buf_clk new_AGEMA_reg_buffer_4875 ( .C (clk), .D (new_AGEMA_signal_10726), .Q (new_AGEMA_signal_10727) ) ;
    buf_clk new_AGEMA_reg_buffer_4879 ( .C (clk), .D (new_AGEMA_signal_10730), .Q (new_AGEMA_signal_10731) ) ;
    buf_clk new_AGEMA_reg_buffer_4883 ( .C (clk), .D (new_AGEMA_signal_10734), .Q (new_AGEMA_signal_10735) ) ;
    buf_clk new_AGEMA_reg_buffer_4887 ( .C (clk), .D (new_AGEMA_signal_10738), .Q (new_AGEMA_signal_10739) ) ;
    buf_clk new_AGEMA_reg_buffer_4891 ( .C (clk), .D (new_AGEMA_signal_10742), .Q (new_AGEMA_signal_10743) ) ;
    buf_clk new_AGEMA_reg_buffer_4895 ( .C (clk), .D (new_AGEMA_signal_10746), .Q (new_AGEMA_signal_10747) ) ;
    buf_clk new_AGEMA_reg_buffer_4899 ( .C (clk), .D (new_AGEMA_signal_10750), .Q (new_AGEMA_signal_10751) ) ;
    buf_clk new_AGEMA_reg_buffer_4903 ( .C (clk), .D (new_AGEMA_signal_10754), .Q (new_AGEMA_signal_10755) ) ;
    buf_clk new_AGEMA_reg_buffer_4907 ( .C (clk), .D (new_AGEMA_signal_10758), .Q (new_AGEMA_signal_10759) ) ;
    buf_clk new_AGEMA_reg_buffer_4911 ( .C (clk), .D (new_AGEMA_signal_10762), .Q (new_AGEMA_signal_10763) ) ;
    buf_clk new_AGEMA_reg_buffer_4915 ( .C (clk), .D (new_AGEMA_signal_10766), .Q (new_AGEMA_signal_10767) ) ;
    buf_clk new_AGEMA_reg_buffer_4919 ( .C (clk), .D (new_AGEMA_signal_10770), .Q (new_AGEMA_signal_10771) ) ;
    buf_clk new_AGEMA_reg_buffer_4923 ( .C (clk), .D (new_AGEMA_signal_10774), .Q (new_AGEMA_signal_10775) ) ;
    buf_clk new_AGEMA_reg_buffer_4927 ( .C (clk), .D (new_AGEMA_signal_10778), .Q (new_AGEMA_signal_10779) ) ;
    buf_clk new_AGEMA_reg_buffer_4931 ( .C (clk), .D (new_AGEMA_signal_10782), .Q (new_AGEMA_signal_10783) ) ;
    buf_clk new_AGEMA_reg_buffer_4935 ( .C (clk), .D (new_AGEMA_signal_10786), .Q (new_AGEMA_signal_10787) ) ;
    buf_clk new_AGEMA_reg_buffer_4939 ( .C (clk), .D (new_AGEMA_signal_10790), .Q (new_AGEMA_signal_10791) ) ;
    buf_clk new_AGEMA_reg_buffer_4943 ( .C (clk), .D (new_AGEMA_signal_10794), .Q (new_AGEMA_signal_10795) ) ;
    buf_clk new_AGEMA_reg_buffer_4947 ( .C (clk), .D (new_AGEMA_signal_10798), .Q (new_AGEMA_signal_10799) ) ;
    buf_clk new_AGEMA_reg_buffer_4951 ( .C (clk), .D (new_AGEMA_signal_10802), .Q (new_AGEMA_signal_10803) ) ;
    buf_clk new_AGEMA_reg_buffer_4955 ( .C (clk), .D (new_AGEMA_signal_10806), .Q (new_AGEMA_signal_10807) ) ;
    buf_clk new_AGEMA_reg_buffer_4959 ( .C (clk), .D (new_AGEMA_signal_10810), .Q (new_AGEMA_signal_10811) ) ;
    buf_clk new_AGEMA_reg_buffer_4963 ( .C (clk), .D (new_AGEMA_signal_10814), .Q (new_AGEMA_signal_10815) ) ;
    buf_clk new_AGEMA_reg_buffer_4967 ( .C (clk), .D (new_AGEMA_signal_10818), .Q (new_AGEMA_signal_10819) ) ;
    buf_clk new_AGEMA_reg_buffer_4971 ( .C (clk), .D (new_AGEMA_signal_10822), .Q (new_AGEMA_signal_10823) ) ;
    buf_clk new_AGEMA_reg_buffer_4975 ( .C (clk), .D (new_AGEMA_signal_10826), .Q (new_AGEMA_signal_10827) ) ;
    buf_clk new_AGEMA_reg_buffer_4979 ( .C (clk), .D (new_AGEMA_signal_10830), .Q (new_AGEMA_signal_10831) ) ;
    buf_clk new_AGEMA_reg_buffer_4983 ( .C (clk), .D (new_AGEMA_signal_10834), .Q (new_AGEMA_signal_10835) ) ;
    buf_clk new_AGEMA_reg_buffer_4987 ( .C (clk), .D (new_AGEMA_signal_10838), .Q (new_AGEMA_signal_10839) ) ;
    buf_clk new_AGEMA_reg_buffer_4991 ( .C (clk), .D (new_AGEMA_signal_10842), .Q (new_AGEMA_signal_10843) ) ;
    buf_clk new_AGEMA_reg_buffer_4995 ( .C (clk), .D (new_AGEMA_signal_10846), .Q (new_AGEMA_signal_10847) ) ;
    buf_clk new_AGEMA_reg_buffer_4999 ( .C (clk), .D (new_AGEMA_signal_10850), .Q (new_AGEMA_signal_10851) ) ;
    buf_clk new_AGEMA_reg_buffer_5003 ( .C (clk), .D (new_AGEMA_signal_10854), .Q (new_AGEMA_signal_10855) ) ;
    buf_clk new_AGEMA_reg_buffer_5007 ( .C (clk), .D (new_AGEMA_signal_10858), .Q (new_AGEMA_signal_10859) ) ;
    buf_clk new_AGEMA_reg_buffer_5011 ( .C (clk), .D (new_AGEMA_signal_10862), .Q (new_AGEMA_signal_10863) ) ;
    buf_clk new_AGEMA_reg_buffer_5015 ( .C (clk), .D (new_AGEMA_signal_10866), .Q (new_AGEMA_signal_10867) ) ;
    buf_clk new_AGEMA_reg_buffer_5019 ( .C (clk), .D (new_AGEMA_signal_10870), .Q (new_AGEMA_signal_10871) ) ;
    buf_clk new_AGEMA_reg_buffer_5023 ( .C (clk), .D (new_AGEMA_signal_10874), .Q (new_AGEMA_signal_10875) ) ;
    buf_clk new_AGEMA_reg_buffer_5027 ( .C (clk), .D (new_AGEMA_signal_10878), .Q (new_AGEMA_signal_10879) ) ;
    buf_clk new_AGEMA_reg_buffer_5031 ( .C (clk), .D (new_AGEMA_signal_10882), .Q (new_AGEMA_signal_10883) ) ;
    buf_clk new_AGEMA_reg_buffer_5035 ( .C (clk), .D (new_AGEMA_signal_10886), .Q (new_AGEMA_signal_10887) ) ;
    buf_clk new_AGEMA_reg_buffer_5039 ( .C (clk), .D (new_AGEMA_signal_10890), .Q (new_AGEMA_signal_10891) ) ;
    buf_clk new_AGEMA_reg_buffer_5043 ( .C (clk), .D (new_AGEMA_signal_10894), .Q (new_AGEMA_signal_10895) ) ;
    buf_clk new_AGEMA_reg_buffer_5047 ( .C (clk), .D (new_AGEMA_signal_10898), .Q (new_AGEMA_signal_10899) ) ;
    buf_clk new_AGEMA_reg_buffer_5051 ( .C (clk), .D (new_AGEMA_signal_10902), .Q (new_AGEMA_signal_10903) ) ;
    buf_clk new_AGEMA_reg_buffer_5055 ( .C (clk), .D (new_AGEMA_signal_10906), .Q (new_AGEMA_signal_10907) ) ;
    buf_clk new_AGEMA_reg_buffer_5059 ( .C (clk), .D (new_AGEMA_signal_10910), .Q (new_AGEMA_signal_10911) ) ;
    buf_clk new_AGEMA_reg_buffer_5063 ( .C (clk), .D (new_AGEMA_signal_10914), .Q (new_AGEMA_signal_10915) ) ;
    buf_clk new_AGEMA_reg_buffer_5067 ( .C (clk), .D (new_AGEMA_signal_10918), .Q (new_AGEMA_signal_10919) ) ;
    buf_clk new_AGEMA_reg_buffer_5071 ( .C (clk), .D (new_AGEMA_signal_10922), .Q (new_AGEMA_signal_10923) ) ;
    buf_clk new_AGEMA_reg_buffer_5075 ( .C (clk), .D (new_AGEMA_signal_10926), .Q (new_AGEMA_signal_10927) ) ;
    buf_clk new_AGEMA_reg_buffer_5079 ( .C (clk), .D (new_AGEMA_signal_10930), .Q (new_AGEMA_signal_10931) ) ;
    buf_clk new_AGEMA_reg_buffer_5083 ( .C (clk), .D (new_AGEMA_signal_10934), .Q (new_AGEMA_signal_10935) ) ;
    buf_clk new_AGEMA_reg_buffer_5087 ( .C (clk), .D (new_AGEMA_signal_10938), .Q (new_AGEMA_signal_10939) ) ;
    buf_clk new_AGEMA_reg_buffer_5091 ( .C (clk), .D (new_AGEMA_signal_10942), .Q (new_AGEMA_signal_10943) ) ;
    buf_clk new_AGEMA_reg_buffer_5095 ( .C (clk), .D (new_AGEMA_signal_10946), .Q (new_AGEMA_signal_10947) ) ;
    buf_clk new_AGEMA_reg_buffer_5099 ( .C (clk), .D (new_AGEMA_signal_10950), .Q (new_AGEMA_signal_10951) ) ;
    buf_clk new_AGEMA_reg_buffer_5103 ( .C (clk), .D (new_AGEMA_signal_10954), .Q (new_AGEMA_signal_10955) ) ;
    buf_clk new_AGEMA_reg_buffer_5107 ( .C (clk), .D (new_AGEMA_signal_10958), .Q (new_AGEMA_signal_10959) ) ;
    buf_clk new_AGEMA_reg_buffer_5111 ( .C (clk), .D (new_AGEMA_signal_10962), .Q (new_AGEMA_signal_10963) ) ;
    buf_clk new_AGEMA_reg_buffer_5115 ( .C (clk), .D (new_AGEMA_signal_10966), .Q (new_AGEMA_signal_10967) ) ;
    buf_clk new_AGEMA_reg_buffer_5119 ( .C (clk), .D (new_AGEMA_signal_10970), .Q (new_AGEMA_signal_10971) ) ;
    buf_clk new_AGEMA_reg_buffer_5123 ( .C (clk), .D (new_AGEMA_signal_10974), .Q (new_AGEMA_signal_10975) ) ;
    buf_clk new_AGEMA_reg_buffer_5127 ( .C (clk), .D (new_AGEMA_signal_10978), .Q (new_AGEMA_signal_10979) ) ;
    buf_clk new_AGEMA_reg_buffer_5131 ( .C (clk), .D (new_AGEMA_signal_10982), .Q (new_AGEMA_signal_10983) ) ;
    buf_clk new_AGEMA_reg_buffer_5135 ( .C (clk), .D (new_AGEMA_signal_10986), .Q (new_AGEMA_signal_10987) ) ;
    buf_clk new_AGEMA_reg_buffer_5139 ( .C (clk), .D (new_AGEMA_signal_10990), .Q (new_AGEMA_signal_10991) ) ;
    buf_clk new_AGEMA_reg_buffer_5143 ( .C (clk), .D (new_AGEMA_signal_10994), .Q (new_AGEMA_signal_10995) ) ;
    buf_clk new_AGEMA_reg_buffer_5147 ( .C (clk), .D (new_AGEMA_signal_10998), .Q (new_AGEMA_signal_10999) ) ;
    buf_clk new_AGEMA_reg_buffer_5151 ( .C (clk), .D (new_AGEMA_signal_11002), .Q (new_AGEMA_signal_11003) ) ;
    buf_clk new_AGEMA_reg_buffer_5155 ( .C (clk), .D (new_AGEMA_signal_11006), .Q (new_AGEMA_signal_11007) ) ;
    buf_clk new_AGEMA_reg_buffer_5159 ( .C (clk), .D (new_AGEMA_signal_11010), .Q (new_AGEMA_signal_11011) ) ;
    buf_clk new_AGEMA_reg_buffer_5163 ( .C (clk), .D (new_AGEMA_signal_11014), .Q (new_AGEMA_signal_11015) ) ;
    buf_clk new_AGEMA_reg_buffer_5167 ( .C (clk), .D (new_AGEMA_signal_11018), .Q (new_AGEMA_signal_11019) ) ;
    buf_clk new_AGEMA_reg_buffer_5171 ( .C (clk), .D (new_AGEMA_signal_11022), .Q (new_AGEMA_signal_11023) ) ;
    buf_clk new_AGEMA_reg_buffer_5175 ( .C (clk), .D (new_AGEMA_signal_11026), .Q (new_AGEMA_signal_11027) ) ;
    buf_clk new_AGEMA_reg_buffer_5179 ( .C (clk), .D (new_AGEMA_signal_11030), .Q (new_AGEMA_signal_11031) ) ;
    buf_clk new_AGEMA_reg_buffer_5183 ( .C (clk), .D (new_AGEMA_signal_11034), .Q (new_AGEMA_signal_11035) ) ;
    buf_clk new_AGEMA_reg_buffer_5187 ( .C (clk), .D (new_AGEMA_signal_11038), .Q (new_AGEMA_signal_11039) ) ;
    buf_clk new_AGEMA_reg_buffer_5191 ( .C (clk), .D (new_AGEMA_signal_11042), .Q (new_AGEMA_signal_11043) ) ;
    buf_clk new_AGEMA_reg_buffer_5195 ( .C (clk), .D (new_AGEMA_signal_11046), .Q (new_AGEMA_signal_11047) ) ;
    buf_clk new_AGEMA_reg_buffer_5199 ( .C (clk), .D (new_AGEMA_signal_11050), .Q (new_AGEMA_signal_11051) ) ;
    buf_clk new_AGEMA_reg_buffer_5203 ( .C (clk), .D (new_AGEMA_signal_11054), .Q (new_AGEMA_signal_11055) ) ;
    buf_clk new_AGEMA_reg_buffer_5207 ( .C (clk), .D (new_AGEMA_signal_11058), .Q (new_AGEMA_signal_11059) ) ;
    buf_clk new_AGEMA_reg_buffer_5211 ( .C (clk), .D (new_AGEMA_signal_11062), .Q (new_AGEMA_signal_11063) ) ;
    buf_clk new_AGEMA_reg_buffer_5215 ( .C (clk), .D (new_AGEMA_signal_11066), .Q (new_AGEMA_signal_11067) ) ;
    buf_clk new_AGEMA_reg_buffer_5219 ( .C (clk), .D (new_AGEMA_signal_11070), .Q (new_AGEMA_signal_11071) ) ;
    buf_clk new_AGEMA_reg_buffer_5223 ( .C (clk), .D (new_AGEMA_signal_11074), .Q (new_AGEMA_signal_11075) ) ;
    buf_clk new_AGEMA_reg_buffer_5227 ( .C (clk), .D (new_AGEMA_signal_11078), .Q (new_AGEMA_signal_11079) ) ;
    buf_clk new_AGEMA_reg_buffer_5231 ( .C (clk), .D (new_AGEMA_signal_11082), .Q (new_AGEMA_signal_11083) ) ;
    buf_clk new_AGEMA_reg_buffer_5235 ( .C (clk), .D (new_AGEMA_signal_11086), .Q (new_AGEMA_signal_11087) ) ;
    buf_clk new_AGEMA_reg_buffer_5239 ( .C (clk), .D (new_AGEMA_signal_11090), .Q (new_AGEMA_signal_11091) ) ;
    buf_clk new_AGEMA_reg_buffer_5243 ( .C (clk), .D (new_AGEMA_signal_11094), .Q (new_AGEMA_signal_11095) ) ;
    buf_clk new_AGEMA_reg_buffer_5247 ( .C (clk), .D (new_AGEMA_signal_11098), .Q (new_AGEMA_signal_11099) ) ;
    buf_clk new_AGEMA_reg_buffer_5251 ( .C (clk), .D (new_AGEMA_signal_11102), .Q (new_AGEMA_signal_11103) ) ;
    buf_clk new_AGEMA_reg_buffer_5255 ( .C (clk), .D (new_AGEMA_signal_11106), .Q (new_AGEMA_signal_11107) ) ;
    buf_clk new_AGEMA_reg_buffer_5259 ( .C (clk), .D (new_AGEMA_signal_11110), .Q (new_AGEMA_signal_11111) ) ;
    buf_clk new_AGEMA_reg_buffer_5263 ( .C (clk), .D (new_AGEMA_signal_11114), .Q (new_AGEMA_signal_11115) ) ;
    buf_clk new_AGEMA_reg_buffer_5267 ( .C (clk), .D (new_AGEMA_signal_11118), .Q (new_AGEMA_signal_11119) ) ;
    buf_clk new_AGEMA_reg_buffer_5271 ( .C (clk), .D (new_AGEMA_signal_11122), .Q (new_AGEMA_signal_11123) ) ;
    buf_clk new_AGEMA_reg_buffer_5275 ( .C (clk), .D (new_AGEMA_signal_11126), .Q (new_AGEMA_signal_11127) ) ;
    buf_clk new_AGEMA_reg_buffer_5279 ( .C (clk), .D (new_AGEMA_signal_11130), .Q (new_AGEMA_signal_11131) ) ;
    buf_clk new_AGEMA_reg_buffer_5283 ( .C (clk), .D (new_AGEMA_signal_11134), .Q (new_AGEMA_signal_11135) ) ;
    buf_clk new_AGEMA_reg_buffer_5287 ( .C (clk), .D (new_AGEMA_signal_11138), .Q (new_AGEMA_signal_11139) ) ;
    buf_clk new_AGEMA_reg_buffer_5291 ( .C (clk), .D (new_AGEMA_signal_11142), .Q (new_AGEMA_signal_11143) ) ;
    buf_clk new_AGEMA_reg_buffer_5295 ( .C (clk), .D (new_AGEMA_signal_11146), .Q (new_AGEMA_signal_11147) ) ;
    buf_clk new_AGEMA_reg_buffer_5299 ( .C (clk), .D (new_AGEMA_signal_11150), .Q (new_AGEMA_signal_11151) ) ;
    buf_clk new_AGEMA_reg_buffer_5303 ( .C (clk), .D (new_AGEMA_signal_11154), .Q (new_AGEMA_signal_11155) ) ;
    buf_clk new_AGEMA_reg_buffer_5307 ( .C (clk), .D (new_AGEMA_signal_11158), .Q (new_AGEMA_signal_11159) ) ;
    buf_clk new_AGEMA_reg_buffer_5311 ( .C (clk), .D (new_AGEMA_signal_11162), .Q (new_AGEMA_signal_11163) ) ;
    buf_clk new_AGEMA_reg_buffer_5315 ( .C (clk), .D (new_AGEMA_signal_11166), .Q (new_AGEMA_signal_11167) ) ;
    buf_clk new_AGEMA_reg_buffer_5319 ( .C (clk), .D (new_AGEMA_signal_11170), .Q (new_AGEMA_signal_11171) ) ;
    buf_clk new_AGEMA_reg_buffer_5323 ( .C (clk), .D (new_AGEMA_signal_11174), .Q (new_AGEMA_signal_11175) ) ;
    buf_clk new_AGEMA_reg_buffer_5327 ( .C (clk), .D (new_AGEMA_signal_11178), .Q (new_AGEMA_signal_11179) ) ;
    buf_clk new_AGEMA_reg_buffer_5331 ( .C (clk), .D (new_AGEMA_signal_11182), .Q (new_AGEMA_signal_11183) ) ;
    buf_clk new_AGEMA_reg_buffer_5335 ( .C (clk), .D (new_AGEMA_signal_11186), .Q (new_AGEMA_signal_11187) ) ;
    buf_clk new_AGEMA_reg_buffer_5339 ( .C (clk), .D (new_AGEMA_signal_11190), .Q (new_AGEMA_signal_11191) ) ;
    buf_clk new_AGEMA_reg_buffer_5343 ( .C (clk), .D (new_AGEMA_signal_11194), .Q (new_AGEMA_signal_11195) ) ;
    buf_clk new_AGEMA_reg_buffer_5347 ( .C (clk), .D (new_AGEMA_signal_11198), .Q (new_AGEMA_signal_11199) ) ;
    buf_clk new_AGEMA_reg_buffer_5351 ( .C (clk), .D (new_AGEMA_signal_11202), .Q (new_AGEMA_signal_11203) ) ;
    buf_clk new_AGEMA_reg_buffer_5355 ( .C (clk), .D (new_AGEMA_signal_11206), .Q (new_AGEMA_signal_11207) ) ;
    buf_clk new_AGEMA_reg_buffer_5359 ( .C (clk), .D (new_AGEMA_signal_11210), .Q (new_AGEMA_signal_11211) ) ;
    buf_clk new_AGEMA_reg_buffer_5363 ( .C (clk), .D (new_AGEMA_signal_11214), .Q (new_AGEMA_signal_11215) ) ;
    buf_clk new_AGEMA_reg_buffer_5367 ( .C (clk), .D (new_AGEMA_signal_11218), .Q (new_AGEMA_signal_11219) ) ;
    buf_clk new_AGEMA_reg_buffer_5371 ( .C (clk), .D (new_AGEMA_signal_11222), .Q (new_AGEMA_signal_11223) ) ;
    buf_clk new_AGEMA_reg_buffer_5375 ( .C (clk), .D (new_AGEMA_signal_11226), .Q (new_AGEMA_signal_11227) ) ;
    buf_clk new_AGEMA_reg_buffer_5379 ( .C (clk), .D (new_AGEMA_signal_11230), .Q (new_AGEMA_signal_11231) ) ;
    buf_clk new_AGEMA_reg_buffer_5383 ( .C (clk), .D (new_AGEMA_signal_11234), .Q (new_AGEMA_signal_11235) ) ;
    buf_clk new_AGEMA_reg_buffer_5387 ( .C (clk), .D (new_AGEMA_signal_11238), .Q (new_AGEMA_signal_11239) ) ;
    buf_clk new_AGEMA_reg_buffer_5391 ( .C (clk), .D (new_AGEMA_signal_11242), .Q (new_AGEMA_signal_11243) ) ;
    buf_clk new_AGEMA_reg_buffer_5395 ( .C (clk), .D (new_AGEMA_signal_11246), .Q (new_AGEMA_signal_11247) ) ;
    buf_clk new_AGEMA_reg_buffer_5399 ( .C (clk), .D (new_AGEMA_signal_11250), .Q (new_AGEMA_signal_11251) ) ;
    buf_clk new_AGEMA_reg_buffer_5403 ( .C (clk), .D (new_AGEMA_signal_11254), .Q (new_AGEMA_signal_11255) ) ;
    buf_clk new_AGEMA_reg_buffer_5407 ( .C (clk), .D (new_AGEMA_signal_11258), .Q (new_AGEMA_signal_11259) ) ;
    buf_clk new_AGEMA_reg_buffer_5411 ( .C (clk), .D (new_AGEMA_signal_11262), .Q (new_AGEMA_signal_11263) ) ;
    buf_clk new_AGEMA_reg_buffer_5415 ( .C (clk), .D (new_AGEMA_signal_11266), .Q (new_AGEMA_signal_11267) ) ;
    buf_clk new_AGEMA_reg_buffer_5419 ( .C (clk), .D (new_AGEMA_signal_11270), .Q (new_AGEMA_signal_11271) ) ;
    buf_clk new_AGEMA_reg_buffer_5423 ( .C (clk), .D (new_AGEMA_signal_11274), .Q (new_AGEMA_signal_11275) ) ;
    buf_clk new_AGEMA_reg_buffer_5427 ( .C (clk), .D (new_AGEMA_signal_11278), .Q (new_AGEMA_signal_11279) ) ;
    buf_clk new_AGEMA_reg_buffer_5431 ( .C (clk), .D (new_AGEMA_signal_11282), .Q (new_AGEMA_signal_11283) ) ;
    buf_clk new_AGEMA_reg_buffer_5435 ( .C (clk), .D (new_AGEMA_signal_11286), .Q (new_AGEMA_signal_11287) ) ;
    buf_clk new_AGEMA_reg_buffer_5439 ( .C (clk), .D (new_AGEMA_signal_11290), .Q (new_AGEMA_signal_11291) ) ;
    buf_clk new_AGEMA_reg_buffer_5443 ( .C (clk), .D (new_AGEMA_signal_11294), .Q (new_AGEMA_signal_11295) ) ;
    buf_clk new_AGEMA_reg_buffer_5447 ( .C (clk), .D (new_AGEMA_signal_11298), .Q (new_AGEMA_signal_11299) ) ;
    buf_clk new_AGEMA_reg_buffer_5451 ( .C (clk), .D (new_AGEMA_signal_11302), .Q (new_AGEMA_signal_11303) ) ;
    buf_clk new_AGEMA_reg_buffer_5455 ( .C (clk), .D (new_AGEMA_signal_11306), .Q (new_AGEMA_signal_11307) ) ;
    buf_clk new_AGEMA_reg_buffer_5459 ( .C (clk), .D (new_AGEMA_signal_11310), .Q (new_AGEMA_signal_11311) ) ;
    buf_clk new_AGEMA_reg_buffer_5463 ( .C (clk), .D (new_AGEMA_signal_11314), .Q (new_AGEMA_signal_11315) ) ;
    buf_clk new_AGEMA_reg_buffer_5467 ( .C (clk), .D (new_AGEMA_signal_11318), .Q (new_AGEMA_signal_11319) ) ;
    buf_clk new_AGEMA_reg_buffer_5471 ( .C (clk), .D (new_AGEMA_signal_11322), .Q (new_AGEMA_signal_11323) ) ;
    buf_clk new_AGEMA_reg_buffer_5475 ( .C (clk), .D (new_AGEMA_signal_11326), .Q (new_AGEMA_signal_11327) ) ;
    buf_clk new_AGEMA_reg_buffer_5479 ( .C (clk), .D (new_AGEMA_signal_11330), .Q (new_AGEMA_signal_11331) ) ;
    buf_clk new_AGEMA_reg_buffer_5483 ( .C (clk), .D (new_AGEMA_signal_11334), .Q (new_AGEMA_signal_11335) ) ;
    buf_clk new_AGEMA_reg_buffer_5487 ( .C (clk), .D (new_AGEMA_signal_11338), .Q (new_AGEMA_signal_11339) ) ;
    buf_clk new_AGEMA_reg_buffer_5491 ( .C (clk), .D (new_AGEMA_signal_11342), .Q (new_AGEMA_signal_11343) ) ;
    buf_clk new_AGEMA_reg_buffer_5495 ( .C (clk), .D (new_AGEMA_signal_11346), .Q (new_AGEMA_signal_11347) ) ;
    buf_clk new_AGEMA_reg_buffer_5499 ( .C (clk), .D (new_AGEMA_signal_11350), .Q (new_AGEMA_signal_11351) ) ;
    buf_clk new_AGEMA_reg_buffer_5503 ( .C (clk), .D (new_AGEMA_signal_11354), .Q (new_AGEMA_signal_11355) ) ;
    buf_clk new_AGEMA_reg_buffer_5507 ( .C (clk), .D (new_AGEMA_signal_11358), .Q (new_AGEMA_signal_11359) ) ;
    buf_clk new_AGEMA_reg_buffer_5511 ( .C (clk), .D (new_AGEMA_signal_11362), .Q (new_AGEMA_signal_11363) ) ;
    buf_clk new_AGEMA_reg_buffer_5515 ( .C (clk), .D (new_AGEMA_signal_11366), .Q (new_AGEMA_signal_11367) ) ;
    buf_clk new_AGEMA_reg_buffer_5519 ( .C (clk), .D (new_AGEMA_signal_11370), .Q (new_AGEMA_signal_11371) ) ;
    buf_clk new_AGEMA_reg_buffer_5523 ( .C (clk), .D (new_AGEMA_signal_11374), .Q (new_AGEMA_signal_11375) ) ;
    buf_clk new_AGEMA_reg_buffer_5527 ( .C (clk), .D (new_AGEMA_signal_11378), .Q (new_AGEMA_signal_11379) ) ;
    buf_clk new_AGEMA_reg_buffer_5531 ( .C (clk), .D (new_AGEMA_signal_11382), .Q (new_AGEMA_signal_11383) ) ;
    buf_clk new_AGEMA_reg_buffer_5535 ( .C (clk), .D (new_AGEMA_signal_11386), .Q (new_AGEMA_signal_11387) ) ;
    buf_clk new_AGEMA_reg_buffer_5539 ( .C (clk), .D (new_AGEMA_signal_11390), .Q (new_AGEMA_signal_11391) ) ;
    buf_clk new_AGEMA_reg_buffer_5543 ( .C (clk), .D (new_AGEMA_signal_11394), .Q (new_AGEMA_signal_11395) ) ;
    buf_clk new_AGEMA_reg_buffer_5547 ( .C (clk), .D (new_AGEMA_signal_11398), .Q (new_AGEMA_signal_11399) ) ;
    buf_clk new_AGEMA_reg_buffer_5551 ( .C (clk), .D (new_AGEMA_signal_11402), .Q (new_AGEMA_signal_11403) ) ;
    buf_clk new_AGEMA_reg_buffer_5555 ( .C (clk), .D (new_AGEMA_signal_11406), .Q (new_AGEMA_signal_11407) ) ;
    buf_clk new_AGEMA_reg_buffer_5559 ( .C (clk), .D (new_AGEMA_signal_11410), .Q (new_AGEMA_signal_11411) ) ;
    buf_clk new_AGEMA_reg_buffer_5563 ( .C (clk), .D (new_AGEMA_signal_11414), .Q (new_AGEMA_signal_11415) ) ;
    buf_clk new_AGEMA_reg_buffer_5567 ( .C (clk), .D (new_AGEMA_signal_11418), .Q (new_AGEMA_signal_11419) ) ;
    buf_clk new_AGEMA_reg_buffer_5571 ( .C (clk), .D (new_AGEMA_signal_11422), .Q (new_AGEMA_signal_11423) ) ;
    buf_clk new_AGEMA_reg_buffer_5575 ( .C (clk), .D (new_AGEMA_signal_11426), .Q (new_AGEMA_signal_11427) ) ;
    buf_clk new_AGEMA_reg_buffer_5579 ( .C (clk), .D (new_AGEMA_signal_11430), .Q (new_AGEMA_signal_11431) ) ;
    buf_clk new_AGEMA_reg_buffer_5583 ( .C (clk), .D (new_AGEMA_signal_11434), .Q (new_AGEMA_signal_11435) ) ;
    buf_clk new_AGEMA_reg_buffer_5587 ( .C (clk), .D (new_AGEMA_signal_11438), .Q (new_AGEMA_signal_11439) ) ;
    buf_clk new_AGEMA_reg_buffer_5591 ( .C (clk), .D (new_AGEMA_signal_11442), .Q (new_AGEMA_signal_11443) ) ;
    buf_clk new_AGEMA_reg_buffer_5595 ( .C (clk), .D (new_AGEMA_signal_11446), .Q (new_AGEMA_signal_11447) ) ;
    buf_clk new_AGEMA_reg_buffer_5599 ( .C (clk), .D (new_AGEMA_signal_11450), .Q (new_AGEMA_signal_11451) ) ;
    buf_clk new_AGEMA_reg_buffer_5603 ( .C (clk), .D (new_AGEMA_signal_11454), .Q (new_AGEMA_signal_11455) ) ;
    buf_clk new_AGEMA_reg_buffer_5607 ( .C (clk), .D (new_AGEMA_signal_11458), .Q (new_AGEMA_signal_11459) ) ;
    buf_clk new_AGEMA_reg_buffer_5611 ( .C (clk), .D (new_AGEMA_signal_11462), .Q (new_AGEMA_signal_11463) ) ;
    buf_clk new_AGEMA_reg_buffer_5615 ( .C (clk), .D (new_AGEMA_signal_11466), .Q (new_AGEMA_signal_11467) ) ;
    buf_clk new_AGEMA_reg_buffer_5619 ( .C (clk), .D (new_AGEMA_signal_11470), .Q (new_AGEMA_signal_11471) ) ;
    buf_clk new_AGEMA_reg_buffer_5623 ( .C (clk), .D (new_AGEMA_signal_11474), .Q (new_AGEMA_signal_11475) ) ;
    buf_clk new_AGEMA_reg_buffer_5627 ( .C (clk), .D (new_AGEMA_signal_11478), .Q (new_AGEMA_signal_11479) ) ;
    buf_clk new_AGEMA_reg_buffer_5631 ( .C (clk), .D (new_AGEMA_signal_11482), .Q (new_AGEMA_signal_11483) ) ;
    buf_clk new_AGEMA_reg_buffer_5635 ( .C (clk), .D (new_AGEMA_signal_11486), .Q (new_AGEMA_signal_11487) ) ;
    buf_clk new_AGEMA_reg_buffer_5639 ( .C (clk), .D (new_AGEMA_signal_11490), .Q (new_AGEMA_signal_11491) ) ;
    buf_clk new_AGEMA_reg_buffer_5643 ( .C (clk), .D (new_AGEMA_signal_11494), .Q (new_AGEMA_signal_11495) ) ;
    buf_clk new_AGEMA_reg_buffer_5647 ( .C (clk), .D (new_AGEMA_signal_11498), .Q (new_AGEMA_signal_11499) ) ;
    buf_clk new_AGEMA_reg_buffer_5651 ( .C (clk), .D (new_AGEMA_signal_11502), .Q (new_AGEMA_signal_11503) ) ;
    buf_clk new_AGEMA_reg_buffer_5655 ( .C (clk), .D (new_AGEMA_signal_11506), .Q (new_AGEMA_signal_11507) ) ;
    buf_clk new_AGEMA_reg_buffer_5659 ( .C (clk), .D (new_AGEMA_signal_11510), .Q (new_AGEMA_signal_11511) ) ;
    buf_clk new_AGEMA_reg_buffer_5663 ( .C (clk), .D (new_AGEMA_signal_11514), .Q (new_AGEMA_signal_11515) ) ;
    buf_clk new_AGEMA_reg_buffer_5667 ( .C (clk), .D (new_AGEMA_signal_11518), .Q (new_AGEMA_signal_11519) ) ;
    buf_clk new_AGEMA_reg_buffer_5671 ( .C (clk), .D (new_AGEMA_signal_11522), .Q (new_AGEMA_signal_11523) ) ;
    buf_clk new_AGEMA_reg_buffer_5675 ( .C (clk), .D (new_AGEMA_signal_11526), .Q (new_AGEMA_signal_11527) ) ;
    buf_clk new_AGEMA_reg_buffer_5679 ( .C (clk), .D (new_AGEMA_signal_11530), .Q (new_AGEMA_signal_11531) ) ;
    buf_clk new_AGEMA_reg_buffer_5683 ( .C (clk), .D (new_AGEMA_signal_11534), .Q (new_AGEMA_signal_11535) ) ;
    buf_clk new_AGEMA_reg_buffer_5687 ( .C (clk), .D (new_AGEMA_signal_11538), .Q (new_AGEMA_signal_11539) ) ;
    buf_clk new_AGEMA_reg_buffer_5691 ( .C (clk), .D (new_AGEMA_signal_11542), .Q (new_AGEMA_signal_11543) ) ;
    buf_clk new_AGEMA_reg_buffer_5695 ( .C (clk), .D (new_AGEMA_signal_11546), .Q (new_AGEMA_signal_11547) ) ;
    buf_clk new_AGEMA_reg_buffer_5699 ( .C (clk), .D (new_AGEMA_signal_11550), .Q (new_AGEMA_signal_11551) ) ;
    buf_clk new_AGEMA_reg_buffer_5703 ( .C (clk), .D (new_AGEMA_signal_11554), .Q (new_AGEMA_signal_11555) ) ;
    buf_clk new_AGEMA_reg_buffer_5707 ( .C (clk), .D (new_AGEMA_signal_11558), .Q (new_AGEMA_signal_11559) ) ;
    buf_clk new_AGEMA_reg_buffer_5711 ( .C (clk), .D (new_AGEMA_signal_11562), .Q (new_AGEMA_signal_11563) ) ;
    buf_clk new_AGEMA_reg_buffer_5715 ( .C (clk), .D (new_AGEMA_signal_11566), .Q (new_AGEMA_signal_11567) ) ;
    buf_clk new_AGEMA_reg_buffer_5719 ( .C (clk), .D (new_AGEMA_signal_11570), .Q (new_AGEMA_signal_11571) ) ;
    buf_clk new_AGEMA_reg_buffer_5723 ( .C (clk), .D (new_AGEMA_signal_11574), .Q (new_AGEMA_signal_11575) ) ;
    buf_clk new_AGEMA_reg_buffer_5727 ( .C (clk), .D (new_AGEMA_signal_11578), .Q (new_AGEMA_signal_11579) ) ;
    buf_clk new_AGEMA_reg_buffer_5731 ( .C (clk), .D (new_AGEMA_signal_11582), .Q (new_AGEMA_signal_11583) ) ;
    buf_clk new_AGEMA_reg_buffer_5735 ( .C (clk), .D (new_AGEMA_signal_11586), .Q (new_AGEMA_signal_11587) ) ;
    buf_clk new_AGEMA_reg_buffer_5739 ( .C (clk), .D (new_AGEMA_signal_11590), .Q (new_AGEMA_signal_11591) ) ;
    buf_clk new_AGEMA_reg_buffer_5743 ( .C (clk), .D (new_AGEMA_signal_11594), .Q (new_AGEMA_signal_11595) ) ;
    buf_clk new_AGEMA_reg_buffer_5747 ( .C (clk), .D (new_AGEMA_signal_11598), .Q (new_AGEMA_signal_11599) ) ;
    buf_clk new_AGEMA_reg_buffer_5750 ( .C (clk), .D (new_AGEMA_signal_11601), .Q (new_AGEMA_signal_11602) ) ;
    buf_clk new_AGEMA_reg_buffer_5753 ( .C (clk), .D (new_AGEMA_signal_11604), .Q (new_AGEMA_signal_11605) ) ;
    buf_clk new_AGEMA_reg_buffer_5756 ( .C (clk), .D (new_AGEMA_signal_11607), .Q (new_AGEMA_signal_11608) ) ;
    buf_clk new_AGEMA_reg_buffer_5759 ( .C (clk), .D (new_AGEMA_signal_11610), .Q (new_AGEMA_signal_11611) ) ;
    buf_clk new_AGEMA_reg_buffer_5762 ( .C (clk), .D (new_AGEMA_signal_11613), .Q (new_AGEMA_signal_11614) ) ;
    buf_clk new_AGEMA_reg_buffer_5765 ( .C (clk), .D (new_AGEMA_signal_11616), .Q (new_AGEMA_signal_11617) ) ;
    buf_clk new_AGEMA_reg_buffer_5768 ( .C (clk), .D (new_AGEMA_signal_11619), .Q (new_AGEMA_signal_11620) ) ;
    buf_clk new_AGEMA_reg_buffer_5771 ( .C (clk), .D (new_AGEMA_signal_11622), .Q (new_AGEMA_signal_11623) ) ;
    buf_clk new_AGEMA_reg_buffer_5774 ( .C (clk), .D (new_AGEMA_signal_11625), .Q (new_AGEMA_signal_11626) ) ;
    buf_clk new_AGEMA_reg_buffer_5777 ( .C (clk), .D (new_AGEMA_signal_11628), .Q (new_AGEMA_signal_11629) ) ;
    buf_clk new_AGEMA_reg_buffer_5780 ( .C (clk), .D (new_AGEMA_signal_11631), .Q (new_AGEMA_signal_11632) ) ;
    buf_clk new_AGEMA_reg_buffer_5783 ( .C (clk), .D (new_AGEMA_signal_11634), .Q (new_AGEMA_signal_11635) ) ;
    buf_clk new_AGEMA_reg_buffer_5786 ( .C (clk), .D (new_AGEMA_signal_11637), .Q (new_AGEMA_signal_11638) ) ;
    buf_clk new_AGEMA_reg_buffer_5789 ( .C (clk), .D (new_AGEMA_signal_11640), .Q (new_AGEMA_signal_11641) ) ;
    buf_clk new_AGEMA_reg_buffer_5792 ( .C (clk), .D (new_AGEMA_signal_11643), .Q (new_AGEMA_signal_11644) ) ;
    buf_clk new_AGEMA_reg_buffer_5795 ( .C (clk), .D (new_AGEMA_signal_11646), .Q (new_AGEMA_signal_11647) ) ;
    buf_clk new_AGEMA_reg_buffer_5798 ( .C (clk), .D (new_AGEMA_signal_11649), .Q (new_AGEMA_signal_11650) ) ;
    buf_clk new_AGEMA_reg_buffer_5801 ( .C (clk), .D (new_AGEMA_signal_11652), .Q (new_AGEMA_signal_11653) ) ;
    buf_clk new_AGEMA_reg_buffer_5804 ( .C (clk), .D (new_AGEMA_signal_11655), .Q (new_AGEMA_signal_11656) ) ;
    buf_clk new_AGEMA_reg_buffer_5807 ( .C (clk), .D (new_AGEMA_signal_11658), .Q (new_AGEMA_signal_11659) ) ;
    buf_clk new_AGEMA_reg_buffer_5810 ( .C (clk), .D (new_AGEMA_signal_11661), .Q (new_AGEMA_signal_11662) ) ;
    buf_clk new_AGEMA_reg_buffer_5813 ( .C (clk), .D (new_AGEMA_signal_11664), .Q (new_AGEMA_signal_11665) ) ;
    buf_clk new_AGEMA_reg_buffer_5816 ( .C (clk), .D (new_AGEMA_signal_11667), .Q (new_AGEMA_signal_11668) ) ;
    buf_clk new_AGEMA_reg_buffer_5819 ( .C (clk), .D (new_AGEMA_signal_11670), .Q (new_AGEMA_signal_11671) ) ;
    buf_clk new_AGEMA_reg_buffer_5822 ( .C (clk), .D (new_AGEMA_signal_11673), .Q (new_AGEMA_signal_11674) ) ;
    buf_clk new_AGEMA_reg_buffer_5825 ( .C (clk), .D (new_AGEMA_signal_11676), .Q (new_AGEMA_signal_11677) ) ;
    buf_clk new_AGEMA_reg_buffer_5828 ( .C (clk), .D (new_AGEMA_signal_11679), .Q (new_AGEMA_signal_11680) ) ;
    buf_clk new_AGEMA_reg_buffer_5831 ( .C (clk), .D (new_AGEMA_signal_11682), .Q (new_AGEMA_signal_11683) ) ;
    buf_clk new_AGEMA_reg_buffer_5834 ( .C (clk), .D (new_AGEMA_signal_11685), .Q (new_AGEMA_signal_11686) ) ;
    buf_clk new_AGEMA_reg_buffer_5837 ( .C (clk), .D (new_AGEMA_signal_11688), .Q (new_AGEMA_signal_11689) ) ;
    buf_clk new_AGEMA_reg_buffer_5840 ( .C (clk), .D (new_AGEMA_signal_11691), .Q (new_AGEMA_signal_11692) ) ;
    buf_clk new_AGEMA_reg_buffer_5843 ( .C (clk), .D (new_AGEMA_signal_11694), .Q (new_AGEMA_signal_11695) ) ;
    buf_clk new_AGEMA_reg_buffer_5846 ( .C (clk), .D (new_AGEMA_signal_11697), .Q (new_AGEMA_signal_11698) ) ;
    buf_clk new_AGEMA_reg_buffer_5849 ( .C (clk), .D (new_AGEMA_signal_11700), .Q (new_AGEMA_signal_11701) ) ;
    buf_clk new_AGEMA_reg_buffer_5852 ( .C (clk), .D (new_AGEMA_signal_11703), .Q (new_AGEMA_signal_11704) ) ;
    buf_clk new_AGEMA_reg_buffer_5855 ( .C (clk), .D (new_AGEMA_signal_11706), .Q (new_AGEMA_signal_11707) ) ;
    buf_clk new_AGEMA_reg_buffer_5858 ( .C (clk), .D (new_AGEMA_signal_11709), .Q (new_AGEMA_signal_11710) ) ;
    buf_clk new_AGEMA_reg_buffer_5861 ( .C (clk), .D (new_AGEMA_signal_11712), .Q (new_AGEMA_signal_11713) ) ;
    buf_clk new_AGEMA_reg_buffer_5864 ( .C (clk), .D (new_AGEMA_signal_11715), .Q (new_AGEMA_signal_11716) ) ;
    buf_clk new_AGEMA_reg_buffer_5867 ( .C (clk), .D (new_AGEMA_signal_11718), .Q (new_AGEMA_signal_11719) ) ;
    buf_clk new_AGEMA_reg_buffer_5870 ( .C (clk), .D (new_AGEMA_signal_11721), .Q (new_AGEMA_signal_11722) ) ;
    buf_clk new_AGEMA_reg_buffer_5873 ( .C (clk), .D (new_AGEMA_signal_11724), .Q (new_AGEMA_signal_11725) ) ;
    buf_clk new_AGEMA_reg_buffer_5876 ( .C (clk), .D (new_AGEMA_signal_11727), .Q (new_AGEMA_signal_11728) ) ;
    buf_clk new_AGEMA_reg_buffer_5879 ( .C (clk), .D (new_AGEMA_signal_11730), .Q (new_AGEMA_signal_11731) ) ;
    buf_clk new_AGEMA_reg_buffer_5882 ( .C (clk), .D (new_AGEMA_signal_11733), .Q (new_AGEMA_signal_11734) ) ;
    buf_clk new_AGEMA_reg_buffer_5885 ( .C (clk), .D (new_AGEMA_signal_11736), .Q (new_AGEMA_signal_11737) ) ;
    buf_clk new_AGEMA_reg_buffer_5888 ( .C (clk), .D (new_AGEMA_signal_11739), .Q (new_AGEMA_signal_11740) ) ;
    buf_clk new_AGEMA_reg_buffer_5891 ( .C (clk), .D (new_AGEMA_signal_11742), .Q (new_AGEMA_signal_11743) ) ;
    buf_clk new_AGEMA_reg_buffer_5894 ( .C (clk), .D (new_AGEMA_signal_11745), .Q (new_AGEMA_signal_11746) ) ;
    buf_clk new_AGEMA_reg_buffer_5897 ( .C (clk), .D (new_AGEMA_signal_11748), .Q (new_AGEMA_signal_11749) ) ;
    buf_clk new_AGEMA_reg_buffer_5900 ( .C (clk), .D (new_AGEMA_signal_11751), .Q (new_AGEMA_signal_11752) ) ;
    buf_clk new_AGEMA_reg_buffer_5903 ( .C (clk), .D (new_AGEMA_signal_11754), .Q (new_AGEMA_signal_11755) ) ;
    buf_clk new_AGEMA_reg_buffer_5906 ( .C (clk), .D (new_AGEMA_signal_11757), .Q (new_AGEMA_signal_11758) ) ;
    buf_clk new_AGEMA_reg_buffer_5909 ( .C (clk), .D (new_AGEMA_signal_11760), .Q (new_AGEMA_signal_11761) ) ;
    buf_clk new_AGEMA_reg_buffer_5912 ( .C (clk), .D (new_AGEMA_signal_11763), .Q (new_AGEMA_signal_11764) ) ;
    buf_clk new_AGEMA_reg_buffer_5915 ( .C (clk), .D (new_AGEMA_signal_11766), .Q (new_AGEMA_signal_11767) ) ;
    buf_clk new_AGEMA_reg_buffer_5918 ( .C (clk), .D (new_AGEMA_signal_11769), .Q (new_AGEMA_signal_11770) ) ;
    buf_clk new_AGEMA_reg_buffer_5921 ( .C (clk), .D (new_AGEMA_signal_11772), .Q (new_AGEMA_signal_11773) ) ;
    buf_clk new_AGEMA_reg_buffer_5924 ( .C (clk), .D (new_AGEMA_signal_11775), .Q (new_AGEMA_signal_11776) ) ;
    buf_clk new_AGEMA_reg_buffer_5927 ( .C (clk), .D (new_AGEMA_signal_11778), .Q (new_AGEMA_signal_11779) ) ;
    buf_clk new_AGEMA_reg_buffer_5930 ( .C (clk), .D (new_AGEMA_signal_11781), .Q (new_AGEMA_signal_11782) ) ;
    buf_clk new_AGEMA_reg_buffer_5933 ( .C (clk), .D (new_AGEMA_signal_11784), .Q (new_AGEMA_signal_11785) ) ;
    buf_clk new_AGEMA_reg_buffer_5936 ( .C (clk), .D (new_AGEMA_signal_11787), .Q (new_AGEMA_signal_11788) ) ;
    buf_clk new_AGEMA_reg_buffer_5939 ( .C (clk), .D (new_AGEMA_signal_11790), .Q (new_AGEMA_signal_11791) ) ;
    buf_clk new_AGEMA_reg_buffer_5942 ( .C (clk), .D (new_AGEMA_signal_11793), .Q (new_AGEMA_signal_11794) ) ;
    buf_clk new_AGEMA_reg_buffer_5945 ( .C (clk), .D (new_AGEMA_signal_11796), .Q (new_AGEMA_signal_11797) ) ;
    buf_clk new_AGEMA_reg_buffer_5948 ( .C (clk), .D (new_AGEMA_signal_11799), .Q (new_AGEMA_signal_11800) ) ;
    buf_clk new_AGEMA_reg_buffer_5951 ( .C (clk), .D (new_AGEMA_signal_11802), .Q (new_AGEMA_signal_11803) ) ;
    buf_clk new_AGEMA_reg_buffer_5954 ( .C (clk), .D (new_AGEMA_signal_11805), .Q (new_AGEMA_signal_11806) ) ;
    buf_clk new_AGEMA_reg_buffer_5957 ( .C (clk), .D (new_AGEMA_signal_11808), .Q (new_AGEMA_signal_11809) ) ;
    buf_clk new_AGEMA_reg_buffer_5960 ( .C (clk), .D (new_AGEMA_signal_11811), .Q (new_AGEMA_signal_11812) ) ;
    buf_clk new_AGEMA_reg_buffer_5963 ( .C (clk), .D (new_AGEMA_signal_11814), .Q (new_AGEMA_signal_11815) ) ;
    buf_clk new_AGEMA_reg_buffer_5966 ( .C (clk), .D (new_AGEMA_signal_11817), .Q (new_AGEMA_signal_11818) ) ;
    buf_clk new_AGEMA_reg_buffer_5969 ( .C (clk), .D (new_AGEMA_signal_11820), .Q (new_AGEMA_signal_11821) ) ;
    buf_clk new_AGEMA_reg_buffer_5972 ( .C (clk), .D (new_AGEMA_signal_11823), .Q (new_AGEMA_signal_11824) ) ;
    buf_clk new_AGEMA_reg_buffer_5975 ( .C (clk), .D (new_AGEMA_signal_11826), .Q (new_AGEMA_signal_11827) ) ;
    buf_clk new_AGEMA_reg_buffer_5978 ( .C (clk), .D (new_AGEMA_signal_11829), .Q (new_AGEMA_signal_11830) ) ;
    buf_clk new_AGEMA_reg_buffer_5981 ( .C (clk), .D (new_AGEMA_signal_11832), .Q (new_AGEMA_signal_11833) ) ;
    buf_clk new_AGEMA_reg_buffer_5984 ( .C (clk), .D (new_AGEMA_signal_11835), .Q (new_AGEMA_signal_11836) ) ;
    buf_clk new_AGEMA_reg_buffer_5987 ( .C (clk), .D (new_AGEMA_signal_11838), .Q (new_AGEMA_signal_11839) ) ;
    buf_clk new_AGEMA_reg_buffer_5990 ( .C (clk), .D (new_AGEMA_signal_11841), .Q (new_AGEMA_signal_11842) ) ;
    buf_clk new_AGEMA_reg_buffer_5993 ( .C (clk), .D (new_AGEMA_signal_11844), .Q (new_AGEMA_signal_11845) ) ;
    buf_clk new_AGEMA_reg_buffer_5996 ( .C (clk), .D (new_AGEMA_signal_11847), .Q (new_AGEMA_signal_11848) ) ;
    buf_clk new_AGEMA_reg_buffer_5999 ( .C (clk), .D (new_AGEMA_signal_11850), .Q (new_AGEMA_signal_11851) ) ;
    buf_clk new_AGEMA_reg_buffer_6002 ( .C (clk), .D (new_AGEMA_signal_11853), .Q (new_AGEMA_signal_11854) ) ;
    buf_clk new_AGEMA_reg_buffer_6005 ( .C (clk), .D (new_AGEMA_signal_11856), .Q (new_AGEMA_signal_11857) ) ;
    buf_clk new_AGEMA_reg_buffer_6008 ( .C (clk), .D (new_AGEMA_signal_11859), .Q (new_AGEMA_signal_11860) ) ;
    buf_clk new_AGEMA_reg_buffer_6011 ( .C (clk), .D (new_AGEMA_signal_11862), .Q (new_AGEMA_signal_11863) ) ;
    buf_clk new_AGEMA_reg_buffer_6014 ( .C (clk), .D (new_AGEMA_signal_11865), .Q (new_AGEMA_signal_11866) ) ;
    buf_clk new_AGEMA_reg_buffer_6017 ( .C (clk), .D (new_AGEMA_signal_11868), .Q (new_AGEMA_signal_11869) ) ;
    buf_clk new_AGEMA_reg_buffer_6020 ( .C (clk), .D (new_AGEMA_signal_11871), .Q (new_AGEMA_signal_11872) ) ;
    buf_clk new_AGEMA_reg_buffer_6023 ( .C (clk), .D (new_AGEMA_signal_11874), .Q (new_AGEMA_signal_11875) ) ;
    buf_clk new_AGEMA_reg_buffer_6026 ( .C (clk), .D (new_AGEMA_signal_11877), .Q (new_AGEMA_signal_11878) ) ;
    buf_clk new_AGEMA_reg_buffer_6029 ( .C (clk), .D (new_AGEMA_signal_11880), .Q (new_AGEMA_signal_11881) ) ;
    buf_clk new_AGEMA_reg_buffer_6032 ( .C (clk), .D (new_AGEMA_signal_11883), .Q (new_AGEMA_signal_11884) ) ;
    buf_clk new_AGEMA_reg_buffer_6035 ( .C (clk), .D (new_AGEMA_signal_11886), .Q (new_AGEMA_signal_11887) ) ;
    buf_clk new_AGEMA_reg_buffer_6038 ( .C (clk), .D (new_AGEMA_signal_11889), .Q (new_AGEMA_signal_11890) ) ;
    buf_clk new_AGEMA_reg_buffer_6041 ( .C (clk), .D (new_AGEMA_signal_11892), .Q (new_AGEMA_signal_11893) ) ;
    buf_clk new_AGEMA_reg_buffer_6044 ( .C (clk), .D (new_AGEMA_signal_11895), .Q (new_AGEMA_signal_11896) ) ;
    buf_clk new_AGEMA_reg_buffer_6047 ( .C (clk), .D (new_AGEMA_signal_11898), .Q (new_AGEMA_signal_11899) ) ;
    buf_clk new_AGEMA_reg_buffer_6050 ( .C (clk), .D (new_AGEMA_signal_11901), .Q (new_AGEMA_signal_11902) ) ;
    buf_clk new_AGEMA_reg_buffer_6053 ( .C (clk), .D (new_AGEMA_signal_11904), .Q (new_AGEMA_signal_11905) ) ;
    buf_clk new_AGEMA_reg_buffer_6056 ( .C (clk), .D (new_AGEMA_signal_11907), .Q (new_AGEMA_signal_11908) ) ;
    buf_clk new_AGEMA_reg_buffer_6059 ( .C (clk), .D (new_AGEMA_signal_11910), .Q (new_AGEMA_signal_11911) ) ;
    buf_clk new_AGEMA_reg_buffer_6062 ( .C (clk), .D (new_AGEMA_signal_11913), .Q (new_AGEMA_signal_11914) ) ;
    buf_clk new_AGEMA_reg_buffer_6065 ( .C (clk), .D (new_AGEMA_signal_11916), .Q (new_AGEMA_signal_11917) ) ;
    buf_clk new_AGEMA_reg_buffer_6068 ( .C (clk), .D (new_AGEMA_signal_11919), .Q (new_AGEMA_signal_11920) ) ;
    buf_clk new_AGEMA_reg_buffer_6071 ( .C (clk), .D (new_AGEMA_signal_11922), .Q (new_AGEMA_signal_11923) ) ;
    buf_clk new_AGEMA_reg_buffer_6074 ( .C (clk), .D (new_AGEMA_signal_11925), .Q (new_AGEMA_signal_11926) ) ;
    buf_clk new_AGEMA_reg_buffer_6077 ( .C (clk), .D (new_AGEMA_signal_11928), .Q (new_AGEMA_signal_11929) ) ;
    buf_clk new_AGEMA_reg_buffer_6080 ( .C (clk), .D (new_AGEMA_signal_11931), .Q (new_AGEMA_signal_11932) ) ;
    buf_clk new_AGEMA_reg_buffer_6083 ( .C (clk), .D (new_AGEMA_signal_11934), .Q (new_AGEMA_signal_11935) ) ;
    buf_clk new_AGEMA_reg_buffer_6086 ( .C (clk), .D (new_AGEMA_signal_11937), .Q (new_AGEMA_signal_11938) ) ;
    buf_clk new_AGEMA_reg_buffer_6089 ( .C (clk), .D (new_AGEMA_signal_11940), .Q (new_AGEMA_signal_11941) ) ;
    buf_clk new_AGEMA_reg_buffer_6092 ( .C (clk), .D (new_AGEMA_signal_11943), .Q (new_AGEMA_signal_11944) ) ;
    buf_clk new_AGEMA_reg_buffer_6095 ( .C (clk), .D (new_AGEMA_signal_11946), .Q (new_AGEMA_signal_11947) ) ;
    buf_clk new_AGEMA_reg_buffer_6098 ( .C (clk), .D (new_AGEMA_signal_11949), .Q (new_AGEMA_signal_11950) ) ;
    buf_clk new_AGEMA_reg_buffer_6101 ( .C (clk), .D (new_AGEMA_signal_11952), .Q (new_AGEMA_signal_11953) ) ;
    buf_clk new_AGEMA_reg_buffer_6104 ( .C (clk), .D (new_AGEMA_signal_11955), .Q (new_AGEMA_signal_11956) ) ;
    buf_clk new_AGEMA_reg_buffer_6107 ( .C (clk), .D (new_AGEMA_signal_11958), .Q (new_AGEMA_signal_11959) ) ;
    buf_clk new_AGEMA_reg_buffer_6110 ( .C (clk), .D (new_AGEMA_signal_11961), .Q (new_AGEMA_signal_11962) ) ;
    buf_clk new_AGEMA_reg_buffer_6113 ( .C (clk), .D (new_AGEMA_signal_11964), .Q (new_AGEMA_signal_11965) ) ;
    buf_clk new_AGEMA_reg_buffer_6116 ( .C (clk), .D (new_AGEMA_signal_11967), .Q (new_AGEMA_signal_11968) ) ;
    buf_clk new_AGEMA_reg_buffer_6119 ( .C (clk), .D (new_AGEMA_signal_11970), .Q (new_AGEMA_signal_11971) ) ;
    buf_clk new_AGEMA_reg_buffer_6122 ( .C (clk), .D (new_AGEMA_signal_11973), .Q (new_AGEMA_signal_11974) ) ;
    buf_clk new_AGEMA_reg_buffer_6125 ( .C (clk), .D (new_AGEMA_signal_11976), .Q (new_AGEMA_signal_11977) ) ;
    buf_clk new_AGEMA_reg_buffer_6128 ( .C (clk), .D (new_AGEMA_signal_11979), .Q (new_AGEMA_signal_11980) ) ;
    buf_clk new_AGEMA_reg_buffer_6131 ( .C (clk), .D (new_AGEMA_signal_11982), .Q (new_AGEMA_signal_11983) ) ;
    buf_clk new_AGEMA_reg_buffer_6134 ( .C (clk), .D (new_AGEMA_signal_11985), .Q (new_AGEMA_signal_11986) ) ;
    buf_clk new_AGEMA_reg_buffer_6137 ( .C (clk), .D (new_AGEMA_signal_11988), .Q (new_AGEMA_signal_11989) ) ;
    buf_clk new_AGEMA_reg_buffer_6140 ( .C (clk), .D (new_AGEMA_signal_11991), .Q (new_AGEMA_signal_11992) ) ;
    buf_clk new_AGEMA_reg_buffer_6143 ( .C (clk), .D (new_AGEMA_signal_11994), .Q (new_AGEMA_signal_11995) ) ;
    buf_clk new_AGEMA_reg_buffer_6146 ( .C (clk), .D (new_AGEMA_signal_11997), .Q (new_AGEMA_signal_11998) ) ;
    buf_clk new_AGEMA_reg_buffer_6149 ( .C (clk), .D (new_AGEMA_signal_12000), .Q (new_AGEMA_signal_12001) ) ;
    buf_clk new_AGEMA_reg_buffer_6152 ( .C (clk), .D (new_AGEMA_signal_12003), .Q (new_AGEMA_signal_12004) ) ;
    buf_clk new_AGEMA_reg_buffer_6155 ( .C (clk), .D (new_AGEMA_signal_12006), .Q (new_AGEMA_signal_12007) ) ;
    buf_clk new_AGEMA_reg_buffer_6158 ( .C (clk), .D (new_AGEMA_signal_12009), .Q (new_AGEMA_signal_12010) ) ;
    buf_clk new_AGEMA_reg_buffer_6161 ( .C (clk), .D (new_AGEMA_signal_12012), .Q (new_AGEMA_signal_12013) ) ;
    buf_clk new_AGEMA_reg_buffer_6164 ( .C (clk), .D (new_AGEMA_signal_12015), .Q (new_AGEMA_signal_12016) ) ;
    buf_clk new_AGEMA_reg_buffer_6167 ( .C (clk), .D (new_AGEMA_signal_12018), .Q (new_AGEMA_signal_12019) ) ;
    buf_clk new_AGEMA_reg_buffer_6170 ( .C (clk), .D (new_AGEMA_signal_12021), .Q (new_AGEMA_signal_12022) ) ;
    buf_clk new_AGEMA_reg_buffer_6173 ( .C (clk), .D (new_AGEMA_signal_12024), .Q (new_AGEMA_signal_12025) ) ;
    buf_clk new_AGEMA_reg_buffer_6176 ( .C (clk), .D (new_AGEMA_signal_12027), .Q (new_AGEMA_signal_12028) ) ;
    buf_clk new_AGEMA_reg_buffer_6179 ( .C (clk), .D (new_AGEMA_signal_12030), .Q (new_AGEMA_signal_12031) ) ;
    buf_clk new_AGEMA_reg_buffer_6182 ( .C (clk), .D (new_AGEMA_signal_12033), .Q (new_AGEMA_signal_12034) ) ;
    buf_clk new_AGEMA_reg_buffer_6185 ( .C (clk), .D (new_AGEMA_signal_12036), .Q (new_AGEMA_signal_12037) ) ;
    buf_clk new_AGEMA_reg_buffer_6188 ( .C (clk), .D (new_AGEMA_signal_12039), .Q (new_AGEMA_signal_12040) ) ;
    buf_clk new_AGEMA_reg_buffer_6191 ( .C (clk), .D (new_AGEMA_signal_12042), .Q (new_AGEMA_signal_12043) ) ;
    buf_clk new_AGEMA_reg_buffer_6194 ( .C (clk), .D (new_AGEMA_signal_12045), .Q (new_AGEMA_signal_12046) ) ;
    buf_clk new_AGEMA_reg_buffer_6197 ( .C (clk), .D (new_AGEMA_signal_12048), .Q (new_AGEMA_signal_12049) ) ;
    buf_clk new_AGEMA_reg_buffer_6200 ( .C (clk), .D (new_AGEMA_signal_12051), .Q (new_AGEMA_signal_12052) ) ;
    buf_clk new_AGEMA_reg_buffer_6203 ( .C (clk), .D (new_AGEMA_signal_12054), .Q (new_AGEMA_signal_12055) ) ;
    buf_clk new_AGEMA_reg_buffer_6206 ( .C (clk), .D (new_AGEMA_signal_12057), .Q (new_AGEMA_signal_12058) ) ;
    buf_clk new_AGEMA_reg_buffer_6209 ( .C (clk), .D (new_AGEMA_signal_12060), .Q (new_AGEMA_signal_12061) ) ;
    buf_clk new_AGEMA_reg_buffer_6212 ( .C (clk), .D (new_AGEMA_signal_12063), .Q (new_AGEMA_signal_12064) ) ;
    buf_clk new_AGEMA_reg_buffer_6215 ( .C (clk), .D (new_AGEMA_signal_12066), .Q (new_AGEMA_signal_12067) ) ;
    buf_clk new_AGEMA_reg_buffer_6218 ( .C (clk), .D (new_AGEMA_signal_12069), .Q (new_AGEMA_signal_12070) ) ;
    buf_clk new_AGEMA_reg_buffer_6221 ( .C (clk), .D (new_AGEMA_signal_12072), .Q (new_AGEMA_signal_12073) ) ;
    buf_clk new_AGEMA_reg_buffer_6224 ( .C (clk), .D (new_AGEMA_signal_12075), .Q (new_AGEMA_signal_12076) ) ;
    buf_clk new_AGEMA_reg_buffer_6227 ( .C (clk), .D (new_AGEMA_signal_12078), .Q (new_AGEMA_signal_12079) ) ;
    buf_clk new_AGEMA_reg_buffer_6230 ( .C (clk), .D (new_AGEMA_signal_12081), .Q (new_AGEMA_signal_12082) ) ;
    buf_clk new_AGEMA_reg_buffer_6233 ( .C (clk), .D (new_AGEMA_signal_12084), .Q (new_AGEMA_signal_12085) ) ;
    buf_clk new_AGEMA_reg_buffer_6236 ( .C (clk), .D (new_AGEMA_signal_12087), .Q (new_AGEMA_signal_12088) ) ;
    buf_clk new_AGEMA_reg_buffer_6239 ( .C (clk), .D (new_AGEMA_signal_12090), .Q (new_AGEMA_signal_12091) ) ;
    buf_clk new_AGEMA_reg_buffer_6242 ( .C (clk), .D (new_AGEMA_signal_12093), .Q (new_AGEMA_signal_12094) ) ;
    buf_clk new_AGEMA_reg_buffer_6245 ( .C (clk), .D (new_AGEMA_signal_12096), .Q (new_AGEMA_signal_12097) ) ;
    buf_clk new_AGEMA_reg_buffer_6248 ( .C (clk), .D (new_AGEMA_signal_12099), .Q (new_AGEMA_signal_12100) ) ;
    buf_clk new_AGEMA_reg_buffer_6251 ( .C (clk), .D (new_AGEMA_signal_12102), .Q (new_AGEMA_signal_12103) ) ;
    buf_clk new_AGEMA_reg_buffer_6254 ( .C (clk), .D (new_AGEMA_signal_12105), .Q (new_AGEMA_signal_12106) ) ;
    buf_clk new_AGEMA_reg_buffer_6257 ( .C (clk), .D (new_AGEMA_signal_12108), .Q (new_AGEMA_signal_12109) ) ;
    buf_clk new_AGEMA_reg_buffer_6260 ( .C (clk), .D (new_AGEMA_signal_12111), .Q (new_AGEMA_signal_12112) ) ;
    buf_clk new_AGEMA_reg_buffer_6263 ( .C (clk), .D (new_AGEMA_signal_12114), .Q (new_AGEMA_signal_12115) ) ;
    buf_clk new_AGEMA_reg_buffer_6266 ( .C (clk), .D (new_AGEMA_signal_12117), .Q (new_AGEMA_signal_12118) ) ;
    buf_clk new_AGEMA_reg_buffer_6269 ( .C (clk), .D (new_AGEMA_signal_12120), .Q (new_AGEMA_signal_12121) ) ;
    buf_clk new_AGEMA_reg_buffer_6272 ( .C (clk), .D (new_AGEMA_signal_12123), .Q (new_AGEMA_signal_12124) ) ;
    buf_clk new_AGEMA_reg_buffer_6275 ( .C (clk), .D (new_AGEMA_signal_12126), .Q (new_AGEMA_signal_12127) ) ;
    buf_clk new_AGEMA_reg_buffer_6278 ( .C (clk), .D (new_AGEMA_signal_12129), .Q (new_AGEMA_signal_12130) ) ;
    buf_clk new_AGEMA_reg_buffer_6281 ( .C (clk), .D (new_AGEMA_signal_12132), .Q (new_AGEMA_signal_12133) ) ;
    buf_clk new_AGEMA_reg_buffer_6284 ( .C (clk), .D (new_AGEMA_signal_12135), .Q (new_AGEMA_signal_12136) ) ;
    buf_clk new_AGEMA_reg_buffer_6287 ( .C (clk), .D (new_AGEMA_signal_12138), .Q (new_AGEMA_signal_12139) ) ;
    buf_clk new_AGEMA_reg_buffer_6290 ( .C (clk), .D (new_AGEMA_signal_12141), .Q (new_AGEMA_signal_12142) ) ;
    buf_clk new_AGEMA_reg_buffer_6293 ( .C (clk), .D (new_AGEMA_signal_12144), .Q (new_AGEMA_signal_12145) ) ;
    buf_clk new_AGEMA_reg_buffer_6296 ( .C (clk), .D (new_AGEMA_signal_12147), .Q (new_AGEMA_signal_12148) ) ;
    buf_clk new_AGEMA_reg_buffer_6299 ( .C (clk), .D (new_AGEMA_signal_12150), .Q (new_AGEMA_signal_12151) ) ;
    buf_clk new_AGEMA_reg_buffer_6302 ( .C (clk), .D (new_AGEMA_signal_12153), .Q (new_AGEMA_signal_12154) ) ;
    buf_clk new_AGEMA_reg_buffer_6305 ( .C (clk), .D (new_AGEMA_signal_12156), .Q (new_AGEMA_signal_12157) ) ;
    buf_clk new_AGEMA_reg_buffer_6308 ( .C (clk), .D (new_AGEMA_signal_12159), .Q (new_AGEMA_signal_12160) ) ;
    buf_clk new_AGEMA_reg_buffer_6311 ( .C (clk), .D (new_AGEMA_signal_12162), .Q (new_AGEMA_signal_12163) ) ;
    buf_clk new_AGEMA_reg_buffer_6314 ( .C (clk), .D (new_AGEMA_signal_12165), .Q (new_AGEMA_signal_12166) ) ;
    buf_clk new_AGEMA_reg_buffer_6317 ( .C (clk), .D (new_AGEMA_signal_12168), .Q (new_AGEMA_signal_12169) ) ;
    buf_clk new_AGEMA_reg_buffer_6320 ( .C (clk), .D (new_AGEMA_signal_12171), .Q (new_AGEMA_signal_12172) ) ;
    buf_clk new_AGEMA_reg_buffer_6323 ( .C (clk), .D (new_AGEMA_signal_12174), .Q (new_AGEMA_signal_12175) ) ;
    buf_clk new_AGEMA_reg_buffer_6326 ( .C (clk), .D (new_AGEMA_signal_12177), .Q (new_AGEMA_signal_12178) ) ;
    buf_clk new_AGEMA_reg_buffer_6329 ( .C (clk), .D (new_AGEMA_signal_12180), .Q (new_AGEMA_signal_12181) ) ;
    buf_clk new_AGEMA_reg_buffer_6332 ( .C (clk), .D (new_AGEMA_signal_12183), .Q (new_AGEMA_signal_12184) ) ;
    buf_clk new_AGEMA_reg_buffer_6335 ( .C (clk), .D (new_AGEMA_signal_12186), .Q (new_AGEMA_signal_12187) ) ;
    buf_clk new_AGEMA_reg_buffer_6338 ( .C (clk), .D (new_AGEMA_signal_12189), .Q (new_AGEMA_signal_12190) ) ;
    buf_clk new_AGEMA_reg_buffer_6341 ( .C (clk), .D (new_AGEMA_signal_12192), .Q (new_AGEMA_signal_12193) ) ;
    buf_clk new_AGEMA_reg_buffer_6344 ( .C (clk), .D (new_AGEMA_signal_12195), .Q (new_AGEMA_signal_12196) ) ;
    buf_clk new_AGEMA_reg_buffer_6347 ( .C (clk), .D (new_AGEMA_signal_12198), .Q (new_AGEMA_signal_12199) ) ;
    buf_clk new_AGEMA_reg_buffer_6350 ( .C (clk), .D (new_AGEMA_signal_12201), .Q (new_AGEMA_signal_12202) ) ;
    buf_clk new_AGEMA_reg_buffer_6353 ( .C (clk), .D (new_AGEMA_signal_12204), .Q (new_AGEMA_signal_12205) ) ;
    buf_clk new_AGEMA_reg_buffer_6356 ( .C (clk), .D (new_AGEMA_signal_12207), .Q (new_AGEMA_signal_12208) ) ;
    buf_clk new_AGEMA_reg_buffer_6359 ( .C (clk), .D (new_AGEMA_signal_12210), .Q (new_AGEMA_signal_12211) ) ;
    buf_clk new_AGEMA_reg_buffer_6362 ( .C (clk), .D (new_AGEMA_signal_12213), .Q (new_AGEMA_signal_12214) ) ;
    buf_clk new_AGEMA_reg_buffer_6365 ( .C (clk), .D (new_AGEMA_signal_12216), .Q (new_AGEMA_signal_12217) ) ;
    buf_clk new_AGEMA_reg_buffer_6368 ( .C (clk), .D (new_AGEMA_signal_12219), .Q (new_AGEMA_signal_12220) ) ;
    buf_clk new_AGEMA_reg_buffer_6371 ( .C (clk), .D (new_AGEMA_signal_12222), .Q (new_AGEMA_signal_12223) ) ;
    buf_clk new_AGEMA_reg_buffer_6374 ( .C (clk), .D (new_AGEMA_signal_12225), .Q (new_AGEMA_signal_12226) ) ;
    buf_clk new_AGEMA_reg_buffer_6377 ( .C (clk), .D (new_AGEMA_signal_12228), .Q (new_AGEMA_signal_12229) ) ;
    buf_clk new_AGEMA_reg_buffer_6380 ( .C (clk), .D (new_AGEMA_signal_12231), .Q (new_AGEMA_signal_12232) ) ;
    buf_clk new_AGEMA_reg_buffer_6383 ( .C (clk), .D (new_AGEMA_signal_12234), .Q (new_AGEMA_signal_12235) ) ;
    buf_clk new_AGEMA_reg_buffer_6386 ( .C (clk), .D (new_AGEMA_signal_12237), .Q (new_AGEMA_signal_12238) ) ;
    buf_clk new_AGEMA_reg_buffer_6389 ( .C (clk), .D (new_AGEMA_signal_12240), .Q (new_AGEMA_signal_12241) ) ;
    buf_clk new_AGEMA_reg_buffer_6392 ( .C (clk), .D (new_AGEMA_signal_12243), .Q (new_AGEMA_signal_12244) ) ;
    buf_clk new_AGEMA_reg_buffer_6395 ( .C (clk), .D (new_AGEMA_signal_12246), .Q (new_AGEMA_signal_12247) ) ;
    buf_clk new_AGEMA_reg_buffer_6398 ( .C (clk), .D (new_AGEMA_signal_12249), .Q (new_AGEMA_signal_12250) ) ;
    buf_clk new_AGEMA_reg_buffer_6401 ( .C (clk), .D (new_AGEMA_signal_12252), .Q (new_AGEMA_signal_12253) ) ;
    buf_clk new_AGEMA_reg_buffer_6404 ( .C (clk), .D (new_AGEMA_signal_12255), .Q (new_AGEMA_signal_12256) ) ;
    buf_clk new_AGEMA_reg_buffer_6407 ( .C (clk), .D (new_AGEMA_signal_12258), .Q (new_AGEMA_signal_12259) ) ;
    buf_clk new_AGEMA_reg_buffer_6410 ( .C (clk), .D (new_AGEMA_signal_12261), .Q (new_AGEMA_signal_12262) ) ;
    buf_clk new_AGEMA_reg_buffer_6413 ( .C (clk), .D (new_AGEMA_signal_12264), .Q (new_AGEMA_signal_12265) ) ;
    buf_clk new_AGEMA_reg_buffer_6416 ( .C (clk), .D (new_AGEMA_signal_12267), .Q (new_AGEMA_signal_12268) ) ;
    buf_clk new_AGEMA_reg_buffer_6419 ( .C (clk), .D (new_AGEMA_signal_12270), .Q (new_AGEMA_signal_12271) ) ;
    buf_clk new_AGEMA_reg_buffer_6422 ( .C (clk), .D (new_AGEMA_signal_12273), .Q (new_AGEMA_signal_12274) ) ;
    buf_clk new_AGEMA_reg_buffer_6425 ( .C (clk), .D (new_AGEMA_signal_12276), .Q (new_AGEMA_signal_12277) ) ;
    buf_clk new_AGEMA_reg_buffer_6428 ( .C (clk), .D (new_AGEMA_signal_12279), .Q (new_AGEMA_signal_12280) ) ;
    buf_clk new_AGEMA_reg_buffer_6431 ( .C (clk), .D (new_AGEMA_signal_12282), .Q (new_AGEMA_signal_12283) ) ;
    buf_clk new_AGEMA_reg_buffer_6434 ( .C (clk), .D (new_AGEMA_signal_12285), .Q (new_AGEMA_signal_12286) ) ;
    buf_clk new_AGEMA_reg_buffer_6437 ( .C (clk), .D (new_AGEMA_signal_12288), .Q (new_AGEMA_signal_12289) ) ;
    buf_clk new_AGEMA_reg_buffer_6440 ( .C (clk), .D (new_AGEMA_signal_12291), .Q (new_AGEMA_signal_12292) ) ;
    buf_clk new_AGEMA_reg_buffer_6443 ( .C (clk), .D (new_AGEMA_signal_12294), .Q (new_AGEMA_signal_12295) ) ;
    buf_clk new_AGEMA_reg_buffer_6446 ( .C (clk), .D (new_AGEMA_signal_12297), .Q (new_AGEMA_signal_12298) ) ;
    buf_clk new_AGEMA_reg_buffer_6449 ( .C (clk), .D (new_AGEMA_signal_12300), .Q (new_AGEMA_signal_12301) ) ;
    buf_clk new_AGEMA_reg_buffer_6452 ( .C (clk), .D (new_AGEMA_signal_12303), .Q (new_AGEMA_signal_12304) ) ;
    buf_clk new_AGEMA_reg_buffer_6455 ( .C (clk), .D (new_AGEMA_signal_12306), .Q (new_AGEMA_signal_12307) ) ;
    buf_clk new_AGEMA_reg_buffer_6458 ( .C (clk), .D (new_AGEMA_signal_12309), .Q (new_AGEMA_signal_12310) ) ;
    buf_clk new_AGEMA_reg_buffer_6461 ( .C (clk), .D (new_AGEMA_signal_12312), .Q (new_AGEMA_signal_12313) ) ;
    buf_clk new_AGEMA_reg_buffer_6464 ( .C (clk), .D (new_AGEMA_signal_12315), .Q (new_AGEMA_signal_12316) ) ;
    buf_clk new_AGEMA_reg_buffer_6467 ( .C (clk), .D (new_AGEMA_signal_12318), .Q (new_AGEMA_signal_12319) ) ;
    buf_clk new_AGEMA_reg_buffer_6470 ( .C (clk), .D (new_AGEMA_signal_12321), .Q (new_AGEMA_signal_12322) ) ;
    buf_clk new_AGEMA_reg_buffer_6473 ( .C (clk), .D (new_AGEMA_signal_12324), .Q (new_AGEMA_signal_12325) ) ;
    buf_clk new_AGEMA_reg_buffer_6476 ( .C (clk), .D (new_AGEMA_signal_12327), .Q (new_AGEMA_signal_12328) ) ;
    buf_clk new_AGEMA_reg_buffer_6479 ( .C (clk), .D (new_AGEMA_signal_12330), .Q (new_AGEMA_signal_12331) ) ;
    buf_clk new_AGEMA_reg_buffer_6482 ( .C (clk), .D (new_AGEMA_signal_12333), .Q (new_AGEMA_signal_12334) ) ;
    buf_clk new_AGEMA_reg_buffer_6485 ( .C (clk), .D (new_AGEMA_signal_12336), .Q (new_AGEMA_signal_12337) ) ;
    buf_clk new_AGEMA_reg_buffer_6488 ( .C (clk), .D (new_AGEMA_signal_12339), .Q (new_AGEMA_signal_12340) ) ;
    buf_clk new_AGEMA_reg_buffer_6491 ( .C (clk), .D (new_AGEMA_signal_12342), .Q (new_AGEMA_signal_12343) ) ;
    buf_clk new_AGEMA_reg_buffer_6494 ( .C (clk), .D (new_AGEMA_signal_12345), .Q (new_AGEMA_signal_12346) ) ;
    buf_clk new_AGEMA_reg_buffer_6497 ( .C (clk), .D (new_AGEMA_signal_12348), .Q (new_AGEMA_signal_12349) ) ;
    buf_clk new_AGEMA_reg_buffer_6500 ( .C (clk), .D (new_AGEMA_signal_12351), .Q (new_AGEMA_signal_12352) ) ;
    buf_clk new_AGEMA_reg_buffer_6503 ( .C (clk), .D (new_AGEMA_signal_12354), .Q (new_AGEMA_signal_12355) ) ;
    buf_clk new_AGEMA_reg_buffer_6506 ( .C (clk), .D (new_AGEMA_signal_12357), .Q (new_AGEMA_signal_12358) ) ;
    buf_clk new_AGEMA_reg_buffer_6509 ( .C (clk), .D (new_AGEMA_signal_12360), .Q (new_AGEMA_signal_12361) ) ;
    buf_clk new_AGEMA_reg_buffer_6512 ( .C (clk), .D (new_AGEMA_signal_12363), .Q (new_AGEMA_signal_12364) ) ;
    buf_clk new_AGEMA_reg_buffer_6515 ( .C (clk), .D (new_AGEMA_signal_12366), .Q (new_AGEMA_signal_12367) ) ;
    buf_clk new_AGEMA_reg_buffer_6518 ( .C (clk), .D (new_AGEMA_signal_12369), .Q (new_AGEMA_signal_12370) ) ;
    buf_clk new_AGEMA_reg_buffer_6521 ( .C (clk), .D (new_AGEMA_signal_12372), .Q (new_AGEMA_signal_12373) ) ;
    buf_clk new_AGEMA_reg_buffer_6524 ( .C (clk), .D (new_AGEMA_signal_12375), .Q (new_AGEMA_signal_12376) ) ;
    buf_clk new_AGEMA_reg_buffer_6527 ( .C (clk), .D (new_AGEMA_signal_12378), .Q (new_AGEMA_signal_12379) ) ;
    buf_clk new_AGEMA_reg_buffer_6530 ( .C (clk), .D (new_AGEMA_signal_12381), .Q (new_AGEMA_signal_12382) ) ;
    buf_clk new_AGEMA_reg_buffer_6533 ( .C (clk), .D (new_AGEMA_signal_12384), .Q (new_AGEMA_signal_12385) ) ;
    buf_clk new_AGEMA_reg_buffer_6536 ( .C (clk), .D (new_AGEMA_signal_12387), .Q (new_AGEMA_signal_12388) ) ;
    buf_clk new_AGEMA_reg_buffer_6539 ( .C (clk), .D (new_AGEMA_signal_12390), .Q (new_AGEMA_signal_12391) ) ;
    buf_clk new_AGEMA_reg_buffer_6542 ( .C (clk), .D (new_AGEMA_signal_12393), .Q (new_AGEMA_signal_12394) ) ;
    buf_clk new_AGEMA_reg_buffer_6545 ( .C (clk), .D (new_AGEMA_signal_12396), .Q (new_AGEMA_signal_12397) ) ;
    buf_clk new_AGEMA_reg_buffer_6548 ( .C (clk), .D (new_AGEMA_signal_12399), .Q (new_AGEMA_signal_12400) ) ;
    buf_clk new_AGEMA_reg_buffer_6551 ( .C (clk), .D (new_AGEMA_signal_12402), .Q (new_AGEMA_signal_12403) ) ;
    buf_clk new_AGEMA_reg_buffer_6554 ( .C (clk), .D (new_AGEMA_signal_12405), .Q (new_AGEMA_signal_12406) ) ;
    buf_clk new_AGEMA_reg_buffer_6557 ( .C (clk), .D (new_AGEMA_signal_12408), .Q (new_AGEMA_signal_12409) ) ;
    buf_clk new_AGEMA_reg_buffer_6560 ( .C (clk), .D (new_AGEMA_signal_12411), .Q (new_AGEMA_signal_12412) ) ;
    buf_clk new_AGEMA_reg_buffer_6563 ( .C (clk), .D (new_AGEMA_signal_12414), .Q (new_AGEMA_signal_12415) ) ;
    buf_clk new_AGEMA_reg_buffer_6566 ( .C (clk), .D (new_AGEMA_signal_12417), .Q (new_AGEMA_signal_12418) ) ;
    buf_clk new_AGEMA_reg_buffer_6569 ( .C (clk), .D (new_AGEMA_signal_12420), .Q (new_AGEMA_signal_12421) ) ;
    buf_clk new_AGEMA_reg_buffer_6572 ( .C (clk), .D (new_AGEMA_signal_12423), .Q (new_AGEMA_signal_12424) ) ;
    buf_clk new_AGEMA_reg_buffer_6575 ( .C (clk), .D (new_AGEMA_signal_12426), .Q (new_AGEMA_signal_12427) ) ;
    buf_clk new_AGEMA_reg_buffer_6578 ( .C (clk), .D (new_AGEMA_signal_12429), .Q (new_AGEMA_signal_12430) ) ;
    buf_clk new_AGEMA_reg_buffer_6581 ( .C (clk), .D (new_AGEMA_signal_12432), .Q (new_AGEMA_signal_12433) ) ;
    buf_clk new_AGEMA_reg_buffer_6584 ( .C (clk), .D (new_AGEMA_signal_12435), .Q (new_AGEMA_signal_12436) ) ;
    buf_clk new_AGEMA_reg_buffer_6587 ( .C (clk), .D (new_AGEMA_signal_12438), .Q (new_AGEMA_signal_12439) ) ;
    buf_clk new_AGEMA_reg_buffer_6590 ( .C (clk), .D (new_AGEMA_signal_12441), .Q (new_AGEMA_signal_12442) ) ;
    buf_clk new_AGEMA_reg_buffer_6593 ( .C (clk), .D (new_AGEMA_signal_12444), .Q (new_AGEMA_signal_12445) ) ;
    buf_clk new_AGEMA_reg_buffer_6596 ( .C (clk), .D (new_AGEMA_signal_12447), .Q (new_AGEMA_signal_12448) ) ;
    buf_clk new_AGEMA_reg_buffer_6599 ( .C (clk), .D (new_AGEMA_signal_12450), .Q (new_AGEMA_signal_12451) ) ;
    buf_clk new_AGEMA_reg_buffer_6602 ( .C (clk), .D (new_AGEMA_signal_12453), .Q (new_AGEMA_signal_12454) ) ;
    buf_clk new_AGEMA_reg_buffer_6605 ( .C (clk), .D (new_AGEMA_signal_12456), .Q (new_AGEMA_signal_12457) ) ;
    buf_clk new_AGEMA_reg_buffer_6608 ( .C (clk), .D (new_AGEMA_signal_12459), .Q (new_AGEMA_signal_12460) ) ;
    buf_clk new_AGEMA_reg_buffer_6611 ( .C (clk), .D (new_AGEMA_signal_12462), .Q (new_AGEMA_signal_12463) ) ;
    buf_clk new_AGEMA_reg_buffer_6614 ( .C (clk), .D (new_AGEMA_signal_12465), .Q (new_AGEMA_signal_12466) ) ;
    buf_clk new_AGEMA_reg_buffer_6617 ( .C (clk), .D (new_AGEMA_signal_12468), .Q (new_AGEMA_signal_12469) ) ;
    buf_clk new_AGEMA_reg_buffer_6620 ( .C (clk), .D (new_AGEMA_signal_12471), .Q (new_AGEMA_signal_12472) ) ;
    buf_clk new_AGEMA_reg_buffer_6623 ( .C (clk), .D (new_AGEMA_signal_12474), .Q (new_AGEMA_signal_12475) ) ;
    buf_clk new_AGEMA_reg_buffer_6626 ( .C (clk), .D (new_AGEMA_signal_12477), .Q (new_AGEMA_signal_12478) ) ;
    buf_clk new_AGEMA_reg_buffer_6629 ( .C (clk), .D (new_AGEMA_signal_12480), .Q (new_AGEMA_signal_12481) ) ;
    buf_clk new_AGEMA_reg_buffer_6632 ( .C (clk), .D (new_AGEMA_signal_12483), .Q (new_AGEMA_signal_12484) ) ;
    buf_clk new_AGEMA_reg_buffer_6635 ( .C (clk), .D (new_AGEMA_signal_12486), .Q (new_AGEMA_signal_12487) ) ;
    buf_clk new_AGEMA_reg_buffer_6638 ( .C (clk), .D (new_AGEMA_signal_12489), .Q (new_AGEMA_signal_12490) ) ;
    buf_clk new_AGEMA_reg_buffer_6641 ( .C (clk), .D (new_AGEMA_signal_12492), .Q (new_AGEMA_signal_12493) ) ;
    buf_clk new_AGEMA_reg_buffer_6644 ( .C (clk), .D (new_AGEMA_signal_12495), .Q (new_AGEMA_signal_12496) ) ;
    buf_clk new_AGEMA_reg_buffer_6647 ( .C (clk), .D (new_AGEMA_signal_12498), .Q (new_AGEMA_signal_12499) ) ;
    buf_clk new_AGEMA_reg_buffer_6650 ( .C (clk), .D (new_AGEMA_signal_12501), .Q (new_AGEMA_signal_12502) ) ;
    buf_clk new_AGEMA_reg_buffer_6653 ( .C (clk), .D (new_AGEMA_signal_12504), .Q (new_AGEMA_signal_12505) ) ;
    buf_clk new_AGEMA_reg_buffer_6656 ( .C (clk), .D (new_AGEMA_signal_12507), .Q (new_AGEMA_signal_12508) ) ;
    buf_clk new_AGEMA_reg_buffer_6659 ( .C (clk), .D (new_AGEMA_signal_12510), .Q (new_AGEMA_signal_12511) ) ;
    buf_clk new_AGEMA_reg_buffer_6662 ( .C (clk), .D (new_AGEMA_signal_12513), .Q (new_AGEMA_signal_12514) ) ;
    buf_clk new_AGEMA_reg_buffer_6665 ( .C (clk), .D (new_AGEMA_signal_12516), .Q (new_AGEMA_signal_12517) ) ;
    buf_clk new_AGEMA_reg_buffer_6668 ( .C (clk), .D (new_AGEMA_signal_12519), .Q (new_AGEMA_signal_12520) ) ;
    buf_clk new_AGEMA_reg_buffer_6671 ( .C (clk), .D (new_AGEMA_signal_12522), .Q (new_AGEMA_signal_12523) ) ;
    buf_clk new_AGEMA_reg_buffer_6674 ( .C (clk), .D (new_AGEMA_signal_12525), .Q (new_AGEMA_signal_12526) ) ;
    buf_clk new_AGEMA_reg_buffer_6677 ( .C (clk), .D (new_AGEMA_signal_12528), .Q (new_AGEMA_signal_12529) ) ;
    buf_clk new_AGEMA_reg_buffer_6680 ( .C (clk), .D (new_AGEMA_signal_12531), .Q (new_AGEMA_signal_12532) ) ;
    buf_clk new_AGEMA_reg_buffer_6683 ( .C (clk), .D (new_AGEMA_signal_12534), .Q (new_AGEMA_signal_12535) ) ;
    buf_clk new_AGEMA_reg_buffer_6686 ( .C (clk), .D (new_AGEMA_signal_12537), .Q (new_AGEMA_signal_12538) ) ;
    buf_clk new_AGEMA_reg_buffer_6689 ( .C (clk), .D (new_AGEMA_signal_12540), .Q (new_AGEMA_signal_12541) ) ;
    buf_clk new_AGEMA_reg_buffer_6692 ( .C (clk), .D (new_AGEMA_signal_12543), .Q (new_AGEMA_signal_12544) ) ;
    buf_clk new_AGEMA_reg_buffer_6695 ( .C (clk), .D (new_AGEMA_signal_12546), .Q (new_AGEMA_signal_12547) ) ;
    buf_clk new_AGEMA_reg_buffer_6698 ( .C (clk), .D (new_AGEMA_signal_12549), .Q (new_AGEMA_signal_12550) ) ;
    buf_clk new_AGEMA_reg_buffer_6701 ( .C (clk), .D (new_AGEMA_signal_12552), .Q (new_AGEMA_signal_12553) ) ;
    buf_clk new_AGEMA_reg_buffer_6704 ( .C (clk), .D (new_AGEMA_signal_12555), .Q (new_AGEMA_signal_12556) ) ;
    buf_clk new_AGEMA_reg_buffer_6707 ( .C (clk), .D (new_AGEMA_signal_12558), .Q (new_AGEMA_signal_12559) ) ;
    buf_clk new_AGEMA_reg_buffer_6710 ( .C (clk), .D (new_AGEMA_signal_12561), .Q (new_AGEMA_signal_12562) ) ;
    buf_clk new_AGEMA_reg_buffer_6713 ( .C (clk), .D (new_AGEMA_signal_12564), .Q (new_AGEMA_signal_12565) ) ;
    buf_clk new_AGEMA_reg_buffer_6716 ( .C (clk), .D (new_AGEMA_signal_12567), .Q (new_AGEMA_signal_12568) ) ;
    buf_clk new_AGEMA_reg_buffer_6719 ( .C (clk), .D (new_AGEMA_signal_12570), .Q (new_AGEMA_signal_12571) ) ;
    buf_clk new_AGEMA_reg_buffer_6722 ( .C (clk), .D (new_AGEMA_signal_12573), .Q (new_AGEMA_signal_12574) ) ;
    buf_clk new_AGEMA_reg_buffer_6725 ( .C (clk), .D (new_AGEMA_signal_12576), .Q (new_AGEMA_signal_12577) ) ;
    buf_clk new_AGEMA_reg_buffer_6728 ( .C (clk), .D (new_AGEMA_signal_12579), .Q (new_AGEMA_signal_12580) ) ;
    buf_clk new_AGEMA_reg_buffer_6731 ( .C (clk), .D (new_AGEMA_signal_12582), .Q (new_AGEMA_signal_12583) ) ;
    buf_clk new_AGEMA_reg_buffer_6734 ( .C (clk), .D (new_AGEMA_signal_12585), .Q (new_AGEMA_signal_12586) ) ;
    buf_clk new_AGEMA_reg_buffer_6737 ( .C (clk), .D (new_AGEMA_signal_12588), .Q (new_AGEMA_signal_12589) ) ;
    buf_clk new_AGEMA_reg_buffer_6740 ( .C (clk), .D (new_AGEMA_signal_12591), .Q (new_AGEMA_signal_12592) ) ;
    buf_clk new_AGEMA_reg_buffer_6743 ( .C (clk), .D (new_AGEMA_signal_12594), .Q (new_AGEMA_signal_12595) ) ;
    buf_clk new_AGEMA_reg_buffer_6746 ( .C (clk), .D (new_AGEMA_signal_12597), .Q (new_AGEMA_signal_12598) ) ;
    buf_clk new_AGEMA_reg_buffer_6749 ( .C (clk), .D (new_AGEMA_signal_12600), .Q (new_AGEMA_signal_12601) ) ;
    buf_clk new_AGEMA_reg_buffer_6752 ( .C (clk), .D (new_AGEMA_signal_12603), .Q (new_AGEMA_signal_12604) ) ;
    buf_clk new_AGEMA_reg_buffer_6755 ( .C (clk), .D (new_AGEMA_signal_12606), .Q (new_AGEMA_signal_12607) ) ;
    buf_clk new_AGEMA_reg_buffer_6758 ( .C (clk), .D (new_AGEMA_signal_12609), .Q (new_AGEMA_signal_12610) ) ;
    buf_clk new_AGEMA_reg_buffer_6761 ( .C (clk), .D (new_AGEMA_signal_12612), .Q (new_AGEMA_signal_12613) ) ;
    buf_clk new_AGEMA_reg_buffer_6764 ( .C (clk), .D (new_AGEMA_signal_12615), .Q (new_AGEMA_signal_12616) ) ;
    buf_clk new_AGEMA_reg_buffer_6767 ( .C (clk), .D (new_AGEMA_signal_12618), .Q (new_AGEMA_signal_12619) ) ;
    buf_clk new_AGEMA_reg_buffer_6770 ( .C (clk), .D (new_AGEMA_signal_12621), .Q (new_AGEMA_signal_12622) ) ;
    buf_clk new_AGEMA_reg_buffer_6773 ( .C (clk), .D (new_AGEMA_signal_12624), .Q (new_AGEMA_signal_12625) ) ;
    buf_clk new_AGEMA_reg_buffer_6776 ( .C (clk), .D (new_AGEMA_signal_12627), .Q (new_AGEMA_signal_12628) ) ;
    buf_clk new_AGEMA_reg_buffer_6779 ( .C (clk), .D (new_AGEMA_signal_12630), .Q (new_AGEMA_signal_12631) ) ;
    buf_clk new_AGEMA_reg_buffer_6782 ( .C (clk), .D (new_AGEMA_signal_12633), .Q (new_AGEMA_signal_12634) ) ;
    buf_clk new_AGEMA_reg_buffer_6785 ( .C (clk), .D (new_AGEMA_signal_12636), .Q (new_AGEMA_signal_12637) ) ;
    buf_clk new_AGEMA_reg_buffer_6788 ( .C (clk), .D (new_AGEMA_signal_12639), .Q (new_AGEMA_signal_12640) ) ;
    buf_clk new_AGEMA_reg_buffer_6791 ( .C (clk), .D (new_AGEMA_signal_12642), .Q (new_AGEMA_signal_12643) ) ;
    buf_clk new_AGEMA_reg_buffer_6794 ( .C (clk), .D (new_AGEMA_signal_12645), .Q (new_AGEMA_signal_12646) ) ;
    buf_clk new_AGEMA_reg_buffer_6797 ( .C (clk), .D (new_AGEMA_signal_12648), .Q (new_AGEMA_signal_12649) ) ;
    buf_clk new_AGEMA_reg_buffer_6800 ( .C (clk), .D (new_AGEMA_signal_12651), .Q (new_AGEMA_signal_12652) ) ;
    buf_clk new_AGEMA_reg_buffer_6803 ( .C (clk), .D (new_AGEMA_signal_12654), .Q (new_AGEMA_signal_12655) ) ;
    buf_clk new_AGEMA_reg_buffer_6806 ( .C (clk), .D (new_AGEMA_signal_12657), .Q (new_AGEMA_signal_12658) ) ;
    buf_clk new_AGEMA_reg_buffer_6809 ( .C (clk), .D (new_AGEMA_signal_12660), .Q (new_AGEMA_signal_12661) ) ;
    buf_clk new_AGEMA_reg_buffer_6812 ( .C (clk), .D (new_AGEMA_signal_12663), .Q (new_AGEMA_signal_12664) ) ;
    buf_clk new_AGEMA_reg_buffer_6815 ( .C (clk), .D (new_AGEMA_signal_12666), .Q (new_AGEMA_signal_12667) ) ;
    buf_clk new_AGEMA_reg_buffer_6818 ( .C (clk), .D (new_AGEMA_signal_12669), .Q (new_AGEMA_signal_12670) ) ;
    buf_clk new_AGEMA_reg_buffer_6821 ( .C (clk), .D (new_AGEMA_signal_12672), .Q (new_AGEMA_signal_12673) ) ;
    buf_clk new_AGEMA_reg_buffer_6824 ( .C (clk), .D (new_AGEMA_signal_12675), .Q (new_AGEMA_signal_12676) ) ;
    buf_clk new_AGEMA_reg_buffer_6827 ( .C (clk), .D (new_AGEMA_signal_12678), .Q (new_AGEMA_signal_12679) ) ;
    buf_clk new_AGEMA_reg_buffer_6830 ( .C (clk), .D (new_AGEMA_signal_12681), .Q (new_AGEMA_signal_12682) ) ;
    buf_clk new_AGEMA_reg_buffer_6833 ( .C (clk), .D (new_AGEMA_signal_12684), .Q (new_AGEMA_signal_12685) ) ;
    buf_clk new_AGEMA_reg_buffer_6836 ( .C (clk), .D (new_AGEMA_signal_12687), .Q (new_AGEMA_signal_12688) ) ;
    buf_clk new_AGEMA_reg_buffer_6839 ( .C (clk), .D (new_AGEMA_signal_12690), .Q (new_AGEMA_signal_12691) ) ;
    buf_clk new_AGEMA_reg_buffer_6842 ( .C (clk), .D (new_AGEMA_signal_12693), .Q (new_AGEMA_signal_12694) ) ;
    buf_clk new_AGEMA_reg_buffer_6845 ( .C (clk), .D (new_AGEMA_signal_12696), .Q (new_AGEMA_signal_12697) ) ;
    buf_clk new_AGEMA_reg_buffer_6848 ( .C (clk), .D (new_AGEMA_signal_12699), .Q (new_AGEMA_signal_12700) ) ;
    buf_clk new_AGEMA_reg_buffer_6851 ( .C (clk), .D (new_AGEMA_signal_12702), .Q (new_AGEMA_signal_12703) ) ;
    buf_clk new_AGEMA_reg_buffer_6854 ( .C (clk), .D (new_AGEMA_signal_12705), .Q (new_AGEMA_signal_12706) ) ;
    buf_clk new_AGEMA_reg_buffer_6857 ( .C (clk), .D (new_AGEMA_signal_12708), .Q (new_AGEMA_signal_12709) ) ;
    buf_clk new_AGEMA_reg_buffer_6860 ( .C (clk), .D (new_AGEMA_signal_12711), .Q (new_AGEMA_signal_12712) ) ;
    buf_clk new_AGEMA_reg_buffer_6863 ( .C (clk), .D (new_AGEMA_signal_12714), .Q (new_AGEMA_signal_12715) ) ;
    buf_clk new_AGEMA_reg_buffer_6866 ( .C (clk), .D (new_AGEMA_signal_12717), .Q (new_AGEMA_signal_12718) ) ;
    buf_clk new_AGEMA_reg_buffer_6869 ( .C (clk), .D (new_AGEMA_signal_12720), .Q (new_AGEMA_signal_12721) ) ;
    buf_clk new_AGEMA_reg_buffer_6872 ( .C (clk), .D (new_AGEMA_signal_12723), .Q (new_AGEMA_signal_12724) ) ;
    buf_clk new_AGEMA_reg_buffer_6875 ( .C (clk), .D (new_AGEMA_signal_12726), .Q (new_AGEMA_signal_12727) ) ;
    buf_clk new_AGEMA_reg_buffer_6878 ( .C (clk), .D (new_AGEMA_signal_12729), .Q (new_AGEMA_signal_12730) ) ;
    buf_clk new_AGEMA_reg_buffer_6881 ( .C (clk), .D (new_AGEMA_signal_12732), .Q (new_AGEMA_signal_12733) ) ;
    buf_clk new_AGEMA_reg_buffer_6884 ( .C (clk), .D (new_AGEMA_signal_12735), .Q (new_AGEMA_signal_12736) ) ;
    buf_clk new_AGEMA_reg_buffer_6887 ( .C (clk), .D (new_AGEMA_signal_12738), .Q (new_AGEMA_signal_12739) ) ;
    buf_clk new_AGEMA_reg_buffer_6890 ( .C (clk), .D (new_AGEMA_signal_12741), .Q (new_AGEMA_signal_12742) ) ;
    buf_clk new_AGEMA_reg_buffer_6893 ( .C (clk), .D (new_AGEMA_signal_12744), .Q (new_AGEMA_signal_12745) ) ;
    buf_clk new_AGEMA_reg_buffer_6896 ( .C (clk), .D (new_AGEMA_signal_12747), .Q (new_AGEMA_signal_12748) ) ;
    buf_clk new_AGEMA_reg_buffer_6899 ( .C (clk), .D (new_AGEMA_signal_12750), .Q (new_AGEMA_signal_12751) ) ;
    buf_clk new_AGEMA_reg_buffer_6902 ( .C (clk), .D (new_AGEMA_signal_12753), .Q (new_AGEMA_signal_12754) ) ;
    buf_clk new_AGEMA_reg_buffer_6905 ( .C (clk), .D (new_AGEMA_signal_12756), .Q (new_AGEMA_signal_12757) ) ;
    buf_clk new_AGEMA_reg_buffer_6908 ( .C (clk), .D (new_AGEMA_signal_12759), .Q (new_AGEMA_signal_12760) ) ;
    buf_clk new_AGEMA_reg_buffer_6911 ( .C (clk), .D (new_AGEMA_signal_12762), .Q (new_AGEMA_signal_12763) ) ;
    buf_clk new_AGEMA_reg_buffer_6914 ( .C (clk), .D (new_AGEMA_signal_12765), .Q (new_AGEMA_signal_12766) ) ;
    buf_clk new_AGEMA_reg_buffer_6917 ( .C (clk), .D (new_AGEMA_signal_12768), .Q (new_AGEMA_signal_12769) ) ;
    buf_clk new_AGEMA_reg_buffer_6920 ( .C (clk), .D (new_AGEMA_signal_12771), .Q (new_AGEMA_signal_12772) ) ;
    buf_clk new_AGEMA_reg_buffer_6923 ( .C (clk), .D (new_AGEMA_signal_12774), .Q (new_AGEMA_signal_12775) ) ;
    buf_clk new_AGEMA_reg_buffer_6926 ( .C (clk), .D (new_AGEMA_signal_12777), .Q (new_AGEMA_signal_12778) ) ;
    buf_clk new_AGEMA_reg_buffer_6929 ( .C (clk), .D (new_AGEMA_signal_12780), .Q (new_AGEMA_signal_12781) ) ;
    buf_clk new_AGEMA_reg_buffer_6932 ( .C (clk), .D (new_AGEMA_signal_12783), .Q (new_AGEMA_signal_12784) ) ;
    buf_clk new_AGEMA_reg_buffer_6935 ( .C (clk), .D (new_AGEMA_signal_12786), .Q (new_AGEMA_signal_12787) ) ;
    buf_clk new_AGEMA_reg_buffer_6938 ( .C (clk), .D (new_AGEMA_signal_12789), .Q (new_AGEMA_signal_12790) ) ;
    buf_clk new_AGEMA_reg_buffer_6941 ( .C (clk), .D (new_AGEMA_signal_12792), .Q (new_AGEMA_signal_12793) ) ;
    buf_clk new_AGEMA_reg_buffer_6944 ( .C (clk), .D (new_AGEMA_signal_12795), .Q (new_AGEMA_signal_12796) ) ;
    buf_clk new_AGEMA_reg_buffer_6947 ( .C (clk), .D (new_AGEMA_signal_12798), .Q (new_AGEMA_signal_12799) ) ;
    buf_clk new_AGEMA_reg_buffer_6950 ( .C (clk), .D (new_AGEMA_signal_12801), .Q (new_AGEMA_signal_12802) ) ;
    buf_clk new_AGEMA_reg_buffer_6953 ( .C (clk), .D (new_AGEMA_signal_12804), .Q (new_AGEMA_signal_12805) ) ;
    buf_clk new_AGEMA_reg_buffer_6956 ( .C (clk), .D (new_AGEMA_signal_12807), .Q (new_AGEMA_signal_12808) ) ;
    buf_clk new_AGEMA_reg_buffer_6959 ( .C (clk), .D (new_AGEMA_signal_12810), .Q (new_AGEMA_signal_12811) ) ;
    buf_clk new_AGEMA_reg_buffer_6962 ( .C (clk), .D (new_AGEMA_signal_12813), .Q (new_AGEMA_signal_12814) ) ;
    buf_clk new_AGEMA_reg_buffer_6965 ( .C (clk), .D (new_AGEMA_signal_12816), .Q (new_AGEMA_signal_12817) ) ;
    buf_clk new_AGEMA_reg_buffer_6968 ( .C (clk), .D (new_AGEMA_signal_12819), .Q (new_AGEMA_signal_12820) ) ;
    buf_clk new_AGEMA_reg_buffer_6971 ( .C (clk), .D (new_AGEMA_signal_12822), .Q (new_AGEMA_signal_12823) ) ;
    buf_clk new_AGEMA_reg_buffer_6974 ( .C (clk), .D (new_AGEMA_signal_12825), .Q (new_AGEMA_signal_12826) ) ;
    buf_clk new_AGEMA_reg_buffer_6977 ( .C (clk), .D (new_AGEMA_signal_12828), .Q (new_AGEMA_signal_12829) ) ;
    buf_clk new_AGEMA_reg_buffer_6980 ( .C (clk), .D (new_AGEMA_signal_12831), .Q (new_AGEMA_signal_12832) ) ;
    buf_clk new_AGEMA_reg_buffer_6983 ( .C (clk), .D (new_AGEMA_signal_12834), .Q (new_AGEMA_signal_12835) ) ;
    buf_clk new_AGEMA_reg_buffer_6986 ( .C (clk), .D (new_AGEMA_signal_12837), .Q (new_AGEMA_signal_12838) ) ;
    buf_clk new_AGEMA_reg_buffer_6989 ( .C (clk), .D (new_AGEMA_signal_12840), .Q (new_AGEMA_signal_12841) ) ;
    buf_clk new_AGEMA_reg_buffer_6992 ( .C (clk), .D (new_AGEMA_signal_12843), .Q (new_AGEMA_signal_12844) ) ;
    buf_clk new_AGEMA_reg_buffer_6995 ( .C (clk), .D (new_AGEMA_signal_12846), .Q (new_AGEMA_signal_12847) ) ;
    buf_clk new_AGEMA_reg_buffer_6998 ( .C (clk), .D (new_AGEMA_signal_12849), .Q (new_AGEMA_signal_12850) ) ;
    buf_clk new_AGEMA_reg_buffer_7001 ( .C (clk), .D (new_AGEMA_signal_12852), .Q (new_AGEMA_signal_12853) ) ;
    buf_clk new_AGEMA_reg_buffer_7004 ( .C (clk), .D (new_AGEMA_signal_12855), .Q (new_AGEMA_signal_12856) ) ;
    buf_clk new_AGEMA_reg_buffer_7007 ( .C (clk), .D (new_AGEMA_signal_12858), .Q (new_AGEMA_signal_12859) ) ;
    buf_clk new_AGEMA_reg_buffer_7010 ( .C (clk), .D (new_AGEMA_signal_12861), .Q (new_AGEMA_signal_12862) ) ;
    buf_clk new_AGEMA_reg_buffer_7013 ( .C (clk), .D (new_AGEMA_signal_12864), .Q (new_AGEMA_signal_12865) ) ;
    buf_clk new_AGEMA_reg_buffer_7016 ( .C (clk), .D (new_AGEMA_signal_12867), .Q (new_AGEMA_signal_12868) ) ;
    buf_clk new_AGEMA_reg_buffer_7019 ( .C (clk), .D (new_AGEMA_signal_12870), .Q (new_AGEMA_signal_12871) ) ;
    buf_clk new_AGEMA_reg_buffer_7022 ( .C (clk), .D (new_AGEMA_signal_12873), .Q (new_AGEMA_signal_12874) ) ;
    buf_clk new_AGEMA_reg_buffer_7025 ( .C (clk), .D (new_AGEMA_signal_12876), .Q (new_AGEMA_signal_12877) ) ;
    buf_clk new_AGEMA_reg_buffer_7028 ( .C (clk), .D (new_AGEMA_signal_12879), .Q (new_AGEMA_signal_12880) ) ;
    buf_clk new_AGEMA_reg_buffer_7031 ( .C (clk), .D (new_AGEMA_signal_12882), .Q (new_AGEMA_signal_12883) ) ;
    buf_clk new_AGEMA_reg_buffer_7034 ( .C (clk), .D (new_AGEMA_signal_12885), .Q (new_AGEMA_signal_12886) ) ;
    buf_clk new_AGEMA_reg_buffer_7037 ( .C (clk), .D (new_AGEMA_signal_12888), .Q (new_AGEMA_signal_12889) ) ;
    buf_clk new_AGEMA_reg_buffer_7040 ( .C (clk), .D (new_AGEMA_signal_12891), .Q (new_AGEMA_signal_12892) ) ;
    buf_clk new_AGEMA_reg_buffer_7043 ( .C (clk), .D (new_AGEMA_signal_12894), .Q (new_AGEMA_signal_12895) ) ;
    buf_clk new_AGEMA_reg_buffer_7046 ( .C (clk), .D (new_AGEMA_signal_12897), .Q (new_AGEMA_signal_12898) ) ;
    buf_clk new_AGEMA_reg_buffer_7049 ( .C (clk), .D (new_AGEMA_signal_12900), .Q (new_AGEMA_signal_12901) ) ;
    buf_clk new_AGEMA_reg_buffer_7052 ( .C (clk), .D (new_AGEMA_signal_12903), .Q (new_AGEMA_signal_12904) ) ;
    buf_clk new_AGEMA_reg_buffer_7055 ( .C (clk), .D (new_AGEMA_signal_12906), .Q (new_AGEMA_signal_12907) ) ;
    buf_clk new_AGEMA_reg_buffer_7058 ( .C (clk), .D (new_AGEMA_signal_12909), .Q (new_AGEMA_signal_12910) ) ;
    buf_clk new_AGEMA_reg_buffer_7061 ( .C (clk), .D (new_AGEMA_signal_12912), .Q (new_AGEMA_signal_12913) ) ;
    buf_clk new_AGEMA_reg_buffer_7064 ( .C (clk), .D (new_AGEMA_signal_12915), .Q (new_AGEMA_signal_12916) ) ;
    buf_clk new_AGEMA_reg_buffer_7067 ( .C (clk), .D (new_AGEMA_signal_12918), .Q (new_AGEMA_signal_12919) ) ;
    buf_clk new_AGEMA_reg_buffer_7070 ( .C (clk), .D (new_AGEMA_signal_12921), .Q (new_AGEMA_signal_12922) ) ;
    buf_clk new_AGEMA_reg_buffer_7073 ( .C (clk), .D (new_AGEMA_signal_12924), .Q (new_AGEMA_signal_12925) ) ;
    buf_clk new_AGEMA_reg_buffer_7076 ( .C (clk), .D (new_AGEMA_signal_12927), .Q (new_AGEMA_signal_12928) ) ;
    buf_clk new_AGEMA_reg_buffer_7079 ( .C (clk), .D (new_AGEMA_signal_12930), .Q (new_AGEMA_signal_12931) ) ;
    buf_clk new_AGEMA_reg_buffer_7082 ( .C (clk), .D (new_AGEMA_signal_12933), .Q (new_AGEMA_signal_12934) ) ;
    buf_clk new_AGEMA_reg_buffer_7085 ( .C (clk), .D (new_AGEMA_signal_12936), .Q (new_AGEMA_signal_12937) ) ;
    buf_clk new_AGEMA_reg_buffer_7088 ( .C (clk), .D (new_AGEMA_signal_12939), .Q (new_AGEMA_signal_12940) ) ;
    buf_clk new_AGEMA_reg_buffer_7091 ( .C (clk), .D (new_AGEMA_signal_12942), .Q (new_AGEMA_signal_12943) ) ;
    buf_clk new_AGEMA_reg_buffer_7094 ( .C (clk), .D (new_AGEMA_signal_12945), .Q (new_AGEMA_signal_12946) ) ;
    buf_clk new_AGEMA_reg_buffer_7097 ( .C (clk), .D (new_AGEMA_signal_12948), .Q (new_AGEMA_signal_12949) ) ;
    buf_clk new_AGEMA_reg_buffer_7100 ( .C (clk), .D (new_AGEMA_signal_12951), .Q (new_AGEMA_signal_12952) ) ;
    buf_clk new_AGEMA_reg_buffer_7103 ( .C (clk), .D (new_AGEMA_signal_12954), .Q (new_AGEMA_signal_12955) ) ;
    buf_clk new_AGEMA_reg_buffer_7106 ( .C (clk), .D (new_AGEMA_signal_12957), .Q (new_AGEMA_signal_12958) ) ;
    buf_clk new_AGEMA_reg_buffer_7109 ( .C (clk), .D (new_AGEMA_signal_12960), .Q (new_AGEMA_signal_12961) ) ;
    buf_clk new_AGEMA_reg_buffer_7112 ( .C (clk), .D (new_AGEMA_signal_12963), .Q (new_AGEMA_signal_12964) ) ;
    buf_clk new_AGEMA_reg_buffer_7115 ( .C (clk), .D (new_AGEMA_signal_12966), .Q (new_AGEMA_signal_12967) ) ;
    buf_clk new_AGEMA_reg_buffer_7118 ( .C (clk), .D (new_AGEMA_signal_12969), .Q (new_AGEMA_signal_12970) ) ;
    buf_clk new_AGEMA_reg_buffer_7121 ( .C (clk), .D (new_AGEMA_signal_12972), .Q (new_AGEMA_signal_12973) ) ;
    buf_clk new_AGEMA_reg_buffer_7124 ( .C (clk), .D (new_AGEMA_signal_12975), .Q (new_AGEMA_signal_12976) ) ;
    buf_clk new_AGEMA_reg_buffer_7127 ( .C (clk), .D (new_AGEMA_signal_12978), .Q (new_AGEMA_signal_12979) ) ;
    buf_clk new_AGEMA_reg_buffer_7130 ( .C (clk), .D (new_AGEMA_signal_12981), .Q (new_AGEMA_signal_12982) ) ;
    buf_clk new_AGEMA_reg_buffer_7133 ( .C (clk), .D (new_AGEMA_signal_12984), .Q (new_AGEMA_signal_12985) ) ;
    buf_clk new_AGEMA_reg_buffer_7136 ( .C (clk), .D (new_AGEMA_signal_12987), .Q (new_AGEMA_signal_12988) ) ;
    buf_clk new_AGEMA_reg_buffer_7139 ( .C (clk), .D (new_AGEMA_signal_12990), .Q (new_AGEMA_signal_12991) ) ;
    buf_clk new_AGEMA_reg_buffer_7142 ( .C (clk), .D (new_AGEMA_signal_12993), .Q (new_AGEMA_signal_12994) ) ;
    buf_clk new_AGEMA_reg_buffer_7145 ( .C (clk), .D (new_AGEMA_signal_12996), .Q (new_AGEMA_signal_12997) ) ;
    buf_clk new_AGEMA_reg_buffer_7148 ( .C (clk), .D (new_AGEMA_signal_12999), .Q (new_AGEMA_signal_13000) ) ;
    buf_clk new_AGEMA_reg_buffer_7151 ( .C (clk), .D (new_AGEMA_signal_13002), .Q (new_AGEMA_signal_13003) ) ;
    buf_clk new_AGEMA_reg_buffer_7154 ( .C (clk), .D (new_AGEMA_signal_13005), .Q (new_AGEMA_signal_13006) ) ;
    buf_clk new_AGEMA_reg_buffer_7157 ( .C (clk), .D (new_AGEMA_signal_13008), .Q (new_AGEMA_signal_13009) ) ;
    buf_clk new_AGEMA_reg_buffer_7160 ( .C (clk), .D (new_AGEMA_signal_13011), .Q (new_AGEMA_signal_13012) ) ;
    buf_clk new_AGEMA_reg_buffer_7163 ( .C (clk), .D (new_AGEMA_signal_13014), .Q (new_AGEMA_signal_13015) ) ;
    buf_clk new_AGEMA_reg_buffer_7166 ( .C (clk), .D (new_AGEMA_signal_13017), .Q (new_AGEMA_signal_13018) ) ;
    buf_clk new_AGEMA_reg_buffer_7169 ( .C (clk), .D (new_AGEMA_signal_13020), .Q (new_AGEMA_signal_13021) ) ;
    buf_clk new_AGEMA_reg_buffer_7172 ( .C (clk), .D (new_AGEMA_signal_13023), .Q (new_AGEMA_signal_13024) ) ;
    buf_clk new_AGEMA_reg_buffer_7175 ( .C (clk), .D (new_AGEMA_signal_13026), .Q (new_AGEMA_signal_13027) ) ;
    buf_clk new_AGEMA_reg_buffer_7178 ( .C (clk), .D (new_AGEMA_signal_13029), .Q (new_AGEMA_signal_13030) ) ;
    buf_clk new_AGEMA_reg_buffer_7181 ( .C (clk), .D (new_AGEMA_signal_13032), .Q (new_AGEMA_signal_13033) ) ;
    buf_clk new_AGEMA_reg_buffer_7184 ( .C (clk), .D (new_AGEMA_signal_13035), .Q (new_AGEMA_signal_13036) ) ;
    buf_clk new_AGEMA_reg_buffer_7187 ( .C (clk), .D (new_AGEMA_signal_13038), .Q (new_AGEMA_signal_13039) ) ;
    buf_clk new_AGEMA_reg_buffer_7190 ( .C (clk), .D (new_AGEMA_signal_13041), .Q (new_AGEMA_signal_13042) ) ;
    buf_clk new_AGEMA_reg_buffer_7193 ( .C (clk), .D (new_AGEMA_signal_13044), .Q (new_AGEMA_signal_13045) ) ;
    buf_clk new_AGEMA_reg_buffer_7196 ( .C (clk), .D (new_AGEMA_signal_13047), .Q (new_AGEMA_signal_13048) ) ;
    buf_clk new_AGEMA_reg_buffer_7199 ( .C (clk), .D (new_AGEMA_signal_13050), .Q (new_AGEMA_signal_13051) ) ;
    buf_clk new_AGEMA_reg_buffer_7202 ( .C (clk), .D (new_AGEMA_signal_13053), .Q (new_AGEMA_signal_13054) ) ;
    buf_clk new_AGEMA_reg_buffer_7205 ( .C (clk), .D (new_AGEMA_signal_13056), .Q (new_AGEMA_signal_13057) ) ;
    buf_clk new_AGEMA_reg_buffer_7208 ( .C (clk), .D (new_AGEMA_signal_13059), .Q (new_AGEMA_signal_13060) ) ;
    buf_clk new_AGEMA_reg_buffer_7211 ( .C (clk), .D (new_AGEMA_signal_13062), .Q (new_AGEMA_signal_13063) ) ;
    buf_clk new_AGEMA_reg_buffer_7214 ( .C (clk), .D (new_AGEMA_signal_13065), .Q (new_AGEMA_signal_13066) ) ;
    buf_clk new_AGEMA_reg_buffer_7217 ( .C (clk), .D (new_AGEMA_signal_13068), .Q (new_AGEMA_signal_13069) ) ;
    buf_clk new_AGEMA_reg_buffer_7220 ( .C (clk), .D (new_AGEMA_signal_13071), .Q (new_AGEMA_signal_13072) ) ;
    buf_clk new_AGEMA_reg_buffer_7223 ( .C (clk), .D (new_AGEMA_signal_13074), .Q (new_AGEMA_signal_13075) ) ;
    buf_clk new_AGEMA_reg_buffer_7226 ( .C (clk), .D (new_AGEMA_signal_13077), .Q (new_AGEMA_signal_13078) ) ;
    buf_clk new_AGEMA_reg_buffer_7229 ( .C (clk), .D (new_AGEMA_signal_13080), .Q (new_AGEMA_signal_13081) ) ;
    buf_clk new_AGEMA_reg_buffer_7232 ( .C (clk), .D (new_AGEMA_signal_13083), .Q (new_AGEMA_signal_13084) ) ;
    buf_clk new_AGEMA_reg_buffer_7235 ( .C (clk), .D (new_AGEMA_signal_13086), .Q (new_AGEMA_signal_13087) ) ;
    buf_clk new_AGEMA_reg_buffer_7238 ( .C (clk), .D (new_AGEMA_signal_13089), .Q (new_AGEMA_signal_13090) ) ;
    buf_clk new_AGEMA_reg_buffer_7241 ( .C (clk), .D (new_AGEMA_signal_13092), .Q (new_AGEMA_signal_13093) ) ;
    buf_clk new_AGEMA_reg_buffer_7244 ( .C (clk), .D (new_AGEMA_signal_13095), .Q (new_AGEMA_signal_13096) ) ;
    buf_clk new_AGEMA_reg_buffer_7247 ( .C (clk), .D (new_AGEMA_signal_13098), .Q (new_AGEMA_signal_13099) ) ;
    buf_clk new_AGEMA_reg_buffer_7250 ( .C (clk), .D (new_AGEMA_signal_13101), .Q (new_AGEMA_signal_13102) ) ;
    buf_clk new_AGEMA_reg_buffer_7253 ( .C (clk), .D (new_AGEMA_signal_13104), .Q (new_AGEMA_signal_13105) ) ;
    buf_clk new_AGEMA_reg_buffer_7256 ( .C (clk), .D (new_AGEMA_signal_13107), .Q (new_AGEMA_signal_13108) ) ;
    buf_clk new_AGEMA_reg_buffer_7259 ( .C (clk), .D (new_AGEMA_signal_13110), .Q (new_AGEMA_signal_13111) ) ;
    buf_clk new_AGEMA_reg_buffer_7262 ( .C (clk), .D (new_AGEMA_signal_13113), .Q (new_AGEMA_signal_13114) ) ;
    buf_clk new_AGEMA_reg_buffer_7265 ( .C (clk), .D (new_AGEMA_signal_13116), .Q (new_AGEMA_signal_13117) ) ;
    buf_clk new_AGEMA_reg_buffer_7268 ( .C (clk), .D (new_AGEMA_signal_13119), .Q (new_AGEMA_signal_13120) ) ;
    buf_clk new_AGEMA_reg_buffer_7271 ( .C (clk), .D (new_AGEMA_signal_13122), .Q (new_AGEMA_signal_13123) ) ;
    buf_clk new_AGEMA_reg_buffer_7274 ( .C (clk), .D (new_AGEMA_signal_13125), .Q (new_AGEMA_signal_13126) ) ;
    buf_clk new_AGEMA_reg_buffer_7277 ( .C (clk), .D (new_AGEMA_signal_13128), .Q (new_AGEMA_signal_13129) ) ;
    buf_clk new_AGEMA_reg_buffer_7280 ( .C (clk), .D (new_AGEMA_signal_13131), .Q (new_AGEMA_signal_13132) ) ;
    buf_clk new_AGEMA_reg_buffer_7283 ( .C (clk), .D (new_AGEMA_signal_13134), .Q (new_AGEMA_signal_13135) ) ;
    buf_clk new_AGEMA_reg_buffer_7286 ( .C (clk), .D (new_AGEMA_signal_13137), .Q (new_AGEMA_signal_13138) ) ;
    buf_clk new_AGEMA_reg_buffer_7289 ( .C (clk), .D (new_AGEMA_signal_13140), .Q (new_AGEMA_signal_13141) ) ;
    buf_clk new_AGEMA_reg_buffer_7292 ( .C (clk), .D (new_AGEMA_signal_13143), .Q (new_AGEMA_signal_13144) ) ;
    buf_clk new_AGEMA_reg_buffer_7295 ( .C (clk), .D (new_AGEMA_signal_13146), .Q (new_AGEMA_signal_13147) ) ;
    buf_clk new_AGEMA_reg_buffer_7298 ( .C (clk), .D (new_AGEMA_signal_13149), .Q (new_AGEMA_signal_13150) ) ;
    buf_clk new_AGEMA_reg_buffer_7301 ( .C (clk), .D (new_AGEMA_signal_13152), .Q (new_AGEMA_signal_13153) ) ;
    buf_clk new_AGEMA_reg_buffer_7304 ( .C (clk), .D (new_AGEMA_signal_13155), .Q (new_AGEMA_signal_13156) ) ;
    buf_clk new_AGEMA_reg_buffer_7307 ( .C (clk), .D (new_AGEMA_signal_13158), .Q (new_AGEMA_signal_13159) ) ;
    buf_clk new_AGEMA_reg_buffer_7310 ( .C (clk), .D (new_AGEMA_signal_13161), .Q (new_AGEMA_signal_13162) ) ;
    buf_clk new_AGEMA_reg_buffer_7313 ( .C (clk), .D (new_AGEMA_signal_13164), .Q (new_AGEMA_signal_13165) ) ;
    buf_clk new_AGEMA_reg_buffer_7316 ( .C (clk), .D (new_AGEMA_signal_13167), .Q (new_AGEMA_signal_13168) ) ;
    buf_clk new_AGEMA_reg_buffer_7319 ( .C (clk), .D (new_AGEMA_signal_13170), .Q (new_AGEMA_signal_13171) ) ;
    buf_clk new_AGEMA_reg_buffer_7322 ( .C (clk), .D (new_AGEMA_signal_13173), .Q (new_AGEMA_signal_13174) ) ;
    buf_clk new_AGEMA_reg_buffer_7325 ( .C (clk), .D (new_AGEMA_signal_13176), .Q (new_AGEMA_signal_13177) ) ;
    buf_clk new_AGEMA_reg_buffer_7328 ( .C (clk), .D (new_AGEMA_signal_13179), .Q (new_AGEMA_signal_13180) ) ;
    buf_clk new_AGEMA_reg_buffer_7331 ( .C (clk), .D (new_AGEMA_signal_13182), .Q (new_AGEMA_signal_13183) ) ;
    buf_clk new_AGEMA_reg_buffer_7334 ( .C (clk), .D (new_AGEMA_signal_13185), .Q (new_AGEMA_signal_13186) ) ;
    buf_clk new_AGEMA_reg_buffer_7337 ( .C (clk), .D (new_AGEMA_signal_13188), .Q (new_AGEMA_signal_13189) ) ;
    buf_clk new_AGEMA_reg_buffer_7340 ( .C (clk), .D (new_AGEMA_signal_13191), .Q (new_AGEMA_signal_13192) ) ;
    buf_clk new_AGEMA_reg_buffer_7343 ( .C (clk), .D (new_AGEMA_signal_13194), .Q (new_AGEMA_signal_13195) ) ;
    buf_clk new_AGEMA_reg_buffer_7346 ( .C (clk), .D (new_AGEMA_signal_13197), .Q (new_AGEMA_signal_13198) ) ;
    buf_clk new_AGEMA_reg_buffer_7349 ( .C (clk), .D (new_AGEMA_signal_13200), .Q (new_AGEMA_signal_13201) ) ;
    buf_clk new_AGEMA_reg_buffer_7352 ( .C (clk), .D (new_AGEMA_signal_13203), .Q (new_AGEMA_signal_13204) ) ;
    buf_clk new_AGEMA_reg_buffer_7355 ( .C (clk), .D (new_AGEMA_signal_13206), .Q (new_AGEMA_signal_13207) ) ;
    buf_clk new_AGEMA_reg_buffer_7358 ( .C (clk), .D (new_AGEMA_signal_13209), .Q (new_AGEMA_signal_13210) ) ;
    buf_clk new_AGEMA_reg_buffer_7361 ( .C (clk), .D (new_AGEMA_signal_13212), .Q (new_AGEMA_signal_13213) ) ;
    buf_clk new_AGEMA_reg_buffer_7364 ( .C (clk), .D (new_AGEMA_signal_13215), .Q (new_AGEMA_signal_13216) ) ;
    buf_clk new_AGEMA_reg_buffer_7367 ( .C (clk), .D (new_AGEMA_signal_13218), .Q (new_AGEMA_signal_13219) ) ;
    buf_clk new_AGEMA_reg_buffer_7370 ( .C (clk), .D (new_AGEMA_signal_13221), .Q (new_AGEMA_signal_13222) ) ;
    buf_clk new_AGEMA_reg_buffer_7373 ( .C (clk), .D (new_AGEMA_signal_13224), .Q (new_AGEMA_signal_13225) ) ;
    buf_clk new_AGEMA_reg_buffer_7376 ( .C (clk), .D (new_AGEMA_signal_13227), .Q (new_AGEMA_signal_13228) ) ;
    buf_clk new_AGEMA_reg_buffer_7379 ( .C (clk), .D (new_AGEMA_signal_13230), .Q (new_AGEMA_signal_13231) ) ;
    buf_clk new_AGEMA_reg_buffer_7382 ( .C (clk), .D (new_AGEMA_signal_13233), .Q (new_AGEMA_signal_13234) ) ;
    buf_clk new_AGEMA_reg_buffer_7385 ( .C (clk), .D (new_AGEMA_signal_13236), .Q (new_AGEMA_signal_13237) ) ;
    buf_clk new_AGEMA_reg_buffer_7388 ( .C (clk), .D (new_AGEMA_signal_13239), .Q (new_AGEMA_signal_13240) ) ;
    buf_clk new_AGEMA_reg_buffer_7391 ( .C (clk), .D (new_AGEMA_signal_13242), .Q (new_AGEMA_signal_13243) ) ;
    buf_clk new_AGEMA_reg_buffer_7394 ( .C (clk), .D (new_AGEMA_signal_13245), .Q (new_AGEMA_signal_13246) ) ;
    buf_clk new_AGEMA_reg_buffer_7397 ( .C (clk), .D (new_AGEMA_signal_13248), .Q (new_AGEMA_signal_13249) ) ;
    buf_clk new_AGEMA_reg_buffer_7400 ( .C (clk), .D (new_AGEMA_signal_13251), .Q (new_AGEMA_signal_13252) ) ;
    buf_clk new_AGEMA_reg_buffer_7403 ( .C (clk), .D (new_AGEMA_signal_13254), .Q (new_AGEMA_signal_13255) ) ;
    buf_clk new_AGEMA_reg_buffer_7406 ( .C (clk), .D (new_AGEMA_signal_13257), .Q (new_AGEMA_signal_13258) ) ;
    buf_clk new_AGEMA_reg_buffer_7409 ( .C (clk), .D (new_AGEMA_signal_13260), .Q (new_AGEMA_signal_13261) ) ;
    buf_clk new_AGEMA_reg_buffer_7412 ( .C (clk), .D (new_AGEMA_signal_13263), .Q (new_AGEMA_signal_13264) ) ;
    buf_clk new_AGEMA_reg_buffer_7415 ( .C (clk), .D (new_AGEMA_signal_13266), .Q (new_AGEMA_signal_13267) ) ;
    buf_clk new_AGEMA_reg_buffer_7418 ( .C (clk), .D (new_AGEMA_signal_13269), .Q (new_AGEMA_signal_13270) ) ;
    buf_clk new_AGEMA_reg_buffer_7421 ( .C (clk), .D (new_AGEMA_signal_13272), .Q (new_AGEMA_signal_13273) ) ;
    buf_clk new_AGEMA_reg_buffer_7424 ( .C (clk), .D (new_AGEMA_signal_13275), .Q (new_AGEMA_signal_13276) ) ;
    buf_clk new_AGEMA_reg_buffer_7427 ( .C (clk), .D (new_AGEMA_signal_13278), .Q (new_AGEMA_signal_13279) ) ;
    buf_clk new_AGEMA_reg_buffer_7430 ( .C (clk), .D (new_AGEMA_signal_13281), .Q (new_AGEMA_signal_13282) ) ;
    buf_clk new_AGEMA_reg_buffer_7433 ( .C (clk), .D (new_AGEMA_signal_13284), .Q (new_AGEMA_signal_13285) ) ;
    buf_clk new_AGEMA_reg_buffer_7436 ( .C (clk), .D (new_AGEMA_signal_13287), .Q (new_AGEMA_signal_13288) ) ;
    buf_clk new_AGEMA_reg_buffer_7439 ( .C (clk), .D (new_AGEMA_signal_13290), .Q (new_AGEMA_signal_13291) ) ;
    buf_clk new_AGEMA_reg_buffer_7442 ( .C (clk), .D (new_AGEMA_signal_13293), .Q (new_AGEMA_signal_13294) ) ;
    buf_clk new_AGEMA_reg_buffer_7445 ( .C (clk), .D (new_AGEMA_signal_13296), .Q (new_AGEMA_signal_13297) ) ;
    buf_clk new_AGEMA_reg_buffer_7448 ( .C (clk), .D (new_AGEMA_signal_13299), .Q (new_AGEMA_signal_13300) ) ;
    buf_clk new_AGEMA_reg_buffer_7451 ( .C (clk), .D (new_AGEMA_signal_13302), .Q (new_AGEMA_signal_13303) ) ;
    buf_clk new_AGEMA_reg_buffer_7454 ( .C (clk), .D (new_AGEMA_signal_13305), .Q (new_AGEMA_signal_13306) ) ;
    buf_clk new_AGEMA_reg_buffer_7457 ( .C (clk), .D (new_AGEMA_signal_13308), .Q (new_AGEMA_signal_13309) ) ;
    buf_clk new_AGEMA_reg_buffer_7460 ( .C (clk), .D (new_AGEMA_signal_13311), .Q (new_AGEMA_signal_13312) ) ;
    buf_clk new_AGEMA_reg_buffer_7463 ( .C (clk), .D (new_AGEMA_signal_13314), .Q (new_AGEMA_signal_13315) ) ;
    buf_clk new_AGEMA_reg_buffer_7466 ( .C (clk), .D (new_AGEMA_signal_13317), .Q (new_AGEMA_signal_13318) ) ;
    buf_clk new_AGEMA_reg_buffer_7469 ( .C (clk), .D (new_AGEMA_signal_13320), .Q (new_AGEMA_signal_13321) ) ;
    buf_clk new_AGEMA_reg_buffer_7472 ( .C (clk), .D (new_AGEMA_signal_13323), .Q (new_AGEMA_signal_13324) ) ;
    buf_clk new_AGEMA_reg_buffer_7475 ( .C (clk), .D (new_AGEMA_signal_13326), .Q (new_AGEMA_signal_13327) ) ;
    buf_clk new_AGEMA_reg_buffer_7479 ( .C (clk), .D (new_AGEMA_signal_13330), .Q (new_AGEMA_signal_13331) ) ;
    buf_clk new_AGEMA_reg_buffer_7483 ( .C (clk), .D (new_AGEMA_signal_13334), .Q (new_AGEMA_signal_13335) ) ;
    buf_clk new_AGEMA_reg_buffer_7487 ( .C (clk), .D (new_AGEMA_signal_13338), .Q (new_AGEMA_signal_13339) ) ;
    buf_clk new_AGEMA_reg_buffer_7491 ( .C (clk), .D (new_AGEMA_signal_13342), .Q (new_AGEMA_signal_13343) ) ;
    buf_clk new_AGEMA_reg_buffer_7495 ( .C (clk), .D (new_AGEMA_signal_13346), .Q (new_AGEMA_signal_13347) ) ;
    buf_clk new_AGEMA_reg_buffer_7499 ( .C (clk), .D (new_AGEMA_signal_13350), .Q (new_AGEMA_signal_13351) ) ;
    buf_clk new_AGEMA_reg_buffer_7503 ( .C (clk), .D (new_AGEMA_signal_13354), .Q (new_AGEMA_signal_13355) ) ;
    buf_clk new_AGEMA_reg_buffer_7507 ( .C (clk), .D (new_AGEMA_signal_13358), .Q (new_AGEMA_signal_13359) ) ;
    buf_clk new_AGEMA_reg_buffer_7511 ( .C (clk), .D (new_AGEMA_signal_13362), .Q (new_AGEMA_signal_13363) ) ;
    buf_clk new_AGEMA_reg_buffer_7515 ( .C (clk), .D (new_AGEMA_signal_13366), .Q (new_AGEMA_signal_13367) ) ;
    buf_clk new_AGEMA_reg_buffer_7519 ( .C (clk), .D (new_AGEMA_signal_13370), .Q (new_AGEMA_signal_13371) ) ;
    buf_clk new_AGEMA_reg_buffer_7523 ( .C (clk), .D (new_AGEMA_signal_13374), .Q (new_AGEMA_signal_13375) ) ;
    buf_clk new_AGEMA_reg_buffer_7527 ( .C (clk), .D (new_AGEMA_signal_13378), .Q (new_AGEMA_signal_13379) ) ;
    buf_clk new_AGEMA_reg_buffer_7531 ( .C (clk), .D (new_AGEMA_signal_13382), .Q (new_AGEMA_signal_13383) ) ;
    buf_clk new_AGEMA_reg_buffer_7535 ( .C (clk), .D (new_AGEMA_signal_13386), .Q (new_AGEMA_signal_13387) ) ;
    buf_clk new_AGEMA_reg_buffer_7539 ( .C (clk), .D (new_AGEMA_signal_13390), .Q (new_AGEMA_signal_13391) ) ;
    buf_clk new_AGEMA_reg_buffer_7543 ( .C (clk), .D (new_AGEMA_signal_13394), .Q (new_AGEMA_signal_13395) ) ;
    buf_clk new_AGEMA_reg_buffer_7547 ( .C (clk), .D (new_AGEMA_signal_13398), .Q (new_AGEMA_signal_13399) ) ;
    buf_clk new_AGEMA_reg_buffer_7551 ( .C (clk), .D (new_AGEMA_signal_13402), .Q (new_AGEMA_signal_13403) ) ;
    buf_clk new_AGEMA_reg_buffer_7555 ( .C (clk), .D (new_AGEMA_signal_13406), .Q (new_AGEMA_signal_13407) ) ;
    buf_clk new_AGEMA_reg_buffer_7559 ( .C (clk), .D (new_AGEMA_signal_13410), .Q (new_AGEMA_signal_13411) ) ;
    buf_clk new_AGEMA_reg_buffer_7563 ( .C (clk), .D (new_AGEMA_signal_13414), .Q (new_AGEMA_signal_13415) ) ;
    buf_clk new_AGEMA_reg_buffer_7567 ( .C (clk), .D (new_AGEMA_signal_13418), .Q (new_AGEMA_signal_13419) ) ;
    buf_clk new_AGEMA_reg_buffer_7571 ( .C (clk), .D (new_AGEMA_signal_13422), .Q (new_AGEMA_signal_13423) ) ;
    buf_clk new_AGEMA_reg_buffer_7575 ( .C (clk), .D (new_AGEMA_signal_13426), .Q (new_AGEMA_signal_13427) ) ;
    buf_clk new_AGEMA_reg_buffer_7579 ( .C (clk), .D (new_AGEMA_signal_13430), .Q (new_AGEMA_signal_13431) ) ;
    buf_clk new_AGEMA_reg_buffer_7583 ( .C (clk), .D (new_AGEMA_signal_13434), .Q (new_AGEMA_signal_13435) ) ;
    buf_clk new_AGEMA_reg_buffer_7587 ( .C (clk), .D (new_AGEMA_signal_13438), .Q (new_AGEMA_signal_13439) ) ;
    buf_clk new_AGEMA_reg_buffer_7591 ( .C (clk), .D (new_AGEMA_signal_13442), .Q (new_AGEMA_signal_13443) ) ;
    buf_clk new_AGEMA_reg_buffer_7595 ( .C (clk), .D (new_AGEMA_signal_13446), .Q (new_AGEMA_signal_13447) ) ;
    buf_clk new_AGEMA_reg_buffer_7599 ( .C (clk), .D (new_AGEMA_signal_13450), .Q (new_AGEMA_signal_13451) ) ;
    buf_clk new_AGEMA_reg_buffer_7603 ( .C (clk), .D (new_AGEMA_signal_13454), .Q (new_AGEMA_signal_13455) ) ;
    buf_clk new_AGEMA_reg_buffer_7607 ( .C (clk), .D (new_AGEMA_signal_13458), .Q (new_AGEMA_signal_13459) ) ;
    buf_clk new_AGEMA_reg_buffer_7611 ( .C (clk), .D (new_AGEMA_signal_13462), .Q (new_AGEMA_signal_13463) ) ;
    buf_clk new_AGEMA_reg_buffer_7615 ( .C (clk), .D (new_AGEMA_signal_13466), .Q (new_AGEMA_signal_13467) ) ;
    buf_clk new_AGEMA_reg_buffer_7619 ( .C (clk), .D (new_AGEMA_signal_13470), .Q (new_AGEMA_signal_13471) ) ;
    buf_clk new_AGEMA_reg_buffer_7623 ( .C (clk), .D (new_AGEMA_signal_13474), .Q (new_AGEMA_signal_13475) ) ;
    buf_clk new_AGEMA_reg_buffer_7627 ( .C (clk), .D (new_AGEMA_signal_13478), .Q (new_AGEMA_signal_13479) ) ;
    buf_clk new_AGEMA_reg_buffer_7631 ( .C (clk), .D (new_AGEMA_signal_13482), .Q (new_AGEMA_signal_13483) ) ;
    buf_clk new_AGEMA_reg_buffer_7635 ( .C (clk), .D (new_AGEMA_signal_13486), .Q (new_AGEMA_signal_13487) ) ;
    buf_clk new_AGEMA_reg_buffer_7639 ( .C (clk), .D (new_AGEMA_signal_13490), .Q (new_AGEMA_signal_13491) ) ;
    buf_clk new_AGEMA_reg_buffer_7643 ( .C (clk), .D (new_AGEMA_signal_13494), .Q (new_AGEMA_signal_13495) ) ;
    buf_clk new_AGEMA_reg_buffer_7647 ( .C (clk), .D (new_AGEMA_signal_13498), .Q (new_AGEMA_signal_13499) ) ;
    buf_clk new_AGEMA_reg_buffer_7651 ( .C (clk), .D (new_AGEMA_signal_13502), .Q (new_AGEMA_signal_13503) ) ;
    buf_clk new_AGEMA_reg_buffer_7655 ( .C (clk), .D (new_AGEMA_signal_13506), .Q (new_AGEMA_signal_13507) ) ;
    buf_clk new_AGEMA_reg_buffer_7659 ( .C (clk), .D (new_AGEMA_signal_13510), .Q (new_AGEMA_signal_13511) ) ;
    buf_clk new_AGEMA_reg_buffer_7663 ( .C (clk), .D (new_AGEMA_signal_13514), .Q (new_AGEMA_signal_13515) ) ;
    buf_clk new_AGEMA_reg_buffer_7667 ( .C (clk), .D (new_AGEMA_signal_13518), .Q (new_AGEMA_signal_13519) ) ;
    buf_clk new_AGEMA_reg_buffer_7671 ( .C (clk), .D (new_AGEMA_signal_13522), .Q (new_AGEMA_signal_13523) ) ;
    buf_clk new_AGEMA_reg_buffer_7675 ( .C (clk), .D (new_AGEMA_signal_13526), .Q (new_AGEMA_signal_13527) ) ;
    buf_clk new_AGEMA_reg_buffer_7679 ( .C (clk), .D (new_AGEMA_signal_13530), .Q (new_AGEMA_signal_13531) ) ;
    buf_clk new_AGEMA_reg_buffer_7683 ( .C (clk), .D (new_AGEMA_signal_13534), .Q (new_AGEMA_signal_13535) ) ;
    buf_clk new_AGEMA_reg_buffer_7687 ( .C (clk), .D (new_AGEMA_signal_13538), .Q (new_AGEMA_signal_13539) ) ;
    buf_clk new_AGEMA_reg_buffer_7691 ( .C (clk), .D (new_AGEMA_signal_13542), .Q (new_AGEMA_signal_13543) ) ;
    buf_clk new_AGEMA_reg_buffer_7695 ( .C (clk), .D (new_AGEMA_signal_13546), .Q (new_AGEMA_signal_13547) ) ;
    buf_clk new_AGEMA_reg_buffer_7699 ( .C (clk), .D (new_AGEMA_signal_13550), .Q (new_AGEMA_signal_13551) ) ;
    buf_clk new_AGEMA_reg_buffer_7703 ( .C (clk), .D (new_AGEMA_signal_13554), .Q (new_AGEMA_signal_13555) ) ;
    buf_clk new_AGEMA_reg_buffer_7707 ( .C (clk), .D (new_AGEMA_signal_13558), .Q (new_AGEMA_signal_13559) ) ;
    buf_clk new_AGEMA_reg_buffer_7711 ( .C (clk), .D (new_AGEMA_signal_13562), .Q (new_AGEMA_signal_13563) ) ;
    buf_clk new_AGEMA_reg_buffer_7715 ( .C (clk), .D (new_AGEMA_signal_13566), .Q (new_AGEMA_signal_13567) ) ;
    buf_clk new_AGEMA_reg_buffer_7719 ( .C (clk), .D (new_AGEMA_signal_13570), .Q (new_AGEMA_signal_13571) ) ;
    buf_clk new_AGEMA_reg_buffer_7723 ( .C (clk), .D (new_AGEMA_signal_13574), .Q (new_AGEMA_signal_13575) ) ;
    buf_clk new_AGEMA_reg_buffer_7727 ( .C (clk), .D (new_AGEMA_signal_13578), .Q (new_AGEMA_signal_13579) ) ;
    buf_clk new_AGEMA_reg_buffer_7731 ( .C (clk), .D (new_AGEMA_signal_13582), .Q (new_AGEMA_signal_13583) ) ;
    buf_clk new_AGEMA_reg_buffer_7735 ( .C (clk), .D (new_AGEMA_signal_13586), .Q (new_AGEMA_signal_13587) ) ;
    buf_clk new_AGEMA_reg_buffer_7739 ( .C (clk), .D (new_AGEMA_signal_13590), .Q (new_AGEMA_signal_13591) ) ;
    buf_clk new_AGEMA_reg_buffer_7743 ( .C (clk), .D (new_AGEMA_signal_13594), .Q (new_AGEMA_signal_13595) ) ;
    buf_clk new_AGEMA_reg_buffer_7747 ( .C (clk), .D (new_AGEMA_signal_13598), .Q (new_AGEMA_signal_13599) ) ;
    buf_clk new_AGEMA_reg_buffer_7751 ( .C (clk), .D (new_AGEMA_signal_13602), .Q (new_AGEMA_signal_13603) ) ;
    buf_clk new_AGEMA_reg_buffer_7755 ( .C (clk), .D (new_AGEMA_signal_13606), .Q (new_AGEMA_signal_13607) ) ;
    buf_clk new_AGEMA_reg_buffer_7759 ( .C (clk), .D (new_AGEMA_signal_13610), .Q (new_AGEMA_signal_13611) ) ;
    buf_clk new_AGEMA_reg_buffer_7763 ( .C (clk), .D (new_AGEMA_signal_13614), .Q (new_AGEMA_signal_13615) ) ;
    buf_clk new_AGEMA_reg_buffer_7767 ( .C (clk), .D (new_AGEMA_signal_13618), .Q (new_AGEMA_signal_13619) ) ;
    buf_clk new_AGEMA_reg_buffer_7771 ( .C (clk), .D (new_AGEMA_signal_13622), .Q (new_AGEMA_signal_13623) ) ;
    buf_clk new_AGEMA_reg_buffer_7775 ( .C (clk), .D (new_AGEMA_signal_13626), .Q (new_AGEMA_signal_13627) ) ;
    buf_clk new_AGEMA_reg_buffer_7779 ( .C (clk), .D (new_AGEMA_signal_13630), .Q (new_AGEMA_signal_13631) ) ;
    buf_clk new_AGEMA_reg_buffer_7783 ( .C (clk), .D (new_AGEMA_signal_13634), .Q (new_AGEMA_signal_13635) ) ;
    buf_clk new_AGEMA_reg_buffer_7787 ( .C (clk), .D (new_AGEMA_signal_13638), .Q (new_AGEMA_signal_13639) ) ;
    buf_clk new_AGEMA_reg_buffer_7791 ( .C (clk), .D (new_AGEMA_signal_13642), .Q (new_AGEMA_signal_13643) ) ;
    buf_clk new_AGEMA_reg_buffer_7795 ( .C (clk), .D (new_AGEMA_signal_13646), .Q (new_AGEMA_signal_13647) ) ;
    buf_clk new_AGEMA_reg_buffer_7799 ( .C (clk), .D (new_AGEMA_signal_13650), .Q (new_AGEMA_signal_13651) ) ;
    buf_clk new_AGEMA_reg_buffer_7803 ( .C (clk), .D (new_AGEMA_signal_13654), .Q (new_AGEMA_signal_13655) ) ;
    buf_clk new_AGEMA_reg_buffer_7807 ( .C (clk), .D (new_AGEMA_signal_13658), .Q (new_AGEMA_signal_13659) ) ;
    buf_clk new_AGEMA_reg_buffer_7811 ( .C (clk), .D (new_AGEMA_signal_13662), .Q (new_AGEMA_signal_13663) ) ;
    buf_clk new_AGEMA_reg_buffer_7815 ( .C (clk), .D (new_AGEMA_signal_13666), .Q (new_AGEMA_signal_13667) ) ;
    buf_clk new_AGEMA_reg_buffer_7819 ( .C (clk), .D (new_AGEMA_signal_13670), .Q (new_AGEMA_signal_13671) ) ;
    buf_clk new_AGEMA_reg_buffer_7823 ( .C (clk), .D (new_AGEMA_signal_13674), .Q (new_AGEMA_signal_13675) ) ;
    buf_clk new_AGEMA_reg_buffer_7827 ( .C (clk), .D (new_AGEMA_signal_13678), .Q (new_AGEMA_signal_13679) ) ;
    buf_clk new_AGEMA_reg_buffer_7831 ( .C (clk), .D (new_AGEMA_signal_13682), .Q (new_AGEMA_signal_13683) ) ;
    buf_clk new_AGEMA_reg_buffer_7835 ( .C (clk), .D (new_AGEMA_signal_13686), .Q (new_AGEMA_signal_13687) ) ;
    buf_clk new_AGEMA_reg_buffer_7839 ( .C (clk), .D (new_AGEMA_signal_13690), .Q (new_AGEMA_signal_13691) ) ;
    buf_clk new_AGEMA_reg_buffer_7843 ( .C (clk), .D (new_AGEMA_signal_13694), .Q (new_AGEMA_signal_13695) ) ;
    buf_clk new_AGEMA_reg_buffer_7847 ( .C (clk), .D (new_AGEMA_signal_13698), .Q (new_AGEMA_signal_13699) ) ;
    buf_clk new_AGEMA_reg_buffer_7851 ( .C (clk), .D (new_AGEMA_signal_13702), .Q (new_AGEMA_signal_13703) ) ;
    buf_clk new_AGEMA_reg_buffer_7855 ( .C (clk), .D (new_AGEMA_signal_13706), .Q (new_AGEMA_signal_13707) ) ;
    buf_clk new_AGEMA_reg_buffer_7859 ( .C (clk), .D (new_AGEMA_signal_13710), .Q (new_AGEMA_signal_13711) ) ;
    buf_clk new_AGEMA_reg_buffer_7863 ( .C (clk), .D (new_AGEMA_signal_13714), .Q (new_AGEMA_signal_13715) ) ;
    buf_clk new_AGEMA_reg_buffer_7867 ( .C (clk), .D (new_AGEMA_signal_13718), .Q (new_AGEMA_signal_13719) ) ;
    buf_clk new_AGEMA_reg_buffer_7871 ( .C (clk), .D (new_AGEMA_signal_13722), .Q (new_AGEMA_signal_13723) ) ;
    buf_clk new_AGEMA_reg_buffer_7875 ( .C (clk), .D (new_AGEMA_signal_13726), .Q (new_AGEMA_signal_13727) ) ;
    buf_clk new_AGEMA_reg_buffer_7879 ( .C (clk), .D (new_AGEMA_signal_13730), .Q (new_AGEMA_signal_13731) ) ;
    buf_clk new_AGEMA_reg_buffer_7883 ( .C (clk), .D (new_AGEMA_signal_13734), .Q (new_AGEMA_signal_13735) ) ;
    buf_clk new_AGEMA_reg_buffer_7887 ( .C (clk), .D (new_AGEMA_signal_13738), .Q (new_AGEMA_signal_13739) ) ;
    buf_clk new_AGEMA_reg_buffer_7891 ( .C (clk), .D (new_AGEMA_signal_13742), .Q (new_AGEMA_signal_13743) ) ;
    buf_clk new_AGEMA_reg_buffer_7895 ( .C (clk), .D (new_AGEMA_signal_13746), .Q (new_AGEMA_signal_13747) ) ;
    buf_clk new_AGEMA_reg_buffer_7899 ( .C (clk), .D (new_AGEMA_signal_13750), .Q (new_AGEMA_signal_13751) ) ;
    buf_clk new_AGEMA_reg_buffer_7903 ( .C (clk), .D (new_AGEMA_signal_13754), .Q (new_AGEMA_signal_13755) ) ;
    buf_clk new_AGEMA_reg_buffer_7907 ( .C (clk), .D (new_AGEMA_signal_13758), .Q (new_AGEMA_signal_13759) ) ;
    buf_clk new_AGEMA_reg_buffer_7911 ( .C (clk), .D (new_AGEMA_signal_13762), .Q (new_AGEMA_signal_13763) ) ;
    buf_clk new_AGEMA_reg_buffer_7915 ( .C (clk), .D (new_AGEMA_signal_13766), .Q (new_AGEMA_signal_13767) ) ;
    buf_clk new_AGEMA_reg_buffer_7919 ( .C (clk), .D (new_AGEMA_signal_13770), .Q (new_AGEMA_signal_13771) ) ;
    buf_clk new_AGEMA_reg_buffer_7923 ( .C (clk), .D (new_AGEMA_signal_13774), .Q (new_AGEMA_signal_13775) ) ;
    buf_clk new_AGEMA_reg_buffer_7927 ( .C (clk), .D (new_AGEMA_signal_13778), .Q (new_AGEMA_signal_13779) ) ;
    buf_clk new_AGEMA_reg_buffer_7931 ( .C (clk), .D (new_AGEMA_signal_13782), .Q (new_AGEMA_signal_13783) ) ;
    buf_clk new_AGEMA_reg_buffer_7935 ( .C (clk), .D (new_AGEMA_signal_13786), .Q (new_AGEMA_signal_13787) ) ;
    buf_clk new_AGEMA_reg_buffer_7939 ( .C (clk), .D (new_AGEMA_signal_13790), .Q (new_AGEMA_signal_13791) ) ;
    buf_clk new_AGEMA_reg_buffer_7943 ( .C (clk), .D (new_AGEMA_signal_13794), .Q (new_AGEMA_signal_13795) ) ;
    buf_clk new_AGEMA_reg_buffer_7947 ( .C (clk), .D (new_AGEMA_signal_13798), .Q (new_AGEMA_signal_13799) ) ;
    buf_clk new_AGEMA_reg_buffer_7951 ( .C (clk), .D (new_AGEMA_signal_13802), .Q (new_AGEMA_signal_13803) ) ;
    buf_clk new_AGEMA_reg_buffer_7955 ( .C (clk), .D (new_AGEMA_signal_13806), .Q (new_AGEMA_signal_13807) ) ;
    buf_clk new_AGEMA_reg_buffer_7959 ( .C (clk), .D (new_AGEMA_signal_13810), .Q (new_AGEMA_signal_13811) ) ;
    buf_clk new_AGEMA_reg_buffer_7963 ( .C (clk), .D (new_AGEMA_signal_13814), .Q (new_AGEMA_signal_13815) ) ;
    buf_clk new_AGEMA_reg_buffer_7967 ( .C (clk), .D (new_AGEMA_signal_13818), .Q (new_AGEMA_signal_13819) ) ;
    buf_clk new_AGEMA_reg_buffer_7971 ( .C (clk), .D (new_AGEMA_signal_13822), .Q (new_AGEMA_signal_13823) ) ;
    buf_clk new_AGEMA_reg_buffer_7975 ( .C (clk), .D (new_AGEMA_signal_13826), .Q (new_AGEMA_signal_13827) ) ;
    buf_clk new_AGEMA_reg_buffer_7979 ( .C (clk), .D (new_AGEMA_signal_13830), .Q (new_AGEMA_signal_13831) ) ;
    buf_clk new_AGEMA_reg_buffer_7983 ( .C (clk), .D (new_AGEMA_signal_13834), .Q (new_AGEMA_signal_13835) ) ;
    buf_clk new_AGEMA_reg_buffer_7987 ( .C (clk), .D (new_AGEMA_signal_13838), .Q (new_AGEMA_signal_13839) ) ;
    buf_clk new_AGEMA_reg_buffer_7991 ( .C (clk), .D (new_AGEMA_signal_13842), .Q (new_AGEMA_signal_13843) ) ;
    buf_clk new_AGEMA_reg_buffer_7995 ( .C (clk), .D (new_AGEMA_signal_13846), .Q (new_AGEMA_signal_13847) ) ;
    buf_clk new_AGEMA_reg_buffer_7999 ( .C (clk), .D (new_AGEMA_signal_13850), .Q (new_AGEMA_signal_13851) ) ;
    buf_clk new_AGEMA_reg_buffer_8003 ( .C (clk), .D (new_AGEMA_signal_13854), .Q (new_AGEMA_signal_13855) ) ;
    buf_clk new_AGEMA_reg_buffer_8007 ( .C (clk), .D (new_AGEMA_signal_13858), .Q (new_AGEMA_signal_13859) ) ;
    buf_clk new_AGEMA_reg_buffer_8011 ( .C (clk), .D (new_AGEMA_signal_13862), .Q (new_AGEMA_signal_13863) ) ;
    buf_clk new_AGEMA_reg_buffer_8015 ( .C (clk), .D (new_AGEMA_signal_13866), .Q (new_AGEMA_signal_13867) ) ;
    buf_clk new_AGEMA_reg_buffer_8019 ( .C (clk), .D (new_AGEMA_signal_13870), .Q (new_AGEMA_signal_13871) ) ;
    buf_clk new_AGEMA_reg_buffer_8023 ( .C (clk), .D (new_AGEMA_signal_13874), .Q (new_AGEMA_signal_13875) ) ;
    buf_clk new_AGEMA_reg_buffer_8027 ( .C (clk), .D (new_AGEMA_signal_13878), .Q (new_AGEMA_signal_13879) ) ;
    buf_clk new_AGEMA_reg_buffer_8031 ( .C (clk), .D (new_AGEMA_signal_13882), .Q (new_AGEMA_signal_13883) ) ;
    buf_clk new_AGEMA_reg_buffer_8035 ( .C (clk), .D (new_AGEMA_signal_13886), .Q (new_AGEMA_signal_13887) ) ;
    buf_clk new_AGEMA_reg_buffer_8039 ( .C (clk), .D (new_AGEMA_signal_13890), .Q (new_AGEMA_signal_13891) ) ;
    buf_clk new_AGEMA_reg_buffer_8043 ( .C (clk), .D (new_AGEMA_signal_13894), .Q (new_AGEMA_signal_13895) ) ;
    buf_clk new_AGEMA_reg_buffer_8047 ( .C (clk), .D (new_AGEMA_signal_13898), .Q (new_AGEMA_signal_13899) ) ;
    buf_clk new_AGEMA_reg_buffer_8051 ( .C (clk), .D (new_AGEMA_signal_13902), .Q (new_AGEMA_signal_13903) ) ;
    buf_clk new_AGEMA_reg_buffer_8055 ( .C (clk), .D (new_AGEMA_signal_13906), .Q (new_AGEMA_signal_13907) ) ;
    buf_clk new_AGEMA_reg_buffer_8059 ( .C (clk), .D (new_AGEMA_signal_13910), .Q (new_AGEMA_signal_13911) ) ;
    buf_clk new_AGEMA_reg_buffer_8063 ( .C (clk), .D (new_AGEMA_signal_13914), .Q (new_AGEMA_signal_13915) ) ;
    buf_clk new_AGEMA_reg_buffer_8067 ( .C (clk), .D (new_AGEMA_signal_13918), .Q (new_AGEMA_signal_13919) ) ;
    buf_clk new_AGEMA_reg_buffer_8071 ( .C (clk), .D (new_AGEMA_signal_13922), .Q (new_AGEMA_signal_13923) ) ;
    buf_clk new_AGEMA_reg_buffer_8075 ( .C (clk), .D (new_AGEMA_signal_13926), .Q (new_AGEMA_signal_13927) ) ;
    buf_clk new_AGEMA_reg_buffer_8079 ( .C (clk), .D (new_AGEMA_signal_13930), .Q (new_AGEMA_signal_13931) ) ;
    buf_clk new_AGEMA_reg_buffer_8083 ( .C (clk), .D (new_AGEMA_signal_13934), .Q (new_AGEMA_signal_13935) ) ;
    buf_clk new_AGEMA_reg_buffer_8087 ( .C (clk), .D (new_AGEMA_signal_13938), .Q (new_AGEMA_signal_13939) ) ;
    buf_clk new_AGEMA_reg_buffer_8091 ( .C (clk), .D (new_AGEMA_signal_13942), .Q (new_AGEMA_signal_13943) ) ;
    buf_clk new_AGEMA_reg_buffer_8095 ( .C (clk), .D (new_AGEMA_signal_13946), .Q (new_AGEMA_signal_13947) ) ;
    buf_clk new_AGEMA_reg_buffer_8099 ( .C (clk), .D (new_AGEMA_signal_13950), .Q (new_AGEMA_signal_13951) ) ;
    buf_clk new_AGEMA_reg_buffer_8103 ( .C (clk), .D (new_AGEMA_signal_13954), .Q (new_AGEMA_signal_13955) ) ;
    buf_clk new_AGEMA_reg_buffer_8107 ( .C (clk), .D (new_AGEMA_signal_13958), .Q (new_AGEMA_signal_13959) ) ;
    buf_clk new_AGEMA_reg_buffer_8111 ( .C (clk), .D (new_AGEMA_signal_13962), .Q (new_AGEMA_signal_13963) ) ;
    buf_clk new_AGEMA_reg_buffer_8115 ( .C (clk), .D (new_AGEMA_signal_13966), .Q (new_AGEMA_signal_13967) ) ;
    buf_clk new_AGEMA_reg_buffer_8119 ( .C (clk), .D (new_AGEMA_signal_13970), .Q (new_AGEMA_signal_13971) ) ;
    buf_clk new_AGEMA_reg_buffer_8123 ( .C (clk), .D (new_AGEMA_signal_13974), .Q (new_AGEMA_signal_13975) ) ;
    buf_clk new_AGEMA_reg_buffer_8127 ( .C (clk), .D (new_AGEMA_signal_13978), .Q (new_AGEMA_signal_13979) ) ;
    buf_clk new_AGEMA_reg_buffer_8131 ( .C (clk), .D (new_AGEMA_signal_13982), .Q (new_AGEMA_signal_13983) ) ;
    buf_clk new_AGEMA_reg_buffer_8135 ( .C (clk), .D (new_AGEMA_signal_13986), .Q (new_AGEMA_signal_13987) ) ;
    buf_clk new_AGEMA_reg_buffer_8139 ( .C (clk), .D (new_AGEMA_signal_13990), .Q (new_AGEMA_signal_13991) ) ;
    buf_clk new_AGEMA_reg_buffer_8143 ( .C (clk), .D (new_AGEMA_signal_13994), .Q (new_AGEMA_signal_13995) ) ;
    buf_clk new_AGEMA_reg_buffer_8147 ( .C (clk), .D (new_AGEMA_signal_13998), .Q (new_AGEMA_signal_13999) ) ;
    buf_clk new_AGEMA_reg_buffer_8151 ( .C (clk), .D (new_AGEMA_signal_14002), .Q (new_AGEMA_signal_14003) ) ;
    buf_clk new_AGEMA_reg_buffer_8155 ( .C (clk), .D (new_AGEMA_signal_14006), .Q (new_AGEMA_signal_14007) ) ;
    buf_clk new_AGEMA_reg_buffer_8159 ( .C (clk), .D (new_AGEMA_signal_14010), .Q (new_AGEMA_signal_14011) ) ;
    buf_clk new_AGEMA_reg_buffer_8163 ( .C (clk), .D (new_AGEMA_signal_14014), .Q (new_AGEMA_signal_14015) ) ;
    buf_clk new_AGEMA_reg_buffer_8167 ( .C (clk), .D (new_AGEMA_signal_14018), .Q (new_AGEMA_signal_14019) ) ;
    buf_clk new_AGEMA_reg_buffer_8171 ( .C (clk), .D (new_AGEMA_signal_14022), .Q (new_AGEMA_signal_14023) ) ;
    buf_clk new_AGEMA_reg_buffer_8175 ( .C (clk), .D (new_AGEMA_signal_14026), .Q (new_AGEMA_signal_14027) ) ;
    buf_clk new_AGEMA_reg_buffer_8179 ( .C (clk), .D (new_AGEMA_signal_14030), .Q (new_AGEMA_signal_14031) ) ;
    buf_clk new_AGEMA_reg_buffer_8183 ( .C (clk), .D (new_AGEMA_signal_14034), .Q (new_AGEMA_signal_14035) ) ;
    buf_clk new_AGEMA_reg_buffer_8187 ( .C (clk), .D (new_AGEMA_signal_14038), .Q (new_AGEMA_signal_14039) ) ;
    buf_clk new_AGEMA_reg_buffer_8191 ( .C (clk), .D (new_AGEMA_signal_14042), .Q (new_AGEMA_signal_14043) ) ;
    buf_clk new_AGEMA_reg_buffer_8195 ( .C (clk), .D (new_AGEMA_signal_14046), .Q (new_AGEMA_signal_14047) ) ;
    buf_clk new_AGEMA_reg_buffer_8199 ( .C (clk), .D (new_AGEMA_signal_14050), .Q (new_AGEMA_signal_14051) ) ;
    buf_clk new_AGEMA_reg_buffer_8203 ( .C (clk), .D (new_AGEMA_signal_14054), .Q (new_AGEMA_signal_14055) ) ;
    buf_clk new_AGEMA_reg_buffer_8207 ( .C (clk), .D (new_AGEMA_signal_14058), .Q (new_AGEMA_signal_14059) ) ;
    buf_clk new_AGEMA_reg_buffer_8211 ( .C (clk), .D (new_AGEMA_signal_14062), .Q (new_AGEMA_signal_14063) ) ;
    buf_clk new_AGEMA_reg_buffer_8215 ( .C (clk), .D (new_AGEMA_signal_14066), .Q (new_AGEMA_signal_14067) ) ;
    buf_clk new_AGEMA_reg_buffer_8219 ( .C (clk), .D (new_AGEMA_signal_14070), .Q (new_AGEMA_signal_14071) ) ;
    buf_clk new_AGEMA_reg_buffer_8223 ( .C (clk), .D (new_AGEMA_signal_14074), .Q (new_AGEMA_signal_14075) ) ;
    buf_clk new_AGEMA_reg_buffer_8227 ( .C (clk), .D (new_AGEMA_signal_14078), .Q (new_AGEMA_signal_14079) ) ;
    buf_clk new_AGEMA_reg_buffer_8231 ( .C (clk), .D (new_AGEMA_signal_14082), .Q (new_AGEMA_signal_14083) ) ;
    buf_clk new_AGEMA_reg_buffer_8235 ( .C (clk), .D (new_AGEMA_signal_14086), .Q (new_AGEMA_signal_14087) ) ;
    buf_clk new_AGEMA_reg_buffer_8239 ( .C (clk), .D (new_AGEMA_signal_14090), .Q (new_AGEMA_signal_14091) ) ;
    buf_clk new_AGEMA_reg_buffer_8243 ( .C (clk), .D (new_AGEMA_signal_14094), .Q (new_AGEMA_signal_14095) ) ;
    buf_clk new_AGEMA_reg_buffer_8247 ( .C (clk), .D (new_AGEMA_signal_14098), .Q (new_AGEMA_signal_14099) ) ;
    buf_clk new_AGEMA_reg_buffer_8251 ( .C (clk), .D (new_AGEMA_signal_14102), .Q (new_AGEMA_signal_14103) ) ;
    buf_clk new_AGEMA_reg_buffer_8255 ( .C (clk), .D (new_AGEMA_signal_14106), .Q (new_AGEMA_signal_14107) ) ;
    buf_clk new_AGEMA_reg_buffer_8259 ( .C (clk), .D (new_AGEMA_signal_14110), .Q (new_AGEMA_signal_14111) ) ;
    buf_clk new_AGEMA_reg_buffer_8263 ( .C (clk), .D (new_AGEMA_signal_14114), .Q (new_AGEMA_signal_14115) ) ;
    buf_clk new_AGEMA_reg_buffer_8267 ( .C (clk), .D (new_AGEMA_signal_14118), .Q (new_AGEMA_signal_14119) ) ;
    buf_clk new_AGEMA_reg_buffer_8271 ( .C (clk), .D (new_AGEMA_signal_14122), .Q (new_AGEMA_signal_14123) ) ;
    buf_clk new_AGEMA_reg_buffer_8275 ( .C (clk), .D (new_AGEMA_signal_14126), .Q (new_AGEMA_signal_14127) ) ;
    buf_clk new_AGEMA_reg_buffer_8279 ( .C (clk), .D (new_AGEMA_signal_14130), .Q (new_AGEMA_signal_14131) ) ;
    buf_clk new_AGEMA_reg_buffer_8283 ( .C (clk), .D (new_AGEMA_signal_14134), .Q (new_AGEMA_signal_14135) ) ;
    buf_clk new_AGEMA_reg_buffer_8287 ( .C (clk), .D (new_AGEMA_signal_14138), .Q (new_AGEMA_signal_14139) ) ;
    buf_clk new_AGEMA_reg_buffer_8291 ( .C (clk), .D (new_AGEMA_signal_14142), .Q (new_AGEMA_signal_14143) ) ;
    buf_clk new_AGEMA_reg_buffer_8295 ( .C (clk), .D (new_AGEMA_signal_14146), .Q (new_AGEMA_signal_14147) ) ;
    buf_clk new_AGEMA_reg_buffer_8299 ( .C (clk), .D (new_AGEMA_signal_14150), .Q (new_AGEMA_signal_14151) ) ;
    buf_clk new_AGEMA_reg_buffer_8303 ( .C (clk), .D (new_AGEMA_signal_14154), .Q (new_AGEMA_signal_14155) ) ;
    buf_clk new_AGEMA_reg_buffer_8307 ( .C (clk), .D (new_AGEMA_signal_14158), .Q (new_AGEMA_signal_14159) ) ;
    buf_clk new_AGEMA_reg_buffer_8311 ( .C (clk), .D (new_AGEMA_signal_14162), .Q (new_AGEMA_signal_14163) ) ;
    buf_clk new_AGEMA_reg_buffer_8315 ( .C (clk), .D (new_AGEMA_signal_14166), .Q (new_AGEMA_signal_14167) ) ;
    buf_clk new_AGEMA_reg_buffer_8319 ( .C (clk), .D (new_AGEMA_signal_14170), .Q (new_AGEMA_signal_14171) ) ;
    buf_clk new_AGEMA_reg_buffer_8323 ( .C (clk), .D (new_AGEMA_signal_14174), .Q (new_AGEMA_signal_14175) ) ;
    buf_clk new_AGEMA_reg_buffer_8327 ( .C (clk), .D (new_AGEMA_signal_14178), .Q (new_AGEMA_signal_14179) ) ;
    buf_clk new_AGEMA_reg_buffer_8331 ( .C (clk), .D (new_AGEMA_signal_14182), .Q (new_AGEMA_signal_14183) ) ;
    buf_clk new_AGEMA_reg_buffer_8335 ( .C (clk), .D (new_AGEMA_signal_14186), .Q (new_AGEMA_signal_14187) ) ;
    buf_clk new_AGEMA_reg_buffer_8339 ( .C (clk), .D (new_AGEMA_signal_14190), .Q (new_AGEMA_signal_14191) ) ;
    buf_clk new_AGEMA_reg_buffer_8343 ( .C (clk), .D (new_AGEMA_signal_14194), .Q (new_AGEMA_signal_14195) ) ;
    buf_clk new_AGEMA_reg_buffer_8347 ( .C (clk), .D (new_AGEMA_signal_14198), .Q (new_AGEMA_signal_14199) ) ;
    buf_clk new_AGEMA_reg_buffer_8351 ( .C (clk), .D (new_AGEMA_signal_14202), .Q (new_AGEMA_signal_14203) ) ;
    buf_clk new_AGEMA_reg_buffer_8355 ( .C (clk), .D (new_AGEMA_signal_14206), .Q (new_AGEMA_signal_14207) ) ;
    buf_clk new_AGEMA_reg_buffer_8359 ( .C (clk), .D (new_AGEMA_signal_14210), .Q (new_AGEMA_signal_14211) ) ;
    buf_clk new_AGEMA_reg_buffer_8363 ( .C (clk), .D (new_AGEMA_signal_14214), .Q (new_AGEMA_signal_14215) ) ;
    buf_clk new_AGEMA_reg_buffer_8367 ( .C (clk), .D (new_AGEMA_signal_14218), .Q (new_AGEMA_signal_14219) ) ;
    buf_clk new_AGEMA_reg_buffer_8371 ( .C (clk), .D (new_AGEMA_signal_14222), .Q (new_AGEMA_signal_14223) ) ;
    buf_clk new_AGEMA_reg_buffer_8375 ( .C (clk), .D (new_AGEMA_signal_14226), .Q (new_AGEMA_signal_14227) ) ;
    buf_clk new_AGEMA_reg_buffer_8379 ( .C (clk), .D (new_AGEMA_signal_14230), .Q (new_AGEMA_signal_14231) ) ;
    buf_clk new_AGEMA_reg_buffer_8383 ( .C (clk), .D (new_AGEMA_signal_14234), .Q (new_AGEMA_signal_14235) ) ;
    buf_clk new_AGEMA_reg_buffer_8387 ( .C (clk), .D (new_AGEMA_signal_14238), .Q (new_AGEMA_signal_14239) ) ;
    buf_clk new_AGEMA_reg_buffer_8391 ( .C (clk), .D (new_AGEMA_signal_14242), .Q (new_AGEMA_signal_14243) ) ;
    buf_clk new_AGEMA_reg_buffer_8395 ( .C (clk), .D (new_AGEMA_signal_14246), .Q (new_AGEMA_signal_14247) ) ;
    buf_clk new_AGEMA_reg_buffer_8399 ( .C (clk), .D (new_AGEMA_signal_14250), .Q (new_AGEMA_signal_14251) ) ;
    buf_clk new_AGEMA_reg_buffer_8403 ( .C (clk), .D (new_AGEMA_signal_14254), .Q (new_AGEMA_signal_14255) ) ;
    buf_clk new_AGEMA_reg_buffer_8407 ( .C (clk), .D (new_AGEMA_signal_14258), .Q (new_AGEMA_signal_14259) ) ;
    buf_clk new_AGEMA_reg_buffer_8411 ( .C (clk), .D (new_AGEMA_signal_14262), .Q (new_AGEMA_signal_14263) ) ;
    buf_clk new_AGEMA_reg_buffer_8415 ( .C (clk), .D (new_AGEMA_signal_14266), .Q (new_AGEMA_signal_14267) ) ;
    buf_clk new_AGEMA_reg_buffer_8419 ( .C (clk), .D (new_AGEMA_signal_14270), .Q (new_AGEMA_signal_14271) ) ;
    buf_clk new_AGEMA_reg_buffer_8423 ( .C (clk), .D (new_AGEMA_signal_14274), .Q (new_AGEMA_signal_14275) ) ;
    buf_clk new_AGEMA_reg_buffer_8427 ( .C (clk), .D (new_AGEMA_signal_14278), .Q (new_AGEMA_signal_14279) ) ;
    buf_clk new_AGEMA_reg_buffer_8431 ( .C (clk), .D (new_AGEMA_signal_14282), .Q (new_AGEMA_signal_14283) ) ;
    buf_clk new_AGEMA_reg_buffer_8435 ( .C (clk), .D (new_AGEMA_signal_14286), .Q (new_AGEMA_signal_14287) ) ;
    buf_clk new_AGEMA_reg_buffer_8439 ( .C (clk), .D (new_AGEMA_signal_14290), .Q (new_AGEMA_signal_14291) ) ;
    buf_clk new_AGEMA_reg_buffer_8443 ( .C (clk), .D (new_AGEMA_signal_14294), .Q (new_AGEMA_signal_14295) ) ;
    buf_clk new_AGEMA_reg_buffer_8447 ( .C (clk), .D (new_AGEMA_signal_14298), .Q (new_AGEMA_signal_14299) ) ;
    buf_clk new_AGEMA_reg_buffer_8451 ( .C (clk), .D (new_AGEMA_signal_14302), .Q (new_AGEMA_signal_14303) ) ;
    buf_clk new_AGEMA_reg_buffer_8455 ( .C (clk), .D (new_AGEMA_signal_14306), .Q (new_AGEMA_signal_14307) ) ;
    buf_clk new_AGEMA_reg_buffer_8459 ( .C (clk), .D (new_AGEMA_signal_14310), .Q (new_AGEMA_signal_14311) ) ;
    buf_clk new_AGEMA_reg_buffer_8463 ( .C (clk), .D (new_AGEMA_signal_14314), .Q (new_AGEMA_signal_14315) ) ;
    buf_clk new_AGEMA_reg_buffer_8467 ( .C (clk), .D (new_AGEMA_signal_14318), .Q (new_AGEMA_signal_14319) ) ;
    buf_clk new_AGEMA_reg_buffer_8471 ( .C (clk), .D (new_AGEMA_signal_14322), .Q (new_AGEMA_signal_14323) ) ;
    buf_clk new_AGEMA_reg_buffer_8475 ( .C (clk), .D (new_AGEMA_signal_14326), .Q (new_AGEMA_signal_14327) ) ;
    buf_clk new_AGEMA_reg_buffer_8479 ( .C (clk), .D (new_AGEMA_signal_14330), .Q (new_AGEMA_signal_14331) ) ;
    buf_clk new_AGEMA_reg_buffer_8483 ( .C (clk), .D (new_AGEMA_signal_14334), .Q (new_AGEMA_signal_14335) ) ;
    buf_clk new_AGEMA_reg_buffer_8487 ( .C (clk), .D (new_AGEMA_signal_14338), .Q (new_AGEMA_signal_14339) ) ;
    buf_clk new_AGEMA_reg_buffer_8491 ( .C (clk), .D (new_AGEMA_signal_14342), .Q (new_AGEMA_signal_14343) ) ;
    buf_clk new_AGEMA_reg_buffer_8495 ( .C (clk), .D (new_AGEMA_signal_14346), .Q (new_AGEMA_signal_14347) ) ;
    buf_clk new_AGEMA_reg_buffer_8499 ( .C (clk), .D (new_AGEMA_signal_14350), .Q (new_AGEMA_signal_14351) ) ;
    buf_clk new_AGEMA_reg_buffer_8503 ( .C (clk), .D (new_AGEMA_signal_14354), .Q (new_AGEMA_signal_14355) ) ;
    buf_clk new_AGEMA_reg_buffer_8507 ( .C (clk), .D (new_AGEMA_signal_14358), .Q (new_AGEMA_signal_14359) ) ;
    buf_clk new_AGEMA_reg_buffer_8511 ( .C (clk), .D (new_AGEMA_signal_14362), .Q (new_AGEMA_signal_14363) ) ;
    buf_clk new_AGEMA_reg_buffer_8515 ( .C (clk), .D (new_AGEMA_signal_14366), .Q (new_AGEMA_signal_14367) ) ;
    buf_clk new_AGEMA_reg_buffer_8519 ( .C (clk), .D (new_AGEMA_signal_14370), .Q (new_AGEMA_signal_14371) ) ;
    buf_clk new_AGEMA_reg_buffer_8523 ( .C (clk), .D (new_AGEMA_signal_14374), .Q (new_AGEMA_signal_14375) ) ;
    buf_clk new_AGEMA_reg_buffer_8527 ( .C (clk), .D (new_AGEMA_signal_14378), .Q (new_AGEMA_signal_14379) ) ;
    buf_clk new_AGEMA_reg_buffer_8531 ( .C (clk), .D (new_AGEMA_signal_14382), .Q (new_AGEMA_signal_14383) ) ;
    buf_clk new_AGEMA_reg_buffer_8535 ( .C (clk), .D (new_AGEMA_signal_14386), .Q (new_AGEMA_signal_14387) ) ;
    buf_clk new_AGEMA_reg_buffer_8539 ( .C (clk), .D (new_AGEMA_signal_14390), .Q (new_AGEMA_signal_14391) ) ;
    buf_clk new_AGEMA_reg_buffer_8543 ( .C (clk), .D (new_AGEMA_signal_14394), .Q (new_AGEMA_signal_14395) ) ;
    buf_clk new_AGEMA_reg_buffer_8547 ( .C (clk), .D (new_AGEMA_signal_14398), .Q (new_AGEMA_signal_14399) ) ;
    buf_clk new_AGEMA_reg_buffer_8551 ( .C (clk), .D (new_AGEMA_signal_14402), .Q (new_AGEMA_signal_14403) ) ;
    buf_clk new_AGEMA_reg_buffer_8555 ( .C (clk), .D (new_AGEMA_signal_14406), .Q (new_AGEMA_signal_14407) ) ;
    buf_clk new_AGEMA_reg_buffer_8559 ( .C (clk), .D (new_AGEMA_signal_14410), .Q (new_AGEMA_signal_14411) ) ;
    buf_clk new_AGEMA_reg_buffer_8563 ( .C (clk), .D (new_AGEMA_signal_14414), .Q (new_AGEMA_signal_14415) ) ;
    buf_clk new_AGEMA_reg_buffer_8567 ( .C (clk), .D (new_AGEMA_signal_14418), .Q (new_AGEMA_signal_14419) ) ;
    buf_clk new_AGEMA_reg_buffer_8571 ( .C (clk), .D (new_AGEMA_signal_14422), .Q (new_AGEMA_signal_14423) ) ;
    buf_clk new_AGEMA_reg_buffer_8575 ( .C (clk), .D (new_AGEMA_signal_14426), .Q (new_AGEMA_signal_14427) ) ;
    buf_clk new_AGEMA_reg_buffer_8579 ( .C (clk), .D (new_AGEMA_signal_14430), .Q (new_AGEMA_signal_14431) ) ;
    buf_clk new_AGEMA_reg_buffer_8583 ( .C (clk), .D (new_AGEMA_signal_14434), .Q (new_AGEMA_signal_14435) ) ;
    buf_clk new_AGEMA_reg_buffer_8587 ( .C (clk), .D (new_AGEMA_signal_14438), .Q (new_AGEMA_signal_14439) ) ;
    buf_clk new_AGEMA_reg_buffer_8591 ( .C (clk), .D (new_AGEMA_signal_14442), .Q (new_AGEMA_signal_14443) ) ;
    buf_clk new_AGEMA_reg_buffer_8595 ( .C (clk), .D (new_AGEMA_signal_14446), .Q (new_AGEMA_signal_14447) ) ;
    buf_clk new_AGEMA_reg_buffer_8599 ( .C (clk), .D (new_AGEMA_signal_14450), .Q (new_AGEMA_signal_14451) ) ;
    buf_clk new_AGEMA_reg_buffer_8603 ( .C (clk), .D (new_AGEMA_signal_14454), .Q (new_AGEMA_signal_14455) ) ;
    buf_clk new_AGEMA_reg_buffer_8607 ( .C (clk), .D (new_AGEMA_signal_14458), .Q (new_AGEMA_signal_14459) ) ;
    buf_clk new_AGEMA_reg_buffer_8611 ( .C (clk), .D (new_AGEMA_signal_14462), .Q (new_AGEMA_signal_14463) ) ;
    buf_clk new_AGEMA_reg_buffer_8615 ( .C (clk), .D (new_AGEMA_signal_14466), .Q (new_AGEMA_signal_14467) ) ;
    buf_clk new_AGEMA_reg_buffer_8619 ( .C (clk), .D (new_AGEMA_signal_14470), .Q (new_AGEMA_signal_14471) ) ;
    buf_clk new_AGEMA_reg_buffer_8623 ( .C (clk), .D (new_AGEMA_signal_14474), .Q (new_AGEMA_signal_14475) ) ;
    buf_clk new_AGEMA_reg_buffer_8627 ( .C (clk), .D (new_AGEMA_signal_14478), .Q (new_AGEMA_signal_14479) ) ;
    buf_clk new_AGEMA_reg_buffer_8631 ( .C (clk), .D (new_AGEMA_signal_14482), .Q (new_AGEMA_signal_14483) ) ;
    buf_clk new_AGEMA_reg_buffer_8635 ( .C (clk), .D (new_AGEMA_signal_14486), .Q (new_AGEMA_signal_14487) ) ;
    buf_clk new_AGEMA_reg_buffer_8639 ( .C (clk), .D (new_AGEMA_signal_14490), .Q (new_AGEMA_signal_14491) ) ;
    buf_clk new_AGEMA_reg_buffer_8643 ( .C (clk), .D (new_AGEMA_signal_14494), .Q (new_AGEMA_signal_14495) ) ;
    buf_clk new_AGEMA_reg_buffer_8647 ( .C (clk), .D (new_AGEMA_signal_14498), .Q (new_AGEMA_signal_14499) ) ;
    buf_clk new_AGEMA_reg_buffer_8651 ( .C (clk), .D (new_AGEMA_signal_14502), .Q (new_AGEMA_signal_14503) ) ;
    buf_clk new_AGEMA_reg_buffer_8655 ( .C (clk), .D (new_AGEMA_signal_14506), .Q (new_AGEMA_signal_14507) ) ;
    buf_clk new_AGEMA_reg_buffer_8659 ( .C (clk), .D (new_AGEMA_signal_14510), .Q (new_AGEMA_signal_14511) ) ;
    buf_clk new_AGEMA_reg_buffer_8663 ( .C (clk), .D (new_AGEMA_signal_14514), .Q (new_AGEMA_signal_14515) ) ;
    buf_clk new_AGEMA_reg_buffer_8667 ( .C (clk), .D (new_AGEMA_signal_14518), .Q (new_AGEMA_signal_14519) ) ;
    buf_clk new_AGEMA_reg_buffer_8671 ( .C (clk), .D (new_AGEMA_signal_14522), .Q (new_AGEMA_signal_14523) ) ;
    buf_clk new_AGEMA_reg_buffer_8675 ( .C (clk), .D (new_AGEMA_signal_14526), .Q (new_AGEMA_signal_14527) ) ;
    buf_clk new_AGEMA_reg_buffer_8679 ( .C (clk), .D (new_AGEMA_signal_14530), .Q (new_AGEMA_signal_14531) ) ;
    buf_clk new_AGEMA_reg_buffer_8683 ( .C (clk), .D (new_AGEMA_signal_14534), .Q (new_AGEMA_signal_14535) ) ;
    buf_clk new_AGEMA_reg_buffer_8687 ( .C (clk), .D (new_AGEMA_signal_14538), .Q (new_AGEMA_signal_14539) ) ;
    buf_clk new_AGEMA_reg_buffer_8691 ( .C (clk), .D (new_AGEMA_signal_14542), .Q (new_AGEMA_signal_14543) ) ;
    buf_clk new_AGEMA_reg_buffer_8695 ( .C (clk), .D (new_AGEMA_signal_14546), .Q (new_AGEMA_signal_14547) ) ;
    buf_clk new_AGEMA_reg_buffer_8699 ( .C (clk), .D (new_AGEMA_signal_14550), .Q (new_AGEMA_signal_14551) ) ;
    buf_clk new_AGEMA_reg_buffer_8703 ( .C (clk), .D (new_AGEMA_signal_14554), .Q (new_AGEMA_signal_14555) ) ;
    buf_clk new_AGEMA_reg_buffer_8707 ( .C (clk), .D (new_AGEMA_signal_14558), .Q (new_AGEMA_signal_14559) ) ;
    buf_clk new_AGEMA_reg_buffer_8711 ( .C (clk), .D (new_AGEMA_signal_14562), .Q (new_AGEMA_signal_14563) ) ;
    buf_clk new_AGEMA_reg_buffer_8715 ( .C (clk), .D (new_AGEMA_signal_14566), .Q (new_AGEMA_signal_14567) ) ;
    buf_clk new_AGEMA_reg_buffer_8719 ( .C (clk), .D (new_AGEMA_signal_14570), .Q (new_AGEMA_signal_14571) ) ;
    buf_clk new_AGEMA_reg_buffer_8723 ( .C (clk), .D (new_AGEMA_signal_14574), .Q (new_AGEMA_signal_14575) ) ;
    buf_clk new_AGEMA_reg_buffer_8727 ( .C (clk), .D (new_AGEMA_signal_14578), .Q (new_AGEMA_signal_14579) ) ;
    buf_clk new_AGEMA_reg_buffer_8731 ( .C (clk), .D (new_AGEMA_signal_14582), .Q (new_AGEMA_signal_14583) ) ;
    buf_clk new_AGEMA_reg_buffer_8735 ( .C (clk), .D (new_AGEMA_signal_14586), .Q (new_AGEMA_signal_14587) ) ;
    buf_clk new_AGEMA_reg_buffer_8739 ( .C (clk), .D (new_AGEMA_signal_14590), .Q (new_AGEMA_signal_14591) ) ;
    buf_clk new_AGEMA_reg_buffer_8743 ( .C (clk), .D (new_AGEMA_signal_14594), .Q (new_AGEMA_signal_14595) ) ;
    buf_clk new_AGEMA_reg_buffer_8747 ( .C (clk), .D (new_AGEMA_signal_14598), .Q (new_AGEMA_signal_14599) ) ;
    buf_clk new_AGEMA_reg_buffer_8751 ( .C (clk), .D (new_AGEMA_signal_14602), .Q (new_AGEMA_signal_14603) ) ;
    buf_clk new_AGEMA_reg_buffer_8755 ( .C (clk), .D (new_AGEMA_signal_14606), .Q (new_AGEMA_signal_14607) ) ;
    buf_clk new_AGEMA_reg_buffer_8759 ( .C (clk), .D (new_AGEMA_signal_14610), .Q (new_AGEMA_signal_14611) ) ;
    buf_clk new_AGEMA_reg_buffer_8763 ( .C (clk), .D (new_AGEMA_signal_14614), .Q (new_AGEMA_signal_14615) ) ;
    buf_clk new_AGEMA_reg_buffer_8767 ( .C (clk), .D (new_AGEMA_signal_14618), .Q (new_AGEMA_signal_14619) ) ;
    buf_clk new_AGEMA_reg_buffer_8771 ( .C (clk), .D (new_AGEMA_signal_14622), .Q (new_AGEMA_signal_14623) ) ;
    buf_clk new_AGEMA_reg_buffer_8775 ( .C (clk), .D (new_AGEMA_signal_14626), .Q (new_AGEMA_signal_14627) ) ;
    buf_clk new_AGEMA_reg_buffer_8779 ( .C (clk), .D (new_AGEMA_signal_14630), .Q (new_AGEMA_signal_14631) ) ;
    buf_clk new_AGEMA_reg_buffer_8783 ( .C (clk), .D (new_AGEMA_signal_14634), .Q (new_AGEMA_signal_14635) ) ;
    buf_clk new_AGEMA_reg_buffer_8787 ( .C (clk), .D (new_AGEMA_signal_14638), .Q (new_AGEMA_signal_14639) ) ;
    buf_clk new_AGEMA_reg_buffer_8791 ( .C (clk), .D (new_AGEMA_signal_14642), .Q (new_AGEMA_signal_14643) ) ;
    buf_clk new_AGEMA_reg_buffer_8795 ( .C (clk), .D (new_AGEMA_signal_14646), .Q (new_AGEMA_signal_14647) ) ;
    buf_clk new_AGEMA_reg_buffer_8799 ( .C (clk), .D (new_AGEMA_signal_14650), .Q (new_AGEMA_signal_14651) ) ;
    buf_clk new_AGEMA_reg_buffer_8803 ( .C (clk), .D (new_AGEMA_signal_14654), .Q (new_AGEMA_signal_14655) ) ;
    buf_clk new_AGEMA_reg_buffer_8807 ( .C (clk), .D (new_AGEMA_signal_14658), .Q (new_AGEMA_signal_14659) ) ;
    buf_clk new_AGEMA_reg_buffer_8811 ( .C (clk), .D (new_AGEMA_signal_14662), .Q (new_AGEMA_signal_14663) ) ;
    buf_clk new_AGEMA_reg_buffer_8815 ( .C (clk), .D (new_AGEMA_signal_14666), .Q (new_AGEMA_signal_14667) ) ;
    buf_clk new_AGEMA_reg_buffer_8819 ( .C (clk), .D (new_AGEMA_signal_14670), .Q (new_AGEMA_signal_14671) ) ;
    buf_clk new_AGEMA_reg_buffer_8823 ( .C (clk), .D (new_AGEMA_signal_14674), .Q (new_AGEMA_signal_14675) ) ;
    buf_clk new_AGEMA_reg_buffer_8827 ( .C (clk), .D (new_AGEMA_signal_14678), .Q (new_AGEMA_signal_14679) ) ;
    buf_clk new_AGEMA_reg_buffer_8831 ( .C (clk), .D (new_AGEMA_signal_14682), .Q (new_AGEMA_signal_14683) ) ;
    buf_clk new_AGEMA_reg_buffer_8835 ( .C (clk), .D (new_AGEMA_signal_14686), .Q (new_AGEMA_signal_14687) ) ;
    buf_clk new_AGEMA_reg_buffer_8839 ( .C (clk), .D (new_AGEMA_signal_14690), .Q (new_AGEMA_signal_14691) ) ;
    buf_clk new_AGEMA_reg_buffer_8843 ( .C (clk), .D (new_AGEMA_signal_14694), .Q (new_AGEMA_signal_14695) ) ;
    buf_clk new_AGEMA_reg_buffer_8847 ( .C (clk), .D (new_AGEMA_signal_14698), .Q (new_AGEMA_signal_14699) ) ;
    buf_clk new_AGEMA_reg_buffer_8851 ( .C (clk), .D (new_AGEMA_signal_14702), .Q (new_AGEMA_signal_14703) ) ;
    buf_clk new_AGEMA_reg_buffer_8855 ( .C (clk), .D (new_AGEMA_signal_14706), .Q (new_AGEMA_signal_14707) ) ;
    buf_clk new_AGEMA_reg_buffer_8859 ( .C (clk), .D (new_AGEMA_signal_14710), .Q (new_AGEMA_signal_14711) ) ;
    buf_clk new_AGEMA_reg_buffer_8863 ( .C (clk), .D (new_AGEMA_signal_14714), .Q (new_AGEMA_signal_14715) ) ;
    buf_clk new_AGEMA_reg_buffer_8867 ( .C (clk), .D (new_AGEMA_signal_14718), .Q (new_AGEMA_signal_14719) ) ;
    buf_clk new_AGEMA_reg_buffer_8871 ( .C (clk), .D (new_AGEMA_signal_14722), .Q (new_AGEMA_signal_14723) ) ;
    buf_clk new_AGEMA_reg_buffer_8875 ( .C (clk), .D (new_AGEMA_signal_14726), .Q (new_AGEMA_signal_14727) ) ;
    buf_clk new_AGEMA_reg_buffer_8879 ( .C (clk), .D (new_AGEMA_signal_14730), .Q (new_AGEMA_signal_14731) ) ;
    buf_clk new_AGEMA_reg_buffer_8883 ( .C (clk), .D (new_AGEMA_signal_14734), .Q (new_AGEMA_signal_14735) ) ;
    buf_clk new_AGEMA_reg_buffer_8887 ( .C (clk), .D (new_AGEMA_signal_14738), .Q (new_AGEMA_signal_14739) ) ;
    buf_clk new_AGEMA_reg_buffer_8891 ( .C (clk), .D (new_AGEMA_signal_14742), .Q (new_AGEMA_signal_14743) ) ;
    buf_clk new_AGEMA_reg_buffer_8895 ( .C (clk), .D (new_AGEMA_signal_14746), .Q (new_AGEMA_signal_14747) ) ;
    buf_clk new_AGEMA_reg_buffer_8899 ( .C (clk), .D (new_AGEMA_signal_14750), .Q (new_AGEMA_signal_14751) ) ;
    buf_clk new_AGEMA_reg_buffer_8903 ( .C (clk), .D (new_AGEMA_signal_14754), .Q (new_AGEMA_signal_14755) ) ;
    buf_clk new_AGEMA_reg_buffer_8907 ( .C (clk), .D (new_AGEMA_signal_14758), .Q (new_AGEMA_signal_14759) ) ;
    buf_clk new_AGEMA_reg_buffer_8911 ( .C (clk), .D (new_AGEMA_signal_14762), .Q (new_AGEMA_signal_14763) ) ;
    buf_clk new_AGEMA_reg_buffer_8915 ( .C (clk), .D (new_AGEMA_signal_14766), .Q (new_AGEMA_signal_14767) ) ;
    buf_clk new_AGEMA_reg_buffer_8919 ( .C (clk), .D (new_AGEMA_signal_14770), .Q (new_AGEMA_signal_14771) ) ;
    buf_clk new_AGEMA_reg_buffer_8923 ( .C (clk), .D (new_AGEMA_signal_14774), .Q (new_AGEMA_signal_14775) ) ;
    buf_clk new_AGEMA_reg_buffer_8927 ( .C (clk), .D (new_AGEMA_signal_14778), .Q (new_AGEMA_signal_14779) ) ;
    buf_clk new_AGEMA_reg_buffer_8931 ( .C (clk), .D (new_AGEMA_signal_14782), .Q (new_AGEMA_signal_14783) ) ;
    buf_clk new_AGEMA_reg_buffer_8935 ( .C (clk), .D (new_AGEMA_signal_14786), .Q (new_AGEMA_signal_14787) ) ;
    buf_clk new_AGEMA_reg_buffer_8939 ( .C (clk), .D (new_AGEMA_signal_14790), .Q (new_AGEMA_signal_14791) ) ;
    buf_clk new_AGEMA_reg_buffer_8943 ( .C (clk), .D (new_AGEMA_signal_14794), .Q (new_AGEMA_signal_14795) ) ;
    buf_clk new_AGEMA_reg_buffer_8947 ( .C (clk), .D (new_AGEMA_signal_14798), .Q (new_AGEMA_signal_14799) ) ;
    buf_clk new_AGEMA_reg_buffer_8951 ( .C (clk), .D (new_AGEMA_signal_14802), .Q (new_AGEMA_signal_14803) ) ;
    buf_clk new_AGEMA_reg_buffer_8955 ( .C (clk), .D (new_AGEMA_signal_14806), .Q (new_AGEMA_signal_14807) ) ;
    buf_clk new_AGEMA_reg_buffer_8959 ( .C (clk), .D (new_AGEMA_signal_14810), .Q (new_AGEMA_signal_14811) ) ;
    buf_clk new_AGEMA_reg_buffer_8963 ( .C (clk), .D (new_AGEMA_signal_14814), .Q (new_AGEMA_signal_14815) ) ;
    buf_clk new_AGEMA_reg_buffer_8967 ( .C (clk), .D (new_AGEMA_signal_14818), .Q (new_AGEMA_signal_14819) ) ;
    buf_clk new_AGEMA_reg_buffer_8971 ( .C (clk), .D (new_AGEMA_signal_14822), .Q (new_AGEMA_signal_14823) ) ;
    buf_clk new_AGEMA_reg_buffer_8975 ( .C (clk), .D (new_AGEMA_signal_14826), .Q (new_AGEMA_signal_14827) ) ;
    buf_clk new_AGEMA_reg_buffer_8979 ( .C (clk), .D (new_AGEMA_signal_14830), .Q (new_AGEMA_signal_14831) ) ;
    buf_clk new_AGEMA_reg_buffer_8983 ( .C (clk), .D (new_AGEMA_signal_14834), .Q (new_AGEMA_signal_14835) ) ;
    buf_clk new_AGEMA_reg_buffer_8987 ( .C (clk), .D (new_AGEMA_signal_14838), .Q (new_AGEMA_signal_14839) ) ;
    buf_clk new_AGEMA_reg_buffer_8991 ( .C (clk), .D (new_AGEMA_signal_14842), .Q (new_AGEMA_signal_14843) ) ;
    buf_clk new_AGEMA_reg_buffer_8995 ( .C (clk), .D (new_AGEMA_signal_14846), .Q (new_AGEMA_signal_14847) ) ;
    buf_clk new_AGEMA_reg_buffer_8999 ( .C (clk), .D (new_AGEMA_signal_14850), .Q (new_AGEMA_signal_14851) ) ;
    buf_clk new_AGEMA_reg_buffer_9003 ( .C (clk), .D (new_AGEMA_signal_14854), .Q (new_AGEMA_signal_14855) ) ;
    buf_clk new_AGEMA_reg_buffer_9007 ( .C (clk), .D (new_AGEMA_signal_14858), .Q (new_AGEMA_signal_14859) ) ;
    buf_clk new_AGEMA_reg_buffer_9011 ( .C (clk), .D (new_AGEMA_signal_14862), .Q (new_AGEMA_signal_14863) ) ;
    buf_clk new_AGEMA_reg_buffer_9015 ( .C (clk), .D (new_AGEMA_signal_14866), .Q (new_AGEMA_signal_14867) ) ;
    buf_clk new_AGEMA_reg_buffer_9019 ( .C (clk), .D (new_AGEMA_signal_14870), .Q (new_AGEMA_signal_14871) ) ;
    buf_clk new_AGEMA_reg_buffer_9023 ( .C (clk), .D (new_AGEMA_signal_14874), .Q (new_AGEMA_signal_14875) ) ;
    buf_clk new_AGEMA_reg_buffer_9027 ( .C (clk), .D (new_AGEMA_signal_14878), .Q (new_AGEMA_signal_14879) ) ;
    buf_clk new_AGEMA_reg_buffer_9031 ( .C (clk), .D (new_AGEMA_signal_14882), .Q (new_AGEMA_signal_14883) ) ;
    buf_clk new_AGEMA_reg_buffer_9035 ( .C (clk), .D (new_AGEMA_signal_14886), .Q (new_AGEMA_signal_14887) ) ;
    buf_clk new_AGEMA_reg_buffer_9039 ( .C (clk), .D (new_AGEMA_signal_14890), .Q (new_AGEMA_signal_14891) ) ;
    buf_clk new_AGEMA_reg_buffer_9043 ( .C (clk), .D (new_AGEMA_signal_14894), .Q (new_AGEMA_signal_14895) ) ;
    buf_clk new_AGEMA_reg_buffer_9047 ( .C (clk), .D (new_AGEMA_signal_14898), .Q (new_AGEMA_signal_14899) ) ;
    buf_clk new_AGEMA_reg_buffer_9051 ( .C (clk), .D (new_AGEMA_signal_14902), .Q (new_AGEMA_signal_14903) ) ;
    buf_clk new_AGEMA_reg_buffer_9055 ( .C (clk), .D (new_AGEMA_signal_14906), .Q (new_AGEMA_signal_14907) ) ;
    buf_clk new_AGEMA_reg_buffer_9059 ( .C (clk), .D (new_AGEMA_signal_14910), .Q (new_AGEMA_signal_14911) ) ;
    buf_clk new_AGEMA_reg_buffer_9063 ( .C (clk), .D (new_AGEMA_signal_14914), .Q (new_AGEMA_signal_14915) ) ;
    buf_clk new_AGEMA_reg_buffer_9067 ( .C (clk), .D (new_AGEMA_signal_14918), .Q (new_AGEMA_signal_14919) ) ;
    buf_clk new_AGEMA_reg_buffer_9071 ( .C (clk), .D (new_AGEMA_signal_14922), .Q (new_AGEMA_signal_14923) ) ;
    buf_clk new_AGEMA_reg_buffer_9075 ( .C (clk), .D (new_AGEMA_signal_14926), .Q (new_AGEMA_signal_14927) ) ;
    buf_clk new_AGEMA_reg_buffer_9079 ( .C (clk), .D (new_AGEMA_signal_14930), .Q (new_AGEMA_signal_14931) ) ;
    buf_clk new_AGEMA_reg_buffer_9083 ( .C (clk), .D (new_AGEMA_signal_14934), .Q (new_AGEMA_signal_14935) ) ;
    buf_clk new_AGEMA_reg_buffer_9087 ( .C (clk), .D (new_AGEMA_signal_14938), .Q (new_AGEMA_signal_14939) ) ;
    buf_clk new_AGEMA_reg_buffer_9091 ( .C (clk), .D (new_AGEMA_signal_14942), .Q (new_AGEMA_signal_14943) ) ;
    buf_clk new_AGEMA_reg_buffer_9095 ( .C (clk), .D (new_AGEMA_signal_14946), .Q (new_AGEMA_signal_14947) ) ;
    buf_clk new_AGEMA_reg_buffer_9099 ( .C (clk), .D (new_AGEMA_signal_14950), .Q (new_AGEMA_signal_14951) ) ;
    buf_clk new_AGEMA_reg_buffer_9103 ( .C (clk), .D (new_AGEMA_signal_14954), .Q (new_AGEMA_signal_14955) ) ;
    buf_clk new_AGEMA_reg_buffer_9107 ( .C (clk), .D (new_AGEMA_signal_14958), .Q (new_AGEMA_signal_14959) ) ;
    buf_clk new_AGEMA_reg_buffer_9111 ( .C (clk), .D (new_AGEMA_signal_14962), .Q (new_AGEMA_signal_14963) ) ;
    buf_clk new_AGEMA_reg_buffer_9115 ( .C (clk), .D (new_AGEMA_signal_14966), .Q (new_AGEMA_signal_14967) ) ;
    buf_clk new_AGEMA_reg_buffer_9119 ( .C (clk), .D (new_AGEMA_signal_14970), .Q (new_AGEMA_signal_14971) ) ;
    buf_clk new_AGEMA_reg_buffer_9123 ( .C (clk), .D (new_AGEMA_signal_14974), .Q (new_AGEMA_signal_14975) ) ;
    buf_clk new_AGEMA_reg_buffer_9127 ( .C (clk), .D (new_AGEMA_signal_14978), .Q (new_AGEMA_signal_14979) ) ;
    buf_clk new_AGEMA_reg_buffer_9131 ( .C (clk), .D (new_AGEMA_signal_14982), .Q (new_AGEMA_signal_14983) ) ;
    buf_clk new_AGEMA_reg_buffer_9135 ( .C (clk), .D (new_AGEMA_signal_14986), .Q (new_AGEMA_signal_14987) ) ;
    buf_clk new_AGEMA_reg_buffer_9139 ( .C (clk), .D (new_AGEMA_signal_14990), .Q (new_AGEMA_signal_14991) ) ;
    buf_clk new_AGEMA_reg_buffer_9143 ( .C (clk), .D (new_AGEMA_signal_14994), .Q (new_AGEMA_signal_14995) ) ;
    buf_clk new_AGEMA_reg_buffer_9147 ( .C (clk), .D (new_AGEMA_signal_14998), .Q (new_AGEMA_signal_14999) ) ;
    buf_clk new_AGEMA_reg_buffer_9151 ( .C (clk), .D (new_AGEMA_signal_15002), .Q (new_AGEMA_signal_15003) ) ;
    buf_clk new_AGEMA_reg_buffer_9155 ( .C (clk), .D (new_AGEMA_signal_15006), .Q (new_AGEMA_signal_15007) ) ;
    buf_clk new_AGEMA_reg_buffer_9159 ( .C (clk), .D (new_AGEMA_signal_15010), .Q (new_AGEMA_signal_15011) ) ;
    buf_clk new_AGEMA_reg_buffer_9163 ( .C (clk), .D (new_AGEMA_signal_15014), .Q (new_AGEMA_signal_15015) ) ;
    buf_clk new_AGEMA_reg_buffer_9167 ( .C (clk), .D (new_AGEMA_signal_15018), .Q (new_AGEMA_signal_15019) ) ;
    buf_clk new_AGEMA_reg_buffer_9171 ( .C (clk), .D (new_AGEMA_signal_15022), .Q (new_AGEMA_signal_15023) ) ;
    buf_clk new_AGEMA_reg_buffer_9175 ( .C (clk), .D (new_AGEMA_signal_15026), .Q (new_AGEMA_signal_15027) ) ;
    buf_clk new_AGEMA_reg_buffer_9179 ( .C (clk), .D (new_AGEMA_signal_15030), .Q (new_AGEMA_signal_15031) ) ;
    buf_clk new_AGEMA_reg_buffer_9183 ( .C (clk), .D (new_AGEMA_signal_15034), .Q (new_AGEMA_signal_15035) ) ;
    buf_clk new_AGEMA_reg_buffer_9187 ( .C (clk), .D (new_AGEMA_signal_15038), .Q (new_AGEMA_signal_15039) ) ;
    buf_clk new_AGEMA_reg_buffer_9191 ( .C (clk), .D (new_AGEMA_signal_15042), .Q (new_AGEMA_signal_15043) ) ;
    buf_clk new_AGEMA_reg_buffer_9195 ( .C (clk), .D (new_AGEMA_signal_15046), .Q (new_AGEMA_signal_15047) ) ;
    buf_clk new_AGEMA_reg_buffer_9199 ( .C (clk), .D (new_AGEMA_signal_15050), .Q (new_AGEMA_signal_15051) ) ;
    buf_clk new_AGEMA_reg_buffer_9203 ( .C (clk), .D (new_AGEMA_signal_15054), .Q (new_AGEMA_signal_15055) ) ;
    buf_clk new_AGEMA_reg_buffer_9207 ( .C (clk), .D (new_AGEMA_signal_15058), .Q (new_AGEMA_signal_15059) ) ;
    buf_clk new_AGEMA_reg_buffer_9211 ( .C (clk), .D (new_AGEMA_signal_15062), .Q (new_AGEMA_signal_15063) ) ;
    buf_clk new_AGEMA_reg_buffer_9215 ( .C (clk), .D (new_AGEMA_signal_15066), .Q (new_AGEMA_signal_15067) ) ;
    buf_clk new_AGEMA_reg_buffer_9219 ( .C (clk), .D (new_AGEMA_signal_15070), .Q (new_AGEMA_signal_15071) ) ;
    buf_clk new_AGEMA_reg_buffer_9223 ( .C (clk), .D (new_AGEMA_signal_15074), .Q (new_AGEMA_signal_15075) ) ;
    buf_clk new_AGEMA_reg_buffer_9227 ( .C (clk), .D (new_AGEMA_signal_15078), .Q (new_AGEMA_signal_15079) ) ;
    buf_clk new_AGEMA_reg_buffer_9231 ( .C (clk), .D (new_AGEMA_signal_15082), .Q (new_AGEMA_signal_15083) ) ;
    buf_clk new_AGEMA_reg_buffer_9235 ( .C (clk), .D (new_AGEMA_signal_15086), .Q (new_AGEMA_signal_15087) ) ;
    buf_clk new_AGEMA_reg_buffer_9239 ( .C (clk), .D (new_AGEMA_signal_15090), .Q (new_AGEMA_signal_15091) ) ;
    buf_clk new_AGEMA_reg_buffer_9243 ( .C (clk), .D (new_AGEMA_signal_15094), .Q (new_AGEMA_signal_15095) ) ;
    buf_clk new_AGEMA_reg_buffer_9247 ( .C (clk), .D (new_AGEMA_signal_15098), .Q (new_AGEMA_signal_15099) ) ;
    buf_clk new_AGEMA_reg_buffer_9251 ( .C (clk), .D (new_AGEMA_signal_15102), .Q (new_AGEMA_signal_15103) ) ;
    buf_clk new_AGEMA_reg_buffer_9255 ( .C (clk), .D (new_AGEMA_signal_15106), .Q (new_AGEMA_signal_15107) ) ;
    buf_clk new_AGEMA_reg_buffer_9259 ( .C (clk), .D (new_AGEMA_signal_15110), .Q (new_AGEMA_signal_15111) ) ;
    buf_clk new_AGEMA_reg_buffer_9263 ( .C (clk), .D (new_AGEMA_signal_15114), .Q (new_AGEMA_signal_15115) ) ;
    buf_clk new_AGEMA_reg_buffer_9267 ( .C (clk), .D (new_AGEMA_signal_15118), .Q (new_AGEMA_signal_15119) ) ;
    buf_clk new_AGEMA_reg_buffer_9271 ( .C (clk), .D (new_AGEMA_signal_15122), .Q (new_AGEMA_signal_15123) ) ;
    buf_clk new_AGEMA_reg_buffer_9275 ( .C (clk), .D (new_AGEMA_signal_15126), .Q (new_AGEMA_signal_15127) ) ;
    buf_clk new_AGEMA_reg_buffer_9279 ( .C (clk), .D (new_AGEMA_signal_15130), .Q (new_AGEMA_signal_15131) ) ;
    buf_clk new_AGEMA_reg_buffer_9283 ( .C (clk), .D (new_AGEMA_signal_15134), .Q (new_AGEMA_signal_15135) ) ;
    buf_clk new_AGEMA_reg_buffer_9287 ( .C (clk), .D (new_AGEMA_signal_15138), .Q (new_AGEMA_signal_15139) ) ;
    buf_clk new_AGEMA_reg_buffer_9291 ( .C (clk), .D (new_AGEMA_signal_15142), .Q (new_AGEMA_signal_15143) ) ;
    buf_clk new_AGEMA_reg_buffer_9295 ( .C (clk), .D (new_AGEMA_signal_15146), .Q (new_AGEMA_signal_15147) ) ;
    buf_clk new_AGEMA_reg_buffer_9299 ( .C (clk), .D (new_AGEMA_signal_15150), .Q (new_AGEMA_signal_15151) ) ;
    buf_clk new_AGEMA_reg_buffer_9303 ( .C (clk), .D (new_AGEMA_signal_15154), .Q (new_AGEMA_signal_15155) ) ;
    buf_clk new_AGEMA_reg_buffer_9307 ( .C (clk), .D (new_AGEMA_signal_15158), .Q (new_AGEMA_signal_15159) ) ;
    buf_clk new_AGEMA_reg_buffer_9311 ( .C (clk), .D (new_AGEMA_signal_15162), .Q (new_AGEMA_signal_15163) ) ;
    buf_clk new_AGEMA_reg_buffer_9315 ( .C (clk), .D (new_AGEMA_signal_15166), .Q (new_AGEMA_signal_15167) ) ;
    buf_clk new_AGEMA_reg_buffer_9319 ( .C (clk), .D (new_AGEMA_signal_15170), .Q (new_AGEMA_signal_15171) ) ;
    buf_clk new_AGEMA_reg_buffer_9323 ( .C (clk), .D (new_AGEMA_signal_15174), .Q (new_AGEMA_signal_15175) ) ;
    buf_clk new_AGEMA_reg_buffer_9327 ( .C (clk), .D (new_AGEMA_signal_15178), .Q (new_AGEMA_signal_15179) ) ;
    buf_clk new_AGEMA_reg_buffer_9331 ( .C (clk), .D (new_AGEMA_signal_15182), .Q (new_AGEMA_signal_15183) ) ;
    buf_clk new_AGEMA_reg_buffer_9335 ( .C (clk), .D (new_AGEMA_signal_15186), .Q (new_AGEMA_signal_15187) ) ;
    buf_clk new_AGEMA_reg_buffer_9339 ( .C (clk), .D (new_AGEMA_signal_15190), .Q (new_AGEMA_signal_15191) ) ;
    buf_clk new_AGEMA_reg_buffer_9343 ( .C (clk), .D (new_AGEMA_signal_15194), .Q (new_AGEMA_signal_15195) ) ;
    buf_clk new_AGEMA_reg_buffer_9347 ( .C (clk), .D (new_AGEMA_signal_15198), .Q (new_AGEMA_signal_15199) ) ;
    buf_clk new_AGEMA_reg_buffer_9351 ( .C (clk), .D (new_AGEMA_signal_15202), .Q (new_AGEMA_signal_15203) ) ;
    buf_clk new_AGEMA_reg_buffer_9355 ( .C (clk), .D (new_AGEMA_signal_15206), .Q (new_AGEMA_signal_15207) ) ;
    buf_clk new_AGEMA_reg_buffer_9359 ( .C (clk), .D (new_AGEMA_signal_15210), .Q (new_AGEMA_signal_15211) ) ;
    buf_clk new_AGEMA_reg_buffer_9363 ( .C (clk), .D (new_AGEMA_signal_15214), .Q (new_AGEMA_signal_15215) ) ;
    buf_clk new_AGEMA_reg_buffer_9367 ( .C (clk), .D (new_AGEMA_signal_15218), .Q (new_AGEMA_signal_15219) ) ;
    buf_clk new_AGEMA_reg_buffer_9371 ( .C (clk), .D (new_AGEMA_signal_15222), .Q (new_AGEMA_signal_15223) ) ;
    buf_clk new_AGEMA_reg_buffer_9375 ( .C (clk), .D (new_AGEMA_signal_15226), .Q (new_AGEMA_signal_15227) ) ;
    buf_clk new_AGEMA_reg_buffer_9379 ( .C (clk), .D (new_AGEMA_signal_15230), .Q (new_AGEMA_signal_15231) ) ;
    buf_clk new_AGEMA_reg_buffer_9383 ( .C (clk), .D (new_AGEMA_signal_15234), .Q (new_AGEMA_signal_15235) ) ;
    buf_clk new_AGEMA_reg_buffer_9387 ( .C (clk), .D (new_AGEMA_signal_15238), .Q (new_AGEMA_signal_15239) ) ;
    buf_clk new_AGEMA_reg_buffer_9391 ( .C (clk), .D (new_AGEMA_signal_15242), .Q (new_AGEMA_signal_15243) ) ;
    buf_clk new_AGEMA_reg_buffer_9395 ( .C (clk), .D (new_AGEMA_signal_15246), .Q (new_AGEMA_signal_15247) ) ;
    buf_clk new_AGEMA_reg_buffer_9399 ( .C (clk), .D (new_AGEMA_signal_15250), .Q (new_AGEMA_signal_15251) ) ;
    buf_clk new_AGEMA_reg_buffer_9403 ( .C (clk), .D (new_AGEMA_signal_15254), .Q (new_AGEMA_signal_15255) ) ;
    buf_clk new_AGEMA_reg_buffer_9407 ( .C (clk), .D (new_AGEMA_signal_15258), .Q (new_AGEMA_signal_15259) ) ;
    buf_clk new_AGEMA_reg_buffer_9411 ( .C (clk), .D (new_AGEMA_signal_15262), .Q (new_AGEMA_signal_15263) ) ;
    buf_clk new_AGEMA_reg_buffer_9415 ( .C (clk), .D (new_AGEMA_signal_15266), .Q (new_AGEMA_signal_15267) ) ;
    buf_clk new_AGEMA_reg_buffer_9419 ( .C (clk), .D (new_AGEMA_signal_15270), .Q (new_AGEMA_signal_15271) ) ;
    buf_clk new_AGEMA_reg_buffer_9423 ( .C (clk), .D (new_AGEMA_signal_15274), .Q (new_AGEMA_signal_15275) ) ;
    buf_clk new_AGEMA_reg_buffer_9427 ( .C (clk), .D (new_AGEMA_signal_15278), .Q (new_AGEMA_signal_15279) ) ;
    buf_clk new_AGEMA_reg_buffer_9431 ( .C (clk), .D (new_AGEMA_signal_15282), .Q (new_AGEMA_signal_15283) ) ;
    buf_clk new_AGEMA_reg_buffer_9435 ( .C (clk), .D (new_AGEMA_signal_15286), .Q (new_AGEMA_signal_15287) ) ;
    buf_clk new_AGEMA_reg_buffer_9439 ( .C (clk), .D (new_AGEMA_signal_15290), .Q (new_AGEMA_signal_15291) ) ;
    buf_clk new_AGEMA_reg_buffer_9443 ( .C (clk), .D (new_AGEMA_signal_15294), .Q (new_AGEMA_signal_15295) ) ;
    buf_clk new_AGEMA_reg_buffer_9447 ( .C (clk), .D (new_AGEMA_signal_15298), .Q (new_AGEMA_signal_15299) ) ;
    buf_clk new_AGEMA_reg_buffer_9451 ( .C (clk), .D (new_AGEMA_signal_15302), .Q (new_AGEMA_signal_15303) ) ;
    buf_clk new_AGEMA_reg_buffer_9455 ( .C (clk), .D (new_AGEMA_signal_15306), .Q (new_AGEMA_signal_15307) ) ;
    buf_clk new_AGEMA_reg_buffer_9459 ( .C (clk), .D (new_AGEMA_signal_15310), .Q (new_AGEMA_signal_15311) ) ;
    buf_clk new_AGEMA_reg_buffer_9463 ( .C (clk), .D (new_AGEMA_signal_15314), .Q (new_AGEMA_signal_15315) ) ;
    buf_clk new_AGEMA_reg_buffer_9467 ( .C (clk), .D (new_AGEMA_signal_15318), .Q (new_AGEMA_signal_15319) ) ;
    buf_clk new_AGEMA_reg_buffer_9471 ( .C (clk), .D (new_AGEMA_signal_15322), .Q (new_AGEMA_signal_15323) ) ;
    buf_clk new_AGEMA_reg_buffer_9475 ( .C (clk), .D (new_AGEMA_signal_15326), .Q (new_AGEMA_signal_15327) ) ;
    buf_clk new_AGEMA_reg_buffer_9479 ( .C (clk), .D (new_AGEMA_signal_15330), .Q (new_AGEMA_signal_15331) ) ;
    buf_clk new_AGEMA_reg_buffer_9483 ( .C (clk), .D (new_AGEMA_signal_15334), .Q (new_AGEMA_signal_15335) ) ;
    buf_clk new_AGEMA_reg_buffer_9487 ( .C (clk), .D (new_AGEMA_signal_15338), .Q (new_AGEMA_signal_15339) ) ;
    buf_clk new_AGEMA_reg_buffer_9491 ( .C (clk), .D (new_AGEMA_signal_15342), .Q (new_AGEMA_signal_15343) ) ;
    buf_clk new_AGEMA_reg_buffer_9495 ( .C (clk), .D (new_AGEMA_signal_15346), .Q (new_AGEMA_signal_15347) ) ;
    buf_clk new_AGEMA_reg_buffer_9499 ( .C (clk), .D (new_AGEMA_signal_15350), .Q (new_AGEMA_signal_15351) ) ;
    buf_clk new_AGEMA_reg_buffer_9503 ( .C (clk), .D (new_AGEMA_signal_15354), .Q (new_AGEMA_signal_15355) ) ;
    buf_clk new_AGEMA_reg_buffer_9507 ( .C (clk), .D (new_AGEMA_signal_15358), .Q (new_AGEMA_signal_15359) ) ;
    buf_clk new_AGEMA_reg_buffer_9511 ( .C (clk), .D (new_AGEMA_signal_15362), .Q (new_AGEMA_signal_15363) ) ;
    buf_clk new_AGEMA_reg_buffer_9515 ( .C (clk), .D (new_AGEMA_signal_15366), .Q (new_AGEMA_signal_15367) ) ;
    buf_clk new_AGEMA_reg_buffer_9519 ( .C (clk), .D (new_AGEMA_signal_15370), .Q (new_AGEMA_signal_15371) ) ;
    buf_clk new_AGEMA_reg_buffer_9523 ( .C (clk), .D (new_AGEMA_signal_15374), .Q (new_AGEMA_signal_15375) ) ;
    buf_clk new_AGEMA_reg_buffer_9527 ( .C (clk), .D (new_AGEMA_signal_15378), .Q (new_AGEMA_signal_15379) ) ;
    buf_clk new_AGEMA_reg_buffer_9531 ( .C (clk), .D (new_AGEMA_signal_15382), .Q (new_AGEMA_signal_15383) ) ;
    buf_clk new_AGEMA_reg_buffer_9535 ( .C (clk), .D (new_AGEMA_signal_15386), .Q (new_AGEMA_signal_15387) ) ;
    buf_clk new_AGEMA_reg_buffer_9539 ( .C (clk), .D (new_AGEMA_signal_15390), .Q (new_AGEMA_signal_15391) ) ;
    buf_clk new_AGEMA_reg_buffer_9543 ( .C (clk), .D (new_AGEMA_signal_15394), .Q (new_AGEMA_signal_15395) ) ;
    buf_clk new_AGEMA_reg_buffer_9547 ( .C (clk), .D (new_AGEMA_signal_15398), .Q (new_AGEMA_signal_15399) ) ;
    buf_clk new_AGEMA_reg_buffer_9551 ( .C (clk), .D (new_AGEMA_signal_15402), .Q (new_AGEMA_signal_15403) ) ;
    buf_clk new_AGEMA_reg_buffer_9555 ( .C (clk), .D (new_AGEMA_signal_15406), .Q (new_AGEMA_signal_15407) ) ;
    buf_clk new_AGEMA_reg_buffer_9558 ( .C (clk), .D (new_AGEMA_signal_15409), .Q (new_AGEMA_signal_15410) ) ;
    buf_clk new_AGEMA_reg_buffer_9561 ( .C (clk), .D (new_AGEMA_signal_15412), .Q (new_AGEMA_signal_15413) ) ;
    buf_clk new_AGEMA_reg_buffer_9564 ( .C (clk), .D (new_AGEMA_signal_15415), .Q (new_AGEMA_signal_15416) ) ;
    buf_clk new_AGEMA_reg_buffer_9567 ( .C (clk), .D (new_AGEMA_signal_15418), .Q (new_AGEMA_signal_15419) ) ;
    buf_clk new_AGEMA_reg_buffer_9570 ( .C (clk), .D (new_AGEMA_signal_15421), .Q (new_AGEMA_signal_15422) ) ;
    buf_clk new_AGEMA_reg_buffer_9573 ( .C (clk), .D (new_AGEMA_signal_15424), .Q (new_AGEMA_signal_15425) ) ;
    buf_clk new_AGEMA_reg_buffer_9576 ( .C (clk), .D (new_AGEMA_signal_15427), .Q (new_AGEMA_signal_15428) ) ;
    buf_clk new_AGEMA_reg_buffer_9579 ( .C (clk), .D (new_AGEMA_signal_15430), .Q (new_AGEMA_signal_15431) ) ;
    buf_clk new_AGEMA_reg_buffer_9582 ( .C (clk), .D (new_AGEMA_signal_15433), .Q (new_AGEMA_signal_15434) ) ;
    buf_clk new_AGEMA_reg_buffer_9585 ( .C (clk), .D (new_AGEMA_signal_15436), .Q (new_AGEMA_signal_15437) ) ;
    buf_clk new_AGEMA_reg_buffer_9588 ( .C (clk), .D (new_AGEMA_signal_15439), .Q (new_AGEMA_signal_15440) ) ;
    buf_clk new_AGEMA_reg_buffer_9591 ( .C (clk), .D (new_AGEMA_signal_15442), .Q (new_AGEMA_signal_15443) ) ;
    buf_clk new_AGEMA_reg_buffer_9594 ( .C (clk), .D (new_AGEMA_signal_15445), .Q (new_AGEMA_signal_15446) ) ;
    buf_clk new_AGEMA_reg_buffer_9597 ( .C (clk), .D (new_AGEMA_signal_15448), .Q (new_AGEMA_signal_15449) ) ;
    buf_clk new_AGEMA_reg_buffer_9600 ( .C (clk), .D (new_AGEMA_signal_15451), .Q (new_AGEMA_signal_15452) ) ;
    buf_clk new_AGEMA_reg_buffer_9603 ( .C (clk), .D (new_AGEMA_signal_15454), .Q (new_AGEMA_signal_15455) ) ;
    buf_clk new_AGEMA_reg_buffer_9606 ( .C (clk), .D (new_AGEMA_signal_15457), .Q (new_AGEMA_signal_15458) ) ;
    buf_clk new_AGEMA_reg_buffer_9609 ( .C (clk), .D (new_AGEMA_signal_15460), .Q (new_AGEMA_signal_15461) ) ;
    buf_clk new_AGEMA_reg_buffer_9612 ( .C (clk), .D (new_AGEMA_signal_15463), .Q (new_AGEMA_signal_15464) ) ;
    buf_clk new_AGEMA_reg_buffer_9615 ( .C (clk), .D (new_AGEMA_signal_15466), .Q (new_AGEMA_signal_15467) ) ;
    buf_clk new_AGEMA_reg_buffer_9618 ( .C (clk), .D (new_AGEMA_signal_15469), .Q (new_AGEMA_signal_15470) ) ;
    buf_clk new_AGEMA_reg_buffer_9621 ( .C (clk), .D (new_AGEMA_signal_15472), .Q (new_AGEMA_signal_15473) ) ;
    buf_clk new_AGEMA_reg_buffer_9624 ( .C (clk), .D (new_AGEMA_signal_15475), .Q (new_AGEMA_signal_15476) ) ;
    buf_clk new_AGEMA_reg_buffer_9627 ( .C (clk), .D (new_AGEMA_signal_15478), .Q (new_AGEMA_signal_15479) ) ;
    buf_clk new_AGEMA_reg_buffer_9630 ( .C (clk), .D (new_AGEMA_signal_15481), .Q (new_AGEMA_signal_15482) ) ;
    buf_clk new_AGEMA_reg_buffer_9633 ( .C (clk), .D (new_AGEMA_signal_15484), .Q (new_AGEMA_signal_15485) ) ;
    buf_clk new_AGEMA_reg_buffer_9636 ( .C (clk), .D (new_AGEMA_signal_15487), .Q (new_AGEMA_signal_15488) ) ;
    buf_clk new_AGEMA_reg_buffer_9639 ( .C (clk), .D (new_AGEMA_signal_15490), .Q (new_AGEMA_signal_15491) ) ;
    buf_clk new_AGEMA_reg_buffer_9642 ( .C (clk), .D (new_AGEMA_signal_15493), .Q (new_AGEMA_signal_15494) ) ;
    buf_clk new_AGEMA_reg_buffer_9645 ( .C (clk), .D (new_AGEMA_signal_15496), .Q (new_AGEMA_signal_15497) ) ;
    buf_clk new_AGEMA_reg_buffer_9648 ( .C (clk), .D (new_AGEMA_signal_15499), .Q (new_AGEMA_signal_15500) ) ;
    buf_clk new_AGEMA_reg_buffer_9651 ( .C (clk), .D (new_AGEMA_signal_15502), .Q (new_AGEMA_signal_15503) ) ;
    buf_clk new_AGEMA_reg_buffer_9654 ( .C (clk), .D (new_AGEMA_signal_15505), .Q (new_AGEMA_signal_15506) ) ;
    buf_clk new_AGEMA_reg_buffer_9657 ( .C (clk), .D (new_AGEMA_signal_15508), .Q (new_AGEMA_signal_15509) ) ;
    buf_clk new_AGEMA_reg_buffer_9660 ( .C (clk), .D (new_AGEMA_signal_15511), .Q (new_AGEMA_signal_15512) ) ;
    buf_clk new_AGEMA_reg_buffer_9663 ( .C (clk), .D (new_AGEMA_signal_15514), .Q (new_AGEMA_signal_15515) ) ;
    buf_clk new_AGEMA_reg_buffer_9666 ( .C (clk), .D (new_AGEMA_signal_15517), .Q (new_AGEMA_signal_15518) ) ;
    buf_clk new_AGEMA_reg_buffer_9669 ( .C (clk), .D (new_AGEMA_signal_15520), .Q (new_AGEMA_signal_15521) ) ;
    buf_clk new_AGEMA_reg_buffer_9672 ( .C (clk), .D (new_AGEMA_signal_15523), .Q (new_AGEMA_signal_15524) ) ;
    buf_clk new_AGEMA_reg_buffer_9675 ( .C (clk), .D (new_AGEMA_signal_15526), .Q (new_AGEMA_signal_15527) ) ;
    buf_clk new_AGEMA_reg_buffer_9678 ( .C (clk), .D (new_AGEMA_signal_15529), .Q (new_AGEMA_signal_15530) ) ;
    buf_clk new_AGEMA_reg_buffer_9681 ( .C (clk), .D (new_AGEMA_signal_15532), .Q (new_AGEMA_signal_15533) ) ;
    buf_clk new_AGEMA_reg_buffer_9684 ( .C (clk), .D (new_AGEMA_signal_15535), .Q (new_AGEMA_signal_15536) ) ;
    buf_clk new_AGEMA_reg_buffer_9687 ( .C (clk), .D (new_AGEMA_signal_15538), .Q (new_AGEMA_signal_15539) ) ;
    buf_clk new_AGEMA_reg_buffer_9690 ( .C (clk), .D (new_AGEMA_signal_15541), .Q (new_AGEMA_signal_15542) ) ;
    buf_clk new_AGEMA_reg_buffer_9693 ( .C (clk), .D (new_AGEMA_signal_15544), .Q (new_AGEMA_signal_15545) ) ;
    buf_clk new_AGEMA_reg_buffer_9696 ( .C (clk), .D (new_AGEMA_signal_15547), .Q (new_AGEMA_signal_15548) ) ;
    buf_clk new_AGEMA_reg_buffer_9699 ( .C (clk), .D (new_AGEMA_signal_15550), .Q (new_AGEMA_signal_15551) ) ;
    buf_clk new_AGEMA_reg_buffer_9702 ( .C (clk), .D (new_AGEMA_signal_15553), .Q (new_AGEMA_signal_15554) ) ;
    buf_clk new_AGEMA_reg_buffer_9705 ( .C (clk), .D (new_AGEMA_signal_15556), .Q (new_AGEMA_signal_15557) ) ;
    buf_clk new_AGEMA_reg_buffer_9708 ( .C (clk), .D (new_AGEMA_signal_15559), .Q (new_AGEMA_signal_15560) ) ;
    buf_clk new_AGEMA_reg_buffer_9711 ( .C (clk), .D (new_AGEMA_signal_15562), .Q (new_AGEMA_signal_15563) ) ;
    buf_clk new_AGEMA_reg_buffer_9714 ( .C (clk), .D (new_AGEMA_signal_15565), .Q (new_AGEMA_signal_15566) ) ;
    buf_clk new_AGEMA_reg_buffer_9717 ( .C (clk), .D (new_AGEMA_signal_15568), .Q (new_AGEMA_signal_15569) ) ;
    buf_clk new_AGEMA_reg_buffer_9720 ( .C (clk), .D (new_AGEMA_signal_15571), .Q (new_AGEMA_signal_15572) ) ;
    buf_clk new_AGEMA_reg_buffer_9723 ( .C (clk), .D (new_AGEMA_signal_15574), .Q (new_AGEMA_signal_15575) ) ;
    buf_clk new_AGEMA_reg_buffer_9726 ( .C (clk), .D (new_AGEMA_signal_15577), .Q (new_AGEMA_signal_15578) ) ;
    buf_clk new_AGEMA_reg_buffer_9729 ( .C (clk), .D (new_AGEMA_signal_15580), .Q (new_AGEMA_signal_15581) ) ;
    buf_clk new_AGEMA_reg_buffer_9732 ( .C (clk), .D (new_AGEMA_signal_15583), .Q (new_AGEMA_signal_15584) ) ;
    buf_clk new_AGEMA_reg_buffer_9735 ( .C (clk), .D (new_AGEMA_signal_15586), .Q (new_AGEMA_signal_15587) ) ;
    buf_clk new_AGEMA_reg_buffer_9738 ( .C (clk), .D (new_AGEMA_signal_15589), .Q (new_AGEMA_signal_15590) ) ;
    buf_clk new_AGEMA_reg_buffer_9741 ( .C (clk), .D (new_AGEMA_signal_15592), .Q (new_AGEMA_signal_15593) ) ;
    buf_clk new_AGEMA_reg_buffer_9744 ( .C (clk), .D (new_AGEMA_signal_15595), .Q (new_AGEMA_signal_15596) ) ;
    buf_clk new_AGEMA_reg_buffer_9747 ( .C (clk), .D (new_AGEMA_signal_15598), .Q (new_AGEMA_signal_15599) ) ;
    buf_clk new_AGEMA_reg_buffer_9750 ( .C (clk), .D (new_AGEMA_signal_15601), .Q (new_AGEMA_signal_15602) ) ;
    buf_clk new_AGEMA_reg_buffer_9753 ( .C (clk), .D (new_AGEMA_signal_15604), .Q (new_AGEMA_signal_15605) ) ;
    buf_clk new_AGEMA_reg_buffer_9756 ( .C (clk), .D (new_AGEMA_signal_15607), .Q (new_AGEMA_signal_15608) ) ;
    buf_clk new_AGEMA_reg_buffer_9759 ( .C (clk), .D (new_AGEMA_signal_15610), .Q (new_AGEMA_signal_15611) ) ;
    buf_clk new_AGEMA_reg_buffer_9762 ( .C (clk), .D (new_AGEMA_signal_15613), .Q (new_AGEMA_signal_15614) ) ;
    buf_clk new_AGEMA_reg_buffer_9765 ( .C (clk), .D (new_AGEMA_signal_15616), .Q (new_AGEMA_signal_15617) ) ;
    buf_clk new_AGEMA_reg_buffer_9768 ( .C (clk), .D (new_AGEMA_signal_15619), .Q (new_AGEMA_signal_15620) ) ;
    buf_clk new_AGEMA_reg_buffer_9771 ( .C (clk), .D (new_AGEMA_signal_15622), .Q (new_AGEMA_signal_15623) ) ;
    buf_clk new_AGEMA_reg_buffer_9774 ( .C (clk), .D (new_AGEMA_signal_15625), .Q (new_AGEMA_signal_15626) ) ;
    buf_clk new_AGEMA_reg_buffer_9777 ( .C (clk), .D (new_AGEMA_signal_15628), .Q (new_AGEMA_signal_15629) ) ;
    buf_clk new_AGEMA_reg_buffer_9780 ( .C (clk), .D (new_AGEMA_signal_15631), .Q (new_AGEMA_signal_15632) ) ;
    buf_clk new_AGEMA_reg_buffer_9783 ( .C (clk), .D (new_AGEMA_signal_15634), .Q (new_AGEMA_signal_15635) ) ;
    buf_clk new_AGEMA_reg_buffer_9786 ( .C (clk), .D (new_AGEMA_signal_15637), .Q (new_AGEMA_signal_15638) ) ;
    buf_clk new_AGEMA_reg_buffer_9789 ( .C (clk), .D (new_AGEMA_signal_15640), .Q (new_AGEMA_signal_15641) ) ;
    buf_clk new_AGEMA_reg_buffer_9792 ( .C (clk), .D (new_AGEMA_signal_15643), .Q (new_AGEMA_signal_15644) ) ;
    buf_clk new_AGEMA_reg_buffer_9795 ( .C (clk), .D (new_AGEMA_signal_15646), .Q (new_AGEMA_signal_15647) ) ;
    buf_clk new_AGEMA_reg_buffer_9798 ( .C (clk), .D (new_AGEMA_signal_15649), .Q (new_AGEMA_signal_15650) ) ;
    buf_clk new_AGEMA_reg_buffer_9801 ( .C (clk), .D (new_AGEMA_signal_15652), .Q (new_AGEMA_signal_15653) ) ;
    buf_clk new_AGEMA_reg_buffer_9804 ( .C (clk), .D (new_AGEMA_signal_15655), .Q (new_AGEMA_signal_15656) ) ;
    buf_clk new_AGEMA_reg_buffer_9807 ( .C (clk), .D (new_AGEMA_signal_15658), .Q (new_AGEMA_signal_15659) ) ;
    buf_clk new_AGEMA_reg_buffer_9810 ( .C (clk), .D (new_AGEMA_signal_15661), .Q (new_AGEMA_signal_15662) ) ;
    buf_clk new_AGEMA_reg_buffer_9813 ( .C (clk), .D (new_AGEMA_signal_15664), .Q (new_AGEMA_signal_15665) ) ;
    buf_clk new_AGEMA_reg_buffer_9816 ( .C (clk), .D (new_AGEMA_signal_15667), .Q (new_AGEMA_signal_15668) ) ;
    buf_clk new_AGEMA_reg_buffer_9819 ( .C (clk), .D (new_AGEMA_signal_15670), .Q (new_AGEMA_signal_15671) ) ;
    buf_clk new_AGEMA_reg_buffer_9822 ( .C (clk), .D (new_AGEMA_signal_15673), .Q (new_AGEMA_signal_15674) ) ;
    buf_clk new_AGEMA_reg_buffer_9825 ( .C (clk), .D (new_AGEMA_signal_15676), .Q (new_AGEMA_signal_15677) ) ;
    buf_clk new_AGEMA_reg_buffer_9828 ( .C (clk), .D (new_AGEMA_signal_15679), .Q (new_AGEMA_signal_15680) ) ;
    buf_clk new_AGEMA_reg_buffer_9831 ( .C (clk), .D (new_AGEMA_signal_15682), .Q (new_AGEMA_signal_15683) ) ;
    buf_clk new_AGEMA_reg_buffer_9834 ( .C (clk), .D (new_AGEMA_signal_15685), .Q (new_AGEMA_signal_15686) ) ;
    buf_clk new_AGEMA_reg_buffer_9837 ( .C (clk), .D (new_AGEMA_signal_15688), .Q (new_AGEMA_signal_15689) ) ;
    buf_clk new_AGEMA_reg_buffer_9840 ( .C (clk), .D (new_AGEMA_signal_15691), .Q (new_AGEMA_signal_15692) ) ;
    buf_clk new_AGEMA_reg_buffer_9843 ( .C (clk), .D (new_AGEMA_signal_15694), .Q (new_AGEMA_signal_15695) ) ;
    buf_clk new_AGEMA_reg_buffer_9846 ( .C (clk), .D (new_AGEMA_signal_15697), .Q (new_AGEMA_signal_15698) ) ;
    buf_clk new_AGEMA_reg_buffer_9849 ( .C (clk), .D (new_AGEMA_signal_15700), .Q (new_AGEMA_signal_15701) ) ;
    buf_clk new_AGEMA_reg_buffer_9852 ( .C (clk), .D (new_AGEMA_signal_15703), .Q (new_AGEMA_signal_15704) ) ;
    buf_clk new_AGEMA_reg_buffer_9855 ( .C (clk), .D (new_AGEMA_signal_15706), .Q (new_AGEMA_signal_15707) ) ;
    buf_clk new_AGEMA_reg_buffer_9858 ( .C (clk), .D (new_AGEMA_signal_15709), .Q (new_AGEMA_signal_15710) ) ;
    buf_clk new_AGEMA_reg_buffer_9861 ( .C (clk), .D (new_AGEMA_signal_15712), .Q (new_AGEMA_signal_15713) ) ;
    buf_clk new_AGEMA_reg_buffer_9864 ( .C (clk), .D (new_AGEMA_signal_15715), .Q (new_AGEMA_signal_15716) ) ;
    buf_clk new_AGEMA_reg_buffer_9867 ( .C (clk), .D (new_AGEMA_signal_15718), .Q (new_AGEMA_signal_15719) ) ;
    buf_clk new_AGEMA_reg_buffer_9870 ( .C (clk), .D (new_AGEMA_signal_15721), .Q (new_AGEMA_signal_15722) ) ;
    buf_clk new_AGEMA_reg_buffer_9873 ( .C (clk), .D (new_AGEMA_signal_15724), .Q (new_AGEMA_signal_15725) ) ;
    buf_clk new_AGEMA_reg_buffer_9876 ( .C (clk), .D (new_AGEMA_signal_15727), .Q (new_AGEMA_signal_15728) ) ;
    buf_clk new_AGEMA_reg_buffer_9879 ( .C (clk), .D (new_AGEMA_signal_15730), .Q (new_AGEMA_signal_15731) ) ;
    buf_clk new_AGEMA_reg_buffer_9882 ( .C (clk), .D (new_AGEMA_signal_15733), .Q (new_AGEMA_signal_15734) ) ;
    buf_clk new_AGEMA_reg_buffer_9885 ( .C (clk), .D (new_AGEMA_signal_15736), .Q (new_AGEMA_signal_15737) ) ;
    buf_clk new_AGEMA_reg_buffer_9888 ( .C (clk), .D (new_AGEMA_signal_15739), .Q (new_AGEMA_signal_15740) ) ;
    buf_clk new_AGEMA_reg_buffer_9891 ( .C (clk), .D (new_AGEMA_signal_15742), .Q (new_AGEMA_signal_15743) ) ;
    buf_clk new_AGEMA_reg_buffer_9894 ( .C (clk), .D (new_AGEMA_signal_15745), .Q (new_AGEMA_signal_15746) ) ;
    buf_clk new_AGEMA_reg_buffer_9897 ( .C (clk), .D (new_AGEMA_signal_15748), .Q (new_AGEMA_signal_15749) ) ;
    buf_clk new_AGEMA_reg_buffer_9900 ( .C (clk), .D (new_AGEMA_signal_15751), .Q (new_AGEMA_signal_15752) ) ;
    buf_clk new_AGEMA_reg_buffer_9903 ( .C (clk), .D (new_AGEMA_signal_15754), .Q (new_AGEMA_signal_15755) ) ;
    buf_clk new_AGEMA_reg_buffer_9906 ( .C (clk), .D (new_AGEMA_signal_15757), .Q (new_AGEMA_signal_15758) ) ;
    buf_clk new_AGEMA_reg_buffer_9909 ( .C (clk), .D (new_AGEMA_signal_15760), .Q (new_AGEMA_signal_15761) ) ;
    buf_clk new_AGEMA_reg_buffer_9912 ( .C (clk), .D (new_AGEMA_signal_15763), .Q (new_AGEMA_signal_15764) ) ;
    buf_clk new_AGEMA_reg_buffer_9915 ( .C (clk), .D (new_AGEMA_signal_15766), .Q (new_AGEMA_signal_15767) ) ;
    buf_clk new_AGEMA_reg_buffer_9918 ( .C (clk), .D (new_AGEMA_signal_15769), .Q (new_AGEMA_signal_15770) ) ;
    buf_clk new_AGEMA_reg_buffer_9921 ( .C (clk), .D (new_AGEMA_signal_15772), .Q (new_AGEMA_signal_15773) ) ;
    buf_clk new_AGEMA_reg_buffer_9924 ( .C (clk), .D (new_AGEMA_signal_15775), .Q (new_AGEMA_signal_15776) ) ;
    buf_clk new_AGEMA_reg_buffer_9927 ( .C (clk), .D (new_AGEMA_signal_15778), .Q (new_AGEMA_signal_15779) ) ;
    buf_clk new_AGEMA_reg_buffer_9930 ( .C (clk), .D (new_AGEMA_signal_15781), .Q (new_AGEMA_signal_15782) ) ;
    buf_clk new_AGEMA_reg_buffer_9933 ( .C (clk), .D (new_AGEMA_signal_15784), .Q (new_AGEMA_signal_15785) ) ;
    buf_clk new_AGEMA_reg_buffer_9936 ( .C (clk), .D (new_AGEMA_signal_15787), .Q (new_AGEMA_signal_15788) ) ;
    buf_clk new_AGEMA_reg_buffer_9939 ( .C (clk), .D (new_AGEMA_signal_15790), .Q (new_AGEMA_signal_15791) ) ;
    buf_clk new_AGEMA_reg_buffer_9942 ( .C (clk), .D (new_AGEMA_signal_15793), .Q (new_AGEMA_signal_15794) ) ;
    buf_clk new_AGEMA_reg_buffer_9945 ( .C (clk), .D (new_AGEMA_signal_15796), .Q (new_AGEMA_signal_15797) ) ;
    buf_clk new_AGEMA_reg_buffer_9948 ( .C (clk), .D (new_AGEMA_signal_15799), .Q (new_AGEMA_signal_15800) ) ;
    buf_clk new_AGEMA_reg_buffer_9951 ( .C (clk), .D (new_AGEMA_signal_15802), .Q (new_AGEMA_signal_15803) ) ;
    buf_clk new_AGEMA_reg_buffer_9954 ( .C (clk), .D (new_AGEMA_signal_15805), .Q (new_AGEMA_signal_15806) ) ;
    buf_clk new_AGEMA_reg_buffer_9957 ( .C (clk), .D (new_AGEMA_signal_15808), .Q (new_AGEMA_signal_15809) ) ;
    buf_clk new_AGEMA_reg_buffer_9960 ( .C (clk), .D (new_AGEMA_signal_15811), .Q (new_AGEMA_signal_15812) ) ;
    buf_clk new_AGEMA_reg_buffer_9963 ( .C (clk), .D (new_AGEMA_signal_15814), .Q (new_AGEMA_signal_15815) ) ;
    buf_clk new_AGEMA_reg_buffer_9967 ( .C (clk), .D (new_AGEMA_signal_15818), .Q (new_AGEMA_signal_15819) ) ;
    buf_clk new_AGEMA_reg_buffer_9971 ( .C (clk), .D (new_AGEMA_signal_15822), .Q (new_AGEMA_signal_15823) ) ;
    buf_clk new_AGEMA_reg_buffer_9975 ( .C (clk), .D (new_AGEMA_signal_15826), .Q (new_AGEMA_signal_15827) ) ;

    /* cells in depth 4 */
    mux2_masked #(.security_order(1), .pipeline(1)) U858 ( .s (new_AGEMA_signal_10544), .b ({new_AGEMA_signal_7231, MixColumnsInput[0]}), .a ({new_AGEMA_signal_8096, MixColumnsOutput[0]}), .c ({new_AGEMA_signal_8190, RoundOutput[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U859 ( .s (new_AGEMA_signal_10544), .b ({new_AGEMA_signal_7388, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]}), .a ({new_AGEMA_signal_8271, MixColumnsOutput[100]}), .c ({new_AGEMA_signal_8383, RoundOutput[100]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U860 ( .s (new_AGEMA_signal_10544), .b ({new_AGEMA_signal_7387, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]}), .a ({new_AGEMA_signal_7973, MixColumnsOutput[101]}), .c ({new_AGEMA_signal_8191, RoundOutput[101]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U861 ( .s (new_AGEMA_signal_10544), .b ({new_AGEMA_signal_7386, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]}), .a ({new_AGEMA_signal_7972, MixColumnsOutput[102]}), .c ({new_AGEMA_signal_8192, RoundOutput[102]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U862 ( .s (new_AGEMA_signal_10544), .b ({new_AGEMA_signal_7385, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .a ({new_AGEMA_signal_7971, MixColumnsOutput[103]}), .c ({new_AGEMA_signal_8193, RoundOutput[103]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U863 ( .s (new_AGEMA_signal_10544), .b ({new_AGEMA_signal_7242, MixColumnsInput[104]}), .a ({new_AGEMA_signal_7970, MixColumnsOutput[104]}), .c ({new_AGEMA_signal_8194, RoundOutput[104]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U864 ( .s (new_AGEMA_signal_10544), .b ({new_AGEMA_signal_7426, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]}), .a ({new_AGEMA_signal_8270, MixColumnsOutput[105]}), .c ({new_AGEMA_signal_8384, RoundOutput[105]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U865 ( .s (new_AGEMA_signal_10544), .b ({new_AGEMA_signal_7425, MixColumnsInput[106]}), .a ({new_AGEMA_signal_7999, MixColumnsOutput[106]}), .c ({new_AGEMA_signal_8195, RoundOutput[106]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U866 ( .s (new_AGEMA_signal_10548), .b ({new_AGEMA_signal_7424, MixColumnsInput[107]}), .a ({new_AGEMA_signal_8281, MixColumnsOutput[107]}), .c ({new_AGEMA_signal_8385, RoundOutput[107]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U867 ( .s (new_AGEMA_signal_10552), .b ({new_AGEMA_signal_7423, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]}), .a ({new_AGEMA_signal_8280, MixColumnsOutput[108]}), .c ({new_AGEMA_signal_8386, RoundOutput[108]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U868 ( .s (new_AGEMA_signal_10556), .b ({new_AGEMA_signal_7422, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]}), .a ({new_AGEMA_signal_7996, MixColumnsOutput[109]}), .c ({new_AGEMA_signal_8196, RoundOutput[109]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U869 ( .s (new_AGEMA_signal_10560), .b ({new_AGEMA_signal_7453, MixColumnsInput[10]}), .a ({new_AGEMA_signal_8095, MixColumnsOutput[10]}), .c ({new_AGEMA_signal_8197, RoundOutput[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U870 ( .s (new_AGEMA_signal_10564), .b ({new_AGEMA_signal_7421, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]}), .a ({new_AGEMA_signal_7995, MixColumnsOutput[110]}), .c ({new_AGEMA_signal_8198, RoundOutput[110]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U871 ( .s (new_AGEMA_signal_10568), .b ({new_AGEMA_signal_7420, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .a ({new_AGEMA_signal_7994, MixColumnsOutput[111]}), .c ({new_AGEMA_signal_8199, RoundOutput[111]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U872 ( .s (new_AGEMA_signal_10564), .b ({new_AGEMA_signal_7297, MixColumnsInput[112]}), .a ({new_AGEMA_signal_7993, MixColumnsOutput[112]}), .c ({new_AGEMA_signal_8200, RoundOutput[112]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U873 ( .s (new_AGEMA_signal_10560), .b ({new_AGEMA_signal_7461, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]}), .a ({new_AGEMA_signal_8279, MixColumnsOutput[113]}), .c ({new_AGEMA_signal_8387, RoundOutput[113]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U874 ( .s (new_AGEMA_signal_10560), .b ({new_AGEMA_signal_7460, MixColumnsInput[114]}), .a ({new_AGEMA_signal_7991, MixColumnsOutput[114]}), .c ({new_AGEMA_signal_8201, RoundOutput[114]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U875 ( .s (new_AGEMA_signal_10548), .b ({new_AGEMA_signal_7459, MixColumnsInput[115]}), .a ({new_AGEMA_signal_8278, MixColumnsOutput[115]}), .c ({new_AGEMA_signal_8388, RoundOutput[115]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U876 ( .s (new_AGEMA_signal_10552), .b ({new_AGEMA_signal_7458, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]}), .a ({new_AGEMA_signal_8276, MixColumnsOutput[116]}), .c ({new_AGEMA_signal_8389, RoundOutput[116]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U877 ( .s (new_AGEMA_signal_10556), .b ({new_AGEMA_signal_7457, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]}), .a ({new_AGEMA_signal_7987, MixColumnsOutput[117]}), .c ({new_AGEMA_signal_8202, RoundOutput[117]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U878 ( .s (new_AGEMA_signal_10564), .b ({new_AGEMA_signal_7456, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]}), .a ({new_AGEMA_signal_7986, MixColumnsOutput[118]}), .c ({new_AGEMA_signal_8203, RoundOutput[118]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U879 ( .s (new_AGEMA_signal_10568), .b ({new_AGEMA_signal_7455, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .a ({new_AGEMA_signal_7985, MixColumnsOutput[119]}), .c ({new_AGEMA_signal_8204, RoundOutput[119]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U880 ( .s (new_AGEMA_signal_10568), .b ({new_AGEMA_signal_7452, MixColumnsInput[11]}), .a ({new_AGEMA_signal_8317, MixColumnsOutput[11]}), .c ({new_AGEMA_signal_8390, RoundOutput[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U881 ( .s (new_AGEMA_signal_10564), .b ({new_AGEMA_signal_7352, MixColumnsInput[120]}), .a ({new_AGEMA_signal_7984, MixColumnsOutput[120]}), .c ({new_AGEMA_signal_8205, RoundOutput[120]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U882 ( .s (new_AGEMA_signal_10560), .b ({new_AGEMA_signal_7496, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]}), .a ({new_AGEMA_signal_8275, MixColumnsOutput[121]}), .c ({new_AGEMA_signal_8391, RoundOutput[121]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U883 ( .s (new_AGEMA_signal_10564), .b ({new_AGEMA_signal_7495, MixColumnsInput[122]}), .a ({new_AGEMA_signal_7982, MixColumnsOutput[122]}), .c ({new_AGEMA_signal_8206, RoundOutput[122]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U884 ( .s (new_AGEMA_signal_10568), .b ({new_AGEMA_signal_7494, MixColumnsInput[123]}), .a ({new_AGEMA_signal_8274, MixColumnsOutput[123]}), .c ({new_AGEMA_signal_8392, RoundOutput[123]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U885 ( .s (new_AGEMA_signal_10552), .b ({new_AGEMA_signal_7493, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]}), .a ({new_AGEMA_signal_8273, MixColumnsOutput[124]}), .c ({new_AGEMA_signal_8393, RoundOutput[124]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U886 ( .s (new_AGEMA_signal_10568), .b ({new_AGEMA_signal_7492, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]}), .a ({new_AGEMA_signal_7979, MixColumnsOutput[125]}), .c ({new_AGEMA_signal_8207, RoundOutput[125]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U887 ( .s (new_AGEMA_signal_10552), .b ({new_AGEMA_signal_7491, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]}), .a ({new_AGEMA_signal_7977, MixColumnsOutput[126]}), .c ({new_AGEMA_signal_8208, RoundOutput[126]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U888 ( .s (new_AGEMA_signal_10556), .b ({new_AGEMA_signal_7490, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .a ({new_AGEMA_signal_7976, MixColumnsOutput[127]}), .c ({new_AGEMA_signal_8209, RoundOutput[127]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U889 ( .s (new_AGEMA_signal_10548), .b ({new_AGEMA_signal_7451, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]}), .a ({new_AGEMA_signal_8316, MixColumnsOutput[12]}), .c ({new_AGEMA_signal_8394, RoundOutput[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U890 ( .s (new_AGEMA_signal_10556), .b ({new_AGEMA_signal_7450, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]}), .a ({new_AGEMA_signal_8092, MixColumnsOutput[13]}), .c ({new_AGEMA_signal_8210, RoundOutput[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U891 ( .s (new_AGEMA_signal_10552), .b ({new_AGEMA_signal_7449, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]}), .a ({new_AGEMA_signal_8091, MixColumnsOutput[14]}), .c ({new_AGEMA_signal_8211, RoundOutput[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U892 ( .s (new_AGEMA_signal_10556), .b ({new_AGEMA_signal_7448, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .a ({new_AGEMA_signal_8090, MixColumnsOutput[15]}), .c ({new_AGEMA_signal_8212, RoundOutput[15]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U893 ( .s (new_AGEMA_signal_10548), .b ({new_AGEMA_signal_7341, MixColumnsInput[16]}), .a ({new_AGEMA_signal_8089, MixColumnsOutput[16]}), .c ({new_AGEMA_signal_8213, RoundOutput[16]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U894 ( .s (new_AGEMA_signal_10560), .b ({new_AGEMA_signal_7489, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]}), .a ({new_AGEMA_signal_8315, MixColumnsOutput[17]}), .c ({new_AGEMA_signal_8395, RoundOutput[17]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U895 ( .s (new_AGEMA_signal_10564), .b ({new_AGEMA_signal_7488, MixColumnsInput[18]}), .a ({new_AGEMA_signal_8087, MixColumnsOutput[18]}), .c ({new_AGEMA_signal_8214, RoundOutput[18]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U896 ( .s (new_AGEMA_signal_10568), .b ({new_AGEMA_signal_7487, MixColumnsInput[19]}), .a ({new_AGEMA_signal_8314, MixColumnsOutput[19]}), .c ({new_AGEMA_signal_8396, RoundOutput[19]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U897 ( .s (new_AGEMA_signal_10560), .b ({new_AGEMA_signal_7419, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]}), .a ({new_AGEMA_signal_8313, MixColumnsOutput[1]}), .c ({new_AGEMA_signal_8397, RoundOutput[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U898 ( .s (new_AGEMA_signal_10564), .b ({new_AGEMA_signal_7486, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]}), .a ({new_AGEMA_signal_8312, MixColumnsOutput[20]}), .c ({new_AGEMA_signal_8398, RoundOutput[20]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U899 ( .s (new_AGEMA_signal_10552), .b ({new_AGEMA_signal_7485, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]}), .a ({new_AGEMA_signal_8083, MixColumnsOutput[21]}), .c ({new_AGEMA_signal_8215, RoundOutput[21]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U900 ( .s (new_AGEMA_signal_10556), .b ({new_AGEMA_signal_7484, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]}), .a ({new_AGEMA_signal_8082, MixColumnsOutput[22]}), .c ({new_AGEMA_signal_8216, RoundOutput[22]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U901 ( .s (new_AGEMA_signal_10548), .b ({new_AGEMA_signal_7483, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .a ({new_AGEMA_signal_8081, MixColumnsOutput[23]}), .c ({new_AGEMA_signal_8217, RoundOutput[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U902 ( .s (new_AGEMA_signal_10568), .b ({new_AGEMA_signal_7220, MixColumnsInput[24]}), .a ({new_AGEMA_signal_8080, MixColumnsOutput[24]}), .c ({new_AGEMA_signal_8218, RoundOutput[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U903 ( .s (new_AGEMA_signal_10560), .b ({new_AGEMA_signal_7412, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]}), .a ({new_AGEMA_signal_8311, MixColumnsOutput[25]}), .c ({new_AGEMA_signal_8399, RoundOutput[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U904 ( .s (new_AGEMA_signal_10552), .b ({new_AGEMA_signal_7411, MixColumnsInput[26]}), .a ({new_AGEMA_signal_8078, MixColumnsOutput[26]}), .c ({new_AGEMA_signal_8219, RoundOutput[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U905 ( .s (new_AGEMA_signal_10556), .b ({new_AGEMA_signal_7410, MixColumnsInput[27]}), .a ({new_AGEMA_signal_8310, MixColumnsOutput[27]}), .c ({new_AGEMA_signal_8400, RoundOutput[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U906 ( .s (new_AGEMA_signal_10548), .b ({new_AGEMA_signal_7409, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]}), .a ({new_AGEMA_signal_8309, MixColumnsOutput[28]}), .c ({new_AGEMA_signal_8401, RoundOutput[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U907 ( .s (new_AGEMA_signal_10564), .b ({new_AGEMA_signal_7408, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]}), .a ({new_AGEMA_signal_8075, MixColumnsOutput[29]}), .c ({new_AGEMA_signal_8220, RoundOutput[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U908 ( .s (new_AGEMA_signal_10548), .b ({new_AGEMA_signal_7418, MixColumnsInput[2]}), .a ({new_AGEMA_signal_8074, MixColumnsOutput[2]}), .c ({new_AGEMA_signal_8221, RoundOutput[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U909 ( .s (new_AGEMA_signal_10568), .b ({new_AGEMA_signal_7407, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]}), .a ({new_AGEMA_signal_8073, MixColumnsOutput[30]}), .c ({new_AGEMA_signal_8222, RoundOutput[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U910 ( .s (new_AGEMA_signal_10560), .b ({new_AGEMA_signal_7406, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .a ({new_AGEMA_signal_8072, MixColumnsOutput[31]}), .c ({new_AGEMA_signal_8223, RoundOutput[31]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U911 ( .s (new_AGEMA_signal_10552), .b ({new_AGEMA_signal_7275, MixColumnsInput[32]}), .a ({new_AGEMA_signal_8064, MixColumnsOutput[32]}), .c ({new_AGEMA_signal_8224, RoundOutput[32]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U912 ( .s (new_AGEMA_signal_10556), .b ({new_AGEMA_signal_7447, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]}), .a ({new_AGEMA_signal_8301, MixColumnsOutput[33]}), .c ({new_AGEMA_signal_8402, RoundOutput[33]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U913 ( .s (new_AGEMA_signal_10548), .b ({new_AGEMA_signal_7446, MixColumnsInput[34]}), .a ({new_AGEMA_signal_8042, MixColumnsOutput[34]}), .c ({new_AGEMA_signal_8225, RoundOutput[34]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U914 ( .s (new_AGEMA_signal_10568), .b ({new_AGEMA_signal_7445, MixColumnsInput[35]}), .a ({new_AGEMA_signal_8296, MixColumnsOutput[35]}), .c ({new_AGEMA_signal_8403, RoundOutput[35]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U915 ( .s (new_AGEMA_signal_10568), .b ({new_AGEMA_signal_7444, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]}), .a ({new_AGEMA_signal_8295, MixColumnsOutput[36]}), .c ({new_AGEMA_signal_8404, RoundOutput[36]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U916 ( .s (new_AGEMA_signal_10568), .b ({new_AGEMA_signal_7443, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]}), .a ({new_AGEMA_signal_8037, MixColumnsOutput[37]}), .c ({new_AGEMA_signal_8226, RoundOutput[37]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U917 ( .s (new_AGEMA_signal_10568), .b ({new_AGEMA_signal_7442, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]}), .a ({new_AGEMA_signal_8036, MixColumnsOutput[38]}), .c ({new_AGEMA_signal_8227, RoundOutput[38]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U918 ( .s (new_AGEMA_signal_10568), .b ({new_AGEMA_signal_7441, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .a ({new_AGEMA_signal_8035, MixColumnsOutput[39]}), .c ({new_AGEMA_signal_8228, RoundOutput[39]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U919 ( .s (new_AGEMA_signal_10568), .b ({new_AGEMA_signal_7417, MixColumnsInput[3]}), .a ({new_AGEMA_signal_8308, MixColumnsOutput[3]}), .c ({new_AGEMA_signal_8405, RoundOutput[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U920 ( .s (new_AGEMA_signal_10568), .b ({new_AGEMA_signal_7330, MixColumnsInput[40]}), .a ({new_AGEMA_signal_8034, MixColumnsOutput[40]}), .c ({new_AGEMA_signal_8229, RoundOutput[40]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U921 ( .s (new_AGEMA_signal_10568), .b ({new_AGEMA_signal_7482, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]}), .a ({new_AGEMA_signal_8294, MixColumnsOutput[41]}), .c ({new_AGEMA_signal_8406, RoundOutput[41]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U922 ( .s (new_AGEMA_signal_10568), .b ({new_AGEMA_signal_7481, MixColumnsInput[42]}), .a ({new_AGEMA_signal_8063, MixColumnsOutput[42]}), .c ({new_AGEMA_signal_8230, RoundOutput[42]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U923 ( .s (new_AGEMA_signal_10568), .b ({new_AGEMA_signal_7480, MixColumnsInput[43]}), .a ({new_AGEMA_signal_8305, MixColumnsOutput[43]}), .c ({new_AGEMA_signal_8407, RoundOutput[43]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U924 ( .s (new_AGEMA_signal_10568), .b ({new_AGEMA_signal_7479, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]}), .a ({new_AGEMA_signal_8304, MixColumnsOutput[44]}), .c ({new_AGEMA_signal_8408, RoundOutput[44]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U925 ( .s (new_AGEMA_signal_10568), .b ({new_AGEMA_signal_7478, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]}), .a ({new_AGEMA_signal_8060, MixColumnsOutput[45]}), .c ({new_AGEMA_signal_8231, RoundOutput[45]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U926 ( .s (new_AGEMA_signal_10564), .b ({new_AGEMA_signal_7477, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]}), .a ({new_AGEMA_signal_8059, MixColumnsOutput[46]}), .c ({new_AGEMA_signal_8232, RoundOutput[46]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U927 ( .s (new_AGEMA_signal_10564), .b ({new_AGEMA_signal_7476, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .a ({new_AGEMA_signal_8058, MixColumnsOutput[47]}), .c ({new_AGEMA_signal_8233, RoundOutput[47]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U928 ( .s (new_AGEMA_signal_10564), .b ({new_AGEMA_signal_7209, MixColumnsInput[48]}), .a ({new_AGEMA_signal_8057, MixColumnsOutput[48]}), .c ({new_AGEMA_signal_8234, RoundOutput[48]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U929 ( .s (new_AGEMA_signal_10564), .b ({new_AGEMA_signal_7405, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]}), .a ({new_AGEMA_signal_8303, MixColumnsOutput[49]}), .c ({new_AGEMA_signal_8409, RoundOutput[49]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U930 ( .s (new_AGEMA_signal_10564), .b ({new_AGEMA_signal_7416, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]}), .a ({new_AGEMA_signal_8307, MixColumnsOutput[4]}), .c ({new_AGEMA_signal_8410, RoundOutput[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U931 ( .s (new_AGEMA_signal_10564), .b ({new_AGEMA_signal_7404, MixColumnsInput[50]}), .a ({new_AGEMA_signal_8055, MixColumnsOutput[50]}), .c ({new_AGEMA_signal_8235, RoundOutput[50]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U932 ( .s (new_AGEMA_signal_10564), .b ({new_AGEMA_signal_7403, MixColumnsInput[51]}), .a ({new_AGEMA_signal_8302, MixColumnsOutput[51]}), .c ({new_AGEMA_signal_8411, RoundOutput[51]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U933 ( .s (new_AGEMA_signal_10564), .b ({new_AGEMA_signal_7402, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]}), .a ({new_AGEMA_signal_8300, MixColumnsOutput[52]}), .c ({new_AGEMA_signal_8412, RoundOutput[52]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U934 ( .s (new_AGEMA_signal_10564), .b ({new_AGEMA_signal_7401, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]}), .a ({new_AGEMA_signal_8051, MixColumnsOutput[53]}), .c ({new_AGEMA_signal_8236, RoundOutput[53]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U935 ( .s (new_AGEMA_signal_10564), .b ({new_AGEMA_signal_7400, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]}), .a ({new_AGEMA_signal_8050, MixColumnsOutput[54]}), .c ({new_AGEMA_signal_8237, RoundOutput[54]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U936 ( .s (new_AGEMA_signal_10564), .b ({new_AGEMA_signal_7399, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .a ({new_AGEMA_signal_8049, MixColumnsOutput[55]}), .c ({new_AGEMA_signal_8238, RoundOutput[55]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U937 ( .s (new_AGEMA_signal_10564), .b ({new_AGEMA_signal_7264, MixColumnsInput[56]}), .a ({new_AGEMA_signal_8048, MixColumnsOutput[56]}), .c ({new_AGEMA_signal_8239, RoundOutput[56]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U938 ( .s (new_AGEMA_signal_10560), .b ({new_AGEMA_signal_7440, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]}), .a ({new_AGEMA_signal_8299, MixColumnsOutput[57]}), .c ({new_AGEMA_signal_8413, RoundOutput[57]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U939 ( .s (new_AGEMA_signal_10560), .b ({new_AGEMA_signal_7439, MixColumnsInput[58]}), .a ({new_AGEMA_signal_8046, MixColumnsOutput[58]}), .c ({new_AGEMA_signal_8240, RoundOutput[58]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U940 ( .s (new_AGEMA_signal_10560), .b ({new_AGEMA_signal_7438, MixColumnsInput[59]}), .a ({new_AGEMA_signal_8298, MixColumnsOutput[59]}), .c ({new_AGEMA_signal_8414, RoundOutput[59]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U941 ( .s (new_AGEMA_signal_10560), .b ({new_AGEMA_signal_7415, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]}), .a ({new_AGEMA_signal_8069, MixColumnsOutput[5]}), .c ({new_AGEMA_signal_8241, RoundOutput[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U942 ( .s (new_AGEMA_signal_10560), .b ({new_AGEMA_signal_7437, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]}), .a ({new_AGEMA_signal_8297, MixColumnsOutput[60]}), .c ({new_AGEMA_signal_8415, RoundOutput[60]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U943 ( .s (new_AGEMA_signal_10560), .b ({new_AGEMA_signal_7436, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]}), .a ({new_AGEMA_signal_8043, MixColumnsOutput[61]}), .c ({new_AGEMA_signal_8242, RoundOutput[61]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U944 ( .s (new_AGEMA_signal_10560), .b ({new_AGEMA_signal_7435, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]}), .a ({new_AGEMA_signal_8041, MixColumnsOutput[62]}), .c ({new_AGEMA_signal_8243, RoundOutput[62]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U945 ( .s (new_AGEMA_signal_10560), .b ({new_AGEMA_signal_7434, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .a ({new_AGEMA_signal_8040, MixColumnsOutput[63]}), .c ({new_AGEMA_signal_8244, RoundOutput[63]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U946 ( .s (new_AGEMA_signal_10560), .b ({new_AGEMA_signal_7319, MixColumnsInput[64]}), .a ({new_AGEMA_signal_8032, MixColumnsOutput[64]}), .c ({new_AGEMA_signal_8245, RoundOutput[64]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U947 ( .s (new_AGEMA_signal_10560), .b ({new_AGEMA_signal_7475, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]}), .a ({new_AGEMA_signal_8289, MixColumnsOutput[65]}), .c ({new_AGEMA_signal_8416, RoundOutput[65]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U948 ( .s (new_AGEMA_signal_10560), .b ({new_AGEMA_signal_7474, MixColumnsInput[66]}), .a ({new_AGEMA_signal_8010, MixColumnsOutput[66]}), .c ({new_AGEMA_signal_8246, RoundOutput[66]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U949 ( .s (new_AGEMA_signal_10560), .b ({new_AGEMA_signal_7473, MixColumnsInput[67]}), .a ({new_AGEMA_signal_8284, MixColumnsOutput[67]}), .c ({new_AGEMA_signal_8417, RoundOutput[67]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U950 ( .s (new_AGEMA_signal_10556), .b ({new_AGEMA_signal_7472, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]}), .a ({new_AGEMA_signal_8283, MixColumnsOutput[68]}), .c ({new_AGEMA_signal_8418, RoundOutput[68]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U951 ( .s (new_AGEMA_signal_10556), .b ({new_AGEMA_signal_7471, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]}), .a ({new_AGEMA_signal_8005, MixColumnsOutput[69]}), .c ({new_AGEMA_signal_8247, RoundOutput[69]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U952 ( .s (new_AGEMA_signal_10556), .b ({new_AGEMA_signal_7414, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]}), .a ({new_AGEMA_signal_8068, MixColumnsOutput[6]}), .c ({new_AGEMA_signal_8248, RoundOutput[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U953 ( .s (new_AGEMA_signal_10556), .b ({new_AGEMA_signal_7470, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]}), .a ({new_AGEMA_signal_8004, MixColumnsOutput[70]}), .c ({new_AGEMA_signal_8249, RoundOutput[70]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U954 ( .s (new_AGEMA_signal_10556), .b ({new_AGEMA_signal_7469, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .a ({new_AGEMA_signal_8003, MixColumnsOutput[71]}), .c ({new_AGEMA_signal_8250, RoundOutput[71]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U955 ( .s (new_AGEMA_signal_10556), .b ({new_AGEMA_signal_7198, MixColumnsInput[72]}), .a ({new_AGEMA_signal_8002, MixColumnsOutput[72]}), .c ({new_AGEMA_signal_8251, RoundOutput[72]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U956 ( .s (new_AGEMA_signal_10556), .b ({new_AGEMA_signal_7398, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]}), .a ({new_AGEMA_signal_8282, MixColumnsOutput[73]}), .c ({new_AGEMA_signal_8419, RoundOutput[73]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U957 ( .s (new_AGEMA_signal_10556), .b ({new_AGEMA_signal_7397, MixColumnsInput[74]}), .a ({new_AGEMA_signal_8031, MixColumnsOutput[74]}), .c ({new_AGEMA_signal_8252, RoundOutput[74]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U958 ( .s (new_AGEMA_signal_10556), .b ({new_AGEMA_signal_7396, MixColumnsInput[75]}), .a ({new_AGEMA_signal_8293, MixColumnsOutput[75]}), .c ({new_AGEMA_signal_8420, RoundOutput[75]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U959 ( .s (new_AGEMA_signal_10556), .b ({new_AGEMA_signal_7395, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]}), .a ({new_AGEMA_signal_8292, MixColumnsOutput[76]}), .c ({new_AGEMA_signal_8421, RoundOutput[76]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U960 ( .s (new_AGEMA_signal_10556), .b ({new_AGEMA_signal_7394, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]}), .a ({new_AGEMA_signal_8028, MixColumnsOutput[77]}), .c ({new_AGEMA_signal_8253, RoundOutput[77]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U961 ( .s (new_AGEMA_signal_10556), .b ({new_AGEMA_signal_7393, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]}), .a ({new_AGEMA_signal_8027, MixColumnsOutput[78]}), .c ({new_AGEMA_signal_8254, RoundOutput[78]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U962 ( .s (new_AGEMA_signal_10552), .b ({new_AGEMA_signal_7392, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .a ({new_AGEMA_signal_8026, MixColumnsOutput[79]}), .c ({new_AGEMA_signal_8255, RoundOutput[79]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U963 ( .s (new_AGEMA_signal_10552), .b ({new_AGEMA_signal_7413, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .a ({new_AGEMA_signal_8067, MixColumnsOutput[7]}), .c ({new_AGEMA_signal_8256, RoundOutput[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U964 ( .s (new_AGEMA_signal_10552), .b ({new_AGEMA_signal_7253, MixColumnsInput[80]}), .a ({new_AGEMA_signal_8025, MixColumnsOutput[80]}), .c ({new_AGEMA_signal_8257, RoundOutput[80]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U965 ( .s (new_AGEMA_signal_10552), .b ({new_AGEMA_signal_7433, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]}), .a ({new_AGEMA_signal_8291, MixColumnsOutput[81]}), .c ({new_AGEMA_signal_8422, RoundOutput[81]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U966 ( .s (new_AGEMA_signal_10552), .b ({new_AGEMA_signal_7432, MixColumnsInput[82]}), .a ({new_AGEMA_signal_8023, MixColumnsOutput[82]}), .c ({new_AGEMA_signal_8258, RoundOutput[82]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U967 ( .s (new_AGEMA_signal_10552), .b ({new_AGEMA_signal_7431, MixColumnsInput[83]}), .a ({new_AGEMA_signal_8290, MixColumnsOutput[83]}), .c ({new_AGEMA_signal_8423, RoundOutput[83]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U968 ( .s (new_AGEMA_signal_10552), .b ({new_AGEMA_signal_7430, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]}), .a ({new_AGEMA_signal_8288, MixColumnsOutput[84]}), .c ({new_AGEMA_signal_8424, RoundOutput[84]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U969 ( .s (new_AGEMA_signal_10552), .b ({new_AGEMA_signal_7429, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]}), .a ({new_AGEMA_signal_8019, MixColumnsOutput[85]}), .c ({new_AGEMA_signal_8259, RoundOutput[85]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U970 ( .s (new_AGEMA_signal_10552), .b ({new_AGEMA_signal_7428, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]}), .a ({new_AGEMA_signal_8018, MixColumnsOutput[86]}), .c ({new_AGEMA_signal_8260, RoundOutput[86]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U971 ( .s (new_AGEMA_signal_10552), .b ({new_AGEMA_signal_7427, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .a ({new_AGEMA_signal_8017, MixColumnsOutput[87]}), .c ({new_AGEMA_signal_8261, RoundOutput[87]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U972 ( .s (new_AGEMA_signal_10552), .b ({new_AGEMA_signal_7308, MixColumnsInput[88]}), .a ({new_AGEMA_signal_8016, MixColumnsOutput[88]}), .c ({new_AGEMA_signal_8262, RoundOutput[88]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U973 ( .s (new_AGEMA_signal_10552), .b ({new_AGEMA_signal_7468, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]}), .a ({new_AGEMA_signal_8287, MixColumnsOutput[89]}), .c ({new_AGEMA_signal_8425, RoundOutput[89]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U974 ( .s (new_AGEMA_signal_10548), .b ({new_AGEMA_signal_7286, MixColumnsInput[8]}), .a ({new_AGEMA_signal_8066, MixColumnsOutput[8]}), .c ({new_AGEMA_signal_8263, RoundOutput[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U975 ( .s (new_AGEMA_signal_10548), .b ({new_AGEMA_signal_7467, MixColumnsInput[90]}), .a ({new_AGEMA_signal_8014, MixColumnsOutput[90]}), .c ({new_AGEMA_signal_8264, RoundOutput[90]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U976 ( .s (new_AGEMA_signal_10548), .b ({new_AGEMA_signal_7466, MixColumnsInput[91]}), .a ({new_AGEMA_signal_8286, MixColumnsOutput[91]}), .c ({new_AGEMA_signal_8426, RoundOutput[91]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U977 ( .s (new_AGEMA_signal_10548), .b ({new_AGEMA_signal_7465, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]}), .a ({new_AGEMA_signal_8285, MixColumnsOutput[92]}), .c ({new_AGEMA_signal_8427, RoundOutput[92]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U978 ( .s (new_AGEMA_signal_10548), .b ({new_AGEMA_signal_7464, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]}), .a ({new_AGEMA_signal_8011, MixColumnsOutput[93]}), .c ({new_AGEMA_signal_8265, RoundOutput[93]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U979 ( .s (new_AGEMA_signal_10548), .b ({new_AGEMA_signal_7463, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]}), .a ({new_AGEMA_signal_8009, MixColumnsOutput[94]}), .c ({new_AGEMA_signal_8266, RoundOutput[94]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U980 ( .s (new_AGEMA_signal_10548), .b ({new_AGEMA_signal_7462, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .a ({new_AGEMA_signal_8008, MixColumnsOutput[95]}), .c ({new_AGEMA_signal_8267, RoundOutput[95]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U981 ( .s (new_AGEMA_signal_10548), .b ({new_AGEMA_signal_7187, MixColumnsInput[96]}), .a ({new_AGEMA_signal_8000, MixColumnsOutput[96]}), .c ({new_AGEMA_signal_8268, RoundOutput[96]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U982 ( .s (new_AGEMA_signal_10548), .b ({new_AGEMA_signal_7391, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]}), .a ({new_AGEMA_signal_8277, MixColumnsOutput[97]}), .c ({new_AGEMA_signal_8428, RoundOutput[97]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U983 ( .s (new_AGEMA_signal_10548), .b ({new_AGEMA_signal_7390, MixColumnsInput[98]}), .a ({new_AGEMA_signal_7978, MixColumnsOutput[98]}), .c ({new_AGEMA_signal_8269, RoundOutput[98]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U984 ( .s (new_AGEMA_signal_10548), .b ({new_AGEMA_signal_7389, MixColumnsInput[99]}), .a ({new_AGEMA_signal_8272, MixColumnsOutput[99]}), .c ({new_AGEMA_signal_8429, RoundOutput[99]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) U985 ( .s (new_AGEMA_signal_10548), .b ({new_AGEMA_signal_7454, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]}), .a ({new_AGEMA_signal_8306, MixColumnsOutput[9]}), .c ({new_AGEMA_signal_8430, RoundOutput[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_0_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8190, RoundOutput[0]}), .a ({new_AGEMA_signal_10580, new_AGEMA_signal_10576}), .c ({new_AGEMA_signal_8432, RoundReg_Inst_ff_SDE_0_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_1_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8397, RoundOutput[1]}), .a ({new_AGEMA_signal_10588, new_AGEMA_signal_10584}), .c ({new_AGEMA_signal_8606, RoundReg_Inst_ff_SDE_1_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_2_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8221, RoundOutput[2]}), .a ({new_AGEMA_signal_10596, new_AGEMA_signal_10592}), .c ({new_AGEMA_signal_8434, RoundReg_Inst_ff_SDE_2_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_3_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8405, RoundOutput[3]}), .a ({new_AGEMA_signal_10604, new_AGEMA_signal_10600}), .c ({new_AGEMA_signal_8608, RoundReg_Inst_ff_SDE_3_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_4_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8410, RoundOutput[4]}), .a ({new_AGEMA_signal_10612, new_AGEMA_signal_10608}), .c ({new_AGEMA_signal_8610, RoundReg_Inst_ff_SDE_4_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_5_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8241, RoundOutput[5]}), .a ({new_AGEMA_signal_10620, new_AGEMA_signal_10616}), .c ({new_AGEMA_signal_8436, RoundReg_Inst_ff_SDE_5_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_6_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8248, RoundOutput[6]}), .a ({new_AGEMA_signal_10628, new_AGEMA_signal_10624}), .c ({new_AGEMA_signal_8438, RoundReg_Inst_ff_SDE_6_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_7_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8256, RoundOutput[7]}), .a ({new_AGEMA_signal_10636, new_AGEMA_signal_10632}), .c ({new_AGEMA_signal_8440, RoundReg_Inst_ff_SDE_7_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_8_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8263, RoundOutput[8]}), .a ({new_AGEMA_signal_10644, new_AGEMA_signal_10640}), .c ({new_AGEMA_signal_8442, RoundReg_Inst_ff_SDE_8_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_9_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8430, RoundOutput[9]}), .a ({new_AGEMA_signal_10652, new_AGEMA_signal_10648}), .c ({new_AGEMA_signal_8612, RoundReg_Inst_ff_SDE_9_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_10_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8197, RoundOutput[10]}), .a ({new_AGEMA_signal_10660, new_AGEMA_signal_10656}), .c ({new_AGEMA_signal_8444, RoundReg_Inst_ff_SDE_10_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_11_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8390, RoundOutput[11]}), .a ({new_AGEMA_signal_10668, new_AGEMA_signal_10664}), .c ({new_AGEMA_signal_8614, RoundReg_Inst_ff_SDE_11_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_12_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8394, RoundOutput[12]}), .a ({new_AGEMA_signal_10676, new_AGEMA_signal_10672}), .c ({new_AGEMA_signal_8616, RoundReg_Inst_ff_SDE_12_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_13_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8210, RoundOutput[13]}), .a ({new_AGEMA_signal_10684, new_AGEMA_signal_10680}), .c ({new_AGEMA_signal_8446, RoundReg_Inst_ff_SDE_13_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_14_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8211, RoundOutput[14]}), .a ({new_AGEMA_signal_10692, new_AGEMA_signal_10688}), .c ({new_AGEMA_signal_8448, RoundReg_Inst_ff_SDE_14_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_15_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8212, RoundOutput[15]}), .a ({new_AGEMA_signal_10700, new_AGEMA_signal_10696}), .c ({new_AGEMA_signal_8450, RoundReg_Inst_ff_SDE_15_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_16_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8213, RoundOutput[16]}), .a ({new_AGEMA_signal_10708, new_AGEMA_signal_10704}), .c ({new_AGEMA_signal_8452, RoundReg_Inst_ff_SDE_16_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_17_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8395, RoundOutput[17]}), .a ({new_AGEMA_signal_10716, new_AGEMA_signal_10712}), .c ({new_AGEMA_signal_8618, RoundReg_Inst_ff_SDE_17_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_18_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8214, RoundOutput[18]}), .a ({new_AGEMA_signal_10724, new_AGEMA_signal_10720}), .c ({new_AGEMA_signal_8454, RoundReg_Inst_ff_SDE_18_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_19_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8396, RoundOutput[19]}), .a ({new_AGEMA_signal_10732, new_AGEMA_signal_10728}), .c ({new_AGEMA_signal_8620, RoundReg_Inst_ff_SDE_19_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_20_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8398, RoundOutput[20]}), .a ({new_AGEMA_signal_10740, new_AGEMA_signal_10736}), .c ({new_AGEMA_signal_8622, RoundReg_Inst_ff_SDE_20_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_21_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8215, RoundOutput[21]}), .a ({new_AGEMA_signal_10748, new_AGEMA_signal_10744}), .c ({new_AGEMA_signal_8456, RoundReg_Inst_ff_SDE_21_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_22_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8216, RoundOutput[22]}), .a ({new_AGEMA_signal_10756, new_AGEMA_signal_10752}), .c ({new_AGEMA_signal_8458, RoundReg_Inst_ff_SDE_22_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_23_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8217, RoundOutput[23]}), .a ({new_AGEMA_signal_10764, new_AGEMA_signal_10760}), .c ({new_AGEMA_signal_8460, RoundReg_Inst_ff_SDE_23_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_24_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8218, RoundOutput[24]}), .a ({new_AGEMA_signal_10772, new_AGEMA_signal_10768}), .c ({new_AGEMA_signal_8462, RoundReg_Inst_ff_SDE_24_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_25_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8399, RoundOutput[25]}), .a ({new_AGEMA_signal_10780, new_AGEMA_signal_10776}), .c ({new_AGEMA_signal_8624, RoundReg_Inst_ff_SDE_25_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_26_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8219, RoundOutput[26]}), .a ({new_AGEMA_signal_10788, new_AGEMA_signal_10784}), .c ({new_AGEMA_signal_8464, RoundReg_Inst_ff_SDE_26_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_27_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8400, RoundOutput[27]}), .a ({new_AGEMA_signal_10796, new_AGEMA_signal_10792}), .c ({new_AGEMA_signal_8626, RoundReg_Inst_ff_SDE_27_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_28_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8401, RoundOutput[28]}), .a ({new_AGEMA_signal_10804, new_AGEMA_signal_10800}), .c ({new_AGEMA_signal_8628, RoundReg_Inst_ff_SDE_28_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_29_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8220, RoundOutput[29]}), .a ({new_AGEMA_signal_10812, new_AGEMA_signal_10808}), .c ({new_AGEMA_signal_8466, RoundReg_Inst_ff_SDE_29_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_30_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8222, RoundOutput[30]}), .a ({new_AGEMA_signal_10820, new_AGEMA_signal_10816}), .c ({new_AGEMA_signal_8468, RoundReg_Inst_ff_SDE_30_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_31_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8223, RoundOutput[31]}), .a ({new_AGEMA_signal_10828, new_AGEMA_signal_10824}), .c ({new_AGEMA_signal_8470, RoundReg_Inst_ff_SDE_31_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_32_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8224, RoundOutput[32]}), .a ({new_AGEMA_signal_10836, new_AGEMA_signal_10832}), .c ({new_AGEMA_signal_8472, RoundReg_Inst_ff_SDE_32_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_33_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8402, RoundOutput[33]}), .a ({new_AGEMA_signal_10844, new_AGEMA_signal_10840}), .c ({new_AGEMA_signal_8630, RoundReg_Inst_ff_SDE_33_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_34_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8225, RoundOutput[34]}), .a ({new_AGEMA_signal_10852, new_AGEMA_signal_10848}), .c ({new_AGEMA_signal_8474, RoundReg_Inst_ff_SDE_34_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_35_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8403, RoundOutput[35]}), .a ({new_AGEMA_signal_10860, new_AGEMA_signal_10856}), .c ({new_AGEMA_signal_8632, RoundReg_Inst_ff_SDE_35_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_36_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8404, RoundOutput[36]}), .a ({new_AGEMA_signal_10868, new_AGEMA_signal_10864}), .c ({new_AGEMA_signal_8634, RoundReg_Inst_ff_SDE_36_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_37_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8226, RoundOutput[37]}), .a ({new_AGEMA_signal_10876, new_AGEMA_signal_10872}), .c ({new_AGEMA_signal_8476, RoundReg_Inst_ff_SDE_37_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_38_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8227, RoundOutput[38]}), .a ({new_AGEMA_signal_10884, new_AGEMA_signal_10880}), .c ({new_AGEMA_signal_8478, RoundReg_Inst_ff_SDE_38_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_39_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8228, RoundOutput[39]}), .a ({new_AGEMA_signal_10892, new_AGEMA_signal_10888}), .c ({new_AGEMA_signal_8480, RoundReg_Inst_ff_SDE_39_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_40_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8229, RoundOutput[40]}), .a ({new_AGEMA_signal_10900, new_AGEMA_signal_10896}), .c ({new_AGEMA_signal_8482, RoundReg_Inst_ff_SDE_40_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_41_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8406, RoundOutput[41]}), .a ({new_AGEMA_signal_10908, new_AGEMA_signal_10904}), .c ({new_AGEMA_signal_8636, RoundReg_Inst_ff_SDE_41_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_42_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8230, RoundOutput[42]}), .a ({new_AGEMA_signal_10916, new_AGEMA_signal_10912}), .c ({new_AGEMA_signal_8484, RoundReg_Inst_ff_SDE_42_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_43_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8407, RoundOutput[43]}), .a ({new_AGEMA_signal_10924, new_AGEMA_signal_10920}), .c ({new_AGEMA_signal_8638, RoundReg_Inst_ff_SDE_43_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_44_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8408, RoundOutput[44]}), .a ({new_AGEMA_signal_10932, new_AGEMA_signal_10928}), .c ({new_AGEMA_signal_8640, RoundReg_Inst_ff_SDE_44_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_45_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8231, RoundOutput[45]}), .a ({new_AGEMA_signal_10940, new_AGEMA_signal_10936}), .c ({new_AGEMA_signal_8486, RoundReg_Inst_ff_SDE_45_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_46_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8232, RoundOutput[46]}), .a ({new_AGEMA_signal_10948, new_AGEMA_signal_10944}), .c ({new_AGEMA_signal_8488, RoundReg_Inst_ff_SDE_46_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_47_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8233, RoundOutput[47]}), .a ({new_AGEMA_signal_10956, new_AGEMA_signal_10952}), .c ({new_AGEMA_signal_8490, RoundReg_Inst_ff_SDE_47_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_48_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8234, RoundOutput[48]}), .a ({new_AGEMA_signal_10964, new_AGEMA_signal_10960}), .c ({new_AGEMA_signal_8492, RoundReg_Inst_ff_SDE_48_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_49_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8409, RoundOutput[49]}), .a ({new_AGEMA_signal_10972, new_AGEMA_signal_10968}), .c ({new_AGEMA_signal_8642, RoundReg_Inst_ff_SDE_49_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_50_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8235, RoundOutput[50]}), .a ({new_AGEMA_signal_10980, new_AGEMA_signal_10976}), .c ({new_AGEMA_signal_8494, RoundReg_Inst_ff_SDE_50_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_51_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8411, RoundOutput[51]}), .a ({new_AGEMA_signal_10988, new_AGEMA_signal_10984}), .c ({new_AGEMA_signal_8644, RoundReg_Inst_ff_SDE_51_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_52_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8412, RoundOutput[52]}), .a ({new_AGEMA_signal_10996, new_AGEMA_signal_10992}), .c ({new_AGEMA_signal_8646, RoundReg_Inst_ff_SDE_52_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_53_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8236, RoundOutput[53]}), .a ({new_AGEMA_signal_11004, new_AGEMA_signal_11000}), .c ({new_AGEMA_signal_8496, RoundReg_Inst_ff_SDE_53_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_54_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8237, RoundOutput[54]}), .a ({new_AGEMA_signal_11012, new_AGEMA_signal_11008}), .c ({new_AGEMA_signal_8498, RoundReg_Inst_ff_SDE_54_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_55_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8238, RoundOutput[55]}), .a ({new_AGEMA_signal_11020, new_AGEMA_signal_11016}), .c ({new_AGEMA_signal_8500, RoundReg_Inst_ff_SDE_55_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_56_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8239, RoundOutput[56]}), .a ({new_AGEMA_signal_11028, new_AGEMA_signal_11024}), .c ({new_AGEMA_signal_8502, RoundReg_Inst_ff_SDE_56_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_57_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8413, RoundOutput[57]}), .a ({new_AGEMA_signal_11036, new_AGEMA_signal_11032}), .c ({new_AGEMA_signal_8648, RoundReg_Inst_ff_SDE_57_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_58_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8240, RoundOutput[58]}), .a ({new_AGEMA_signal_11044, new_AGEMA_signal_11040}), .c ({new_AGEMA_signal_8504, RoundReg_Inst_ff_SDE_58_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_59_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8414, RoundOutput[59]}), .a ({new_AGEMA_signal_11052, new_AGEMA_signal_11048}), .c ({new_AGEMA_signal_8650, RoundReg_Inst_ff_SDE_59_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_60_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8415, RoundOutput[60]}), .a ({new_AGEMA_signal_11060, new_AGEMA_signal_11056}), .c ({new_AGEMA_signal_8652, RoundReg_Inst_ff_SDE_60_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_61_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8242, RoundOutput[61]}), .a ({new_AGEMA_signal_11068, new_AGEMA_signal_11064}), .c ({new_AGEMA_signal_8506, RoundReg_Inst_ff_SDE_61_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_62_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8243, RoundOutput[62]}), .a ({new_AGEMA_signal_11076, new_AGEMA_signal_11072}), .c ({new_AGEMA_signal_8508, RoundReg_Inst_ff_SDE_62_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_63_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8244, RoundOutput[63]}), .a ({new_AGEMA_signal_11084, new_AGEMA_signal_11080}), .c ({new_AGEMA_signal_8510, RoundReg_Inst_ff_SDE_63_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_64_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8245, RoundOutput[64]}), .a ({new_AGEMA_signal_11092, new_AGEMA_signal_11088}), .c ({new_AGEMA_signal_8512, RoundReg_Inst_ff_SDE_64_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_65_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8416, RoundOutput[65]}), .a ({new_AGEMA_signal_11100, new_AGEMA_signal_11096}), .c ({new_AGEMA_signal_8654, RoundReg_Inst_ff_SDE_65_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_66_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8246, RoundOutput[66]}), .a ({new_AGEMA_signal_11108, new_AGEMA_signal_11104}), .c ({new_AGEMA_signal_8514, RoundReg_Inst_ff_SDE_66_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_67_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8417, RoundOutput[67]}), .a ({new_AGEMA_signal_11116, new_AGEMA_signal_11112}), .c ({new_AGEMA_signal_8656, RoundReg_Inst_ff_SDE_67_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_68_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8418, RoundOutput[68]}), .a ({new_AGEMA_signal_11124, new_AGEMA_signal_11120}), .c ({new_AGEMA_signal_8658, RoundReg_Inst_ff_SDE_68_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_69_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8247, RoundOutput[69]}), .a ({new_AGEMA_signal_11132, new_AGEMA_signal_11128}), .c ({new_AGEMA_signal_8516, RoundReg_Inst_ff_SDE_69_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_70_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8249, RoundOutput[70]}), .a ({new_AGEMA_signal_11140, new_AGEMA_signal_11136}), .c ({new_AGEMA_signal_8518, RoundReg_Inst_ff_SDE_70_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_71_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8250, RoundOutput[71]}), .a ({new_AGEMA_signal_11148, new_AGEMA_signal_11144}), .c ({new_AGEMA_signal_8520, RoundReg_Inst_ff_SDE_71_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_72_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8251, RoundOutput[72]}), .a ({new_AGEMA_signal_11156, new_AGEMA_signal_11152}), .c ({new_AGEMA_signal_8522, RoundReg_Inst_ff_SDE_72_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_73_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8419, RoundOutput[73]}), .a ({new_AGEMA_signal_11164, new_AGEMA_signal_11160}), .c ({new_AGEMA_signal_8660, RoundReg_Inst_ff_SDE_73_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_74_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8252, RoundOutput[74]}), .a ({new_AGEMA_signal_11172, new_AGEMA_signal_11168}), .c ({new_AGEMA_signal_8524, RoundReg_Inst_ff_SDE_74_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_75_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8420, RoundOutput[75]}), .a ({new_AGEMA_signal_11180, new_AGEMA_signal_11176}), .c ({new_AGEMA_signal_8662, RoundReg_Inst_ff_SDE_75_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_76_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8421, RoundOutput[76]}), .a ({new_AGEMA_signal_11188, new_AGEMA_signal_11184}), .c ({new_AGEMA_signal_8664, RoundReg_Inst_ff_SDE_76_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_77_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8253, RoundOutput[77]}), .a ({new_AGEMA_signal_11196, new_AGEMA_signal_11192}), .c ({new_AGEMA_signal_8526, RoundReg_Inst_ff_SDE_77_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_78_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8254, RoundOutput[78]}), .a ({new_AGEMA_signal_11204, new_AGEMA_signal_11200}), .c ({new_AGEMA_signal_8528, RoundReg_Inst_ff_SDE_78_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_79_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8255, RoundOutput[79]}), .a ({new_AGEMA_signal_11212, new_AGEMA_signal_11208}), .c ({new_AGEMA_signal_8530, RoundReg_Inst_ff_SDE_79_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_80_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8257, RoundOutput[80]}), .a ({new_AGEMA_signal_11220, new_AGEMA_signal_11216}), .c ({new_AGEMA_signal_8532, RoundReg_Inst_ff_SDE_80_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_81_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8422, RoundOutput[81]}), .a ({new_AGEMA_signal_11228, new_AGEMA_signal_11224}), .c ({new_AGEMA_signal_8666, RoundReg_Inst_ff_SDE_81_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_82_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8258, RoundOutput[82]}), .a ({new_AGEMA_signal_11236, new_AGEMA_signal_11232}), .c ({new_AGEMA_signal_8534, RoundReg_Inst_ff_SDE_82_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_83_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8423, RoundOutput[83]}), .a ({new_AGEMA_signal_11244, new_AGEMA_signal_11240}), .c ({new_AGEMA_signal_8668, RoundReg_Inst_ff_SDE_83_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_84_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8424, RoundOutput[84]}), .a ({new_AGEMA_signal_11252, new_AGEMA_signal_11248}), .c ({new_AGEMA_signal_8670, RoundReg_Inst_ff_SDE_84_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_85_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8259, RoundOutput[85]}), .a ({new_AGEMA_signal_11260, new_AGEMA_signal_11256}), .c ({new_AGEMA_signal_8536, RoundReg_Inst_ff_SDE_85_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_86_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8260, RoundOutput[86]}), .a ({new_AGEMA_signal_11268, new_AGEMA_signal_11264}), .c ({new_AGEMA_signal_8538, RoundReg_Inst_ff_SDE_86_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_87_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8261, RoundOutput[87]}), .a ({new_AGEMA_signal_11276, new_AGEMA_signal_11272}), .c ({new_AGEMA_signal_8540, RoundReg_Inst_ff_SDE_87_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_88_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8262, RoundOutput[88]}), .a ({new_AGEMA_signal_11284, new_AGEMA_signal_11280}), .c ({new_AGEMA_signal_8542, RoundReg_Inst_ff_SDE_88_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_89_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8425, RoundOutput[89]}), .a ({new_AGEMA_signal_11292, new_AGEMA_signal_11288}), .c ({new_AGEMA_signal_8672, RoundReg_Inst_ff_SDE_89_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_90_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8264, RoundOutput[90]}), .a ({new_AGEMA_signal_11300, new_AGEMA_signal_11296}), .c ({new_AGEMA_signal_8544, RoundReg_Inst_ff_SDE_90_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_91_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8426, RoundOutput[91]}), .a ({new_AGEMA_signal_11308, new_AGEMA_signal_11304}), .c ({new_AGEMA_signal_8674, RoundReg_Inst_ff_SDE_91_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_92_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8427, RoundOutput[92]}), .a ({new_AGEMA_signal_11316, new_AGEMA_signal_11312}), .c ({new_AGEMA_signal_8676, RoundReg_Inst_ff_SDE_92_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_93_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8265, RoundOutput[93]}), .a ({new_AGEMA_signal_11324, new_AGEMA_signal_11320}), .c ({new_AGEMA_signal_8546, RoundReg_Inst_ff_SDE_93_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_94_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8266, RoundOutput[94]}), .a ({new_AGEMA_signal_11332, new_AGEMA_signal_11328}), .c ({new_AGEMA_signal_8548, RoundReg_Inst_ff_SDE_94_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_95_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8267, RoundOutput[95]}), .a ({new_AGEMA_signal_11340, new_AGEMA_signal_11336}), .c ({new_AGEMA_signal_8550, RoundReg_Inst_ff_SDE_95_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_96_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8268, RoundOutput[96]}), .a ({new_AGEMA_signal_11348, new_AGEMA_signal_11344}), .c ({new_AGEMA_signal_8552, RoundReg_Inst_ff_SDE_96_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_97_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8428, RoundOutput[97]}), .a ({new_AGEMA_signal_11356, new_AGEMA_signal_11352}), .c ({new_AGEMA_signal_8678, RoundReg_Inst_ff_SDE_97_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_98_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8269, RoundOutput[98]}), .a ({new_AGEMA_signal_11364, new_AGEMA_signal_11360}), .c ({new_AGEMA_signal_8554, RoundReg_Inst_ff_SDE_98_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_99_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8429, RoundOutput[99]}), .a ({new_AGEMA_signal_11372, new_AGEMA_signal_11368}), .c ({new_AGEMA_signal_8680, RoundReg_Inst_ff_SDE_99_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_100_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8383, RoundOutput[100]}), .a ({new_AGEMA_signal_11380, new_AGEMA_signal_11376}), .c ({new_AGEMA_signal_8682, RoundReg_Inst_ff_SDE_100_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_101_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8191, RoundOutput[101]}), .a ({new_AGEMA_signal_11388, new_AGEMA_signal_11384}), .c ({new_AGEMA_signal_8556, RoundReg_Inst_ff_SDE_101_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_102_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8192, RoundOutput[102]}), .a ({new_AGEMA_signal_11396, new_AGEMA_signal_11392}), .c ({new_AGEMA_signal_8558, RoundReg_Inst_ff_SDE_102_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_103_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8193, RoundOutput[103]}), .a ({new_AGEMA_signal_11404, new_AGEMA_signal_11400}), .c ({new_AGEMA_signal_8560, RoundReg_Inst_ff_SDE_103_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_104_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8194, RoundOutput[104]}), .a ({new_AGEMA_signal_11412, new_AGEMA_signal_11408}), .c ({new_AGEMA_signal_8562, RoundReg_Inst_ff_SDE_104_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_105_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8384, RoundOutput[105]}), .a ({new_AGEMA_signal_11420, new_AGEMA_signal_11416}), .c ({new_AGEMA_signal_8684, RoundReg_Inst_ff_SDE_105_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_106_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8195, RoundOutput[106]}), .a ({new_AGEMA_signal_11428, new_AGEMA_signal_11424}), .c ({new_AGEMA_signal_8564, RoundReg_Inst_ff_SDE_106_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_107_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8385, RoundOutput[107]}), .a ({new_AGEMA_signal_11436, new_AGEMA_signal_11432}), .c ({new_AGEMA_signal_8686, RoundReg_Inst_ff_SDE_107_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_108_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8386, RoundOutput[108]}), .a ({new_AGEMA_signal_11444, new_AGEMA_signal_11440}), .c ({new_AGEMA_signal_8688, RoundReg_Inst_ff_SDE_108_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_109_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8196, RoundOutput[109]}), .a ({new_AGEMA_signal_11452, new_AGEMA_signal_11448}), .c ({new_AGEMA_signal_8566, RoundReg_Inst_ff_SDE_109_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_110_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8198, RoundOutput[110]}), .a ({new_AGEMA_signal_11460, new_AGEMA_signal_11456}), .c ({new_AGEMA_signal_8568, RoundReg_Inst_ff_SDE_110_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_111_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8199, RoundOutput[111]}), .a ({new_AGEMA_signal_11468, new_AGEMA_signal_11464}), .c ({new_AGEMA_signal_8570, RoundReg_Inst_ff_SDE_111_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_112_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8200, RoundOutput[112]}), .a ({new_AGEMA_signal_11476, new_AGEMA_signal_11472}), .c ({new_AGEMA_signal_8572, RoundReg_Inst_ff_SDE_112_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_113_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8387, RoundOutput[113]}), .a ({new_AGEMA_signal_11484, new_AGEMA_signal_11480}), .c ({new_AGEMA_signal_8690, RoundReg_Inst_ff_SDE_113_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_114_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8201, RoundOutput[114]}), .a ({new_AGEMA_signal_11492, new_AGEMA_signal_11488}), .c ({new_AGEMA_signal_8574, RoundReg_Inst_ff_SDE_114_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_115_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8388, RoundOutput[115]}), .a ({new_AGEMA_signal_11500, new_AGEMA_signal_11496}), .c ({new_AGEMA_signal_8692, RoundReg_Inst_ff_SDE_115_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_116_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8389, RoundOutput[116]}), .a ({new_AGEMA_signal_11508, new_AGEMA_signal_11504}), .c ({new_AGEMA_signal_8694, RoundReg_Inst_ff_SDE_116_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_117_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8202, RoundOutput[117]}), .a ({new_AGEMA_signal_11516, new_AGEMA_signal_11512}), .c ({new_AGEMA_signal_8576, RoundReg_Inst_ff_SDE_117_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_118_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8203, RoundOutput[118]}), .a ({new_AGEMA_signal_11524, new_AGEMA_signal_11520}), .c ({new_AGEMA_signal_8578, RoundReg_Inst_ff_SDE_118_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_119_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8204, RoundOutput[119]}), .a ({new_AGEMA_signal_11532, new_AGEMA_signal_11528}), .c ({new_AGEMA_signal_8580, RoundReg_Inst_ff_SDE_119_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_120_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8205, RoundOutput[120]}), .a ({new_AGEMA_signal_11540, new_AGEMA_signal_11536}), .c ({new_AGEMA_signal_8582, RoundReg_Inst_ff_SDE_120_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_121_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8391, RoundOutput[121]}), .a ({new_AGEMA_signal_11548, new_AGEMA_signal_11544}), .c ({new_AGEMA_signal_8696, RoundReg_Inst_ff_SDE_121_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_122_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8206, RoundOutput[122]}), .a ({new_AGEMA_signal_11556, new_AGEMA_signal_11552}), .c ({new_AGEMA_signal_8584, RoundReg_Inst_ff_SDE_122_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_123_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8392, RoundOutput[123]}), .a ({new_AGEMA_signal_11564, new_AGEMA_signal_11560}), .c ({new_AGEMA_signal_8698, RoundReg_Inst_ff_SDE_123_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_124_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8393, RoundOutput[124]}), .a ({new_AGEMA_signal_11572, new_AGEMA_signal_11568}), .c ({new_AGEMA_signal_8700, RoundReg_Inst_ff_SDE_124_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_125_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8207, RoundOutput[125]}), .a ({new_AGEMA_signal_11580, new_AGEMA_signal_11576}), .c ({new_AGEMA_signal_8586, RoundReg_Inst_ff_SDE_125_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_126_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8208, RoundOutput[126]}), .a ({new_AGEMA_signal_11588, new_AGEMA_signal_11584}), .c ({new_AGEMA_signal_8588, RoundReg_Inst_ff_SDE_126_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_127_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8209, RoundOutput[127]}), .a ({new_AGEMA_signal_11596, new_AGEMA_signal_11592}), .c ({new_AGEMA_signal_8590, RoundReg_Inst_ff_SDE_127_next_state}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M46_U1 ( .a ({new_AGEMA_signal_6324, SubBytesIns_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_11602, new_AGEMA_signal_11599}), .clk (clk), .r ({Fresh[641], Fresh[640]}), .c ({new_AGEMA_signal_6562, SubBytesIns_Inst_Sbox_0_M46}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M47_U1 ( .a ({new_AGEMA_signal_6212, SubBytesIns_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_11608, new_AGEMA_signal_11605}), .clk (clk), .r ({Fresh[643], Fresh[642]}), .c ({new_AGEMA_signal_6325, SubBytesIns_Inst_Sbox_0_M47}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M48_U1 ( .a ({new_AGEMA_signal_6211, SubBytesIns_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_11614, new_AGEMA_signal_11611}), .clk (clk), .r ({Fresh[645], Fresh[644]}), .c ({new_AGEMA_signal_6326, SubBytesIns_Inst_Sbox_0_M48}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M49_U1 ( .a ({new_AGEMA_signal_6323, SubBytesIns_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_11620, new_AGEMA_signal_11617}), .clk (clk), .r ({Fresh[647], Fresh[646]}), .c ({new_AGEMA_signal_6563, SubBytesIns_Inst_Sbox_0_M49}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M50_U1 ( .a ({new_AGEMA_signal_6210, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_11626, new_AGEMA_signal_11623}), .clk (clk), .r ({Fresh[649], Fresh[648]}), .c ({new_AGEMA_signal_6327, SubBytesIns_Inst_Sbox_0_M50}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M51_U1 ( .a ({new_AGEMA_signal_6209, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_11632, new_AGEMA_signal_11629}), .clk (clk), .r ({Fresh[651], Fresh[650]}), .c ({new_AGEMA_signal_6328, SubBytesIns_Inst_Sbox_0_M51}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M52_U1 ( .a ({new_AGEMA_signal_6322, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_11638, new_AGEMA_signal_11635}), .clk (clk), .r ({Fresh[653], Fresh[652]}), .c ({new_AGEMA_signal_6564, SubBytesIns_Inst_Sbox_0_M52}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M53_U1 ( .a ({new_AGEMA_signal_6561, SubBytesIns_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_11644, new_AGEMA_signal_11641}), .clk (clk), .r ({Fresh[655], Fresh[654]}), .c ({new_AGEMA_signal_6793, SubBytesIns_Inst_Sbox_0_M53}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M54_U1 ( .a ({new_AGEMA_signal_6321, SubBytesIns_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_11650, new_AGEMA_signal_11647}), .clk (clk), .r ({Fresh[657], Fresh[656]}), .c ({new_AGEMA_signal_6565, SubBytesIns_Inst_Sbox_0_M54}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M55_U1 ( .a ({new_AGEMA_signal_6324, SubBytesIns_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_11656, new_AGEMA_signal_11653}), .clk (clk), .r ({Fresh[659], Fresh[658]}), .c ({new_AGEMA_signal_6566, SubBytesIns_Inst_Sbox_0_M55}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M56_U1 ( .a ({new_AGEMA_signal_6212, SubBytesIns_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_11662, new_AGEMA_signal_11659}), .clk (clk), .r ({Fresh[661], Fresh[660]}), .c ({new_AGEMA_signal_6329, SubBytesIns_Inst_Sbox_0_M56}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M57_U1 ( .a ({new_AGEMA_signal_6211, SubBytesIns_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_11668, new_AGEMA_signal_11665}), .clk (clk), .r ({Fresh[663], Fresh[662]}), .c ({new_AGEMA_signal_6330, SubBytesIns_Inst_Sbox_0_M57}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M58_U1 ( .a ({new_AGEMA_signal_6323, SubBytesIns_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_11674, new_AGEMA_signal_11671}), .clk (clk), .r ({Fresh[665], Fresh[664]}), .c ({new_AGEMA_signal_6567, SubBytesIns_Inst_Sbox_0_M58}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M59_U1 ( .a ({new_AGEMA_signal_6210, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_11680, new_AGEMA_signal_11677}), .clk (clk), .r ({Fresh[667], Fresh[666]}), .c ({new_AGEMA_signal_6331, SubBytesIns_Inst_Sbox_0_M59}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M60_U1 ( .a ({new_AGEMA_signal_6209, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_11686, new_AGEMA_signal_11683}), .clk (clk), .r ({Fresh[669], Fresh[668]}), .c ({new_AGEMA_signal_6332, SubBytesIns_Inst_Sbox_0_M60}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M61_U1 ( .a ({new_AGEMA_signal_6322, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_11692, new_AGEMA_signal_11689}), .clk (clk), .r ({Fresh[671], Fresh[670]}), .c ({new_AGEMA_signal_6568, SubBytesIns_Inst_Sbox_0_M61}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M62_U1 ( .a ({new_AGEMA_signal_6561, SubBytesIns_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_11698, new_AGEMA_signal_11695}), .clk (clk), .r ({Fresh[673], Fresh[672]}), .c ({new_AGEMA_signal_6794, SubBytesIns_Inst_Sbox_0_M62}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M63_U1 ( .a ({new_AGEMA_signal_6321, SubBytesIns_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_11704, new_AGEMA_signal_11701}), .clk (clk), .r ({Fresh[675], Fresh[674]}), .c ({new_AGEMA_signal_6569, SubBytesIns_Inst_Sbox_0_M63}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L0_U1 ( .a ({new_AGEMA_signal_6568, SubBytesIns_Inst_Sbox_0_M61}), .b ({new_AGEMA_signal_6794, SubBytesIns_Inst_Sbox_0_M62}), .c ({new_AGEMA_signal_6989, SubBytesIns_Inst_Sbox_0_L0}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L1_U1 ( .a ({new_AGEMA_signal_6327, SubBytesIns_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_6329, SubBytesIns_Inst_Sbox_0_M56}), .c ({new_AGEMA_signal_6570, SubBytesIns_Inst_Sbox_0_L1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L2_U1 ( .a ({new_AGEMA_signal_6562, SubBytesIns_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_6326, SubBytesIns_Inst_Sbox_0_M48}), .c ({new_AGEMA_signal_6795, SubBytesIns_Inst_Sbox_0_L2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L3_U1 ( .a ({new_AGEMA_signal_6325, SubBytesIns_Inst_Sbox_0_M47}), .b ({new_AGEMA_signal_6566, SubBytesIns_Inst_Sbox_0_M55}), .c ({new_AGEMA_signal_6796, SubBytesIns_Inst_Sbox_0_L3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L4_U1 ( .a ({new_AGEMA_signal_6565, SubBytesIns_Inst_Sbox_0_M54}), .b ({new_AGEMA_signal_6567, SubBytesIns_Inst_Sbox_0_M58}), .c ({new_AGEMA_signal_6797, SubBytesIns_Inst_Sbox_0_L4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L5_U1 ( .a ({new_AGEMA_signal_6563, SubBytesIns_Inst_Sbox_0_M49}), .b ({new_AGEMA_signal_6568, SubBytesIns_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_6798, SubBytesIns_Inst_Sbox_0_L5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L6_U1 ( .a ({new_AGEMA_signal_6794, SubBytesIns_Inst_Sbox_0_M62}), .b ({new_AGEMA_signal_6798, SubBytesIns_Inst_Sbox_0_L5}), .c ({new_AGEMA_signal_6990, SubBytesIns_Inst_Sbox_0_L6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L7_U1 ( .a ({new_AGEMA_signal_6562, SubBytesIns_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_6796, SubBytesIns_Inst_Sbox_0_L3}), .c ({new_AGEMA_signal_6991, SubBytesIns_Inst_Sbox_0_L7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L8_U1 ( .a ({new_AGEMA_signal_6328, SubBytesIns_Inst_Sbox_0_M51}), .b ({new_AGEMA_signal_6331, SubBytesIns_Inst_Sbox_0_M59}), .c ({new_AGEMA_signal_6571, SubBytesIns_Inst_Sbox_0_L8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L9_U1 ( .a ({new_AGEMA_signal_6564, SubBytesIns_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_6793, SubBytesIns_Inst_Sbox_0_M53}), .c ({new_AGEMA_signal_6992, SubBytesIns_Inst_Sbox_0_L9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L10_U1 ( .a ({new_AGEMA_signal_6793, SubBytesIns_Inst_Sbox_0_M53}), .b ({new_AGEMA_signal_6797, SubBytesIns_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_6993, SubBytesIns_Inst_Sbox_0_L10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L11_U1 ( .a ({new_AGEMA_signal_6332, SubBytesIns_Inst_Sbox_0_M60}), .b ({new_AGEMA_signal_6795, SubBytesIns_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_6994, SubBytesIns_Inst_Sbox_0_L11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L12_U1 ( .a ({new_AGEMA_signal_6326, SubBytesIns_Inst_Sbox_0_M48}), .b ({new_AGEMA_signal_6328, SubBytesIns_Inst_Sbox_0_M51}), .c ({new_AGEMA_signal_6572, SubBytesIns_Inst_Sbox_0_L12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L13_U1 ( .a ({new_AGEMA_signal_6327, SubBytesIns_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_6989, SubBytesIns_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_7177, SubBytesIns_Inst_Sbox_0_L13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L14_U1 ( .a ({new_AGEMA_signal_6564, SubBytesIns_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_6568, SubBytesIns_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_6799, SubBytesIns_Inst_Sbox_0_L14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L15_U1 ( .a ({new_AGEMA_signal_6566, SubBytesIns_Inst_Sbox_0_M55}), .b ({new_AGEMA_signal_6570, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_6800, SubBytesIns_Inst_Sbox_0_L15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L16_U1 ( .a ({new_AGEMA_signal_6329, SubBytesIns_Inst_Sbox_0_M56}), .b ({new_AGEMA_signal_6989, SubBytesIns_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_7178, SubBytesIns_Inst_Sbox_0_L16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L17_U1 ( .a ({new_AGEMA_signal_6330, SubBytesIns_Inst_Sbox_0_M57}), .b ({new_AGEMA_signal_6570, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_6801, SubBytesIns_Inst_Sbox_0_L17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L18_U1 ( .a ({new_AGEMA_signal_6567, SubBytesIns_Inst_Sbox_0_M58}), .b ({new_AGEMA_signal_6571, SubBytesIns_Inst_Sbox_0_L8}), .c ({new_AGEMA_signal_6802, SubBytesIns_Inst_Sbox_0_L18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L19_U1 ( .a ({new_AGEMA_signal_6569, SubBytesIns_Inst_Sbox_0_M63}), .b ({new_AGEMA_signal_6797, SubBytesIns_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_6995, SubBytesIns_Inst_Sbox_0_L19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L20_U1 ( .a ({new_AGEMA_signal_6989, SubBytesIns_Inst_Sbox_0_L0}), .b ({new_AGEMA_signal_6570, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_7179, SubBytesIns_Inst_Sbox_0_L20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L21_U1 ( .a ({new_AGEMA_signal_6570, SubBytesIns_Inst_Sbox_0_L1}), .b ({new_AGEMA_signal_6991, SubBytesIns_Inst_Sbox_0_L7}), .c ({new_AGEMA_signal_7180, SubBytesIns_Inst_Sbox_0_L21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L22_U1 ( .a ({new_AGEMA_signal_6796, SubBytesIns_Inst_Sbox_0_L3}), .b ({new_AGEMA_signal_6572, SubBytesIns_Inst_Sbox_0_L12}), .c ({new_AGEMA_signal_6996, SubBytesIns_Inst_Sbox_0_L22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L23_U1 ( .a ({new_AGEMA_signal_6802, SubBytesIns_Inst_Sbox_0_L18}), .b ({new_AGEMA_signal_6795, SubBytesIns_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_6997, SubBytesIns_Inst_Sbox_0_L23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L24_U1 ( .a ({new_AGEMA_signal_6800, SubBytesIns_Inst_Sbox_0_L15}), .b ({new_AGEMA_signal_6992, SubBytesIns_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_7181, SubBytesIns_Inst_Sbox_0_L24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L25_U1 ( .a ({new_AGEMA_signal_6990, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_6993, SubBytesIns_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_7182, SubBytesIns_Inst_Sbox_0_L25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L26_U1 ( .a ({new_AGEMA_signal_6991, SubBytesIns_Inst_Sbox_0_L7}), .b ({new_AGEMA_signal_6992, SubBytesIns_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_7183, SubBytesIns_Inst_Sbox_0_L26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L27_U1 ( .a ({new_AGEMA_signal_6571, SubBytesIns_Inst_Sbox_0_L8}), .b ({new_AGEMA_signal_6993, SubBytesIns_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_7184, SubBytesIns_Inst_Sbox_0_L27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L28_U1 ( .a ({new_AGEMA_signal_6994, SubBytesIns_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_6799, SubBytesIns_Inst_Sbox_0_L14}), .c ({new_AGEMA_signal_7185, SubBytesIns_Inst_Sbox_0_L28}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L29_U1 ( .a ({new_AGEMA_signal_6994, SubBytesIns_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_6801, SubBytesIns_Inst_Sbox_0_L17}), .c ({new_AGEMA_signal_7186, SubBytesIns_Inst_Sbox_0_L29}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S0_U1 ( .a ({new_AGEMA_signal_6990, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_7181, SubBytesIns_Inst_Sbox_0_L24}), .c ({new_AGEMA_signal_7385, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S1_U1 ( .a ({new_AGEMA_signal_7178, SubBytesIns_Inst_Sbox_0_L16}), .b ({new_AGEMA_signal_7183, SubBytesIns_Inst_Sbox_0_L26}), .c ({new_AGEMA_signal_7386, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S2_U1 ( .a ({new_AGEMA_signal_6995, SubBytesIns_Inst_Sbox_0_L19}), .b ({new_AGEMA_signal_7185, SubBytesIns_Inst_Sbox_0_L28}), .c ({new_AGEMA_signal_7387, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S3_U1 ( .a ({new_AGEMA_signal_6990, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_7180, SubBytesIns_Inst_Sbox_0_L21}), .c ({new_AGEMA_signal_7388, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S4_U1 ( .a ({new_AGEMA_signal_7179, SubBytesIns_Inst_Sbox_0_L20}), .b ({new_AGEMA_signal_6996, SubBytesIns_Inst_Sbox_0_L22}), .c ({new_AGEMA_signal_7389, MixColumnsInput[99]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S5_U1 ( .a ({new_AGEMA_signal_7182, SubBytesIns_Inst_Sbox_0_L25}), .b ({new_AGEMA_signal_7186, SubBytesIns_Inst_Sbox_0_L29}), .c ({new_AGEMA_signal_7390, MixColumnsInput[98]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S6_U1 ( .a ({new_AGEMA_signal_7177, SubBytesIns_Inst_Sbox_0_L13}), .b ({new_AGEMA_signal_7184, SubBytesIns_Inst_Sbox_0_L27}), .c ({new_AGEMA_signal_7391, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S7_U1 ( .a ({new_AGEMA_signal_6990, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_6997, SubBytesIns_Inst_Sbox_0_L23}), .c ({new_AGEMA_signal_7187, MixColumnsInput[96]}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M46_U1 ( .a ({new_AGEMA_signal_6336, SubBytesIns_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_11710, new_AGEMA_signal_11707}), .clk (clk), .r ({Fresh[677], Fresh[676]}), .c ({new_AGEMA_signal_6574, SubBytesIns_Inst_Sbox_1_M46}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M47_U1 ( .a ({new_AGEMA_signal_6216, SubBytesIns_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_11716, new_AGEMA_signal_11713}), .clk (clk), .r ({Fresh[679], Fresh[678]}), .c ({new_AGEMA_signal_6337, SubBytesIns_Inst_Sbox_1_M47}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M48_U1 ( .a ({new_AGEMA_signal_6215, SubBytesIns_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_11722, new_AGEMA_signal_11719}), .clk (clk), .r ({Fresh[681], Fresh[680]}), .c ({new_AGEMA_signal_6338, SubBytesIns_Inst_Sbox_1_M48}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M49_U1 ( .a ({new_AGEMA_signal_6335, SubBytesIns_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_11728, new_AGEMA_signal_11725}), .clk (clk), .r ({Fresh[683], Fresh[682]}), .c ({new_AGEMA_signal_6575, SubBytesIns_Inst_Sbox_1_M49}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M50_U1 ( .a ({new_AGEMA_signal_6214, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_11734, new_AGEMA_signal_11731}), .clk (clk), .r ({Fresh[685], Fresh[684]}), .c ({new_AGEMA_signal_6339, SubBytesIns_Inst_Sbox_1_M50}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M51_U1 ( .a ({new_AGEMA_signal_6213, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_11740, new_AGEMA_signal_11737}), .clk (clk), .r ({Fresh[687], Fresh[686]}), .c ({new_AGEMA_signal_6340, SubBytesIns_Inst_Sbox_1_M51}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M52_U1 ( .a ({new_AGEMA_signal_6334, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_11746, new_AGEMA_signal_11743}), .clk (clk), .r ({Fresh[689], Fresh[688]}), .c ({new_AGEMA_signal_6576, SubBytesIns_Inst_Sbox_1_M52}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M53_U1 ( .a ({new_AGEMA_signal_6573, SubBytesIns_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_11752, new_AGEMA_signal_11749}), .clk (clk), .r ({Fresh[691], Fresh[690]}), .c ({new_AGEMA_signal_6803, SubBytesIns_Inst_Sbox_1_M53}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M54_U1 ( .a ({new_AGEMA_signal_6333, SubBytesIns_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_11758, new_AGEMA_signal_11755}), .clk (clk), .r ({Fresh[693], Fresh[692]}), .c ({new_AGEMA_signal_6577, SubBytesIns_Inst_Sbox_1_M54}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M55_U1 ( .a ({new_AGEMA_signal_6336, SubBytesIns_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_11764, new_AGEMA_signal_11761}), .clk (clk), .r ({Fresh[695], Fresh[694]}), .c ({new_AGEMA_signal_6578, SubBytesIns_Inst_Sbox_1_M55}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M56_U1 ( .a ({new_AGEMA_signal_6216, SubBytesIns_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_11770, new_AGEMA_signal_11767}), .clk (clk), .r ({Fresh[697], Fresh[696]}), .c ({new_AGEMA_signal_6341, SubBytesIns_Inst_Sbox_1_M56}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M57_U1 ( .a ({new_AGEMA_signal_6215, SubBytesIns_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_11776, new_AGEMA_signal_11773}), .clk (clk), .r ({Fresh[699], Fresh[698]}), .c ({new_AGEMA_signal_6342, SubBytesIns_Inst_Sbox_1_M57}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M58_U1 ( .a ({new_AGEMA_signal_6335, SubBytesIns_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_11782, new_AGEMA_signal_11779}), .clk (clk), .r ({Fresh[701], Fresh[700]}), .c ({new_AGEMA_signal_6579, SubBytesIns_Inst_Sbox_1_M58}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M59_U1 ( .a ({new_AGEMA_signal_6214, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_11788, new_AGEMA_signal_11785}), .clk (clk), .r ({Fresh[703], Fresh[702]}), .c ({new_AGEMA_signal_6343, SubBytesIns_Inst_Sbox_1_M59}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M60_U1 ( .a ({new_AGEMA_signal_6213, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_11794, new_AGEMA_signal_11791}), .clk (clk), .r ({Fresh[705], Fresh[704]}), .c ({new_AGEMA_signal_6344, SubBytesIns_Inst_Sbox_1_M60}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M61_U1 ( .a ({new_AGEMA_signal_6334, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_11800, new_AGEMA_signal_11797}), .clk (clk), .r ({Fresh[707], Fresh[706]}), .c ({new_AGEMA_signal_6580, SubBytesIns_Inst_Sbox_1_M61}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M62_U1 ( .a ({new_AGEMA_signal_6573, SubBytesIns_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_11806, new_AGEMA_signal_11803}), .clk (clk), .r ({Fresh[709], Fresh[708]}), .c ({new_AGEMA_signal_6804, SubBytesIns_Inst_Sbox_1_M62}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M63_U1 ( .a ({new_AGEMA_signal_6333, SubBytesIns_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_11812, new_AGEMA_signal_11809}), .clk (clk), .r ({Fresh[711], Fresh[710]}), .c ({new_AGEMA_signal_6581, SubBytesIns_Inst_Sbox_1_M63}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L0_U1 ( .a ({new_AGEMA_signal_6580, SubBytesIns_Inst_Sbox_1_M61}), .b ({new_AGEMA_signal_6804, SubBytesIns_Inst_Sbox_1_M62}), .c ({new_AGEMA_signal_6998, SubBytesIns_Inst_Sbox_1_L0}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L1_U1 ( .a ({new_AGEMA_signal_6339, SubBytesIns_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_6341, SubBytesIns_Inst_Sbox_1_M56}), .c ({new_AGEMA_signal_6582, SubBytesIns_Inst_Sbox_1_L1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L2_U1 ( .a ({new_AGEMA_signal_6574, SubBytesIns_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_6338, SubBytesIns_Inst_Sbox_1_M48}), .c ({new_AGEMA_signal_6805, SubBytesIns_Inst_Sbox_1_L2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L3_U1 ( .a ({new_AGEMA_signal_6337, SubBytesIns_Inst_Sbox_1_M47}), .b ({new_AGEMA_signal_6578, SubBytesIns_Inst_Sbox_1_M55}), .c ({new_AGEMA_signal_6806, SubBytesIns_Inst_Sbox_1_L3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L4_U1 ( .a ({new_AGEMA_signal_6577, SubBytesIns_Inst_Sbox_1_M54}), .b ({new_AGEMA_signal_6579, SubBytesIns_Inst_Sbox_1_M58}), .c ({new_AGEMA_signal_6807, SubBytesIns_Inst_Sbox_1_L4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L5_U1 ( .a ({new_AGEMA_signal_6575, SubBytesIns_Inst_Sbox_1_M49}), .b ({new_AGEMA_signal_6580, SubBytesIns_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_6808, SubBytesIns_Inst_Sbox_1_L5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L6_U1 ( .a ({new_AGEMA_signal_6804, SubBytesIns_Inst_Sbox_1_M62}), .b ({new_AGEMA_signal_6808, SubBytesIns_Inst_Sbox_1_L5}), .c ({new_AGEMA_signal_6999, SubBytesIns_Inst_Sbox_1_L6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L7_U1 ( .a ({new_AGEMA_signal_6574, SubBytesIns_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_6806, SubBytesIns_Inst_Sbox_1_L3}), .c ({new_AGEMA_signal_7000, SubBytesIns_Inst_Sbox_1_L7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L8_U1 ( .a ({new_AGEMA_signal_6340, SubBytesIns_Inst_Sbox_1_M51}), .b ({new_AGEMA_signal_6343, SubBytesIns_Inst_Sbox_1_M59}), .c ({new_AGEMA_signal_6583, SubBytesIns_Inst_Sbox_1_L8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L9_U1 ( .a ({new_AGEMA_signal_6576, SubBytesIns_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_6803, SubBytesIns_Inst_Sbox_1_M53}), .c ({new_AGEMA_signal_7001, SubBytesIns_Inst_Sbox_1_L9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L10_U1 ( .a ({new_AGEMA_signal_6803, SubBytesIns_Inst_Sbox_1_M53}), .b ({new_AGEMA_signal_6807, SubBytesIns_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_7002, SubBytesIns_Inst_Sbox_1_L10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L11_U1 ( .a ({new_AGEMA_signal_6344, SubBytesIns_Inst_Sbox_1_M60}), .b ({new_AGEMA_signal_6805, SubBytesIns_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_7003, SubBytesIns_Inst_Sbox_1_L11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L12_U1 ( .a ({new_AGEMA_signal_6338, SubBytesIns_Inst_Sbox_1_M48}), .b ({new_AGEMA_signal_6340, SubBytesIns_Inst_Sbox_1_M51}), .c ({new_AGEMA_signal_6584, SubBytesIns_Inst_Sbox_1_L12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L13_U1 ( .a ({new_AGEMA_signal_6339, SubBytesIns_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_6998, SubBytesIns_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_7188, SubBytesIns_Inst_Sbox_1_L13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L14_U1 ( .a ({new_AGEMA_signal_6576, SubBytesIns_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_6580, SubBytesIns_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_6809, SubBytesIns_Inst_Sbox_1_L14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L15_U1 ( .a ({new_AGEMA_signal_6578, SubBytesIns_Inst_Sbox_1_M55}), .b ({new_AGEMA_signal_6582, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_6810, SubBytesIns_Inst_Sbox_1_L15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L16_U1 ( .a ({new_AGEMA_signal_6341, SubBytesIns_Inst_Sbox_1_M56}), .b ({new_AGEMA_signal_6998, SubBytesIns_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_7189, SubBytesIns_Inst_Sbox_1_L16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L17_U1 ( .a ({new_AGEMA_signal_6342, SubBytesIns_Inst_Sbox_1_M57}), .b ({new_AGEMA_signal_6582, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_6811, SubBytesIns_Inst_Sbox_1_L17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L18_U1 ( .a ({new_AGEMA_signal_6579, SubBytesIns_Inst_Sbox_1_M58}), .b ({new_AGEMA_signal_6583, SubBytesIns_Inst_Sbox_1_L8}), .c ({new_AGEMA_signal_6812, SubBytesIns_Inst_Sbox_1_L18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L19_U1 ( .a ({new_AGEMA_signal_6581, SubBytesIns_Inst_Sbox_1_M63}), .b ({new_AGEMA_signal_6807, SubBytesIns_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_7004, SubBytesIns_Inst_Sbox_1_L19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L20_U1 ( .a ({new_AGEMA_signal_6998, SubBytesIns_Inst_Sbox_1_L0}), .b ({new_AGEMA_signal_6582, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_7190, SubBytesIns_Inst_Sbox_1_L20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L21_U1 ( .a ({new_AGEMA_signal_6582, SubBytesIns_Inst_Sbox_1_L1}), .b ({new_AGEMA_signal_7000, SubBytesIns_Inst_Sbox_1_L7}), .c ({new_AGEMA_signal_7191, SubBytesIns_Inst_Sbox_1_L21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L22_U1 ( .a ({new_AGEMA_signal_6806, SubBytesIns_Inst_Sbox_1_L3}), .b ({new_AGEMA_signal_6584, SubBytesIns_Inst_Sbox_1_L12}), .c ({new_AGEMA_signal_7005, SubBytesIns_Inst_Sbox_1_L22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L23_U1 ( .a ({new_AGEMA_signal_6812, SubBytesIns_Inst_Sbox_1_L18}), .b ({new_AGEMA_signal_6805, SubBytesIns_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_7006, SubBytesIns_Inst_Sbox_1_L23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L24_U1 ( .a ({new_AGEMA_signal_6810, SubBytesIns_Inst_Sbox_1_L15}), .b ({new_AGEMA_signal_7001, SubBytesIns_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_7192, SubBytesIns_Inst_Sbox_1_L24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L25_U1 ( .a ({new_AGEMA_signal_6999, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_7002, SubBytesIns_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_7193, SubBytesIns_Inst_Sbox_1_L25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L26_U1 ( .a ({new_AGEMA_signal_7000, SubBytesIns_Inst_Sbox_1_L7}), .b ({new_AGEMA_signal_7001, SubBytesIns_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_7194, SubBytesIns_Inst_Sbox_1_L26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L27_U1 ( .a ({new_AGEMA_signal_6583, SubBytesIns_Inst_Sbox_1_L8}), .b ({new_AGEMA_signal_7002, SubBytesIns_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_7195, SubBytesIns_Inst_Sbox_1_L27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L28_U1 ( .a ({new_AGEMA_signal_7003, SubBytesIns_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_6809, SubBytesIns_Inst_Sbox_1_L14}), .c ({new_AGEMA_signal_7196, SubBytesIns_Inst_Sbox_1_L28}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L29_U1 ( .a ({new_AGEMA_signal_7003, SubBytesIns_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_6811, SubBytesIns_Inst_Sbox_1_L17}), .c ({new_AGEMA_signal_7197, SubBytesIns_Inst_Sbox_1_L29}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S0_U1 ( .a ({new_AGEMA_signal_6999, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_7192, SubBytesIns_Inst_Sbox_1_L24}), .c ({new_AGEMA_signal_7392, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S1_U1 ( .a ({new_AGEMA_signal_7189, SubBytesIns_Inst_Sbox_1_L16}), .b ({new_AGEMA_signal_7194, SubBytesIns_Inst_Sbox_1_L26}), .c ({new_AGEMA_signal_7393, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S2_U1 ( .a ({new_AGEMA_signal_7004, SubBytesIns_Inst_Sbox_1_L19}), .b ({new_AGEMA_signal_7196, SubBytesIns_Inst_Sbox_1_L28}), .c ({new_AGEMA_signal_7394, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S3_U1 ( .a ({new_AGEMA_signal_6999, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_7191, SubBytesIns_Inst_Sbox_1_L21}), .c ({new_AGEMA_signal_7395, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S4_U1 ( .a ({new_AGEMA_signal_7190, SubBytesIns_Inst_Sbox_1_L20}), .b ({new_AGEMA_signal_7005, SubBytesIns_Inst_Sbox_1_L22}), .c ({new_AGEMA_signal_7396, MixColumnsInput[75]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S5_U1 ( .a ({new_AGEMA_signal_7193, SubBytesIns_Inst_Sbox_1_L25}), .b ({new_AGEMA_signal_7197, SubBytesIns_Inst_Sbox_1_L29}), .c ({new_AGEMA_signal_7397, MixColumnsInput[74]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S6_U1 ( .a ({new_AGEMA_signal_7188, SubBytesIns_Inst_Sbox_1_L13}), .b ({new_AGEMA_signal_7195, SubBytesIns_Inst_Sbox_1_L27}), .c ({new_AGEMA_signal_7398, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S7_U1 ( .a ({new_AGEMA_signal_6999, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_7006, SubBytesIns_Inst_Sbox_1_L23}), .c ({new_AGEMA_signal_7198, MixColumnsInput[72]}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M46_U1 ( .a ({new_AGEMA_signal_6348, SubBytesIns_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_11818, new_AGEMA_signal_11815}), .clk (clk), .r ({Fresh[713], Fresh[712]}), .c ({new_AGEMA_signal_6586, SubBytesIns_Inst_Sbox_2_M46}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M47_U1 ( .a ({new_AGEMA_signal_6220, SubBytesIns_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_11824, new_AGEMA_signal_11821}), .clk (clk), .r ({Fresh[715], Fresh[714]}), .c ({new_AGEMA_signal_6349, SubBytesIns_Inst_Sbox_2_M47}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M48_U1 ( .a ({new_AGEMA_signal_6219, SubBytesIns_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_11830, new_AGEMA_signal_11827}), .clk (clk), .r ({Fresh[717], Fresh[716]}), .c ({new_AGEMA_signal_6350, SubBytesIns_Inst_Sbox_2_M48}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M49_U1 ( .a ({new_AGEMA_signal_6347, SubBytesIns_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_11836, new_AGEMA_signal_11833}), .clk (clk), .r ({Fresh[719], Fresh[718]}), .c ({new_AGEMA_signal_6587, SubBytesIns_Inst_Sbox_2_M49}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M50_U1 ( .a ({new_AGEMA_signal_6218, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_11842, new_AGEMA_signal_11839}), .clk (clk), .r ({Fresh[721], Fresh[720]}), .c ({new_AGEMA_signal_6351, SubBytesIns_Inst_Sbox_2_M50}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M51_U1 ( .a ({new_AGEMA_signal_6217, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_11848, new_AGEMA_signal_11845}), .clk (clk), .r ({Fresh[723], Fresh[722]}), .c ({new_AGEMA_signal_6352, SubBytesIns_Inst_Sbox_2_M51}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M52_U1 ( .a ({new_AGEMA_signal_6346, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_11854, new_AGEMA_signal_11851}), .clk (clk), .r ({Fresh[725], Fresh[724]}), .c ({new_AGEMA_signal_6588, SubBytesIns_Inst_Sbox_2_M52}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M53_U1 ( .a ({new_AGEMA_signal_6585, SubBytesIns_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_11860, new_AGEMA_signal_11857}), .clk (clk), .r ({Fresh[727], Fresh[726]}), .c ({new_AGEMA_signal_6813, SubBytesIns_Inst_Sbox_2_M53}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M54_U1 ( .a ({new_AGEMA_signal_6345, SubBytesIns_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_11866, new_AGEMA_signal_11863}), .clk (clk), .r ({Fresh[729], Fresh[728]}), .c ({new_AGEMA_signal_6589, SubBytesIns_Inst_Sbox_2_M54}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M55_U1 ( .a ({new_AGEMA_signal_6348, SubBytesIns_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_11872, new_AGEMA_signal_11869}), .clk (clk), .r ({Fresh[731], Fresh[730]}), .c ({new_AGEMA_signal_6590, SubBytesIns_Inst_Sbox_2_M55}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M56_U1 ( .a ({new_AGEMA_signal_6220, SubBytesIns_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_11878, new_AGEMA_signal_11875}), .clk (clk), .r ({Fresh[733], Fresh[732]}), .c ({new_AGEMA_signal_6353, SubBytesIns_Inst_Sbox_2_M56}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M57_U1 ( .a ({new_AGEMA_signal_6219, SubBytesIns_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_11884, new_AGEMA_signal_11881}), .clk (clk), .r ({Fresh[735], Fresh[734]}), .c ({new_AGEMA_signal_6354, SubBytesIns_Inst_Sbox_2_M57}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M58_U1 ( .a ({new_AGEMA_signal_6347, SubBytesIns_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_11890, new_AGEMA_signal_11887}), .clk (clk), .r ({Fresh[737], Fresh[736]}), .c ({new_AGEMA_signal_6591, SubBytesIns_Inst_Sbox_2_M58}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M59_U1 ( .a ({new_AGEMA_signal_6218, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_11896, new_AGEMA_signal_11893}), .clk (clk), .r ({Fresh[739], Fresh[738]}), .c ({new_AGEMA_signal_6355, SubBytesIns_Inst_Sbox_2_M59}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M60_U1 ( .a ({new_AGEMA_signal_6217, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_11902, new_AGEMA_signal_11899}), .clk (clk), .r ({Fresh[741], Fresh[740]}), .c ({new_AGEMA_signal_6356, SubBytesIns_Inst_Sbox_2_M60}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M61_U1 ( .a ({new_AGEMA_signal_6346, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_11908, new_AGEMA_signal_11905}), .clk (clk), .r ({Fresh[743], Fresh[742]}), .c ({new_AGEMA_signal_6592, SubBytesIns_Inst_Sbox_2_M61}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M62_U1 ( .a ({new_AGEMA_signal_6585, SubBytesIns_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_11914, new_AGEMA_signal_11911}), .clk (clk), .r ({Fresh[745], Fresh[744]}), .c ({new_AGEMA_signal_6814, SubBytesIns_Inst_Sbox_2_M62}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M63_U1 ( .a ({new_AGEMA_signal_6345, SubBytesIns_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_11920, new_AGEMA_signal_11917}), .clk (clk), .r ({Fresh[747], Fresh[746]}), .c ({new_AGEMA_signal_6593, SubBytesIns_Inst_Sbox_2_M63}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L0_U1 ( .a ({new_AGEMA_signal_6592, SubBytesIns_Inst_Sbox_2_M61}), .b ({new_AGEMA_signal_6814, SubBytesIns_Inst_Sbox_2_M62}), .c ({new_AGEMA_signal_7007, SubBytesIns_Inst_Sbox_2_L0}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L1_U1 ( .a ({new_AGEMA_signal_6351, SubBytesIns_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_6353, SubBytesIns_Inst_Sbox_2_M56}), .c ({new_AGEMA_signal_6594, SubBytesIns_Inst_Sbox_2_L1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L2_U1 ( .a ({new_AGEMA_signal_6586, SubBytesIns_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_6350, SubBytesIns_Inst_Sbox_2_M48}), .c ({new_AGEMA_signal_6815, SubBytesIns_Inst_Sbox_2_L2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L3_U1 ( .a ({new_AGEMA_signal_6349, SubBytesIns_Inst_Sbox_2_M47}), .b ({new_AGEMA_signal_6590, SubBytesIns_Inst_Sbox_2_M55}), .c ({new_AGEMA_signal_6816, SubBytesIns_Inst_Sbox_2_L3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L4_U1 ( .a ({new_AGEMA_signal_6589, SubBytesIns_Inst_Sbox_2_M54}), .b ({new_AGEMA_signal_6591, SubBytesIns_Inst_Sbox_2_M58}), .c ({new_AGEMA_signal_6817, SubBytesIns_Inst_Sbox_2_L4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L5_U1 ( .a ({new_AGEMA_signal_6587, SubBytesIns_Inst_Sbox_2_M49}), .b ({new_AGEMA_signal_6592, SubBytesIns_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_6818, SubBytesIns_Inst_Sbox_2_L5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L6_U1 ( .a ({new_AGEMA_signal_6814, SubBytesIns_Inst_Sbox_2_M62}), .b ({new_AGEMA_signal_6818, SubBytesIns_Inst_Sbox_2_L5}), .c ({new_AGEMA_signal_7008, SubBytesIns_Inst_Sbox_2_L6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L7_U1 ( .a ({new_AGEMA_signal_6586, SubBytesIns_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_6816, SubBytesIns_Inst_Sbox_2_L3}), .c ({new_AGEMA_signal_7009, SubBytesIns_Inst_Sbox_2_L7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L8_U1 ( .a ({new_AGEMA_signal_6352, SubBytesIns_Inst_Sbox_2_M51}), .b ({new_AGEMA_signal_6355, SubBytesIns_Inst_Sbox_2_M59}), .c ({new_AGEMA_signal_6595, SubBytesIns_Inst_Sbox_2_L8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L9_U1 ( .a ({new_AGEMA_signal_6588, SubBytesIns_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_6813, SubBytesIns_Inst_Sbox_2_M53}), .c ({new_AGEMA_signal_7010, SubBytesIns_Inst_Sbox_2_L9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L10_U1 ( .a ({new_AGEMA_signal_6813, SubBytesIns_Inst_Sbox_2_M53}), .b ({new_AGEMA_signal_6817, SubBytesIns_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_7011, SubBytesIns_Inst_Sbox_2_L10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L11_U1 ( .a ({new_AGEMA_signal_6356, SubBytesIns_Inst_Sbox_2_M60}), .b ({new_AGEMA_signal_6815, SubBytesIns_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_7012, SubBytesIns_Inst_Sbox_2_L11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L12_U1 ( .a ({new_AGEMA_signal_6350, SubBytesIns_Inst_Sbox_2_M48}), .b ({new_AGEMA_signal_6352, SubBytesIns_Inst_Sbox_2_M51}), .c ({new_AGEMA_signal_6596, SubBytesIns_Inst_Sbox_2_L12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L13_U1 ( .a ({new_AGEMA_signal_6351, SubBytesIns_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_7007, SubBytesIns_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_7199, SubBytesIns_Inst_Sbox_2_L13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L14_U1 ( .a ({new_AGEMA_signal_6588, SubBytesIns_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_6592, SubBytesIns_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_6819, SubBytesIns_Inst_Sbox_2_L14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L15_U1 ( .a ({new_AGEMA_signal_6590, SubBytesIns_Inst_Sbox_2_M55}), .b ({new_AGEMA_signal_6594, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_6820, SubBytesIns_Inst_Sbox_2_L15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L16_U1 ( .a ({new_AGEMA_signal_6353, SubBytesIns_Inst_Sbox_2_M56}), .b ({new_AGEMA_signal_7007, SubBytesIns_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_7200, SubBytesIns_Inst_Sbox_2_L16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L17_U1 ( .a ({new_AGEMA_signal_6354, SubBytesIns_Inst_Sbox_2_M57}), .b ({new_AGEMA_signal_6594, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_6821, SubBytesIns_Inst_Sbox_2_L17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L18_U1 ( .a ({new_AGEMA_signal_6591, SubBytesIns_Inst_Sbox_2_M58}), .b ({new_AGEMA_signal_6595, SubBytesIns_Inst_Sbox_2_L8}), .c ({new_AGEMA_signal_6822, SubBytesIns_Inst_Sbox_2_L18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L19_U1 ( .a ({new_AGEMA_signal_6593, SubBytesIns_Inst_Sbox_2_M63}), .b ({new_AGEMA_signal_6817, SubBytesIns_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_7013, SubBytesIns_Inst_Sbox_2_L19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L20_U1 ( .a ({new_AGEMA_signal_7007, SubBytesIns_Inst_Sbox_2_L0}), .b ({new_AGEMA_signal_6594, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_7201, SubBytesIns_Inst_Sbox_2_L20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L21_U1 ( .a ({new_AGEMA_signal_6594, SubBytesIns_Inst_Sbox_2_L1}), .b ({new_AGEMA_signal_7009, SubBytesIns_Inst_Sbox_2_L7}), .c ({new_AGEMA_signal_7202, SubBytesIns_Inst_Sbox_2_L21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L22_U1 ( .a ({new_AGEMA_signal_6816, SubBytesIns_Inst_Sbox_2_L3}), .b ({new_AGEMA_signal_6596, SubBytesIns_Inst_Sbox_2_L12}), .c ({new_AGEMA_signal_7014, SubBytesIns_Inst_Sbox_2_L22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L23_U1 ( .a ({new_AGEMA_signal_6822, SubBytesIns_Inst_Sbox_2_L18}), .b ({new_AGEMA_signal_6815, SubBytesIns_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_7015, SubBytesIns_Inst_Sbox_2_L23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L24_U1 ( .a ({new_AGEMA_signal_6820, SubBytesIns_Inst_Sbox_2_L15}), .b ({new_AGEMA_signal_7010, SubBytesIns_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_7203, SubBytesIns_Inst_Sbox_2_L24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L25_U1 ( .a ({new_AGEMA_signal_7008, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_7011, SubBytesIns_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_7204, SubBytesIns_Inst_Sbox_2_L25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L26_U1 ( .a ({new_AGEMA_signal_7009, SubBytesIns_Inst_Sbox_2_L7}), .b ({new_AGEMA_signal_7010, SubBytesIns_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_7205, SubBytesIns_Inst_Sbox_2_L26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L27_U1 ( .a ({new_AGEMA_signal_6595, SubBytesIns_Inst_Sbox_2_L8}), .b ({new_AGEMA_signal_7011, SubBytesIns_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_7206, SubBytesIns_Inst_Sbox_2_L27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L28_U1 ( .a ({new_AGEMA_signal_7012, SubBytesIns_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_6819, SubBytesIns_Inst_Sbox_2_L14}), .c ({new_AGEMA_signal_7207, SubBytesIns_Inst_Sbox_2_L28}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L29_U1 ( .a ({new_AGEMA_signal_7012, SubBytesIns_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_6821, SubBytesIns_Inst_Sbox_2_L17}), .c ({new_AGEMA_signal_7208, SubBytesIns_Inst_Sbox_2_L29}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S0_U1 ( .a ({new_AGEMA_signal_7008, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_7203, SubBytesIns_Inst_Sbox_2_L24}), .c ({new_AGEMA_signal_7399, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S1_U1 ( .a ({new_AGEMA_signal_7200, SubBytesIns_Inst_Sbox_2_L16}), .b ({new_AGEMA_signal_7205, SubBytesIns_Inst_Sbox_2_L26}), .c ({new_AGEMA_signal_7400, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S2_U1 ( .a ({new_AGEMA_signal_7013, SubBytesIns_Inst_Sbox_2_L19}), .b ({new_AGEMA_signal_7207, SubBytesIns_Inst_Sbox_2_L28}), .c ({new_AGEMA_signal_7401, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S3_U1 ( .a ({new_AGEMA_signal_7008, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_7202, SubBytesIns_Inst_Sbox_2_L21}), .c ({new_AGEMA_signal_7402, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S4_U1 ( .a ({new_AGEMA_signal_7201, SubBytesIns_Inst_Sbox_2_L20}), .b ({new_AGEMA_signal_7014, SubBytesIns_Inst_Sbox_2_L22}), .c ({new_AGEMA_signal_7403, MixColumnsInput[51]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S5_U1 ( .a ({new_AGEMA_signal_7204, SubBytesIns_Inst_Sbox_2_L25}), .b ({new_AGEMA_signal_7208, SubBytesIns_Inst_Sbox_2_L29}), .c ({new_AGEMA_signal_7404, MixColumnsInput[50]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S6_U1 ( .a ({new_AGEMA_signal_7199, SubBytesIns_Inst_Sbox_2_L13}), .b ({new_AGEMA_signal_7206, SubBytesIns_Inst_Sbox_2_L27}), .c ({new_AGEMA_signal_7405, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S7_U1 ( .a ({new_AGEMA_signal_7008, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_7015, SubBytesIns_Inst_Sbox_2_L23}), .c ({new_AGEMA_signal_7209, MixColumnsInput[48]}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M46_U1 ( .a ({new_AGEMA_signal_6360, SubBytesIns_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_11926, new_AGEMA_signal_11923}), .clk (clk), .r ({Fresh[749], Fresh[748]}), .c ({new_AGEMA_signal_6598, SubBytesIns_Inst_Sbox_3_M46}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M47_U1 ( .a ({new_AGEMA_signal_6224, SubBytesIns_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_11932, new_AGEMA_signal_11929}), .clk (clk), .r ({Fresh[751], Fresh[750]}), .c ({new_AGEMA_signal_6361, SubBytesIns_Inst_Sbox_3_M47}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M48_U1 ( .a ({new_AGEMA_signal_6223, SubBytesIns_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_11938, new_AGEMA_signal_11935}), .clk (clk), .r ({Fresh[753], Fresh[752]}), .c ({new_AGEMA_signal_6362, SubBytesIns_Inst_Sbox_3_M48}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M49_U1 ( .a ({new_AGEMA_signal_6359, SubBytesIns_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_11944, new_AGEMA_signal_11941}), .clk (clk), .r ({Fresh[755], Fresh[754]}), .c ({new_AGEMA_signal_6599, SubBytesIns_Inst_Sbox_3_M49}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M50_U1 ( .a ({new_AGEMA_signal_6222, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_11950, new_AGEMA_signal_11947}), .clk (clk), .r ({Fresh[757], Fresh[756]}), .c ({new_AGEMA_signal_6363, SubBytesIns_Inst_Sbox_3_M50}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M51_U1 ( .a ({new_AGEMA_signal_6221, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_11956, new_AGEMA_signal_11953}), .clk (clk), .r ({Fresh[759], Fresh[758]}), .c ({new_AGEMA_signal_6364, SubBytesIns_Inst_Sbox_3_M51}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M52_U1 ( .a ({new_AGEMA_signal_6358, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_11962, new_AGEMA_signal_11959}), .clk (clk), .r ({Fresh[761], Fresh[760]}), .c ({new_AGEMA_signal_6600, SubBytesIns_Inst_Sbox_3_M52}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M53_U1 ( .a ({new_AGEMA_signal_6597, SubBytesIns_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_11968, new_AGEMA_signal_11965}), .clk (clk), .r ({Fresh[763], Fresh[762]}), .c ({new_AGEMA_signal_6823, SubBytesIns_Inst_Sbox_3_M53}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M54_U1 ( .a ({new_AGEMA_signal_6357, SubBytesIns_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_11974, new_AGEMA_signal_11971}), .clk (clk), .r ({Fresh[765], Fresh[764]}), .c ({new_AGEMA_signal_6601, SubBytesIns_Inst_Sbox_3_M54}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M55_U1 ( .a ({new_AGEMA_signal_6360, SubBytesIns_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_11980, new_AGEMA_signal_11977}), .clk (clk), .r ({Fresh[767], Fresh[766]}), .c ({new_AGEMA_signal_6602, SubBytesIns_Inst_Sbox_3_M55}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M56_U1 ( .a ({new_AGEMA_signal_6224, SubBytesIns_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_11986, new_AGEMA_signal_11983}), .clk (clk), .r ({Fresh[769], Fresh[768]}), .c ({new_AGEMA_signal_6365, SubBytesIns_Inst_Sbox_3_M56}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M57_U1 ( .a ({new_AGEMA_signal_6223, SubBytesIns_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_11992, new_AGEMA_signal_11989}), .clk (clk), .r ({Fresh[771], Fresh[770]}), .c ({new_AGEMA_signal_6366, SubBytesIns_Inst_Sbox_3_M57}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M58_U1 ( .a ({new_AGEMA_signal_6359, SubBytesIns_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_11998, new_AGEMA_signal_11995}), .clk (clk), .r ({Fresh[773], Fresh[772]}), .c ({new_AGEMA_signal_6603, SubBytesIns_Inst_Sbox_3_M58}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M59_U1 ( .a ({new_AGEMA_signal_6222, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_12004, new_AGEMA_signal_12001}), .clk (clk), .r ({Fresh[775], Fresh[774]}), .c ({new_AGEMA_signal_6367, SubBytesIns_Inst_Sbox_3_M59}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M60_U1 ( .a ({new_AGEMA_signal_6221, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_12010, new_AGEMA_signal_12007}), .clk (clk), .r ({Fresh[777], Fresh[776]}), .c ({new_AGEMA_signal_6368, SubBytesIns_Inst_Sbox_3_M60}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M61_U1 ( .a ({new_AGEMA_signal_6358, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_12016, new_AGEMA_signal_12013}), .clk (clk), .r ({Fresh[779], Fresh[778]}), .c ({new_AGEMA_signal_6604, SubBytesIns_Inst_Sbox_3_M61}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M62_U1 ( .a ({new_AGEMA_signal_6597, SubBytesIns_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_12022, new_AGEMA_signal_12019}), .clk (clk), .r ({Fresh[781], Fresh[780]}), .c ({new_AGEMA_signal_6824, SubBytesIns_Inst_Sbox_3_M62}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M63_U1 ( .a ({new_AGEMA_signal_6357, SubBytesIns_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_12028, new_AGEMA_signal_12025}), .clk (clk), .r ({Fresh[783], Fresh[782]}), .c ({new_AGEMA_signal_6605, SubBytesIns_Inst_Sbox_3_M63}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L0_U1 ( .a ({new_AGEMA_signal_6604, SubBytesIns_Inst_Sbox_3_M61}), .b ({new_AGEMA_signal_6824, SubBytesIns_Inst_Sbox_3_M62}), .c ({new_AGEMA_signal_7016, SubBytesIns_Inst_Sbox_3_L0}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L1_U1 ( .a ({new_AGEMA_signal_6363, SubBytesIns_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_6365, SubBytesIns_Inst_Sbox_3_M56}), .c ({new_AGEMA_signal_6606, SubBytesIns_Inst_Sbox_3_L1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L2_U1 ( .a ({new_AGEMA_signal_6598, SubBytesIns_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_6362, SubBytesIns_Inst_Sbox_3_M48}), .c ({new_AGEMA_signal_6825, SubBytesIns_Inst_Sbox_3_L2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L3_U1 ( .a ({new_AGEMA_signal_6361, SubBytesIns_Inst_Sbox_3_M47}), .b ({new_AGEMA_signal_6602, SubBytesIns_Inst_Sbox_3_M55}), .c ({new_AGEMA_signal_6826, SubBytesIns_Inst_Sbox_3_L3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L4_U1 ( .a ({new_AGEMA_signal_6601, SubBytesIns_Inst_Sbox_3_M54}), .b ({new_AGEMA_signal_6603, SubBytesIns_Inst_Sbox_3_M58}), .c ({new_AGEMA_signal_6827, SubBytesIns_Inst_Sbox_3_L4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L5_U1 ( .a ({new_AGEMA_signal_6599, SubBytesIns_Inst_Sbox_3_M49}), .b ({new_AGEMA_signal_6604, SubBytesIns_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_6828, SubBytesIns_Inst_Sbox_3_L5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L6_U1 ( .a ({new_AGEMA_signal_6824, SubBytesIns_Inst_Sbox_3_M62}), .b ({new_AGEMA_signal_6828, SubBytesIns_Inst_Sbox_3_L5}), .c ({new_AGEMA_signal_7017, SubBytesIns_Inst_Sbox_3_L6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L7_U1 ( .a ({new_AGEMA_signal_6598, SubBytesIns_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_6826, SubBytesIns_Inst_Sbox_3_L3}), .c ({new_AGEMA_signal_7018, SubBytesIns_Inst_Sbox_3_L7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L8_U1 ( .a ({new_AGEMA_signal_6364, SubBytesIns_Inst_Sbox_3_M51}), .b ({new_AGEMA_signal_6367, SubBytesIns_Inst_Sbox_3_M59}), .c ({new_AGEMA_signal_6607, SubBytesIns_Inst_Sbox_3_L8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L9_U1 ( .a ({new_AGEMA_signal_6600, SubBytesIns_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_6823, SubBytesIns_Inst_Sbox_3_M53}), .c ({new_AGEMA_signal_7019, SubBytesIns_Inst_Sbox_3_L9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L10_U1 ( .a ({new_AGEMA_signal_6823, SubBytesIns_Inst_Sbox_3_M53}), .b ({new_AGEMA_signal_6827, SubBytesIns_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_7020, SubBytesIns_Inst_Sbox_3_L10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L11_U1 ( .a ({new_AGEMA_signal_6368, SubBytesIns_Inst_Sbox_3_M60}), .b ({new_AGEMA_signal_6825, SubBytesIns_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_7021, SubBytesIns_Inst_Sbox_3_L11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L12_U1 ( .a ({new_AGEMA_signal_6362, SubBytesIns_Inst_Sbox_3_M48}), .b ({new_AGEMA_signal_6364, SubBytesIns_Inst_Sbox_3_M51}), .c ({new_AGEMA_signal_6608, SubBytesIns_Inst_Sbox_3_L12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L13_U1 ( .a ({new_AGEMA_signal_6363, SubBytesIns_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_7016, SubBytesIns_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_7210, SubBytesIns_Inst_Sbox_3_L13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L14_U1 ( .a ({new_AGEMA_signal_6600, SubBytesIns_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_6604, SubBytesIns_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_6829, SubBytesIns_Inst_Sbox_3_L14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L15_U1 ( .a ({new_AGEMA_signal_6602, SubBytesIns_Inst_Sbox_3_M55}), .b ({new_AGEMA_signal_6606, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_6830, SubBytesIns_Inst_Sbox_3_L15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L16_U1 ( .a ({new_AGEMA_signal_6365, SubBytesIns_Inst_Sbox_3_M56}), .b ({new_AGEMA_signal_7016, SubBytesIns_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_7211, SubBytesIns_Inst_Sbox_3_L16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L17_U1 ( .a ({new_AGEMA_signal_6366, SubBytesIns_Inst_Sbox_3_M57}), .b ({new_AGEMA_signal_6606, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_6831, SubBytesIns_Inst_Sbox_3_L17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L18_U1 ( .a ({new_AGEMA_signal_6603, SubBytesIns_Inst_Sbox_3_M58}), .b ({new_AGEMA_signal_6607, SubBytesIns_Inst_Sbox_3_L8}), .c ({new_AGEMA_signal_6832, SubBytesIns_Inst_Sbox_3_L18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L19_U1 ( .a ({new_AGEMA_signal_6605, SubBytesIns_Inst_Sbox_3_M63}), .b ({new_AGEMA_signal_6827, SubBytesIns_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_7022, SubBytesIns_Inst_Sbox_3_L19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L20_U1 ( .a ({new_AGEMA_signal_7016, SubBytesIns_Inst_Sbox_3_L0}), .b ({new_AGEMA_signal_6606, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_7212, SubBytesIns_Inst_Sbox_3_L20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L21_U1 ( .a ({new_AGEMA_signal_6606, SubBytesIns_Inst_Sbox_3_L1}), .b ({new_AGEMA_signal_7018, SubBytesIns_Inst_Sbox_3_L7}), .c ({new_AGEMA_signal_7213, SubBytesIns_Inst_Sbox_3_L21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L22_U1 ( .a ({new_AGEMA_signal_6826, SubBytesIns_Inst_Sbox_3_L3}), .b ({new_AGEMA_signal_6608, SubBytesIns_Inst_Sbox_3_L12}), .c ({new_AGEMA_signal_7023, SubBytesIns_Inst_Sbox_3_L22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L23_U1 ( .a ({new_AGEMA_signal_6832, SubBytesIns_Inst_Sbox_3_L18}), .b ({new_AGEMA_signal_6825, SubBytesIns_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_7024, SubBytesIns_Inst_Sbox_3_L23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L24_U1 ( .a ({new_AGEMA_signal_6830, SubBytesIns_Inst_Sbox_3_L15}), .b ({new_AGEMA_signal_7019, SubBytesIns_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_7214, SubBytesIns_Inst_Sbox_3_L24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L25_U1 ( .a ({new_AGEMA_signal_7017, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_7020, SubBytesIns_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_7215, SubBytesIns_Inst_Sbox_3_L25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L26_U1 ( .a ({new_AGEMA_signal_7018, SubBytesIns_Inst_Sbox_3_L7}), .b ({new_AGEMA_signal_7019, SubBytesIns_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_7216, SubBytesIns_Inst_Sbox_3_L26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L27_U1 ( .a ({new_AGEMA_signal_6607, SubBytesIns_Inst_Sbox_3_L8}), .b ({new_AGEMA_signal_7020, SubBytesIns_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_7217, SubBytesIns_Inst_Sbox_3_L27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L28_U1 ( .a ({new_AGEMA_signal_7021, SubBytesIns_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_6829, SubBytesIns_Inst_Sbox_3_L14}), .c ({new_AGEMA_signal_7218, SubBytesIns_Inst_Sbox_3_L28}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L29_U1 ( .a ({new_AGEMA_signal_7021, SubBytesIns_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_6831, SubBytesIns_Inst_Sbox_3_L17}), .c ({new_AGEMA_signal_7219, SubBytesIns_Inst_Sbox_3_L29}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S0_U1 ( .a ({new_AGEMA_signal_7017, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_7214, SubBytesIns_Inst_Sbox_3_L24}), .c ({new_AGEMA_signal_7406, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S1_U1 ( .a ({new_AGEMA_signal_7211, SubBytesIns_Inst_Sbox_3_L16}), .b ({new_AGEMA_signal_7216, SubBytesIns_Inst_Sbox_3_L26}), .c ({new_AGEMA_signal_7407, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S2_U1 ( .a ({new_AGEMA_signal_7022, SubBytesIns_Inst_Sbox_3_L19}), .b ({new_AGEMA_signal_7218, SubBytesIns_Inst_Sbox_3_L28}), .c ({new_AGEMA_signal_7408, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S3_U1 ( .a ({new_AGEMA_signal_7017, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_7213, SubBytesIns_Inst_Sbox_3_L21}), .c ({new_AGEMA_signal_7409, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S4_U1 ( .a ({new_AGEMA_signal_7212, SubBytesIns_Inst_Sbox_3_L20}), .b ({new_AGEMA_signal_7023, SubBytesIns_Inst_Sbox_3_L22}), .c ({new_AGEMA_signal_7410, MixColumnsInput[27]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S5_U1 ( .a ({new_AGEMA_signal_7215, SubBytesIns_Inst_Sbox_3_L25}), .b ({new_AGEMA_signal_7219, SubBytesIns_Inst_Sbox_3_L29}), .c ({new_AGEMA_signal_7411, MixColumnsInput[26]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S6_U1 ( .a ({new_AGEMA_signal_7210, SubBytesIns_Inst_Sbox_3_L13}), .b ({new_AGEMA_signal_7217, SubBytesIns_Inst_Sbox_3_L27}), .c ({new_AGEMA_signal_7412, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S7_U1 ( .a ({new_AGEMA_signal_7017, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_7024, SubBytesIns_Inst_Sbox_3_L23}), .c ({new_AGEMA_signal_7220, MixColumnsInput[24]}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M46_U1 ( .a ({new_AGEMA_signal_6372, SubBytesIns_Inst_Sbox_4_M44}), .b ({new_AGEMA_signal_12034, new_AGEMA_signal_12031}), .clk (clk), .r ({Fresh[785], Fresh[784]}), .c ({new_AGEMA_signal_6610, SubBytesIns_Inst_Sbox_4_M46}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M47_U1 ( .a ({new_AGEMA_signal_6228, SubBytesIns_Inst_Sbox_4_M40}), .b ({new_AGEMA_signal_12040, new_AGEMA_signal_12037}), .clk (clk), .r ({Fresh[787], Fresh[786]}), .c ({new_AGEMA_signal_6373, SubBytesIns_Inst_Sbox_4_M47}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M48_U1 ( .a ({new_AGEMA_signal_6227, SubBytesIns_Inst_Sbox_4_M39}), .b ({new_AGEMA_signal_12046, new_AGEMA_signal_12043}), .clk (clk), .r ({Fresh[789], Fresh[788]}), .c ({new_AGEMA_signal_6374, SubBytesIns_Inst_Sbox_4_M48}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M49_U1 ( .a ({new_AGEMA_signal_6371, SubBytesIns_Inst_Sbox_4_M43}), .b ({new_AGEMA_signal_12052, new_AGEMA_signal_12049}), .clk (clk), .r ({Fresh[791], Fresh[790]}), .c ({new_AGEMA_signal_6611, SubBytesIns_Inst_Sbox_4_M49}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M50_U1 ( .a ({new_AGEMA_signal_6226, SubBytesIns_Inst_Sbox_4_M38}), .b ({new_AGEMA_signal_12058, new_AGEMA_signal_12055}), .clk (clk), .r ({Fresh[793], Fresh[792]}), .c ({new_AGEMA_signal_6375, SubBytesIns_Inst_Sbox_4_M50}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M51_U1 ( .a ({new_AGEMA_signal_6225, SubBytesIns_Inst_Sbox_4_M37}), .b ({new_AGEMA_signal_12064, new_AGEMA_signal_12061}), .clk (clk), .r ({Fresh[795], Fresh[794]}), .c ({new_AGEMA_signal_6376, SubBytesIns_Inst_Sbox_4_M51}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M52_U1 ( .a ({new_AGEMA_signal_6370, SubBytesIns_Inst_Sbox_4_M42}), .b ({new_AGEMA_signal_12070, new_AGEMA_signal_12067}), .clk (clk), .r ({Fresh[797], Fresh[796]}), .c ({new_AGEMA_signal_6612, SubBytesIns_Inst_Sbox_4_M52}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M53_U1 ( .a ({new_AGEMA_signal_6609, SubBytesIns_Inst_Sbox_4_M45}), .b ({new_AGEMA_signal_12076, new_AGEMA_signal_12073}), .clk (clk), .r ({Fresh[799], Fresh[798]}), .c ({new_AGEMA_signal_6833, SubBytesIns_Inst_Sbox_4_M53}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M54_U1 ( .a ({new_AGEMA_signal_6369, SubBytesIns_Inst_Sbox_4_M41}), .b ({new_AGEMA_signal_12082, new_AGEMA_signal_12079}), .clk (clk), .r ({Fresh[801], Fresh[800]}), .c ({new_AGEMA_signal_6613, SubBytesIns_Inst_Sbox_4_M54}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M55_U1 ( .a ({new_AGEMA_signal_6372, SubBytesIns_Inst_Sbox_4_M44}), .b ({new_AGEMA_signal_12088, new_AGEMA_signal_12085}), .clk (clk), .r ({Fresh[803], Fresh[802]}), .c ({new_AGEMA_signal_6614, SubBytesIns_Inst_Sbox_4_M55}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M56_U1 ( .a ({new_AGEMA_signal_6228, SubBytesIns_Inst_Sbox_4_M40}), .b ({new_AGEMA_signal_12094, new_AGEMA_signal_12091}), .clk (clk), .r ({Fresh[805], Fresh[804]}), .c ({new_AGEMA_signal_6377, SubBytesIns_Inst_Sbox_4_M56}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M57_U1 ( .a ({new_AGEMA_signal_6227, SubBytesIns_Inst_Sbox_4_M39}), .b ({new_AGEMA_signal_12100, new_AGEMA_signal_12097}), .clk (clk), .r ({Fresh[807], Fresh[806]}), .c ({new_AGEMA_signal_6378, SubBytesIns_Inst_Sbox_4_M57}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M58_U1 ( .a ({new_AGEMA_signal_6371, SubBytesIns_Inst_Sbox_4_M43}), .b ({new_AGEMA_signal_12106, new_AGEMA_signal_12103}), .clk (clk), .r ({Fresh[809], Fresh[808]}), .c ({new_AGEMA_signal_6615, SubBytesIns_Inst_Sbox_4_M58}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M59_U1 ( .a ({new_AGEMA_signal_6226, SubBytesIns_Inst_Sbox_4_M38}), .b ({new_AGEMA_signal_12112, new_AGEMA_signal_12109}), .clk (clk), .r ({Fresh[811], Fresh[810]}), .c ({new_AGEMA_signal_6379, SubBytesIns_Inst_Sbox_4_M59}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M60_U1 ( .a ({new_AGEMA_signal_6225, SubBytesIns_Inst_Sbox_4_M37}), .b ({new_AGEMA_signal_12118, new_AGEMA_signal_12115}), .clk (clk), .r ({Fresh[813], Fresh[812]}), .c ({new_AGEMA_signal_6380, SubBytesIns_Inst_Sbox_4_M60}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M61_U1 ( .a ({new_AGEMA_signal_6370, SubBytesIns_Inst_Sbox_4_M42}), .b ({new_AGEMA_signal_12124, new_AGEMA_signal_12121}), .clk (clk), .r ({Fresh[815], Fresh[814]}), .c ({new_AGEMA_signal_6616, SubBytesIns_Inst_Sbox_4_M61}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M62_U1 ( .a ({new_AGEMA_signal_6609, SubBytesIns_Inst_Sbox_4_M45}), .b ({new_AGEMA_signal_12130, new_AGEMA_signal_12127}), .clk (clk), .r ({Fresh[817], Fresh[816]}), .c ({new_AGEMA_signal_6834, SubBytesIns_Inst_Sbox_4_M62}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M63_U1 ( .a ({new_AGEMA_signal_6369, SubBytesIns_Inst_Sbox_4_M41}), .b ({new_AGEMA_signal_12136, new_AGEMA_signal_12133}), .clk (clk), .r ({Fresh[819], Fresh[818]}), .c ({new_AGEMA_signal_6617, SubBytesIns_Inst_Sbox_4_M63}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L0_U1 ( .a ({new_AGEMA_signal_6616, SubBytesIns_Inst_Sbox_4_M61}), .b ({new_AGEMA_signal_6834, SubBytesIns_Inst_Sbox_4_M62}), .c ({new_AGEMA_signal_7025, SubBytesIns_Inst_Sbox_4_L0}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L1_U1 ( .a ({new_AGEMA_signal_6375, SubBytesIns_Inst_Sbox_4_M50}), .b ({new_AGEMA_signal_6377, SubBytesIns_Inst_Sbox_4_M56}), .c ({new_AGEMA_signal_6618, SubBytesIns_Inst_Sbox_4_L1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L2_U1 ( .a ({new_AGEMA_signal_6610, SubBytesIns_Inst_Sbox_4_M46}), .b ({new_AGEMA_signal_6374, SubBytesIns_Inst_Sbox_4_M48}), .c ({new_AGEMA_signal_6835, SubBytesIns_Inst_Sbox_4_L2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L3_U1 ( .a ({new_AGEMA_signal_6373, SubBytesIns_Inst_Sbox_4_M47}), .b ({new_AGEMA_signal_6614, SubBytesIns_Inst_Sbox_4_M55}), .c ({new_AGEMA_signal_6836, SubBytesIns_Inst_Sbox_4_L3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L4_U1 ( .a ({new_AGEMA_signal_6613, SubBytesIns_Inst_Sbox_4_M54}), .b ({new_AGEMA_signal_6615, SubBytesIns_Inst_Sbox_4_M58}), .c ({new_AGEMA_signal_6837, SubBytesIns_Inst_Sbox_4_L4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L5_U1 ( .a ({new_AGEMA_signal_6611, SubBytesIns_Inst_Sbox_4_M49}), .b ({new_AGEMA_signal_6616, SubBytesIns_Inst_Sbox_4_M61}), .c ({new_AGEMA_signal_6838, SubBytesIns_Inst_Sbox_4_L5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L6_U1 ( .a ({new_AGEMA_signal_6834, SubBytesIns_Inst_Sbox_4_M62}), .b ({new_AGEMA_signal_6838, SubBytesIns_Inst_Sbox_4_L5}), .c ({new_AGEMA_signal_7026, SubBytesIns_Inst_Sbox_4_L6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L7_U1 ( .a ({new_AGEMA_signal_6610, SubBytesIns_Inst_Sbox_4_M46}), .b ({new_AGEMA_signal_6836, SubBytesIns_Inst_Sbox_4_L3}), .c ({new_AGEMA_signal_7027, SubBytesIns_Inst_Sbox_4_L7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L8_U1 ( .a ({new_AGEMA_signal_6376, SubBytesIns_Inst_Sbox_4_M51}), .b ({new_AGEMA_signal_6379, SubBytesIns_Inst_Sbox_4_M59}), .c ({new_AGEMA_signal_6619, SubBytesIns_Inst_Sbox_4_L8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L9_U1 ( .a ({new_AGEMA_signal_6612, SubBytesIns_Inst_Sbox_4_M52}), .b ({new_AGEMA_signal_6833, SubBytesIns_Inst_Sbox_4_M53}), .c ({new_AGEMA_signal_7028, SubBytesIns_Inst_Sbox_4_L9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L10_U1 ( .a ({new_AGEMA_signal_6833, SubBytesIns_Inst_Sbox_4_M53}), .b ({new_AGEMA_signal_6837, SubBytesIns_Inst_Sbox_4_L4}), .c ({new_AGEMA_signal_7029, SubBytesIns_Inst_Sbox_4_L10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L11_U1 ( .a ({new_AGEMA_signal_6380, SubBytesIns_Inst_Sbox_4_M60}), .b ({new_AGEMA_signal_6835, SubBytesIns_Inst_Sbox_4_L2}), .c ({new_AGEMA_signal_7030, SubBytesIns_Inst_Sbox_4_L11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L12_U1 ( .a ({new_AGEMA_signal_6374, SubBytesIns_Inst_Sbox_4_M48}), .b ({new_AGEMA_signal_6376, SubBytesIns_Inst_Sbox_4_M51}), .c ({new_AGEMA_signal_6620, SubBytesIns_Inst_Sbox_4_L12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L13_U1 ( .a ({new_AGEMA_signal_6375, SubBytesIns_Inst_Sbox_4_M50}), .b ({new_AGEMA_signal_7025, SubBytesIns_Inst_Sbox_4_L0}), .c ({new_AGEMA_signal_7221, SubBytesIns_Inst_Sbox_4_L13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L14_U1 ( .a ({new_AGEMA_signal_6612, SubBytesIns_Inst_Sbox_4_M52}), .b ({new_AGEMA_signal_6616, SubBytesIns_Inst_Sbox_4_M61}), .c ({new_AGEMA_signal_6839, SubBytesIns_Inst_Sbox_4_L14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L15_U1 ( .a ({new_AGEMA_signal_6614, SubBytesIns_Inst_Sbox_4_M55}), .b ({new_AGEMA_signal_6618, SubBytesIns_Inst_Sbox_4_L1}), .c ({new_AGEMA_signal_6840, SubBytesIns_Inst_Sbox_4_L15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L16_U1 ( .a ({new_AGEMA_signal_6377, SubBytesIns_Inst_Sbox_4_M56}), .b ({new_AGEMA_signal_7025, SubBytesIns_Inst_Sbox_4_L0}), .c ({new_AGEMA_signal_7222, SubBytesIns_Inst_Sbox_4_L16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L17_U1 ( .a ({new_AGEMA_signal_6378, SubBytesIns_Inst_Sbox_4_M57}), .b ({new_AGEMA_signal_6618, SubBytesIns_Inst_Sbox_4_L1}), .c ({new_AGEMA_signal_6841, SubBytesIns_Inst_Sbox_4_L17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L18_U1 ( .a ({new_AGEMA_signal_6615, SubBytesIns_Inst_Sbox_4_M58}), .b ({new_AGEMA_signal_6619, SubBytesIns_Inst_Sbox_4_L8}), .c ({new_AGEMA_signal_6842, SubBytesIns_Inst_Sbox_4_L18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L19_U1 ( .a ({new_AGEMA_signal_6617, SubBytesIns_Inst_Sbox_4_M63}), .b ({new_AGEMA_signal_6837, SubBytesIns_Inst_Sbox_4_L4}), .c ({new_AGEMA_signal_7031, SubBytesIns_Inst_Sbox_4_L19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L20_U1 ( .a ({new_AGEMA_signal_7025, SubBytesIns_Inst_Sbox_4_L0}), .b ({new_AGEMA_signal_6618, SubBytesIns_Inst_Sbox_4_L1}), .c ({new_AGEMA_signal_7223, SubBytesIns_Inst_Sbox_4_L20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L21_U1 ( .a ({new_AGEMA_signal_6618, SubBytesIns_Inst_Sbox_4_L1}), .b ({new_AGEMA_signal_7027, SubBytesIns_Inst_Sbox_4_L7}), .c ({new_AGEMA_signal_7224, SubBytesIns_Inst_Sbox_4_L21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L22_U1 ( .a ({new_AGEMA_signal_6836, SubBytesIns_Inst_Sbox_4_L3}), .b ({new_AGEMA_signal_6620, SubBytesIns_Inst_Sbox_4_L12}), .c ({new_AGEMA_signal_7032, SubBytesIns_Inst_Sbox_4_L22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L23_U1 ( .a ({new_AGEMA_signal_6842, SubBytesIns_Inst_Sbox_4_L18}), .b ({new_AGEMA_signal_6835, SubBytesIns_Inst_Sbox_4_L2}), .c ({new_AGEMA_signal_7033, SubBytesIns_Inst_Sbox_4_L23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L24_U1 ( .a ({new_AGEMA_signal_6840, SubBytesIns_Inst_Sbox_4_L15}), .b ({new_AGEMA_signal_7028, SubBytesIns_Inst_Sbox_4_L9}), .c ({new_AGEMA_signal_7225, SubBytesIns_Inst_Sbox_4_L24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L25_U1 ( .a ({new_AGEMA_signal_7026, SubBytesIns_Inst_Sbox_4_L6}), .b ({new_AGEMA_signal_7029, SubBytesIns_Inst_Sbox_4_L10}), .c ({new_AGEMA_signal_7226, SubBytesIns_Inst_Sbox_4_L25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L26_U1 ( .a ({new_AGEMA_signal_7027, SubBytesIns_Inst_Sbox_4_L7}), .b ({new_AGEMA_signal_7028, SubBytesIns_Inst_Sbox_4_L9}), .c ({new_AGEMA_signal_7227, SubBytesIns_Inst_Sbox_4_L26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L27_U1 ( .a ({new_AGEMA_signal_6619, SubBytesIns_Inst_Sbox_4_L8}), .b ({new_AGEMA_signal_7029, SubBytesIns_Inst_Sbox_4_L10}), .c ({new_AGEMA_signal_7228, SubBytesIns_Inst_Sbox_4_L27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L28_U1 ( .a ({new_AGEMA_signal_7030, SubBytesIns_Inst_Sbox_4_L11}), .b ({new_AGEMA_signal_6839, SubBytesIns_Inst_Sbox_4_L14}), .c ({new_AGEMA_signal_7229, SubBytesIns_Inst_Sbox_4_L28}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L29_U1 ( .a ({new_AGEMA_signal_7030, SubBytesIns_Inst_Sbox_4_L11}), .b ({new_AGEMA_signal_6841, SubBytesIns_Inst_Sbox_4_L17}), .c ({new_AGEMA_signal_7230, SubBytesIns_Inst_Sbox_4_L29}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_S0_U1 ( .a ({new_AGEMA_signal_7026, SubBytesIns_Inst_Sbox_4_L6}), .b ({new_AGEMA_signal_7225, SubBytesIns_Inst_Sbox_4_L24}), .c ({new_AGEMA_signal_7413, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_S1_U1 ( .a ({new_AGEMA_signal_7222, SubBytesIns_Inst_Sbox_4_L16}), .b ({new_AGEMA_signal_7227, SubBytesIns_Inst_Sbox_4_L26}), .c ({new_AGEMA_signal_7414, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_S2_U1 ( .a ({new_AGEMA_signal_7031, SubBytesIns_Inst_Sbox_4_L19}), .b ({new_AGEMA_signal_7229, SubBytesIns_Inst_Sbox_4_L28}), .c ({new_AGEMA_signal_7415, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_S3_U1 ( .a ({new_AGEMA_signal_7026, SubBytesIns_Inst_Sbox_4_L6}), .b ({new_AGEMA_signal_7224, SubBytesIns_Inst_Sbox_4_L21}), .c ({new_AGEMA_signal_7416, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_S4_U1 ( .a ({new_AGEMA_signal_7223, SubBytesIns_Inst_Sbox_4_L20}), .b ({new_AGEMA_signal_7032, SubBytesIns_Inst_Sbox_4_L22}), .c ({new_AGEMA_signal_7417, MixColumnsInput[3]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_S5_U1 ( .a ({new_AGEMA_signal_7226, SubBytesIns_Inst_Sbox_4_L25}), .b ({new_AGEMA_signal_7230, SubBytesIns_Inst_Sbox_4_L29}), .c ({new_AGEMA_signal_7418, MixColumnsInput[2]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_S6_U1 ( .a ({new_AGEMA_signal_7221, SubBytesIns_Inst_Sbox_4_L13}), .b ({new_AGEMA_signal_7228, SubBytesIns_Inst_Sbox_4_L27}), .c ({new_AGEMA_signal_7419, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_S7_U1 ( .a ({new_AGEMA_signal_7026, SubBytesIns_Inst_Sbox_4_L6}), .b ({new_AGEMA_signal_7033, SubBytesIns_Inst_Sbox_4_L23}), .c ({new_AGEMA_signal_7231, MixColumnsInput[0]}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M46_U1 ( .a ({new_AGEMA_signal_6384, SubBytesIns_Inst_Sbox_5_M44}), .b ({new_AGEMA_signal_12142, new_AGEMA_signal_12139}), .clk (clk), .r ({Fresh[821], Fresh[820]}), .c ({new_AGEMA_signal_6622, SubBytesIns_Inst_Sbox_5_M46}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M47_U1 ( .a ({new_AGEMA_signal_6232, SubBytesIns_Inst_Sbox_5_M40}), .b ({new_AGEMA_signal_12148, new_AGEMA_signal_12145}), .clk (clk), .r ({Fresh[823], Fresh[822]}), .c ({new_AGEMA_signal_6385, SubBytesIns_Inst_Sbox_5_M47}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M48_U1 ( .a ({new_AGEMA_signal_6231, SubBytesIns_Inst_Sbox_5_M39}), .b ({new_AGEMA_signal_12154, new_AGEMA_signal_12151}), .clk (clk), .r ({Fresh[825], Fresh[824]}), .c ({new_AGEMA_signal_6386, SubBytesIns_Inst_Sbox_5_M48}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M49_U1 ( .a ({new_AGEMA_signal_6383, SubBytesIns_Inst_Sbox_5_M43}), .b ({new_AGEMA_signal_12160, new_AGEMA_signal_12157}), .clk (clk), .r ({Fresh[827], Fresh[826]}), .c ({new_AGEMA_signal_6623, SubBytesIns_Inst_Sbox_5_M49}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M50_U1 ( .a ({new_AGEMA_signal_6230, SubBytesIns_Inst_Sbox_5_M38}), .b ({new_AGEMA_signal_12166, new_AGEMA_signal_12163}), .clk (clk), .r ({Fresh[829], Fresh[828]}), .c ({new_AGEMA_signal_6387, SubBytesIns_Inst_Sbox_5_M50}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M51_U1 ( .a ({new_AGEMA_signal_6229, SubBytesIns_Inst_Sbox_5_M37}), .b ({new_AGEMA_signal_12172, new_AGEMA_signal_12169}), .clk (clk), .r ({Fresh[831], Fresh[830]}), .c ({new_AGEMA_signal_6388, SubBytesIns_Inst_Sbox_5_M51}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M52_U1 ( .a ({new_AGEMA_signal_6382, SubBytesIns_Inst_Sbox_5_M42}), .b ({new_AGEMA_signal_12178, new_AGEMA_signal_12175}), .clk (clk), .r ({Fresh[833], Fresh[832]}), .c ({new_AGEMA_signal_6624, SubBytesIns_Inst_Sbox_5_M52}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M53_U1 ( .a ({new_AGEMA_signal_6621, SubBytesIns_Inst_Sbox_5_M45}), .b ({new_AGEMA_signal_12184, new_AGEMA_signal_12181}), .clk (clk), .r ({Fresh[835], Fresh[834]}), .c ({new_AGEMA_signal_6843, SubBytesIns_Inst_Sbox_5_M53}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M54_U1 ( .a ({new_AGEMA_signal_6381, SubBytesIns_Inst_Sbox_5_M41}), .b ({new_AGEMA_signal_12190, new_AGEMA_signal_12187}), .clk (clk), .r ({Fresh[837], Fresh[836]}), .c ({new_AGEMA_signal_6625, SubBytesIns_Inst_Sbox_5_M54}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M55_U1 ( .a ({new_AGEMA_signal_6384, SubBytesIns_Inst_Sbox_5_M44}), .b ({new_AGEMA_signal_12196, new_AGEMA_signal_12193}), .clk (clk), .r ({Fresh[839], Fresh[838]}), .c ({new_AGEMA_signal_6626, SubBytesIns_Inst_Sbox_5_M55}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M56_U1 ( .a ({new_AGEMA_signal_6232, SubBytesIns_Inst_Sbox_5_M40}), .b ({new_AGEMA_signal_12202, new_AGEMA_signal_12199}), .clk (clk), .r ({Fresh[841], Fresh[840]}), .c ({new_AGEMA_signal_6389, SubBytesIns_Inst_Sbox_5_M56}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M57_U1 ( .a ({new_AGEMA_signal_6231, SubBytesIns_Inst_Sbox_5_M39}), .b ({new_AGEMA_signal_12208, new_AGEMA_signal_12205}), .clk (clk), .r ({Fresh[843], Fresh[842]}), .c ({new_AGEMA_signal_6390, SubBytesIns_Inst_Sbox_5_M57}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M58_U1 ( .a ({new_AGEMA_signal_6383, SubBytesIns_Inst_Sbox_5_M43}), .b ({new_AGEMA_signal_12214, new_AGEMA_signal_12211}), .clk (clk), .r ({Fresh[845], Fresh[844]}), .c ({new_AGEMA_signal_6627, SubBytesIns_Inst_Sbox_5_M58}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M59_U1 ( .a ({new_AGEMA_signal_6230, SubBytesIns_Inst_Sbox_5_M38}), .b ({new_AGEMA_signal_12220, new_AGEMA_signal_12217}), .clk (clk), .r ({Fresh[847], Fresh[846]}), .c ({new_AGEMA_signal_6391, SubBytesIns_Inst_Sbox_5_M59}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M60_U1 ( .a ({new_AGEMA_signal_6229, SubBytesIns_Inst_Sbox_5_M37}), .b ({new_AGEMA_signal_12226, new_AGEMA_signal_12223}), .clk (clk), .r ({Fresh[849], Fresh[848]}), .c ({new_AGEMA_signal_6392, SubBytesIns_Inst_Sbox_5_M60}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M61_U1 ( .a ({new_AGEMA_signal_6382, SubBytesIns_Inst_Sbox_5_M42}), .b ({new_AGEMA_signal_12232, new_AGEMA_signal_12229}), .clk (clk), .r ({Fresh[851], Fresh[850]}), .c ({new_AGEMA_signal_6628, SubBytesIns_Inst_Sbox_5_M61}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M62_U1 ( .a ({new_AGEMA_signal_6621, SubBytesIns_Inst_Sbox_5_M45}), .b ({new_AGEMA_signal_12238, new_AGEMA_signal_12235}), .clk (clk), .r ({Fresh[853], Fresh[852]}), .c ({new_AGEMA_signal_6844, SubBytesIns_Inst_Sbox_5_M62}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M63_U1 ( .a ({new_AGEMA_signal_6381, SubBytesIns_Inst_Sbox_5_M41}), .b ({new_AGEMA_signal_12244, new_AGEMA_signal_12241}), .clk (clk), .r ({Fresh[855], Fresh[854]}), .c ({new_AGEMA_signal_6629, SubBytesIns_Inst_Sbox_5_M63}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L0_U1 ( .a ({new_AGEMA_signal_6628, SubBytesIns_Inst_Sbox_5_M61}), .b ({new_AGEMA_signal_6844, SubBytesIns_Inst_Sbox_5_M62}), .c ({new_AGEMA_signal_7034, SubBytesIns_Inst_Sbox_5_L0}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L1_U1 ( .a ({new_AGEMA_signal_6387, SubBytesIns_Inst_Sbox_5_M50}), .b ({new_AGEMA_signal_6389, SubBytesIns_Inst_Sbox_5_M56}), .c ({new_AGEMA_signal_6630, SubBytesIns_Inst_Sbox_5_L1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L2_U1 ( .a ({new_AGEMA_signal_6622, SubBytesIns_Inst_Sbox_5_M46}), .b ({new_AGEMA_signal_6386, SubBytesIns_Inst_Sbox_5_M48}), .c ({new_AGEMA_signal_6845, SubBytesIns_Inst_Sbox_5_L2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L3_U1 ( .a ({new_AGEMA_signal_6385, SubBytesIns_Inst_Sbox_5_M47}), .b ({new_AGEMA_signal_6626, SubBytesIns_Inst_Sbox_5_M55}), .c ({new_AGEMA_signal_6846, SubBytesIns_Inst_Sbox_5_L3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L4_U1 ( .a ({new_AGEMA_signal_6625, SubBytesIns_Inst_Sbox_5_M54}), .b ({new_AGEMA_signal_6627, SubBytesIns_Inst_Sbox_5_M58}), .c ({new_AGEMA_signal_6847, SubBytesIns_Inst_Sbox_5_L4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L5_U1 ( .a ({new_AGEMA_signal_6623, SubBytesIns_Inst_Sbox_5_M49}), .b ({new_AGEMA_signal_6628, SubBytesIns_Inst_Sbox_5_M61}), .c ({new_AGEMA_signal_6848, SubBytesIns_Inst_Sbox_5_L5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L6_U1 ( .a ({new_AGEMA_signal_6844, SubBytesIns_Inst_Sbox_5_M62}), .b ({new_AGEMA_signal_6848, SubBytesIns_Inst_Sbox_5_L5}), .c ({new_AGEMA_signal_7035, SubBytesIns_Inst_Sbox_5_L6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L7_U1 ( .a ({new_AGEMA_signal_6622, SubBytesIns_Inst_Sbox_5_M46}), .b ({new_AGEMA_signal_6846, SubBytesIns_Inst_Sbox_5_L3}), .c ({new_AGEMA_signal_7036, SubBytesIns_Inst_Sbox_5_L7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L8_U1 ( .a ({new_AGEMA_signal_6388, SubBytesIns_Inst_Sbox_5_M51}), .b ({new_AGEMA_signal_6391, SubBytesIns_Inst_Sbox_5_M59}), .c ({new_AGEMA_signal_6631, SubBytesIns_Inst_Sbox_5_L8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L9_U1 ( .a ({new_AGEMA_signal_6624, SubBytesIns_Inst_Sbox_5_M52}), .b ({new_AGEMA_signal_6843, SubBytesIns_Inst_Sbox_5_M53}), .c ({new_AGEMA_signal_7037, SubBytesIns_Inst_Sbox_5_L9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L10_U1 ( .a ({new_AGEMA_signal_6843, SubBytesIns_Inst_Sbox_5_M53}), .b ({new_AGEMA_signal_6847, SubBytesIns_Inst_Sbox_5_L4}), .c ({new_AGEMA_signal_7038, SubBytesIns_Inst_Sbox_5_L10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L11_U1 ( .a ({new_AGEMA_signal_6392, SubBytesIns_Inst_Sbox_5_M60}), .b ({new_AGEMA_signal_6845, SubBytesIns_Inst_Sbox_5_L2}), .c ({new_AGEMA_signal_7039, SubBytesIns_Inst_Sbox_5_L11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L12_U1 ( .a ({new_AGEMA_signal_6386, SubBytesIns_Inst_Sbox_5_M48}), .b ({new_AGEMA_signal_6388, SubBytesIns_Inst_Sbox_5_M51}), .c ({new_AGEMA_signal_6632, SubBytesIns_Inst_Sbox_5_L12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L13_U1 ( .a ({new_AGEMA_signal_6387, SubBytesIns_Inst_Sbox_5_M50}), .b ({new_AGEMA_signal_7034, SubBytesIns_Inst_Sbox_5_L0}), .c ({new_AGEMA_signal_7232, SubBytesIns_Inst_Sbox_5_L13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L14_U1 ( .a ({new_AGEMA_signal_6624, SubBytesIns_Inst_Sbox_5_M52}), .b ({new_AGEMA_signal_6628, SubBytesIns_Inst_Sbox_5_M61}), .c ({new_AGEMA_signal_6849, SubBytesIns_Inst_Sbox_5_L14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L15_U1 ( .a ({new_AGEMA_signal_6626, SubBytesIns_Inst_Sbox_5_M55}), .b ({new_AGEMA_signal_6630, SubBytesIns_Inst_Sbox_5_L1}), .c ({new_AGEMA_signal_6850, SubBytesIns_Inst_Sbox_5_L15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L16_U1 ( .a ({new_AGEMA_signal_6389, SubBytesIns_Inst_Sbox_5_M56}), .b ({new_AGEMA_signal_7034, SubBytesIns_Inst_Sbox_5_L0}), .c ({new_AGEMA_signal_7233, SubBytesIns_Inst_Sbox_5_L16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L17_U1 ( .a ({new_AGEMA_signal_6390, SubBytesIns_Inst_Sbox_5_M57}), .b ({new_AGEMA_signal_6630, SubBytesIns_Inst_Sbox_5_L1}), .c ({new_AGEMA_signal_6851, SubBytesIns_Inst_Sbox_5_L17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L18_U1 ( .a ({new_AGEMA_signal_6627, SubBytesIns_Inst_Sbox_5_M58}), .b ({new_AGEMA_signal_6631, SubBytesIns_Inst_Sbox_5_L8}), .c ({new_AGEMA_signal_6852, SubBytesIns_Inst_Sbox_5_L18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L19_U1 ( .a ({new_AGEMA_signal_6629, SubBytesIns_Inst_Sbox_5_M63}), .b ({new_AGEMA_signal_6847, SubBytesIns_Inst_Sbox_5_L4}), .c ({new_AGEMA_signal_7040, SubBytesIns_Inst_Sbox_5_L19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L20_U1 ( .a ({new_AGEMA_signal_7034, SubBytesIns_Inst_Sbox_5_L0}), .b ({new_AGEMA_signal_6630, SubBytesIns_Inst_Sbox_5_L1}), .c ({new_AGEMA_signal_7234, SubBytesIns_Inst_Sbox_5_L20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L21_U1 ( .a ({new_AGEMA_signal_6630, SubBytesIns_Inst_Sbox_5_L1}), .b ({new_AGEMA_signal_7036, SubBytesIns_Inst_Sbox_5_L7}), .c ({new_AGEMA_signal_7235, SubBytesIns_Inst_Sbox_5_L21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L22_U1 ( .a ({new_AGEMA_signal_6846, SubBytesIns_Inst_Sbox_5_L3}), .b ({new_AGEMA_signal_6632, SubBytesIns_Inst_Sbox_5_L12}), .c ({new_AGEMA_signal_7041, SubBytesIns_Inst_Sbox_5_L22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L23_U1 ( .a ({new_AGEMA_signal_6852, SubBytesIns_Inst_Sbox_5_L18}), .b ({new_AGEMA_signal_6845, SubBytesIns_Inst_Sbox_5_L2}), .c ({new_AGEMA_signal_7042, SubBytesIns_Inst_Sbox_5_L23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L24_U1 ( .a ({new_AGEMA_signal_6850, SubBytesIns_Inst_Sbox_5_L15}), .b ({new_AGEMA_signal_7037, SubBytesIns_Inst_Sbox_5_L9}), .c ({new_AGEMA_signal_7236, SubBytesIns_Inst_Sbox_5_L24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L25_U1 ( .a ({new_AGEMA_signal_7035, SubBytesIns_Inst_Sbox_5_L6}), .b ({new_AGEMA_signal_7038, SubBytesIns_Inst_Sbox_5_L10}), .c ({new_AGEMA_signal_7237, SubBytesIns_Inst_Sbox_5_L25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L26_U1 ( .a ({new_AGEMA_signal_7036, SubBytesIns_Inst_Sbox_5_L7}), .b ({new_AGEMA_signal_7037, SubBytesIns_Inst_Sbox_5_L9}), .c ({new_AGEMA_signal_7238, SubBytesIns_Inst_Sbox_5_L26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L27_U1 ( .a ({new_AGEMA_signal_6631, SubBytesIns_Inst_Sbox_5_L8}), .b ({new_AGEMA_signal_7038, SubBytesIns_Inst_Sbox_5_L10}), .c ({new_AGEMA_signal_7239, SubBytesIns_Inst_Sbox_5_L27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L28_U1 ( .a ({new_AGEMA_signal_7039, SubBytesIns_Inst_Sbox_5_L11}), .b ({new_AGEMA_signal_6849, SubBytesIns_Inst_Sbox_5_L14}), .c ({new_AGEMA_signal_7240, SubBytesIns_Inst_Sbox_5_L28}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L29_U1 ( .a ({new_AGEMA_signal_7039, SubBytesIns_Inst_Sbox_5_L11}), .b ({new_AGEMA_signal_6851, SubBytesIns_Inst_Sbox_5_L17}), .c ({new_AGEMA_signal_7241, SubBytesIns_Inst_Sbox_5_L29}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_S0_U1 ( .a ({new_AGEMA_signal_7035, SubBytesIns_Inst_Sbox_5_L6}), .b ({new_AGEMA_signal_7236, SubBytesIns_Inst_Sbox_5_L24}), .c ({new_AGEMA_signal_7420, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_S1_U1 ( .a ({new_AGEMA_signal_7233, SubBytesIns_Inst_Sbox_5_L16}), .b ({new_AGEMA_signal_7238, SubBytesIns_Inst_Sbox_5_L26}), .c ({new_AGEMA_signal_7421, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_S2_U1 ( .a ({new_AGEMA_signal_7040, SubBytesIns_Inst_Sbox_5_L19}), .b ({new_AGEMA_signal_7240, SubBytesIns_Inst_Sbox_5_L28}), .c ({new_AGEMA_signal_7422, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_S3_U1 ( .a ({new_AGEMA_signal_7035, SubBytesIns_Inst_Sbox_5_L6}), .b ({new_AGEMA_signal_7235, SubBytesIns_Inst_Sbox_5_L21}), .c ({new_AGEMA_signal_7423, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_S4_U1 ( .a ({new_AGEMA_signal_7234, SubBytesIns_Inst_Sbox_5_L20}), .b ({new_AGEMA_signal_7041, SubBytesIns_Inst_Sbox_5_L22}), .c ({new_AGEMA_signal_7424, MixColumnsInput[107]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_S5_U1 ( .a ({new_AGEMA_signal_7237, SubBytesIns_Inst_Sbox_5_L25}), .b ({new_AGEMA_signal_7241, SubBytesIns_Inst_Sbox_5_L29}), .c ({new_AGEMA_signal_7425, MixColumnsInput[106]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_S6_U1 ( .a ({new_AGEMA_signal_7232, SubBytesIns_Inst_Sbox_5_L13}), .b ({new_AGEMA_signal_7239, SubBytesIns_Inst_Sbox_5_L27}), .c ({new_AGEMA_signal_7426, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_S7_U1 ( .a ({new_AGEMA_signal_7035, SubBytesIns_Inst_Sbox_5_L6}), .b ({new_AGEMA_signal_7042, SubBytesIns_Inst_Sbox_5_L23}), .c ({new_AGEMA_signal_7242, MixColumnsInput[104]}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M46_U1 ( .a ({new_AGEMA_signal_6396, SubBytesIns_Inst_Sbox_6_M44}), .b ({new_AGEMA_signal_12250, new_AGEMA_signal_12247}), .clk (clk), .r ({Fresh[857], Fresh[856]}), .c ({new_AGEMA_signal_6634, SubBytesIns_Inst_Sbox_6_M46}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M47_U1 ( .a ({new_AGEMA_signal_6236, SubBytesIns_Inst_Sbox_6_M40}), .b ({new_AGEMA_signal_12256, new_AGEMA_signal_12253}), .clk (clk), .r ({Fresh[859], Fresh[858]}), .c ({new_AGEMA_signal_6397, SubBytesIns_Inst_Sbox_6_M47}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M48_U1 ( .a ({new_AGEMA_signal_6235, SubBytesIns_Inst_Sbox_6_M39}), .b ({new_AGEMA_signal_12262, new_AGEMA_signal_12259}), .clk (clk), .r ({Fresh[861], Fresh[860]}), .c ({new_AGEMA_signal_6398, SubBytesIns_Inst_Sbox_6_M48}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M49_U1 ( .a ({new_AGEMA_signal_6395, SubBytesIns_Inst_Sbox_6_M43}), .b ({new_AGEMA_signal_12268, new_AGEMA_signal_12265}), .clk (clk), .r ({Fresh[863], Fresh[862]}), .c ({new_AGEMA_signal_6635, SubBytesIns_Inst_Sbox_6_M49}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M50_U1 ( .a ({new_AGEMA_signal_6234, SubBytesIns_Inst_Sbox_6_M38}), .b ({new_AGEMA_signal_12274, new_AGEMA_signal_12271}), .clk (clk), .r ({Fresh[865], Fresh[864]}), .c ({new_AGEMA_signal_6399, SubBytesIns_Inst_Sbox_6_M50}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M51_U1 ( .a ({new_AGEMA_signal_6233, SubBytesIns_Inst_Sbox_6_M37}), .b ({new_AGEMA_signal_12280, new_AGEMA_signal_12277}), .clk (clk), .r ({Fresh[867], Fresh[866]}), .c ({new_AGEMA_signal_6400, SubBytesIns_Inst_Sbox_6_M51}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M52_U1 ( .a ({new_AGEMA_signal_6394, SubBytesIns_Inst_Sbox_6_M42}), .b ({new_AGEMA_signal_12286, new_AGEMA_signal_12283}), .clk (clk), .r ({Fresh[869], Fresh[868]}), .c ({new_AGEMA_signal_6636, SubBytesIns_Inst_Sbox_6_M52}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M53_U1 ( .a ({new_AGEMA_signal_6633, SubBytesIns_Inst_Sbox_6_M45}), .b ({new_AGEMA_signal_12292, new_AGEMA_signal_12289}), .clk (clk), .r ({Fresh[871], Fresh[870]}), .c ({new_AGEMA_signal_6853, SubBytesIns_Inst_Sbox_6_M53}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M54_U1 ( .a ({new_AGEMA_signal_6393, SubBytesIns_Inst_Sbox_6_M41}), .b ({new_AGEMA_signal_12298, new_AGEMA_signal_12295}), .clk (clk), .r ({Fresh[873], Fresh[872]}), .c ({new_AGEMA_signal_6637, SubBytesIns_Inst_Sbox_6_M54}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M55_U1 ( .a ({new_AGEMA_signal_6396, SubBytesIns_Inst_Sbox_6_M44}), .b ({new_AGEMA_signal_12304, new_AGEMA_signal_12301}), .clk (clk), .r ({Fresh[875], Fresh[874]}), .c ({new_AGEMA_signal_6638, SubBytesIns_Inst_Sbox_6_M55}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M56_U1 ( .a ({new_AGEMA_signal_6236, SubBytesIns_Inst_Sbox_6_M40}), .b ({new_AGEMA_signal_12310, new_AGEMA_signal_12307}), .clk (clk), .r ({Fresh[877], Fresh[876]}), .c ({new_AGEMA_signal_6401, SubBytesIns_Inst_Sbox_6_M56}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M57_U1 ( .a ({new_AGEMA_signal_6235, SubBytesIns_Inst_Sbox_6_M39}), .b ({new_AGEMA_signal_12316, new_AGEMA_signal_12313}), .clk (clk), .r ({Fresh[879], Fresh[878]}), .c ({new_AGEMA_signal_6402, SubBytesIns_Inst_Sbox_6_M57}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M58_U1 ( .a ({new_AGEMA_signal_6395, SubBytesIns_Inst_Sbox_6_M43}), .b ({new_AGEMA_signal_12322, new_AGEMA_signal_12319}), .clk (clk), .r ({Fresh[881], Fresh[880]}), .c ({new_AGEMA_signal_6639, SubBytesIns_Inst_Sbox_6_M58}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M59_U1 ( .a ({new_AGEMA_signal_6234, SubBytesIns_Inst_Sbox_6_M38}), .b ({new_AGEMA_signal_12328, new_AGEMA_signal_12325}), .clk (clk), .r ({Fresh[883], Fresh[882]}), .c ({new_AGEMA_signal_6403, SubBytesIns_Inst_Sbox_6_M59}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M60_U1 ( .a ({new_AGEMA_signal_6233, SubBytesIns_Inst_Sbox_6_M37}), .b ({new_AGEMA_signal_12334, new_AGEMA_signal_12331}), .clk (clk), .r ({Fresh[885], Fresh[884]}), .c ({new_AGEMA_signal_6404, SubBytesIns_Inst_Sbox_6_M60}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M61_U1 ( .a ({new_AGEMA_signal_6394, SubBytesIns_Inst_Sbox_6_M42}), .b ({new_AGEMA_signal_12340, new_AGEMA_signal_12337}), .clk (clk), .r ({Fresh[887], Fresh[886]}), .c ({new_AGEMA_signal_6640, SubBytesIns_Inst_Sbox_6_M61}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M62_U1 ( .a ({new_AGEMA_signal_6633, SubBytesIns_Inst_Sbox_6_M45}), .b ({new_AGEMA_signal_12346, new_AGEMA_signal_12343}), .clk (clk), .r ({Fresh[889], Fresh[888]}), .c ({new_AGEMA_signal_6854, SubBytesIns_Inst_Sbox_6_M62}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M63_U1 ( .a ({new_AGEMA_signal_6393, SubBytesIns_Inst_Sbox_6_M41}), .b ({new_AGEMA_signal_12352, new_AGEMA_signal_12349}), .clk (clk), .r ({Fresh[891], Fresh[890]}), .c ({new_AGEMA_signal_6641, SubBytesIns_Inst_Sbox_6_M63}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L0_U1 ( .a ({new_AGEMA_signal_6640, SubBytesIns_Inst_Sbox_6_M61}), .b ({new_AGEMA_signal_6854, SubBytesIns_Inst_Sbox_6_M62}), .c ({new_AGEMA_signal_7043, SubBytesIns_Inst_Sbox_6_L0}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L1_U1 ( .a ({new_AGEMA_signal_6399, SubBytesIns_Inst_Sbox_6_M50}), .b ({new_AGEMA_signal_6401, SubBytesIns_Inst_Sbox_6_M56}), .c ({new_AGEMA_signal_6642, SubBytesIns_Inst_Sbox_6_L1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L2_U1 ( .a ({new_AGEMA_signal_6634, SubBytesIns_Inst_Sbox_6_M46}), .b ({new_AGEMA_signal_6398, SubBytesIns_Inst_Sbox_6_M48}), .c ({new_AGEMA_signal_6855, SubBytesIns_Inst_Sbox_6_L2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L3_U1 ( .a ({new_AGEMA_signal_6397, SubBytesIns_Inst_Sbox_6_M47}), .b ({new_AGEMA_signal_6638, SubBytesIns_Inst_Sbox_6_M55}), .c ({new_AGEMA_signal_6856, SubBytesIns_Inst_Sbox_6_L3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L4_U1 ( .a ({new_AGEMA_signal_6637, SubBytesIns_Inst_Sbox_6_M54}), .b ({new_AGEMA_signal_6639, SubBytesIns_Inst_Sbox_6_M58}), .c ({new_AGEMA_signal_6857, SubBytesIns_Inst_Sbox_6_L4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L5_U1 ( .a ({new_AGEMA_signal_6635, SubBytesIns_Inst_Sbox_6_M49}), .b ({new_AGEMA_signal_6640, SubBytesIns_Inst_Sbox_6_M61}), .c ({new_AGEMA_signal_6858, SubBytesIns_Inst_Sbox_6_L5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L6_U1 ( .a ({new_AGEMA_signal_6854, SubBytesIns_Inst_Sbox_6_M62}), .b ({new_AGEMA_signal_6858, SubBytesIns_Inst_Sbox_6_L5}), .c ({new_AGEMA_signal_7044, SubBytesIns_Inst_Sbox_6_L6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L7_U1 ( .a ({new_AGEMA_signal_6634, SubBytesIns_Inst_Sbox_6_M46}), .b ({new_AGEMA_signal_6856, SubBytesIns_Inst_Sbox_6_L3}), .c ({new_AGEMA_signal_7045, SubBytesIns_Inst_Sbox_6_L7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L8_U1 ( .a ({new_AGEMA_signal_6400, SubBytesIns_Inst_Sbox_6_M51}), .b ({new_AGEMA_signal_6403, SubBytesIns_Inst_Sbox_6_M59}), .c ({new_AGEMA_signal_6643, SubBytesIns_Inst_Sbox_6_L8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L9_U1 ( .a ({new_AGEMA_signal_6636, SubBytesIns_Inst_Sbox_6_M52}), .b ({new_AGEMA_signal_6853, SubBytesIns_Inst_Sbox_6_M53}), .c ({new_AGEMA_signal_7046, SubBytesIns_Inst_Sbox_6_L9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L10_U1 ( .a ({new_AGEMA_signal_6853, SubBytesIns_Inst_Sbox_6_M53}), .b ({new_AGEMA_signal_6857, SubBytesIns_Inst_Sbox_6_L4}), .c ({new_AGEMA_signal_7047, SubBytesIns_Inst_Sbox_6_L10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L11_U1 ( .a ({new_AGEMA_signal_6404, SubBytesIns_Inst_Sbox_6_M60}), .b ({new_AGEMA_signal_6855, SubBytesIns_Inst_Sbox_6_L2}), .c ({new_AGEMA_signal_7048, SubBytesIns_Inst_Sbox_6_L11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L12_U1 ( .a ({new_AGEMA_signal_6398, SubBytesIns_Inst_Sbox_6_M48}), .b ({new_AGEMA_signal_6400, SubBytesIns_Inst_Sbox_6_M51}), .c ({new_AGEMA_signal_6644, SubBytesIns_Inst_Sbox_6_L12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L13_U1 ( .a ({new_AGEMA_signal_6399, SubBytesIns_Inst_Sbox_6_M50}), .b ({new_AGEMA_signal_7043, SubBytesIns_Inst_Sbox_6_L0}), .c ({new_AGEMA_signal_7243, SubBytesIns_Inst_Sbox_6_L13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L14_U1 ( .a ({new_AGEMA_signal_6636, SubBytesIns_Inst_Sbox_6_M52}), .b ({new_AGEMA_signal_6640, SubBytesIns_Inst_Sbox_6_M61}), .c ({new_AGEMA_signal_6859, SubBytesIns_Inst_Sbox_6_L14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L15_U1 ( .a ({new_AGEMA_signal_6638, SubBytesIns_Inst_Sbox_6_M55}), .b ({new_AGEMA_signal_6642, SubBytesIns_Inst_Sbox_6_L1}), .c ({new_AGEMA_signal_6860, SubBytesIns_Inst_Sbox_6_L15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L16_U1 ( .a ({new_AGEMA_signal_6401, SubBytesIns_Inst_Sbox_6_M56}), .b ({new_AGEMA_signal_7043, SubBytesIns_Inst_Sbox_6_L0}), .c ({new_AGEMA_signal_7244, SubBytesIns_Inst_Sbox_6_L16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L17_U1 ( .a ({new_AGEMA_signal_6402, SubBytesIns_Inst_Sbox_6_M57}), .b ({new_AGEMA_signal_6642, SubBytesIns_Inst_Sbox_6_L1}), .c ({new_AGEMA_signal_6861, SubBytesIns_Inst_Sbox_6_L17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L18_U1 ( .a ({new_AGEMA_signal_6639, SubBytesIns_Inst_Sbox_6_M58}), .b ({new_AGEMA_signal_6643, SubBytesIns_Inst_Sbox_6_L8}), .c ({new_AGEMA_signal_6862, SubBytesIns_Inst_Sbox_6_L18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L19_U1 ( .a ({new_AGEMA_signal_6641, SubBytesIns_Inst_Sbox_6_M63}), .b ({new_AGEMA_signal_6857, SubBytesIns_Inst_Sbox_6_L4}), .c ({new_AGEMA_signal_7049, SubBytesIns_Inst_Sbox_6_L19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L20_U1 ( .a ({new_AGEMA_signal_7043, SubBytesIns_Inst_Sbox_6_L0}), .b ({new_AGEMA_signal_6642, SubBytesIns_Inst_Sbox_6_L1}), .c ({new_AGEMA_signal_7245, SubBytesIns_Inst_Sbox_6_L20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L21_U1 ( .a ({new_AGEMA_signal_6642, SubBytesIns_Inst_Sbox_6_L1}), .b ({new_AGEMA_signal_7045, SubBytesIns_Inst_Sbox_6_L7}), .c ({new_AGEMA_signal_7246, SubBytesIns_Inst_Sbox_6_L21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L22_U1 ( .a ({new_AGEMA_signal_6856, SubBytesIns_Inst_Sbox_6_L3}), .b ({new_AGEMA_signal_6644, SubBytesIns_Inst_Sbox_6_L12}), .c ({new_AGEMA_signal_7050, SubBytesIns_Inst_Sbox_6_L22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L23_U1 ( .a ({new_AGEMA_signal_6862, SubBytesIns_Inst_Sbox_6_L18}), .b ({new_AGEMA_signal_6855, SubBytesIns_Inst_Sbox_6_L2}), .c ({new_AGEMA_signal_7051, SubBytesIns_Inst_Sbox_6_L23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L24_U1 ( .a ({new_AGEMA_signal_6860, SubBytesIns_Inst_Sbox_6_L15}), .b ({new_AGEMA_signal_7046, SubBytesIns_Inst_Sbox_6_L9}), .c ({new_AGEMA_signal_7247, SubBytesIns_Inst_Sbox_6_L24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L25_U1 ( .a ({new_AGEMA_signal_7044, SubBytesIns_Inst_Sbox_6_L6}), .b ({new_AGEMA_signal_7047, SubBytesIns_Inst_Sbox_6_L10}), .c ({new_AGEMA_signal_7248, SubBytesIns_Inst_Sbox_6_L25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L26_U1 ( .a ({new_AGEMA_signal_7045, SubBytesIns_Inst_Sbox_6_L7}), .b ({new_AGEMA_signal_7046, SubBytesIns_Inst_Sbox_6_L9}), .c ({new_AGEMA_signal_7249, SubBytesIns_Inst_Sbox_6_L26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L27_U1 ( .a ({new_AGEMA_signal_6643, SubBytesIns_Inst_Sbox_6_L8}), .b ({new_AGEMA_signal_7047, SubBytesIns_Inst_Sbox_6_L10}), .c ({new_AGEMA_signal_7250, SubBytesIns_Inst_Sbox_6_L27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L28_U1 ( .a ({new_AGEMA_signal_7048, SubBytesIns_Inst_Sbox_6_L11}), .b ({new_AGEMA_signal_6859, SubBytesIns_Inst_Sbox_6_L14}), .c ({new_AGEMA_signal_7251, SubBytesIns_Inst_Sbox_6_L28}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L29_U1 ( .a ({new_AGEMA_signal_7048, SubBytesIns_Inst_Sbox_6_L11}), .b ({new_AGEMA_signal_6861, SubBytesIns_Inst_Sbox_6_L17}), .c ({new_AGEMA_signal_7252, SubBytesIns_Inst_Sbox_6_L29}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_S0_U1 ( .a ({new_AGEMA_signal_7044, SubBytesIns_Inst_Sbox_6_L6}), .b ({new_AGEMA_signal_7247, SubBytesIns_Inst_Sbox_6_L24}), .c ({new_AGEMA_signal_7427, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_S1_U1 ( .a ({new_AGEMA_signal_7244, SubBytesIns_Inst_Sbox_6_L16}), .b ({new_AGEMA_signal_7249, SubBytesIns_Inst_Sbox_6_L26}), .c ({new_AGEMA_signal_7428, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_S2_U1 ( .a ({new_AGEMA_signal_7049, SubBytesIns_Inst_Sbox_6_L19}), .b ({new_AGEMA_signal_7251, SubBytesIns_Inst_Sbox_6_L28}), .c ({new_AGEMA_signal_7429, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_S3_U1 ( .a ({new_AGEMA_signal_7044, SubBytesIns_Inst_Sbox_6_L6}), .b ({new_AGEMA_signal_7246, SubBytesIns_Inst_Sbox_6_L21}), .c ({new_AGEMA_signal_7430, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_S4_U1 ( .a ({new_AGEMA_signal_7245, SubBytesIns_Inst_Sbox_6_L20}), .b ({new_AGEMA_signal_7050, SubBytesIns_Inst_Sbox_6_L22}), .c ({new_AGEMA_signal_7431, MixColumnsInput[83]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_S5_U1 ( .a ({new_AGEMA_signal_7248, SubBytesIns_Inst_Sbox_6_L25}), .b ({new_AGEMA_signal_7252, SubBytesIns_Inst_Sbox_6_L29}), .c ({new_AGEMA_signal_7432, MixColumnsInput[82]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_S6_U1 ( .a ({new_AGEMA_signal_7243, SubBytesIns_Inst_Sbox_6_L13}), .b ({new_AGEMA_signal_7250, SubBytesIns_Inst_Sbox_6_L27}), .c ({new_AGEMA_signal_7433, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_S7_U1 ( .a ({new_AGEMA_signal_7044, SubBytesIns_Inst_Sbox_6_L6}), .b ({new_AGEMA_signal_7051, SubBytesIns_Inst_Sbox_6_L23}), .c ({new_AGEMA_signal_7253, MixColumnsInput[80]}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M46_U1 ( .a ({new_AGEMA_signal_6408, SubBytesIns_Inst_Sbox_7_M44}), .b ({new_AGEMA_signal_12358, new_AGEMA_signal_12355}), .clk (clk), .r ({Fresh[893], Fresh[892]}), .c ({new_AGEMA_signal_6646, SubBytesIns_Inst_Sbox_7_M46}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M47_U1 ( .a ({new_AGEMA_signal_6240, SubBytesIns_Inst_Sbox_7_M40}), .b ({new_AGEMA_signal_12364, new_AGEMA_signal_12361}), .clk (clk), .r ({Fresh[895], Fresh[894]}), .c ({new_AGEMA_signal_6409, SubBytesIns_Inst_Sbox_7_M47}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M48_U1 ( .a ({new_AGEMA_signal_6239, SubBytesIns_Inst_Sbox_7_M39}), .b ({new_AGEMA_signal_12370, new_AGEMA_signal_12367}), .clk (clk), .r ({Fresh[897], Fresh[896]}), .c ({new_AGEMA_signal_6410, SubBytesIns_Inst_Sbox_7_M48}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M49_U1 ( .a ({new_AGEMA_signal_6407, SubBytesIns_Inst_Sbox_7_M43}), .b ({new_AGEMA_signal_12376, new_AGEMA_signal_12373}), .clk (clk), .r ({Fresh[899], Fresh[898]}), .c ({new_AGEMA_signal_6647, SubBytesIns_Inst_Sbox_7_M49}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M50_U1 ( .a ({new_AGEMA_signal_6238, SubBytesIns_Inst_Sbox_7_M38}), .b ({new_AGEMA_signal_12382, new_AGEMA_signal_12379}), .clk (clk), .r ({Fresh[901], Fresh[900]}), .c ({new_AGEMA_signal_6411, SubBytesIns_Inst_Sbox_7_M50}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M51_U1 ( .a ({new_AGEMA_signal_6237, SubBytesIns_Inst_Sbox_7_M37}), .b ({new_AGEMA_signal_12388, new_AGEMA_signal_12385}), .clk (clk), .r ({Fresh[903], Fresh[902]}), .c ({new_AGEMA_signal_6412, SubBytesIns_Inst_Sbox_7_M51}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M52_U1 ( .a ({new_AGEMA_signal_6406, SubBytesIns_Inst_Sbox_7_M42}), .b ({new_AGEMA_signal_12394, new_AGEMA_signal_12391}), .clk (clk), .r ({Fresh[905], Fresh[904]}), .c ({new_AGEMA_signal_6648, SubBytesIns_Inst_Sbox_7_M52}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M53_U1 ( .a ({new_AGEMA_signal_6645, SubBytesIns_Inst_Sbox_7_M45}), .b ({new_AGEMA_signal_12400, new_AGEMA_signal_12397}), .clk (clk), .r ({Fresh[907], Fresh[906]}), .c ({new_AGEMA_signal_6863, SubBytesIns_Inst_Sbox_7_M53}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M54_U1 ( .a ({new_AGEMA_signal_6405, SubBytesIns_Inst_Sbox_7_M41}), .b ({new_AGEMA_signal_12406, new_AGEMA_signal_12403}), .clk (clk), .r ({Fresh[909], Fresh[908]}), .c ({new_AGEMA_signal_6649, SubBytesIns_Inst_Sbox_7_M54}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M55_U1 ( .a ({new_AGEMA_signal_6408, SubBytesIns_Inst_Sbox_7_M44}), .b ({new_AGEMA_signal_12412, new_AGEMA_signal_12409}), .clk (clk), .r ({Fresh[911], Fresh[910]}), .c ({new_AGEMA_signal_6650, SubBytesIns_Inst_Sbox_7_M55}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M56_U1 ( .a ({new_AGEMA_signal_6240, SubBytesIns_Inst_Sbox_7_M40}), .b ({new_AGEMA_signal_12418, new_AGEMA_signal_12415}), .clk (clk), .r ({Fresh[913], Fresh[912]}), .c ({new_AGEMA_signal_6413, SubBytesIns_Inst_Sbox_7_M56}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M57_U1 ( .a ({new_AGEMA_signal_6239, SubBytesIns_Inst_Sbox_7_M39}), .b ({new_AGEMA_signal_12424, new_AGEMA_signal_12421}), .clk (clk), .r ({Fresh[915], Fresh[914]}), .c ({new_AGEMA_signal_6414, SubBytesIns_Inst_Sbox_7_M57}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M58_U1 ( .a ({new_AGEMA_signal_6407, SubBytesIns_Inst_Sbox_7_M43}), .b ({new_AGEMA_signal_12430, new_AGEMA_signal_12427}), .clk (clk), .r ({Fresh[917], Fresh[916]}), .c ({new_AGEMA_signal_6651, SubBytesIns_Inst_Sbox_7_M58}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M59_U1 ( .a ({new_AGEMA_signal_6238, SubBytesIns_Inst_Sbox_7_M38}), .b ({new_AGEMA_signal_12436, new_AGEMA_signal_12433}), .clk (clk), .r ({Fresh[919], Fresh[918]}), .c ({new_AGEMA_signal_6415, SubBytesIns_Inst_Sbox_7_M59}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M60_U1 ( .a ({new_AGEMA_signal_6237, SubBytesIns_Inst_Sbox_7_M37}), .b ({new_AGEMA_signal_12442, new_AGEMA_signal_12439}), .clk (clk), .r ({Fresh[921], Fresh[920]}), .c ({new_AGEMA_signal_6416, SubBytesIns_Inst_Sbox_7_M60}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M61_U1 ( .a ({new_AGEMA_signal_6406, SubBytesIns_Inst_Sbox_7_M42}), .b ({new_AGEMA_signal_12448, new_AGEMA_signal_12445}), .clk (clk), .r ({Fresh[923], Fresh[922]}), .c ({new_AGEMA_signal_6652, SubBytesIns_Inst_Sbox_7_M61}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M62_U1 ( .a ({new_AGEMA_signal_6645, SubBytesIns_Inst_Sbox_7_M45}), .b ({new_AGEMA_signal_12454, new_AGEMA_signal_12451}), .clk (clk), .r ({Fresh[925], Fresh[924]}), .c ({new_AGEMA_signal_6864, SubBytesIns_Inst_Sbox_7_M62}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M63_U1 ( .a ({new_AGEMA_signal_6405, SubBytesIns_Inst_Sbox_7_M41}), .b ({new_AGEMA_signal_12460, new_AGEMA_signal_12457}), .clk (clk), .r ({Fresh[927], Fresh[926]}), .c ({new_AGEMA_signal_6653, SubBytesIns_Inst_Sbox_7_M63}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L0_U1 ( .a ({new_AGEMA_signal_6652, SubBytesIns_Inst_Sbox_7_M61}), .b ({new_AGEMA_signal_6864, SubBytesIns_Inst_Sbox_7_M62}), .c ({new_AGEMA_signal_7052, SubBytesIns_Inst_Sbox_7_L0}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L1_U1 ( .a ({new_AGEMA_signal_6411, SubBytesIns_Inst_Sbox_7_M50}), .b ({new_AGEMA_signal_6413, SubBytesIns_Inst_Sbox_7_M56}), .c ({new_AGEMA_signal_6654, SubBytesIns_Inst_Sbox_7_L1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L2_U1 ( .a ({new_AGEMA_signal_6646, SubBytesIns_Inst_Sbox_7_M46}), .b ({new_AGEMA_signal_6410, SubBytesIns_Inst_Sbox_7_M48}), .c ({new_AGEMA_signal_6865, SubBytesIns_Inst_Sbox_7_L2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L3_U1 ( .a ({new_AGEMA_signal_6409, SubBytesIns_Inst_Sbox_7_M47}), .b ({new_AGEMA_signal_6650, SubBytesIns_Inst_Sbox_7_M55}), .c ({new_AGEMA_signal_6866, SubBytesIns_Inst_Sbox_7_L3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L4_U1 ( .a ({new_AGEMA_signal_6649, SubBytesIns_Inst_Sbox_7_M54}), .b ({new_AGEMA_signal_6651, SubBytesIns_Inst_Sbox_7_M58}), .c ({new_AGEMA_signal_6867, SubBytesIns_Inst_Sbox_7_L4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L5_U1 ( .a ({new_AGEMA_signal_6647, SubBytesIns_Inst_Sbox_7_M49}), .b ({new_AGEMA_signal_6652, SubBytesIns_Inst_Sbox_7_M61}), .c ({new_AGEMA_signal_6868, SubBytesIns_Inst_Sbox_7_L5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L6_U1 ( .a ({new_AGEMA_signal_6864, SubBytesIns_Inst_Sbox_7_M62}), .b ({new_AGEMA_signal_6868, SubBytesIns_Inst_Sbox_7_L5}), .c ({new_AGEMA_signal_7053, SubBytesIns_Inst_Sbox_7_L6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L7_U1 ( .a ({new_AGEMA_signal_6646, SubBytesIns_Inst_Sbox_7_M46}), .b ({new_AGEMA_signal_6866, SubBytesIns_Inst_Sbox_7_L3}), .c ({new_AGEMA_signal_7054, SubBytesIns_Inst_Sbox_7_L7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L8_U1 ( .a ({new_AGEMA_signal_6412, SubBytesIns_Inst_Sbox_7_M51}), .b ({new_AGEMA_signal_6415, SubBytesIns_Inst_Sbox_7_M59}), .c ({new_AGEMA_signal_6655, SubBytesIns_Inst_Sbox_7_L8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L9_U1 ( .a ({new_AGEMA_signal_6648, SubBytesIns_Inst_Sbox_7_M52}), .b ({new_AGEMA_signal_6863, SubBytesIns_Inst_Sbox_7_M53}), .c ({new_AGEMA_signal_7055, SubBytesIns_Inst_Sbox_7_L9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L10_U1 ( .a ({new_AGEMA_signal_6863, SubBytesIns_Inst_Sbox_7_M53}), .b ({new_AGEMA_signal_6867, SubBytesIns_Inst_Sbox_7_L4}), .c ({new_AGEMA_signal_7056, SubBytesIns_Inst_Sbox_7_L10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L11_U1 ( .a ({new_AGEMA_signal_6416, SubBytesIns_Inst_Sbox_7_M60}), .b ({new_AGEMA_signal_6865, SubBytesIns_Inst_Sbox_7_L2}), .c ({new_AGEMA_signal_7057, SubBytesIns_Inst_Sbox_7_L11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L12_U1 ( .a ({new_AGEMA_signal_6410, SubBytesIns_Inst_Sbox_7_M48}), .b ({new_AGEMA_signal_6412, SubBytesIns_Inst_Sbox_7_M51}), .c ({new_AGEMA_signal_6656, SubBytesIns_Inst_Sbox_7_L12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L13_U1 ( .a ({new_AGEMA_signal_6411, SubBytesIns_Inst_Sbox_7_M50}), .b ({new_AGEMA_signal_7052, SubBytesIns_Inst_Sbox_7_L0}), .c ({new_AGEMA_signal_7254, SubBytesIns_Inst_Sbox_7_L13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L14_U1 ( .a ({new_AGEMA_signal_6648, SubBytesIns_Inst_Sbox_7_M52}), .b ({new_AGEMA_signal_6652, SubBytesIns_Inst_Sbox_7_M61}), .c ({new_AGEMA_signal_6869, SubBytesIns_Inst_Sbox_7_L14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L15_U1 ( .a ({new_AGEMA_signal_6650, SubBytesIns_Inst_Sbox_7_M55}), .b ({new_AGEMA_signal_6654, SubBytesIns_Inst_Sbox_7_L1}), .c ({new_AGEMA_signal_6870, SubBytesIns_Inst_Sbox_7_L15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L16_U1 ( .a ({new_AGEMA_signal_6413, SubBytesIns_Inst_Sbox_7_M56}), .b ({new_AGEMA_signal_7052, SubBytesIns_Inst_Sbox_7_L0}), .c ({new_AGEMA_signal_7255, SubBytesIns_Inst_Sbox_7_L16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L17_U1 ( .a ({new_AGEMA_signal_6414, SubBytesIns_Inst_Sbox_7_M57}), .b ({new_AGEMA_signal_6654, SubBytesIns_Inst_Sbox_7_L1}), .c ({new_AGEMA_signal_6871, SubBytesIns_Inst_Sbox_7_L17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L18_U1 ( .a ({new_AGEMA_signal_6651, SubBytesIns_Inst_Sbox_7_M58}), .b ({new_AGEMA_signal_6655, SubBytesIns_Inst_Sbox_7_L8}), .c ({new_AGEMA_signal_6872, SubBytesIns_Inst_Sbox_7_L18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L19_U1 ( .a ({new_AGEMA_signal_6653, SubBytesIns_Inst_Sbox_7_M63}), .b ({new_AGEMA_signal_6867, SubBytesIns_Inst_Sbox_7_L4}), .c ({new_AGEMA_signal_7058, SubBytesIns_Inst_Sbox_7_L19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L20_U1 ( .a ({new_AGEMA_signal_7052, SubBytesIns_Inst_Sbox_7_L0}), .b ({new_AGEMA_signal_6654, SubBytesIns_Inst_Sbox_7_L1}), .c ({new_AGEMA_signal_7256, SubBytesIns_Inst_Sbox_7_L20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L21_U1 ( .a ({new_AGEMA_signal_6654, SubBytesIns_Inst_Sbox_7_L1}), .b ({new_AGEMA_signal_7054, SubBytesIns_Inst_Sbox_7_L7}), .c ({new_AGEMA_signal_7257, SubBytesIns_Inst_Sbox_7_L21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L22_U1 ( .a ({new_AGEMA_signal_6866, SubBytesIns_Inst_Sbox_7_L3}), .b ({new_AGEMA_signal_6656, SubBytesIns_Inst_Sbox_7_L12}), .c ({new_AGEMA_signal_7059, SubBytesIns_Inst_Sbox_7_L22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L23_U1 ( .a ({new_AGEMA_signal_6872, SubBytesIns_Inst_Sbox_7_L18}), .b ({new_AGEMA_signal_6865, SubBytesIns_Inst_Sbox_7_L2}), .c ({new_AGEMA_signal_7060, SubBytesIns_Inst_Sbox_7_L23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L24_U1 ( .a ({new_AGEMA_signal_6870, SubBytesIns_Inst_Sbox_7_L15}), .b ({new_AGEMA_signal_7055, SubBytesIns_Inst_Sbox_7_L9}), .c ({new_AGEMA_signal_7258, SubBytesIns_Inst_Sbox_7_L24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L25_U1 ( .a ({new_AGEMA_signal_7053, SubBytesIns_Inst_Sbox_7_L6}), .b ({new_AGEMA_signal_7056, SubBytesIns_Inst_Sbox_7_L10}), .c ({new_AGEMA_signal_7259, SubBytesIns_Inst_Sbox_7_L25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L26_U1 ( .a ({new_AGEMA_signal_7054, SubBytesIns_Inst_Sbox_7_L7}), .b ({new_AGEMA_signal_7055, SubBytesIns_Inst_Sbox_7_L9}), .c ({new_AGEMA_signal_7260, SubBytesIns_Inst_Sbox_7_L26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L27_U1 ( .a ({new_AGEMA_signal_6655, SubBytesIns_Inst_Sbox_7_L8}), .b ({new_AGEMA_signal_7056, SubBytesIns_Inst_Sbox_7_L10}), .c ({new_AGEMA_signal_7261, SubBytesIns_Inst_Sbox_7_L27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L28_U1 ( .a ({new_AGEMA_signal_7057, SubBytesIns_Inst_Sbox_7_L11}), .b ({new_AGEMA_signal_6869, SubBytesIns_Inst_Sbox_7_L14}), .c ({new_AGEMA_signal_7262, SubBytesIns_Inst_Sbox_7_L28}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L29_U1 ( .a ({new_AGEMA_signal_7057, SubBytesIns_Inst_Sbox_7_L11}), .b ({new_AGEMA_signal_6871, SubBytesIns_Inst_Sbox_7_L17}), .c ({new_AGEMA_signal_7263, SubBytesIns_Inst_Sbox_7_L29}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_S0_U1 ( .a ({new_AGEMA_signal_7053, SubBytesIns_Inst_Sbox_7_L6}), .b ({new_AGEMA_signal_7258, SubBytesIns_Inst_Sbox_7_L24}), .c ({new_AGEMA_signal_7434, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_S1_U1 ( .a ({new_AGEMA_signal_7255, SubBytesIns_Inst_Sbox_7_L16}), .b ({new_AGEMA_signal_7260, SubBytesIns_Inst_Sbox_7_L26}), .c ({new_AGEMA_signal_7435, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_S2_U1 ( .a ({new_AGEMA_signal_7058, SubBytesIns_Inst_Sbox_7_L19}), .b ({new_AGEMA_signal_7262, SubBytesIns_Inst_Sbox_7_L28}), .c ({new_AGEMA_signal_7436, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_S3_U1 ( .a ({new_AGEMA_signal_7053, SubBytesIns_Inst_Sbox_7_L6}), .b ({new_AGEMA_signal_7257, SubBytesIns_Inst_Sbox_7_L21}), .c ({new_AGEMA_signal_7437, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_S4_U1 ( .a ({new_AGEMA_signal_7256, SubBytesIns_Inst_Sbox_7_L20}), .b ({new_AGEMA_signal_7059, SubBytesIns_Inst_Sbox_7_L22}), .c ({new_AGEMA_signal_7438, MixColumnsInput[59]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_S5_U1 ( .a ({new_AGEMA_signal_7259, SubBytesIns_Inst_Sbox_7_L25}), .b ({new_AGEMA_signal_7263, SubBytesIns_Inst_Sbox_7_L29}), .c ({new_AGEMA_signal_7439, MixColumnsInput[58]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_S6_U1 ( .a ({new_AGEMA_signal_7254, SubBytesIns_Inst_Sbox_7_L13}), .b ({new_AGEMA_signal_7261, SubBytesIns_Inst_Sbox_7_L27}), .c ({new_AGEMA_signal_7440, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_S7_U1 ( .a ({new_AGEMA_signal_7053, SubBytesIns_Inst_Sbox_7_L6}), .b ({new_AGEMA_signal_7060, SubBytesIns_Inst_Sbox_7_L23}), .c ({new_AGEMA_signal_7264, MixColumnsInput[56]}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M46_U1 ( .a ({new_AGEMA_signal_6420, SubBytesIns_Inst_Sbox_8_M44}), .b ({new_AGEMA_signal_12466, new_AGEMA_signal_12463}), .clk (clk), .r ({Fresh[929], Fresh[928]}), .c ({new_AGEMA_signal_6658, SubBytesIns_Inst_Sbox_8_M46}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M47_U1 ( .a ({new_AGEMA_signal_6244, SubBytesIns_Inst_Sbox_8_M40}), .b ({new_AGEMA_signal_12472, new_AGEMA_signal_12469}), .clk (clk), .r ({Fresh[931], Fresh[930]}), .c ({new_AGEMA_signal_6421, SubBytesIns_Inst_Sbox_8_M47}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M48_U1 ( .a ({new_AGEMA_signal_6243, SubBytesIns_Inst_Sbox_8_M39}), .b ({new_AGEMA_signal_12478, new_AGEMA_signal_12475}), .clk (clk), .r ({Fresh[933], Fresh[932]}), .c ({new_AGEMA_signal_6422, SubBytesIns_Inst_Sbox_8_M48}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M49_U1 ( .a ({new_AGEMA_signal_6419, SubBytesIns_Inst_Sbox_8_M43}), .b ({new_AGEMA_signal_12484, new_AGEMA_signal_12481}), .clk (clk), .r ({Fresh[935], Fresh[934]}), .c ({new_AGEMA_signal_6659, SubBytesIns_Inst_Sbox_8_M49}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M50_U1 ( .a ({new_AGEMA_signal_6242, SubBytesIns_Inst_Sbox_8_M38}), .b ({new_AGEMA_signal_12490, new_AGEMA_signal_12487}), .clk (clk), .r ({Fresh[937], Fresh[936]}), .c ({new_AGEMA_signal_6423, SubBytesIns_Inst_Sbox_8_M50}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M51_U1 ( .a ({new_AGEMA_signal_6241, SubBytesIns_Inst_Sbox_8_M37}), .b ({new_AGEMA_signal_12496, new_AGEMA_signal_12493}), .clk (clk), .r ({Fresh[939], Fresh[938]}), .c ({new_AGEMA_signal_6424, SubBytesIns_Inst_Sbox_8_M51}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M52_U1 ( .a ({new_AGEMA_signal_6418, SubBytesIns_Inst_Sbox_8_M42}), .b ({new_AGEMA_signal_12502, new_AGEMA_signal_12499}), .clk (clk), .r ({Fresh[941], Fresh[940]}), .c ({new_AGEMA_signal_6660, SubBytesIns_Inst_Sbox_8_M52}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M53_U1 ( .a ({new_AGEMA_signal_6657, SubBytesIns_Inst_Sbox_8_M45}), .b ({new_AGEMA_signal_12508, new_AGEMA_signal_12505}), .clk (clk), .r ({Fresh[943], Fresh[942]}), .c ({new_AGEMA_signal_6873, SubBytesIns_Inst_Sbox_8_M53}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M54_U1 ( .a ({new_AGEMA_signal_6417, SubBytesIns_Inst_Sbox_8_M41}), .b ({new_AGEMA_signal_12514, new_AGEMA_signal_12511}), .clk (clk), .r ({Fresh[945], Fresh[944]}), .c ({new_AGEMA_signal_6661, SubBytesIns_Inst_Sbox_8_M54}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M55_U1 ( .a ({new_AGEMA_signal_6420, SubBytesIns_Inst_Sbox_8_M44}), .b ({new_AGEMA_signal_12520, new_AGEMA_signal_12517}), .clk (clk), .r ({Fresh[947], Fresh[946]}), .c ({new_AGEMA_signal_6662, SubBytesIns_Inst_Sbox_8_M55}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M56_U1 ( .a ({new_AGEMA_signal_6244, SubBytesIns_Inst_Sbox_8_M40}), .b ({new_AGEMA_signal_12526, new_AGEMA_signal_12523}), .clk (clk), .r ({Fresh[949], Fresh[948]}), .c ({new_AGEMA_signal_6425, SubBytesIns_Inst_Sbox_8_M56}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M57_U1 ( .a ({new_AGEMA_signal_6243, SubBytesIns_Inst_Sbox_8_M39}), .b ({new_AGEMA_signal_12532, new_AGEMA_signal_12529}), .clk (clk), .r ({Fresh[951], Fresh[950]}), .c ({new_AGEMA_signal_6426, SubBytesIns_Inst_Sbox_8_M57}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M58_U1 ( .a ({new_AGEMA_signal_6419, SubBytesIns_Inst_Sbox_8_M43}), .b ({new_AGEMA_signal_12538, new_AGEMA_signal_12535}), .clk (clk), .r ({Fresh[953], Fresh[952]}), .c ({new_AGEMA_signal_6663, SubBytesIns_Inst_Sbox_8_M58}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M59_U1 ( .a ({new_AGEMA_signal_6242, SubBytesIns_Inst_Sbox_8_M38}), .b ({new_AGEMA_signal_12544, new_AGEMA_signal_12541}), .clk (clk), .r ({Fresh[955], Fresh[954]}), .c ({new_AGEMA_signal_6427, SubBytesIns_Inst_Sbox_8_M59}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M60_U1 ( .a ({new_AGEMA_signal_6241, SubBytesIns_Inst_Sbox_8_M37}), .b ({new_AGEMA_signal_12550, new_AGEMA_signal_12547}), .clk (clk), .r ({Fresh[957], Fresh[956]}), .c ({new_AGEMA_signal_6428, SubBytesIns_Inst_Sbox_8_M60}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M61_U1 ( .a ({new_AGEMA_signal_6418, SubBytesIns_Inst_Sbox_8_M42}), .b ({new_AGEMA_signal_12556, new_AGEMA_signal_12553}), .clk (clk), .r ({Fresh[959], Fresh[958]}), .c ({new_AGEMA_signal_6664, SubBytesIns_Inst_Sbox_8_M61}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M62_U1 ( .a ({new_AGEMA_signal_6657, SubBytesIns_Inst_Sbox_8_M45}), .b ({new_AGEMA_signal_12562, new_AGEMA_signal_12559}), .clk (clk), .r ({Fresh[961], Fresh[960]}), .c ({new_AGEMA_signal_6874, SubBytesIns_Inst_Sbox_8_M62}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M63_U1 ( .a ({new_AGEMA_signal_6417, SubBytesIns_Inst_Sbox_8_M41}), .b ({new_AGEMA_signal_12568, new_AGEMA_signal_12565}), .clk (clk), .r ({Fresh[963], Fresh[962]}), .c ({new_AGEMA_signal_6665, SubBytesIns_Inst_Sbox_8_M63}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L0_U1 ( .a ({new_AGEMA_signal_6664, SubBytesIns_Inst_Sbox_8_M61}), .b ({new_AGEMA_signal_6874, SubBytesIns_Inst_Sbox_8_M62}), .c ({new_AGEMA_signal_7061, SubBytesIns_Inst_Sbox_8_L0}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L1_U1 ( .a ({new_AGEMA_signal_6423, SubBytesIns_Inst_Sbox_8_M50}), .b ({new_AGEMA_signal_6425, SubBytesIns_Inst_Sbox_8_M56}), .c ({new_AGEMA_signal_6666, SubBytesIns_Inst_Sbox_8_L1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L2_U1 ( .a ({new_AGEMA_signal_6658, SubBytesIns_Inst_Sbox_8_M46}), .b ({new_AGEMA_signal_6422, SubBytesIns_Inst_Sbox_8_M48}), .c ({new_AGEMA_signal_6875, SubBytesIns_Inst_Sbox_8_L2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L3_U1 ( .a ({new_AGEMA_signal_6421, SubBytesIns_Inst_Sbox_8_M47}), .b ({new_AGEMA_signal_6662, SubBytesIns_Inst_Sbox_8_M55}), .c ({new_AGEMA_signal_6876, SubBytesIns_Inst_Sbox_8_L3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L4_U1 ( .a ({new_AGEMA_signal_6661, SubBytesIns_Inst_Sbox_8_M54}), .b ({new_AGEMA_signal_6663, SubBytesIns_Inst_Sbox_8_M58}), .c ({new_AGEMA_signal_6877, SubBytesIns_Inst_Sbox_8_L4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L5_U1 ( .a ({new_AGEMA_signal_6659, SubBytesIns_Inst_Sbox_8_M49}), .b ({new_AGEMA_signal_6664, SubBytesIns_Inst_Sbox_8_M61}), .c ({new_AGEMA_signal_6878, SubBytesIns_Inst_Sbox_8_L5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L6_U1 ( .a ({new_AGEMA_signal_6874, SubBytesIns_Inst_Sbox_8_M62}), .b ({new_AGEMA_signal_6878, SubBytesIns_Inst_Sbox_8_L5}), .c ({new_AGEMA_signal_7062, SubBytesIns_Inst_Sbox_8_L6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L7_U1 ( .a ({new_AGEMA_signal_6658, SubBytesIns_Inst_Sbox_8_M46}), .b ({new_AGEMA_signal_6876, SubBytesIns_Inst_Sbox_8_L3}), .c ({new_AGEMA_signal_7063, SubBytesIns_Inst_Sbox_8_L7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L8_U1 ( .a ({new_AGEMA_signal_6424, SubBytesIns_Inst_Sbox_8_M51}), .b ({new_AGEMA_signal_6427, SubBytesIns_Inst_Sbox_8_M59}), .c ({new_AGEMA_signal_6667, SubBytesIns_Inst_Sbox_8_L8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L9_U1 ( .a ({new_AGEMA_signal_6660, SubBytesIns_Inst_Sbox_8_M52}), .b ({new_AGEMA_signal_6873, SubBytesIns_Inst_Sbox_8_M53}), .c ({new_AGEMA_signal_7064, SubBytesIns_Inst_Sbox_8_L9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L10_U1 ( .a ({new_AGEMA_signal_6873, SubBytesIns_Inst_Sbox_8_M53}), .b ({new_AGEMA_signal_6877, SubBytesIns_Inst_Sbox_8_L4}), .c ({new_AGEMA_signal_7065, SubBytesIns_Inst_Sbox_8_L10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L11_U1 ( .a ({new_AGEMA_signal_6428, SubBytesIns_Inst_Sbox_8_M60}), .b ({new_AGEMA_signal_6875, SubBytesIns_Inst_Sbox_8_L2}), .c ({new_AGEMA_signal_7066, SubBytesIns_Inst_Sbox_8_L11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L12_U1 ( .a ({new_AGEMA_signal_6422, SubBytesIns_Inst_Sbox_8_M48}), .b ({new_AGEMA_signal_6424, SubBytesIns_Inst_Sbox_8_M51}), .c ({new_AGEMA_signal_6668, SubBytesIns_Inst_Sbox_8_L12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L13_U1 ( .a ({new_AGEMA_signal_6423, SubBytesIns_Inst_Sbox_8_M50}), .b ({new_AGEMA_signal_7061, SubBytesIns_Inst_Sbox_8_L0}), .c ({new_AGEMA_signal_7265, SubBytesIns_Inst_Sbox_8_L13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L14_U1 ( .a ({new_AGEMA_signal_6660, SubBytesIns_Inst_Sbox_8_M52}), .b ({new_AGEMA_signal_6664, SubBytesIns_Inst_Sbox_8_M61}), .c ({new_AGEMA_signal_6879, SubBytesIns_Inst_Sbox_8_L14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L15_U1 ( .a ({new_AGEMA_signal_6662, SubBytesIns_Inst_Sbox_8_M55}), .b ({new_AGEMA_signal_6666, SubBytesIns_Inst_Sbox_8_L1}), .c ({new_AGEMA_signal_6880, SubBytesIns_Inst_Sbox_8_L15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L16_U1 ( .a ({new_AGEMA_signal_6425, SubBytesIns_Inst_Sbox_8_M56}), .b ({new_AGEMA_signal_7061, SubBytesIns_Inst_Sbox_8_L0}), .c ({new_AGEMA_signal_7266, SubBytesIns_Inst_Sbox_8_L16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L17_U1 ( .a ({new_AGEMA_signal_6426, SubBytesIns_Inst_Sbox_8_M57}), .b ({new_AGEMA_signal_6666, SubBytesIns_Inst_Sbox_8_L1}), .c ({new_AGEMA_signal_6881, SubBytesIns_Inst_Sbox_8_L17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L18_U1 ( .a ({new_AGEMA_signal_6663, SubBytesIns_Inst_Sbox_8_M58}), .b ({new_AGEMA_signal_6667, SubBytesIns_Inst_Sbox_8_L8}), .c ({new_AGEMA_signal_6882, SubBytesIns_Inst_Sbox_8_L18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L19_U1 ( .a ({new_AGEMA_signal_6665, SubBytesIns_Inst_Sbox_8_M63}), .b ({new_AGEMA_signal_6877, SubBytesIns_Inst_Sbox_8_L4}), .c ({new_AGEMA_signal_7067, SubBytesIns_Inst_Sbox_8_L19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L20_U1 ( .a ({new_AGEMA_signal_7061, SubBytesIns_Inst_Sbox_8_L0}), .b ({new_AGEMA_signal_6666, SubBytesIns_Inst_Sbox_8_L1}), .c ({new_AGEMA_signal_7267, SubBytesIns_Inst_Sbox_8_L20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L21_U1 ( .a ({new_AGEMA_signal_6666, SubBytesIns_Inst_Sbox_8_L1}), .b ({new_AGEMA_signal_7063, SubBytesIns_Inst_Sbox_8_L7}), .c ({new_AGEMA_signal_7268, SubBytesIns_Inst_Sbox_8_L21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L22_U1 ( .a ({new_AGEMA_signal_6876, SubBytesIns_Inst_Sbox_8_L3}), .b ({new_AGEMA_signal_6668, SubBytesIns_Inst_Sbox_8_L12}), .c ({new_AGEMA_signal_7068, SubBytesIns_Inst_Sbox_8_L22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L23_U1 ( .a ({new_AGEMA_signal_6882, SubBytesIns_Inst_Sbox_8_L18}), .b ({new_AGEMA_signal_6875, SubBytesIns_Inst_Sbox_8_L2}), .c ({new_AGEMA_signal_7069, SubBytesIns_Inst_Sbox_8_L23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L24_U1 ( .a ({new_AGEMA_signal_6880, SubBytesIns_Inst_Sbox_8_L15}), .b ({new_AGEMA_signal_7064, SubBytesIns_Inst_Sbox_8_L9}), .c ({new_AGEMA_signal_7269, SubBytesIns_Inst_Sbox_8_L24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L25_U1 ( .a ({new_AGEMA_signal_7062, SubBytesIns_Inst_Sbox_8_L6}), .b ({new_AGEMA_signal_7065, SubBytesIns_Inst_Sbox_8_L10}), .c ({new_AGEMA_signal_7270, SubBytesIns_Inst_Sbox_8_L25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L26_U1 ( .a ({new_AGEMA_signal_7063, SubBytesIns_Inst_Sbox_8_L7}), .b ({new_AGEMA_signal_7064, SubBytesIns_Inst_Sbox_8_L9}), .c ({new_AGEMA_signal_7271, SubBytesIns_Inst_Sbox_8_L26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L27_U1 ( .a ({new_AGEMA_signal_6667, SubBytesIns_Inst_Sbox_8_L8}), .b ({new_AGEMA_signal_7065, SubBytesIns_Inst_Sbox_8_L10}), .c ({new_AGEMA_signal_7272, SubBytesIns_Inst_Sbox_8_L27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L28_U1 ( .a ({new_AGEMA_signal_7066, SubBytesIns_Inst_Sbox_8_L11}), .b ({new_AGEMA_signal_6879, SubBytesIns_Inst_Sbox_8_L14}), .c ({new_AGEMA_signal_7273, SubBytesIns_Inst_Sbox_8_L28}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L29_U1 ( .a ({new_AGEMA_signal_7066, SubBytesIns_Inst_Sbox_8_L11}), .b ({new_AGEMA_signal_6881, SubBytesIns_Inst_Sbox_8_L17}), .c ({new_AGEMA_signal_7274, SubBytesIns_Inst_Sbox_8_L29}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_S0_U1 ( .a ({new_AGEMA_signal_7062, SubBytesIns_Inst_Sbox_8_L6}), .b ({new_AGEMA_signal_7269, SubBytesIns_Inst_Sbox_8_L24}), .c ({new_AGEMA_signal_7441, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_S1_U1 ( .a ({new_AGEMA_signal_7266, SubBytesIns_Inst_Sbox_8_L16}), .b ({new_AGEMA_signal_7271, SubBytesIns_Inst_Sbox_8_L26}), .c ({new_AGEMA_signal_7442, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_S2_U1 ( .a ({new_AGEMA_signal_7067, SubBytesIns_Inst_Sbox_8_L19}), .b ({new_AGEMA_signal_7273, SubBytesIns_Inst_Sbox_8_L28}), .c ({new_AGEMA_signal_7443, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_S3_U1 ( .a ({new_AGEMA_signal_7062, SubBytesIns_Inst_Sbox_8_L6}), .b ({new_AGEMA_signal_7268, SubBytesIns_Inst_Sbox_8_L21}), .c ({new_AGEMA_signal_7444, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_S4_U1 ( .a ({new_AGEMA_signal_7267, SubBytesIns_Inst_Sbox_8_L20}), .b ({new_AGEMA_signal_7068, SubBytesIns_Inst_Sbox_8_L22}), .c ({new_AGEMA_signal_7445, MixColumnsInput[35]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_S5_U1 ( .a ({new_AGEMA_signal_7270, SubBytesIns_Inst_Sbox_8_L25}), .b ({new_AGEMA_signal_7274, SubBytesIns_Inst_Sbox_8_L29}), .c ({new_AGEMA_signal_7446, MixColumnsInput[34]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_S6_U1 ( .a ({new_AGEMA_signal_7265, SubBytesIns_Inst_Sbox_8_L13}), .b ({new_AGEMA_signal_7272, SubBytesIns_Inst_Sbox_8_L27}), .c ({new_AGEMA_signal_7447, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_S7_U1 ( .a ({new_AGEMA_signal_7062, SubBytesIns_Inst_Sbox_8_L6}), .b ({new_AGEMA_signal_7069, SubBytesIns_Inst_Sbox_8_L23}), .c ({new_AGEMA_signal_7275, MixColumnsInput[32]}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M46_U1 ( .a ({new_AGEMA_signal_6432, SubBytesIns_Inst_Sbox_9_M44}), .b ({new_AGEMA_signal_12574, new_AGEMA_signal_12571}), .clk (clk), .r ({Fresh[965], Fresh[964]}), .c ({new_AGEMA_signal_6670, SubBytesIns_Inst_Sbox_9_M46}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M47_U1 ( .a ({new_AGEMA_signal_6248, SubBytesIns_Inst_Sbox_9_M40}), .b ({new_AGEMA_signal_12580, new_AGEMA_signal_12577}), .clk (clk), .r ({Fresh[967], Fresh[966]}), .c ({new_AGEMA_signal_6433, SubBytesIns_Inst_Sbox_9_M47}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M48_U1 ( .a ({new_AGEMA_signal_6247, SubBytesIns_Inst_Sbox_9_M39}), .b ({new_AGEMA_signal_12586, new_AGEMA_signal_12583}), .clk (clk), .r ({Fresh[969], Fresh[968]}), .c ({new_AGEMA_signal_6434, SubBytesIns_Inst_Sbox_9_M48}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M49_U1 ( .a ({new_AGEMA_signal_6431, SubBytesIns_Inst_Sbox_9_M43}), .b ({new_AGEMA_signal_12592, new_AGEMA_signal_12589}), .clk (clk), .r ({Fresh[971], Fresh[970]}), .c ({new_AGEMA_signal_6671, SubBytesIns_Inst_Sbox_9_M49}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M50_U1 ( .a ({new_AGEMA_signal_6246, SubBytesIns_Inst_Sbox_9_M38}), .b ({new_AGEMA_signal_12598, new_AGEMA_signal_12595}), .clk (clk), .r ({Fresh[973], Fresh[972]}), .c ({new_AGEMA_signal_6435, SubBytesIns_Inst_Sbox_9_M50}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M51_U1 ( .a ({new_AGEMA_signal_6245, SubBytesIns_Inst_Sbox_9_M37}), .b ({new_AGEMA_signal_12604, new_AGEMA_signal_12601}), .clk (clk), .r ({Fresh[975], Fresh[974]}), .c ({new_AGEMA_signal_6436, SubBytesIns_Inst_Sbox_9_M51}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M52_U1 ( .a ({new_AGEMA_signal_6430, SubBytesIns_Inst_Sbox_9_M42}), .b ({new_AGEMA_signal_12610, new_AGEMA_signal_12607}), .clk (clk), .r ({Fresh[977], Fresh[976]}), .c ({new_AGEMA_signal_6672, SubBytesIns_Inst_Sbox_9_M52}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M53_U1 ( .a ({new_AGEMA_signal_6669, SubBytesIns_Inst_Sbox_9_M45}), .b ({new_AGEMA_signal_12616, new_AGEMA_signal_12613}), .clk (clk), .r ({Fresh[979], Fresh[978]}), .c ({new_AGEMA_signal_6883, SubBytesIns_Inst_Sbox_9_M53}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M54_U1 ( .a ({new_AGEMA_signal_6429, SubBytesIns_Inst_Sbox_9_M41}), .b ({new_AGEMA_signal_12622, new_AGEMA_signal_12619}), .clk (clk), .r ({Fresh[981], Fresh[980]}), .c ({new_AGEMA_signal_6673, SubBytesIns_Inst_Sbox_9_M54}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M55_U1 ( .a ({new_AGEMA_signal_6432, SubBytesIns_Inst_Sbox_9_M44}), .b ({new_AGEMA_signal_12628, new_AGEMA_signal_12625}), .clk (clk), .r ({Fresh[983], Fresh[982]}), .c ({new_AGEMA_signal_6674, SubBytesIns_Inst_Sbox_9_M55}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M56_U1 ( .a ({new_AGEMA_signal_6248, SubBytesIns_Inst_Sbox_9_M40}), .b ({new_AGEMA_signal_12634, new_AGEMA_signal_12631}), .clk (clk), .r ({Fresh[985], Fresh[984]}), .c ({new_AGEMA_signal_6437, SubBytesIns_Inst_Sbox_9_M56}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M57_U1 ( .a ({new_AGEMA_signal_6247, SubBytesIns_Inst_Sbox_9_M39}), .b ({new_AGEMA_signal_12640, new_AGEMA_signal_12637}), .clk (clk), .r ({Fresh[987], Fresh[986]}), .c ({new_AGEMA_signal_6438, SubBytesIns_Inst_Sbox_9_M57}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M58_U1 ( .a ({new_AGEMA_signal_6431, SubBytesIns_Inst_Sbox_9_M43}), .b ({new_AGEMA_signal_12646, new_AGEMA_signal_12643}), .clk (clk), .r ({Fresh[989], Fresh[988]}), .c ({new_AGEMA_signal_6675, SubBytesIns_Inst_Sbox_9_M58}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M59_U1 ( .a ({new_AGEMA_signal_6246, SubBytesIns_Inst_Sbox_9_M38}), .b ({new_AGEMA_signal_12652, new_AGEMA_signal_12649}), .clk (clk), .r ({Fresh[991], Fresh[990]}), .c ({new_AGEMA_signal_6439, SubBytesIns_Inst_Sbox_9_M59}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M60_U1 ( .a ({new_AGEMA_signal_6245, SubBytesIns_Inst_Sbox_9_M37}), .b ({new_AGEMA_signal_12658, new_AGEMA_signal_12655}), .clk (clk), .r ({Fresh[993], Fresh[992]}), .c ({new_AGEMA_signal_6440, SubBytesIns_Inst_Sbox_9_M60}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M61_U1 ( .a ({new_AGEMA_signal_6430, SubBytesIns_Inst_Sbox_9_M42}), .b ({new_AGEMA_signal_12664, new_AGEMA_signal_12661}), .clk (clk), .r ({Fresh[995], Fresh[994]}), .c ({new_AGEMA_signal_6676, SubBytesIns_Inst_Sbox_9_M61}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M62_U1 ( .a ({new_AGEMA_signal_6669, SubBytesIns_Inst_Sbox_9_M45}), .b ({new_AGEMA_signal_12670, new_AGEMA_signal_12667}), .clk (clk), .r ({Fresh[997], Fresh[996]}), .c ({new_AGEMA_signal_6884, SubBytesIns_Inst_Sbox_9_M62}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M63_U1 ( .a ({new_AGEMA_signal_6429, SubBytesIns_Inst_Sbox_9_M41}), .b ({new_AGEMA_signal_12676, new_AGEMA_signal_12673}), .clk (clk), .r ({Fresh[999], Fresh[998]}), .c ({new_AGEMA_signal_6677, SubBytesIns_Inst_Sbox_9_M63}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L0_U1 ( .a ({new_AGEMA_signal_6676, SubBytesIns_Inst_Sbox_9_M61}), .b ({new_AGEMA_signal_6884, SubBytesIns_Inst_Sbox_9_M62}), .c ({new_AGEMA_signal_7070, SubBytesIns_Inst_Sbox_9_L0}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L1_U1 ( .a ({new_AGEMA_signal_6435, SubBytesIns_Inst_Sbox_9_M50}), .b ({new_AGEMA_signal_6437, SubBytesIns_Inst_Sbox_9_M56}), .c ({new_AGEMA_signal_6678, SubBytesIns_Inst_Sbox_9_L1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L2_U1 ( .a ({new_AGEMA_signal_6670, SubBytesIns_Inst_Sbox_9_M46}), .b ({new_AGEMA_signal_6434, SubBytesIns_Inst_Sbox_9_M48}), .c ({new_AGEMA_signal_6885, SubBytesIns_Inst_Sbox_9_L2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L3_U1 ( .a ({new_AGEMA_signal_6433, SubBytesIns_Inst_Sbox_9_M47}), .b ({new_AGEMA_signal_6674, SubBytesIns_Inst_Sbox_9_M55}), .c ({new_AGEMA_signal_6886, SubBytesIns_Inst_Sbox_9_L3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L4_U1 ( .a ({new_AGEMA_signal_6673, SubBytesIns_Inst_Sbox_9_M54}), .b ({new_AGEMA_signal_6675, SubBytesIns_Inst_Sbox_9_M58}), .c ({new_AGEMA_signal_6887, SubBytesIns_Inst_Sbox_9_L4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L5_U1 ( .a ({new_AGEMA_signal_6671, SubBytesIns_Inst_Sbox_9_M49}), .b ({new_AGEMA_signal_6676, SubBytesIns_Inst_Sbox_9_M61}), .c ({new_AGEMA_signal_6888, SubBytesIns_Inst_Sbox_9_L5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L6_U1 ( .a ({new_AGEMA_signal_6884, SubBytesIns_Inst_Sbox_9_M62}), .b ({new_AGEMA_signal_6888, SubBytesIns_Inst_Sbox_9_L5}), .c ({new_AGEMA_signal_7071, SubBytesIns_Inst_Sbox_9_L6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L7_U1 ( .a ({new_AGEMA_signal_6670, SubBytesIns_Inst_Sbox_9_M46}), .b ({new_AGEMA_signal_6886, SubBytesIns_Inst_Sbox_9_L3}), .c ({new_AGEMA_signal_7072, SubBytesIns_Inst_Sbox_9_L7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L8_U1 ( .a ({new_AGEMA_signal_6436, SubBytesIns_Inst_Sbox_9_M51}), .b ({new_AGEMA_signal_6439, SubBytesIns_Inst_Sbox_9_M59}), .c ({new_AGEMA_signal_6679, SubBytesIns_Inst_Sbox_9_L8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L9_U1 ( .a ({new_AGEMA_signal_6672, SubBytesIns_Inst_Sbox_9_M52}), .b ({new_AGEMA_signal_6883, SubBytesIns_Inst_Sbox_9_M53}), .c ({new_AGEMA_signal_7073, SubBytesIns_Inst_Sbox_9_L9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L10_U1 ( .a ({new_AGEMA_signal_6883, SubBytesIns_Inst_Sbox_9_M53}), .b ({new_AGEMA_signal_6887, SubBytesIns_Inst_Sbox_9_L4}), .c ({new_AGEMA_signal_7074, SubBytesIns_Inst_Sbox_9_L10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L11_U1 ( .a ({new_AGEMA_signal_6440, SubBytesIns_Inst_Sbox_9_M60}), .b ({new_AGEMA_signal_6885, SubBytesIns_Inst_Sbox_9_L2}), .c ({new_AGEMA_signal_7075, SubBytesIns_Inst_Sbox_9_L11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L12_U1 ( .a ({new_AGEMA_signal_6434, SubBytesIns_Inst_Sbox_9_M48}), .b ({new_AGEMA_signal_6436, SubBytesIns_Inst_Sbox_9_M51}), .c ({new_AGEMA_signal_6680, SubBytesIns_Inst_Sbox_9_L12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L13_U1 ( .a ({new_AGEMA_signal_6435, SubBytesIns_Inst_Sbox_9_M50}), .b ({new_AGEMA_signal_7070, SubBytesIns_Inst_Sbox_9_L0}), .c ({new_AGEMA_signal_7276, SubBytesIns_Inst_Sbox_9_L13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L14_U1 ( .a ({new_AGEMA_signal_6672, SubBytesIns_Inst_Sbox_9_M52}), .b ({new_AGEMA_signal_6676, SubBytesIns_Inst_Sbox_9_M61}), .c ({new_AGEMA_signal_6889, SubBytesIns_Inst_Sbox_9_L14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L15_U1 ( .a ({new_AGEMA_signal_6674, SubBytesIns_Inst_Sbox_9_M55}), .b ({new_AGEMA_signal_6678, SubBytesIns_Inst_Sbox_9_L1}), .c ({new_AGEMA_signal_6890, SubBytesIns_Inst_Sbox_9_L15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L16_U1 ( .a ({new_AGEMA_signal_6437, SubBytesIns_Inst_Sbox_9_M56}), .b ({new_AGEMA_signal_7070, SubBytesIns_Inst_Sbox_9_L0}), .c ({new_AGEMA_signal_7277, SubBytesIns_Inst_Sbox_9_L16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L17_U1 ( .a ({new_AGEMA_signal_6438, SubBytesIns_Inst_Sbox_9_M57}), .b ({new_AGEMA_signal_6678, SubBytesIns_Inst_Sbox_9_L1}), .c ({new_AGEMA_signal_6891, SubBytesIns_Inst_Sbox_9_L17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L18_U1 ( .a ({new_AGEMA_signal_6675, SubBytesIns_Inst_Sbox_9_M58}), .b ({new_AGEMA_signal_6679, SubBytesIns_Inst_Sbox_9_L8}), .c ({new_AGEMA_signal_6892, SubBytesIns_Inst_Sbox_9_L18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L19_U1 ( .a ({new_AGEMA_signal_6677, SubBytesIns_Inst_Sbox_9_M63}), .b ({new_AGEMA_signal_6887, SubBytesIns_Inst_Sbox_9_L4}), .c ({new_AGEMA_signal_7076, SubBytesIns_Inst_Sbox_9_L19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L20_U1 ( .a ({new_AGEMA_signal_7070, SubBytesIns_Inst_Sbox_9_L0}), .b ({new_AGEMA_signal_6678, SubBytesIns_Inst_Sbox_9_L1}), .c ({new_AGEMA_signal_7278, SubBytesIns_Inst_Sbox_9_L20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L21_U1 ( .a ({new_AGEMA_signal_6678, SubBytesIns_Inst_Sbox_9_L1}), .b ({new_AGEMA_signal_7072, SubBytesIns_Inst_Sbox_9_L7}), .c ({new_AGEMA_signal_7279, SubBytesIns_Inst_Sbox_9_L21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L22_U1 ( .a ({new_AGEMA_signal_6886, SubBytesIns_Inst_Sbox_9_L3}), .b ({new_AGEMA_signal_6680, SubBytesIns_Inst_Sbox_9_L12}), .c ({new_AGEMA_signal_7077, SubBytesIns_Inst_Sbox_9_L22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L23_U1 ( .a ({new_AGEMA_signal_6892, SubBytesIns_Inst_Sbox_9_L18}), .b ({new_AGEMA_signal_6885, SubBytesIns_Inst_Sbox_9_L2}), .c ({new_AGEMA_signal_7078, SubBytesIns_Inst_Sbox_9_L23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L24_U1 ( .a ({new_AGEMA_signal_6890, SubBytesIns_Inst_Sbox_9_L15}), .b ({new_AGEMA_signal_7073, SubBytesIns_Inst_Sbox_9_L9}), .c ({new_AGEMA_signal_7280, SubBytesIns_Inst_Sbox_9_L24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L25_U1 ( .a ({new_AGEMA_signal_7071, SubBytesIns_Inst_Sbox_9_L6}), .b ({new_AGEMA_signal_7074, SubBytesIns_Inst_Sbox_9_L10}), .c ({new_AGEMA_signal_7281, SubBytesIns_Inst_Sbox_9_L25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L26_U1 ( .a ({new_AGEMA_signal_7072, SubBytesIns_Inst_Sbox_9_L7}), .b ({new_AGEMA_signal_7073, SubBytesIns_Inst_Sbox_9_L9}), .c ({new_AGEMA_signal_7282, SubBytesIns_Inst_Sbox_9_L26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L27_U1 ( .a ({new_AGEMA_signal_6679, SubBytesIns_Inst_Sbox_9_L8}), .b ({new_AGEMA_signal_7074, SubBytesIns_Inst_Sbox_9_L10}), .c ({new_AGEMA_signal_7283, SubBytesIns_Inst_Sbox_9_L27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L28_U1 ( .a ({new_AGEMA_signal_7075, SubBytesIns_Inst_Sbox_9_L11}), .b ({new_AGEMA_signal_6889, SubBytesIns_Inst_Sbox_9_L14}), .c ({new_AGEMA_signal_7284, SubBytesIns_Inst_Sbox_9_L28}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L29_U1 ( .a ({new_AGEMA_signal_7075, SubBytesIns_Inst_Sbox_9_L11}), .b ({new_AGEMA_signal_6891, SubBytesIns_Inst_Sbox_9_L17}), .c ({new_AGEMA_signal_7285, SubBytesIns_Inst_Sbox_9_L29}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_S0_U1 ( .a ({new_AGEMA_signal_7071, SubBytesIns_Inst_Sbox_9_L6}), .b ({new_AGEMA_signal_7280, SubBytesIns_Inst_Sbox_9_L24}), .c ({new_AGEMA_signal_7448, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_S1_U1 ( .a ({new_AGEMA_signal_7277, SubBytesIns_Inst_Sbox_9_L16}), .b ({new_AGEMA_signal_7282, SubBytesIns_Inst_Sbox_9_L26}), .c ({new_AGEMA_signal_7449, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_S2_U1 ( .a ({new_AGEMA_signal_7076, SubBytesIns_Inst_Sbox_9_L19}), .b ({new_AGEMA_signal_7284, SubBytesIns_Inst_Sbox_9_L28}), .c ({new_AGEMA_signal_7450, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_S3_U1 ( .a ({new_AGEMA_signal_7071, SubBytesIns_Inst_Sbox_9_L6}), .b ({new_AGEMA_signal_7279, SubBytesIns_Inst_Sbox_9_L21}), .c ({new_AGEMA_signal_7451, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_S4_U1 ( .a ({new_AGEMA_signal_7278, SubBytesIns_Inst_Sbox_9_L20}), .b ({new_AGEMA_signal_7077, SubBytesIns_Inst_Sbox_9_L22}), .c ({new_AGEMA_signal_7452, MixColumnsInput[11]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_S5_U1 ( .a ({new_AGEMA_signal_7281, SubBytesIns_Inst_Sbox_9_L25}), .b ({new_AGEMA_signal_7285, SubBytesIns_Inst_Sbox_9_L29}), .c ({new_AGEMA_signal_7453, MixColumnsInput[10]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_S6_U1 ( .a ({new_AGEMA_signal_7276, SubBytesIns_Inst_Sbox_9_L13}), .b ({new_AGEMA_signal_7283, SubBytesIns_Inst_Sbox_9_L27}), .c ({new_AGEMA_signal_7454, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_S7_U1 ( .a ({new_AGEMA_signal_7071, SubBytesIns_Inst_Sbox_9_L6}), .b ({new_AGEMA_signal_7078, SubBytesIns_Inst_Sbox_9_L23}), .c ({new_AGEMA_signal_7286, MixColumnsInput[8]}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M46_U1 ( .a ({new_AGEMA_signal_6444, SubBytesIns_Inst_Sbox_10_M44}), .b ({new_AGEMA_signal_12682, new_AGEMA_signal_12679}), .clk (clk), .r ({Fresh[1001], Fresh[1000]}), .c ({new_AGEMA_signal_6682, SubBytesIns_Inst_Sbox_10_M46}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M47_U1 ( .a ({new_AGEMA_signal_6252, SubBytesIns_Inst_Sbox_10_M40}), .b ({new_AGEMA_signal_12688, new_AGEMA_signal_12685}), .clk (clk), .r ({Fresh[1003], Fresh[1002]}), .c ({new_AGEMA_signal_6445, SubBytesIns_Inst_Sbox_10_M47}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M48_U1 ( .a ({new_AGEMA_signal_6251, SubBytesIns_Inst_Sbox_10_M39}), .b ({new_AGEMA_signal_12694, new_AGEMA_signal_12691}), .clk (clk), .r ({Fresh[1005], Fresh[1004]}), .c ({new_AGEMA_signal_6446, SubBytesIns_Inst_Sbox_10_M48}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M49_U1 ( .a ({new_AGEMA_signal_6443, SubBytesIns_Inst_Sbox_10_M43}), .b ({new_AGEMA_signal_12700, new_AGEMA_signal_12697}), .clk (clk), .r ({Fresh[1007], Fresh[1006]}), .c ({new_AGEMA_signal_6683, SubBytesIns_Inst_Sbox_10_M49}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M50_U1 ( .a ({new_AGEMA_signal_6250, SubBytesIns_Inst_Sbox_10_M38}), .b ({new_AGEMA_signal_12706, new_AGEMA_signal_12703}), .clk (clk), .r ({Fresh[1009], Fresh[1008]}), .c ({new_AGEMA_signal_6447, SubBytesIns_Inst_Sbox_10_M50}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M51_U1 ( .a ({new_AGEMA_signal_6249, SubBytesIns_Inst_Sbox_10_M37}), .b ({new_AGEMA_signal_12712, new_AGEMA_signal_12709}), .clk (clk), .r ({Fresh[1011], Fresh[1010]}), .c ({new_AGEMA_signal_6448, SubBytesIns_Inst_Sbox_10_M51}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M52_U1 ( .a ({new_AGEMA_signal_6442, SubBytesIns_Inst_Sbox_10_M42}), .b ({new_AGEMA_signal_12718, new_AGEMA_signal_12715}), .clk (clk), .r ({Fresh[1013], Fresh[1012]}), .c ({new_AGEMA_signal_6684, SubBytesIns_Inst_Sbox_10_M52}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M53_U1 ( .a ({new_AGEMA_signal_6681, SubBytesIns_Inst_Sbox_10_M45}), .b ({new_AGEMA_signal_12724, new_AGEMA_signal_12721}), .clk (clk), .r ({Fresh[1015], Fresh[1014]}), .c ({new_AGEMA_signal_6893, SubBytesIns_Inst_Sbox_10_M53}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M54_U1 ( .a ({new_AGEMA_signal_6441, SubBytesIns_Inst_Sbox_10_M41}), .b ({new_AGEMA_signal_12730, new_AGEMA_signal_12727}), .clk (clk), .r ({Fresh[1017], Fresh[1016]}), .c ({new_AGEMA_signal_6685, SubBytesIns_Inst_Sbox_10_M54}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M55_U1 ( .a ({new_AGEMA_signal_6444, SubBytesIns_Inst_Sbox_10_M44}), .b ({new_AGEMA_signal_12736, new_AGEMA_signal_12733}), .clk (clk), .r ({Fresh[1019], Fresh[1018]}), .c ({new_AGEMA_signal_6686, SubBytesIns_Inst_Sbox_10_M55}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M56_U1 ( .a ({new_AGEMA_signal_6252, SubBytesIns_Inst_Sbox_10_M40}), .b ({new_AGEMA_signal_12742, new_AGEMA_signal_12739}), .clk (clk), .r ({Fresh[1021], Fresh[1020]}), .c ({new_AGEMA_signal_6449, SubBytesIns_Inst_Sbox_10_M56}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M57_U1 ( .a ({new_AGEMA_signal_6251, SubBytesIns_Inst_Sbox_10_M39}), .b ({new_AGEMA_signal_12748, new_AGEMA_signal_12745}), .clk (clk), .r ({Fresh[1023], Fresh[1022]}), .c ({new_AGEMA_signal_6450, SubBytesIns_Inst_Sbox_10_M57}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M58_U1 ( .a ({new_AGEMA_signal_6443, SubBytesIns_Inst_Sbox_10_M43}), .b ({new_AGEMA_signal_12754, new_AGEMA_signal_12751}), .clk (clk), .r ({Fresh[1025], Fresh[1024]}), .c ({new_AGEMA_signal_6687, SubBytesIns_Inst_Sbox_10_M58}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M59_U1 ( .a ({new_AGEMA_signal_6250, SubBytesIns_Inst_Sbox_10_M38}), .b ({new_AGEMA_signal_12760, new_AGEMA_signal_12757}), .clk (clk), .r ({Fresh[1027], Fresh[1026]}), .c ({new_AGEMA_signal_6451, SubBytesIns_Inst_Sbox_10_M59}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M60_U1 ( .a ({new_AGEMA_signal_6249, SubBytesIns_Inst_Sbox_10_M37}), .b ({new_AGEMA_signal_12766, new_AGEMA_signal_12763}), .clk (clk), .r ({Fresh[1029], Fresh[1028]}), .c ({new_AGEMA_signal_6452, SubBytesIns_Inst_Sbox_10_M60}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M61_U1 ( .a ({new_AGEMA_signal_6442, SubBytesIns_Inst_Sbox_10_M42}), .b ({new_AGEMA_signal_12772, new_AGEMA_signal_12769}), .clk (clk), .r ({Fresh[1031], Fresh[1030]}), .c ({new_AGEMA_signal_6688, SubBytesIns_Inst_Sbox_10_M61}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M62_U1 ( .a ({new_AGEMA_signal_6681, SubBytesIns_Inst_Sbox_10_M45}), .b ({new_AGEMA_signal_12778, new_AGEMA_signal_12775}), .clk (clk), .r ({Fresh[1033], Fresh[1032]}), .c ({new_AGEMA_signal_6894, SubBytesIns_Inst_Sbox_10_M62}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M63_U1 ( .a ({new_AGEMA_signal_6441, SubBytesIns_Inst_Sbox_10_M41}), .b ({new_AGEMA_signal_12784, new_AGEMA_signal_12781}), .clk (clk), .r ({Fresh[1035], Fresh[1034]}), .c ({new_AGEMA_signal_6689, SubBytesIns_Inst_Sbox_10_M63}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L0_U1 ( .a ({new_AGEMA_signal_6688, SubBytesIns_Inst_Sbox_10_M61}), .b ({new_AGEMA_signal_6894, SubBytesIns_Inst_Sbox_10_M62}), .c ({new_AGEMA_signal_7079, SubBytesIns_Inst_Sbox_10_L0}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L1_U1 ( .a ({new_AGEMA_signal_6447, SubBytesIns_Inst_Sbox_10_M50}), .b ({new_AGEMA_signal_6449, SubBytesIns_Inst_Sbox_10_M56}), .c ({new_AGEMA_signal_6690, SubBytesIns_Inst_Sbox_10_L1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L2_U1 ( .a ({new_AGEMA_signal_6682, SubBytesIns_Inst_Sbox_10_M46}), .b ({new_AGEMA_signal_6446, SubBytesIns_Inst_Sbox_10_M48}), .c ({new_AGEMA_signal_6895, SubBytesIns_Inst_Sbox_10_L2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L3_U1 ( .a ({new_AGEMA_signal_6445, SubBytesIns_Inst_Sbox_10_M47}), .b ({new_AGEMA_signal_6686, SubBytesIns_Inst_Sbox_10_M55}), .c ({new_AGEMA_signal_6896, SubBytesIns_Inst_Sbox_10_L3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L4_U1 ( .a ({new_AGEMA_signal_6685, SubBytesIns_Inst_Sbox_10_M54}), .b ({new_AGEMA_signal_6687, SubBytesIns_Inst_Sbox_10_M58}), .c ({new_AGEMA_signal_6897, SubBytesIns_Inst_Sbox_10_L4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L5_U1 ( .a ({new_AGEMA_signal_6683, SubBytesIns_Inst_Sbox_10_M49}), .b ({new_AGEMA_signal_6688, SubBytesIns_Inst_Sbox_10_M61}), .c ({new_AGEMA_signal_6898, SubBytesIns_Inst_Sbox_10_L5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L6_U1 ( .a ({new_AGEMA_signal_6894, SubBytesIns_Inst_Sbox_10_M62}), .b ({new_AGEMA_signal_6898, SubBytesIns_Inst_Sbox_10_L5}), .c ({new_AGEMA_signal_7080, SubBytesIns_Inst_Sbox_10_L6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L7_U1 ( .a ({new_AGEMA_signal_6682, SubBytesIns_Inst_Sbox_10_M46}), .b ({new_AGEMA_signal_6896, SubBytesIns_Inst_Sbox_10_L3}), .c ({new_AGEMA_signal_7081, SubBytesIns_Inst_Sbox_10_L7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L8_U1 ( .a ({new_AGEMA_signal_6448, SubBytesIns_Inst_Sbox_10_M51}), .b ({new_AGEMA_signal_6451, SubBytesIns_Inst_Sbox_10_M59}), .c ({new_AGEMA_signal_6691, SubBytesIns_Inst_Sbox_10_L8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L9_U1 ( .a ({new_AGEMA_signal_6684, SubBytesIns_Inst_Sbox_10_M52}), .b ({new_AGEMA_signal_6893, SubBytesIns_Inst_Sbox_10_M53}), .c ({new_AGEMA_signal_7082, SubBytesIns_Inst_Sbox_10_L9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L10_U1 ( .a ({new_AGEMA_signal_6893, SubBytesIns_Inst_Sbox_10_M53}), .b ({new_AGEMA_signal_6897, SubBytesIns_Inst_Sbox_10_L4}), .c ({new_AGEMA_signal_7083, SubBytesIns_Inst_Sbox_10_L10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L11_U1 ( .a ({new_AGEMA_signal_6452, SubBytesIns_Inst_Sbox_10_M60}), .b ({new_AGEMA_signal_6895, SubBytesIns_Inst_Sbox_10_L2}), .c ({new_AGEMA_signal_7084, SubBytesIns_Inst_Sbox_10_L11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L12_U1 ( .a ({new_AGEMA_signal_6446, SubBytesIns_Inst_Sbox_10_M48}), .b ({new_AGEMA_signal_6448, SubBytesIns_Inst_Sbox_10_M51}), .c ({new_AGEMA_signal_6692, SubBytesIns_Inst_Sbox_10_L12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L13_U1 ( .a ({new_AGEMA_signal_6447, SubBytesIns_Inst_Sbox_10_M50}), .b ({new_AGEMA_signal_7079, SubBytesIns_Inst_Sbox_10_L0}), .c ({new_AGEMA_signal_7287, SubBytesIns_Inst_Sbox_10_L13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L14_U1 ( .a ({new_AGEMA_signal_6684, SubBytesIns_Inst_Sbox_10_M52}), .b ({new_AGEMA_signal_6688, SubBytesIns_Inst_Sbox_10_M61}), .c ({new_AGEMA_signal_6899, SubBytesIns_Inst_Sbox_10_L14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L15_U1 ( .a ({new_AGEMA_signal_6686, SubBytesIns_Inst_Sbox_10_M55}), .b ({new_AGEMA_signal_6690, SubBytesIns_Inst_Sbox_10_L1}), .c ({new_AGEMA_signal_6900, SubBytesIns_Inst_Sbox_10_L15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L16_U1 ( .a ({new_AGEMA_signal_6449, SubBytesIns_Inst_Sbox_10_M56}), .b ({new_AGEMA_signal_7079, SubBytesIns_Inst_Sbox_10_L0}), .c ({new_AGEMA_signal_7288, SubBytesIns_Inst_Sbox_10_L16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L17_U1 ( .a ({new_AGEMA_signal_6450, SubBytesIns_Inst_Sbox_10_M57}), .b ({new_AGEMA_signal_6690, SubBytesIns_Inst_Sbox_10_L1}), .c ({new_AGEMA_signal_6901, SubBytesIns_Inst_Sbox_10_L17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L18_U1 ( .a ({new_AGEMA_signal_6687, SubBytesIns_Inst_Sbox_10_M58}), .b ({new_AGEMA_signal_6691, SubBytesIns_Inst_Sbox_10_L8}), .c ({new_AGEMA_signal_6902, SubBytesIns_Inst_Sbox_10_L18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L19_U1 ( .a ({new_AGEMA_signal_6689, SubBytesIns_Inst_Sbox_10_M63}), .b ({new_AGEMA_signal_6897, SubBytesIns_Inst_Sbox_10_L4}), .c ({new_AGEMA_signal_7085, SubBytesIns_Inst_Sbox_10_L19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L20_U1 ( .a ({new_AGEMA_signal_7079, SubBytesIns_Inst_Sbox_10_L0}), .b ({new_AGEMA_signal_6690, SubBytesIns_Inst_Sbox_10_L1}), .c ({new_AGEMA_signal_7289, SubBytesIns_Inst_Sbox_10_L20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L21_U1 ( .a ({new_AGEMA_signal_6690, SubBytesIns_Inst_Sbox_10_L1}), .b ({new_AGEMA_signal_7081, SubBytesIns_Inst_Sbox_10_L7}), .c ({new_AGEMA_signal_7290, SubBytesIns_Inst_Sbox_10_L21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L22_U1 ( .a ({new_AGEMA_signal_6896, SubBytesIns_Inst_Sbox_10_L3}), .b ({new_AGEMA_signal_6692, SubBytesIns_Inst_Sbox_10_L12}), .c ({new_AGEMA_signal_7086, SubBytesIns_Inst_Sbox_10_L22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L23_U1 ( .a ({new_AGEMA_signal_6902, SubBytesIns_Inst_Sbox_10_L18}), .b ({new_AGEMA_signal_6895, SubBytesIns_Inst_Sbox_10_L2}), .c ({new_AGEMA_signal_7087, SubBytesIns_Inst_Sbox_10_L23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L24_U1 ( .a ({new_AGEMA_signal_6900, SubBytesIns_Inst_Sbox_10_L15}), .b ({new_AGEMA_signal_7082, SubBytesIns_Inst_Sbox_10_L9}), .c ({new_AGEMA_signal_7291, SubBytesIns_Inst_Sbox_10_L24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L25_U1 ( .a ({new_AGEMA_signal_7080, SubBytesIns_Inst_Sbox_10_L6}), .b ({new_AGEMA_signal_7083, SubBytesIns_Inst_Sbox_10_L10}), .c ({new_AGEMA_signal_7292, SubBytesIns_Inst_Sbox_10_L25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L26_U1 ( .a ({new_AGEMA_signal_7081, SubBytesIns_Inst_Sbox_10_L7}), .b ({new_AGEMA_signal_7082, SubBytesIns_Inst_Sbox_10_L9}), .c ({new_AGEMA_signal_7293, SubBytesIns_Inst_Sbox_10_L26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L27_U1 ( .a ({new_AGEMA_signal_6691, SubBytesIns_Inst_Sbox_10_L8}), .b ({new_AGEMA_signal_7083, SubBytesIns_Inst_Sbox_10_L10}), .c ({new_AGEMA_signal_7294, SubBytesIns_Inst_Sbox_10_L27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L28_U1 ( .a ({new_AGEMA_signal_7084, SubBytesIns_Inst_Sbox_10_L11}), .b ({new_AGEMA_signal_6899, SubBytesIns_Inst_Sbox_10_L14}), .c ({new_AGEMA_signal_7295, SubBytesIns_Inst_Sbox_10_L28}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L29_U1 ( .a ({new_AGEMA_signal_7084, SubBytesIns_Inst_Sbox_10_L11}), .b ({new_AGEMA_signal_6901, SubBytesIns_Inst_Sbox_10_L17}), .c ({new_AGEMA_signal_7296, SubBytesIns_Inst_Sbox_10_L29}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_S0_U1 ( .a ({new_AGEMA_signal_7080, SubBytesIns_Inst_Sbox_10_L6}), .b ({new_AGEMA_signal_7291, SubBytesIns_Inst_Sbox_10_L24}), .c ({new_AGEMA_signal_7455, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_S1_U1 ( .a ({new_AGEMA_signal_7288, SubBytesIns_Inst_Sbox_10_L16}), .b ({new_AGEMA_signal_7293, SubBytesIns_Inst_Sbox_10_L26}), .c ({new_AGEMA_signal_7456, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_S2_U1 ( .a ({new_AGEMA_signal_7085, SubBytesIns_Inst_Sbox_10_L19}), .b ({new_AGEMA_signal_7295, SubBytesIns_Inst_Sbox_10_L28}), .c ({new_AGEMA_signal_7457, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_S3_U1 ( .a ({new_AGEMA_signal_7080, SubBytesIns_Inst_Sbox_10_L6}), .b ({new_AGEMA_signal_7290, SubBytesIns_Inst_Sbox_10_L21}), .c ({new_AGEMA_signal_7458, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_S4_U1 ( .a ({new_AGEMA_signal_7289, SubBytesIns_Inst_Sbox_10_L20}), .b ({new_AGEMA_signal_7086, SubBytesIns_Inst_Sbox_10_L22}), .c ({new_AGEMA_signal_7459, MixColumnsInput[115]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_S5_U1 ( .a ({new_AGEMA_signal_7292, SubBytesIns_Inst_Sbox_10_L25}), .b ({new_AGEMA_signal_7296, SubBytesIns_Inst_Sbox_10_L29}), .c ({new_AGEMA_signal_7460, MixColumnsInput[114]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_S6_U1 ( .a ({new_AGEMA_signal_7287, SubBytesIns_Inst_Sbox_10_L13}), .b ({new_AGEMA_signal_7294, SubBytesIns_Inst_Sbox_10_L27}), .c ({new_AGEMA_signal_7461, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_S7_U1 ( .a ({new_AGEMA_signal_7080, SubBytesIns_Inst_Sbox_10_L6}), .b ({new_AGEMA_signal_7087, SubBytesIns_Inst_Sbox_10_L23}), .c ({new_AGEMA_signal_7297, MixColumnsInput[112]}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M46_U1 ( .a ({new_AGEMA_signal_6456, SubBytesIns_Inst_Sbox_11_M44}), .b ({new_AGEMA_signal_12790, new_AGEMA_signal_12787}), .clk (clk), .r ({Fresh[1037], Fresh[1036]}), .c ({new_AGEMA_signal_6694, SubBytesIns_Inst_Sbox_11_M46}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M47_U1 ( .a ({new_AGEMA_signal_6256, SubBytesIns_Inst_Sbox_11_M40}), .b ({new_AGEMA_signal_12796, new_AGEMA_signal_12793}), .clk (clk), .r ({Fresh[1039], Fresh[1038]}), .c ({new_AGEMA_signal_6457, SubBytesIns_Inst_Sbox_11_M47}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M48_U1 ( .a ({new_AGEMA_signal_6255, SubBytesIns_Inst_Sbox_11_M39}), .b ({new_AGEMA_signal_12802, new_AGEMA_signal_12799}), .clk (clk), .r ({Fresh[1041], Fresh[1040]}), .c ({new_AGEMA_signal_6458, SubBytesIns_Inst_Sbox_11_M48}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M49_U1 ( .a ({new_AGEMA_signal_6455, SubBytesIns_Inst_Sbox_11_M43}), .b ({new_AGEMA_signal_12808, new_AGEMA_signal_12805}), .clk (clk), .r ({Fresh[1043], Fresh[1042]}), .c ({new_AGEMA_signal_6695, SubBytesIns_Inst_Sbox_11_M49}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M50_U1 ( .a ({new_AGEMA_signal_6254, SubBytesIns_Inst_Sbox_11_M38}), .b ({new_AGEMA_signal_12814, new_AGEMA_signal_12811}), .clk (clk), .r ({Fresh[1045], Fresh[1044]}), .c ({new_AGEMA_signal_6459, SubBytesIns_Inst_Sbox_11_M50}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M51_U1 ( .a ({new_AGEMA_signal_6253, SubBytesIns_Inst_Sbox_11_M37}), .b ({new_AGEMA_signal_12820, new_AGEMA_signal_12817}), .clk (clk), .r ({Fresh[1047], Fresh[1046]}), .c ({new_AGEMA_signal_6460, SubBytesIns_Inst_Sbox_11_M51}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M52_U1 ( .a ({new_AGEMA_signal_6454, SubBytesIns_Inst_Sbox_11_M42}), .b ({new_AGEMA_signal_12826, new_AGEMA_signal_12823}), .clk (clk), .r ({Fresh[1049], Fresh[1048]}), .c ({new_AGEMA_signal_6696, SubBytesIns_Inst_Sbox_11_M52}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M53_U1 ( .a ({new_AGEMA_signal_6693, SubBytesIns_Inst_Sbox_11_M45}), .b ({new_AGEMA_signal_12832, new_AGEMA_signal_12829}), .clk (clk), .r ({Fresh[1051], Fresh[1050]}), .c ({new_AGEMA_signal_6903, SubBytesIns_Inst_Sbox_11_M53}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M54_U1 ( .a ({new_AGEMA_signal_6453, SubBytesIns_Inst_Sbox_11_M41}), .b ({new_AGEMA_signal_12838, new_AGEMA_signal_12835}), .clk (clk), .r ({Fresh[1053], Fresh[1052]}), .c ({new_AGEMA_signal_6697, SubBytesIns_Inst_Sbox_11_M54}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M55_U1 ( .a ({new_AGEMA_signal_6456, SubBytesIns_Inst_Sbox_11_M44}), .b ({new_AGEMA_signal_12844, new_AGEMA_signal_12841}), .clk (clk), .r ({Fresh[1055], Fresh[1054]}), .c ({new_AGEMA_signal_6698, SubBytesIns_Inst_Sbox_11_M55}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M56_U1 ( .a ({new_AGEMA_signal_6256, SubBytesIns_Inst_Sbox_11_M40}), .b ({new_AGEMA_signal_12850, new_AGEMA_signal_12847}), .clk (clk), .r ({Fresh[1057], Fresh[1056]}), .c ({new_AGEMA_signal_6461, SubBytesIns_Inst_Sbox_11_M56}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M57_U1 ( .a ({new_AGEMA_signal_6255, SubBytesIns_Inst_Sbox_11_M39}), .b ({new_AGEMA_signal_12856, new_AGEMA_signal_12853}), .clk (clk), .r ({Fresh[1059], Fresh[1058]}), .c ({new_AGEMA_signal_6462, SubBytesIns_Inst_Sbox_11_M57}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M58_U1 ( .a ({new_AGEMA_signal_6455, SubBytesIns_Inst_Sbox_11_M43}), .b ({new_AGEMA_signal_12862, new_AGEMA_signal_12859}), .clk (clk), .r ({Fresh[1061], Fresh[1060]}), .c ({new_AGEMA_signal_6699, SubBytesIns_Inst_Sbox_11_M58}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M59_U1 ( .a ({new_AGEMA_signal_6254, SubBytesIns_Inst_Sbox_11_M38}), .b ({new_AGEMA_signal_12868, new_AGEMA_signal_12865}), .clk (clk), .r ({Fresh[1063], Fresh[1062]}), .c ({new_AGEMA_signal_6463, SubBytesIns_Inst_Sbox_11_M59}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M60_U1 ( .a ({new_AGEMA_signal_6253, SubBytesIns_Inst_Sbox_11_M37}), .b ({new_AGEMA_signal_12874, new_AGEMA_signal_12871}), .clk (clk), .r ({Fresh[1065], Fresh[1064]}), .c ({new_AGEMA_signal_6464, SubBytesIns_Inst_Sbox_11_M60}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M61_U1 ( .a ({new_AGEMA_signal_6454, SubBytesIns_Inst_Sbox_11_M42}), .b ({new_AGEMA_signal_12880, new_AGEMA_signal_12877}), .clk (clk), .r ({Fresh[1067], Fresh[1066]}), .c ({new_AGEMA_signal_6700, SubBytesIns_Inst_Sbox_11_M61}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M62_U1 ( .a ({new_AGEMA_signal_6693, SubBytesIns_Inst_Sbox_11_M45}), .b ({new_AGEMA_signal_12886, new_AGEMA_signal_12883}), .clk (clk), .r ({Fresh[1069], Fresh[1068]}), .c ({new_AGEMA_signal_6904, SubBytesIns_Inst_Sbox_11_M62}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M63_U1 ( .a ({new_AGEMA_signal_6453, SubBytesIns_Inst_Sbox_11_M41}), .b ({new_AGEMA_signal_12892, new_AGEMA_signal_12889}), .clk (clk), .r ({Fresh[1071], Fresh[1070]}), .c ({new_AGEMA_signal_6701, SubBytesIns_Inst_Sbox_11_M63}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L0_U1 ( .a ({new_AGEMA_signal_6700, SubBytesIns_Inst_Sbox_11_M61}), .b ({new_AGEMA_signal_6904, SubBytesIns_Inst_Sbox_11_M62}), .c ({new_AGEMA_signal_7088, SubBytesIns_Inst_Sbox_11_L0}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L1_U1 ( .a ({new_AGEMA_signal_6459, SubBytesIns_Inst_Sbox_11_M50}), .b ({new_AGEMA_signal_6461, SubBytesIns_Inst_Sbox_11_M56}), .c ({new_AGEMA_signal_6702, SubBytesIns_Inst_Sbox_11_L1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L2_U1 ( .a ({new_AGEMA_signal_6694, SubBytesIns_Inst_Sbox_11_M46}), .b ({new_AGEMA_signal_6458, SubBytesIns_Inst_Sbox_11_M48}), .c ({new_AGEMA_signal_6905, SubBytesIns_Inst_Sbox_11_L2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L3_U1 ( .a ({new_AGEMA_signal_6457, SubBytesIns_Inst_Sbox_11_M47}), .b ({new_AGEMA_signal_6698, SubBytesIns_Inst_Sbox_11_M55}), .c ({new_AGEMA_signal_6906, SubBytesIns_Inst_Sbox_11_L3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L4_U1 ( .a ({new_AGEMA_signal_6697, SubBytesIns_Inst_Sbox_11_M54}), .b ({new_AGEMA_signal_6699, SubBytesIns_Inst_Sbox_11_M58}), .c ({new_AGEMA_signal_6907, SubBytesIns_Inst_Sbox_11_L4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L5_U1 ( .a ({new_AGEMA_signal_6695, SubBytesIns_Inst_Sbox_11_M49}), .b ({new_AGEMA_signal_6700, SubBytesIns_Inst_Sbox_11_M61}), .c ({new_AGEMA_signal_6908, SubBytesIns_Inst_Sbox_11_L5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L6_U1 ( .a ({new_AGEMA_signal_6904, SubBytesIns_Inst_Sbox_11_M62}), .b ({new_AGEMA_signal_6908, SubBytesIns_Inst_Sbox_11_L5}), .c ({new_AGEMA_signal_7089, SubBytesIns_Inst_Sbox_11_L6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L7_U1 ( .a ({new_AGEMA_signal_6694, SubBytesIns_Inst_Sbox_11_M46}), .b ({new_AGEMA_signal_6906, SubBytesIns_Inst_Sbox_11_L3}), .c ({new_AGEMA_signal_7090, SubBytesIns_Inst_Sbox_11_L7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L8_U1 ( .a ({new_AGEMA_signal_6460, SubBytesIns_Inst_Sbox_11_M51}), .b ({new_AGEMA_signal_6463, SubBytesIns_Inst_Sbox_11_M59}), .c ({new_AGEMA_signal_6703, SubBytesIns_Inst_Sbox_11_L8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L9_U1 ( .a ({new_AGEMA_signal_6696, SubBytesIns_Inst_Sbox_11_M52}), .b ({new_AGEMA_signal_6903, SubBytesIns_Inst_Sbox_11_M53}), .c ({new_AGEMA_signal_7091, SubBytesIns_Inst_Sbox_11_L9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L10_U1 ( .a ({new_AGEMA_signal_6903, SubBytesIns_Inst_Sbox_11_M53}), .b ({new_AGEMA_signal_6907, SubBytesIns_Inst_Sbox_11_L4}), .c ({new_AGEMA_signal_7092, SubBytesIns_Inst_Sbox_11_L10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L11_U1 ( .a ({new_AGEMA_signal_6464, SubBytesIns_Inst_Sbox_11_M60}), .b ({new_AGEMA_signal_6905, SubBytesIns_Inst_Sbox_11_L2}), .c ({new_AGEMA_signal_7093, SubBytesIns_Inst_Sbox_11_L11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L12_U1 ( .a ({new_AGEMA_signal_6458, SubBytesIns_Inst_Sbox_11_M48}), .b ({new_AGEMA_signal_6460, SubBytesIns_Inst_Sbox_11_M51}), .c ({new_AGEMA_signal_6704, SubBytesIns_Inst_Sbox_11_L12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L13_U1 ( .a ({new_AGEMA_signal_6459, SubBytesIns_Inst_Sbox_11_M50}), .b ({new_AGEMA_signal_7088, SubBytesIns_Inst_Sbox_11_L0}), .c ({new_AGEMA_signal_7298, SubBytesIns_Inst_Sbox_11_L13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L14_U1 ( .a ({new_AGEMA_signal_6696, SubBytesIns_Inst_Sbox_11_M52}), .b ({new_AGEMA_signal_6700, SubBytesIns_Inst_Sbox_11_M61}), .c ({new_AGEMA_signal_6909, SubBytesIns_Inst_Sbox_11_L14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L15_U1 ( .a ({new_AGEMA_signal_6698, SubBytesIns_Inst_Sbox_11_M55}), .b ({new_AGEMA_signal_6702, SubBytesIns_Inst_Sbox_11_L1}), .c ({new_AGEMA_signal_6910, SubBytesIns_Inst_Sbox_11_L15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L16_U1 ( .a ({new_AGEMA_signal_6461, SubBytesIns_Inst_Sbox_11_M56}), .b ({new_AGEMA_signal_7088, SubBytesIns_Inst_Sbox_11_L0}), .c ({new_AGEMA_signal_7299, SubBytesIns_Inst_Sbox_11_L16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L17_U1 ( .a ({new_AGEMA_signal_6462, SubBytesIns_Inst_Sbox_11_M57}), .b ({new_AGEMA_signal_6702, SubBytesIns_Inst_Sbox_11_L1}), .c ({new_AGEMA_signal_6911, SubBytesIns_Inst_Sbox_11_L17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L18_U1 ( .a ({new_AGEMA_signal_6699, SubBytesIns_Inst_Sbox_11_M58}), .b ({new_AGEMA_signal_6703, SubBytesIns_Inst_Sbox_11_L8}), .c ({new_AGEMA_signal_6912, SubBytesIns_Inst_Sbox_11_L18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L19_U1 ( .a ({new_AGEMA_signal_6701, SubBytesIns_Inst_Sbox_11_M63}), .b ({new_AGEMA_signal_6907, SubBytesIns_Inst_Sbox_11_L4}), .c ({new_AGEMA_signal_7094, SubBytesIns_Inst_Sbox_11_L19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L20_U1 ( .a ({new_AGEMA_signal_7088, SubBytesIns_Inst_Sbox_11_L0}), .b ({new_AGEMA_signal_6702, SubBytesIns_Inst_Sbox_11_L1}), .c ({new_AGEMA_signal_7300, SubBytesIns_Inst_Sbox_11_L20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L21_U1 ( .a ({new_AGEMA_signal_6702, SubBytesIns_Inst_Sbox_11_L1}), .b ({new_AGEMA_signal_7090, SubBytesIns_Inst_Sbox_11_L7}), .c ({new_AGEMA_signal_7301, SubBytesIns_Inst_Sbox_11_L21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L22_U1 ( .a ({new_AGEMA_signal_6906, SubBytesIns_Inst_Sbox_11_L3}), .b ({new_AGEMA_signal_6704, SubBytesIns_Inst_Sbox_11_L12}), .c ({new_AGEMA_signal_7095, SubBytesIns_Inst_Sbox_11_L22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L23_U1 ( .a ({new_AGEMA_signal_6912, SubBytesIns_Inst_Sbox_11_L18}), .b ({new_AGEMA_signal_6905, SubBytesIns_Inst_Sbox_11_L2}), .c ({new_AGEMA_signal_7096, SubBytesIns_Inst_Sbox_11_L23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L24_U1 ( .a ({new_AGEMA_signal_6910, SubBytesIns_Inst_Sbox_11_L15}), .b ({new_AGEMA_signal_7091, SubBytesIns_Inst_Sbox_11_L9}), .c ({new_AGEMA_signal_7302, SubBytesIns_Inst_Sbox_11_L24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L25_U1 ( .a ({new_AGEMA_signal_7089, SubBytesIns_Inst_Sbox_11_L6}), .b ({new_AGEMA_signal_7092, SubBytesIns_Inst_Sbox_11_L10}), .c ({new_AGEMA_signal_7303, SubBytesIns_Inst_Sbox_11_L25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L26_U1 ( .a ({new_AGEMA_signal_7090, SubBytesIns_Inst_Sbox_11_L7}), .b ({new_AGEMA_signal_7091, SubBytesIns_Inst_Sbox_11_L9}), .c ({new_AGEMA_signal_7304, SubBytesIns_Inst_Sbox_11_L26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L27_U1 ( .a ({new_AGEMA_signal_6703, SubBytesIns_Inst_Sbox_11_L8}), .b ({new_AGEMA_signal_7092, SubBytesIns_Inst_Sbox_11_L10}), .c ({new_AGEMA_signal_7305, SubBytesIns_Inst_Sbox_11_L27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L28_U1 ( .a ({new_AGEMA_signal_7093, SubBytesIns_Inst_Sbox_11_L11}), .b ({new_AGEMA_signal_6909, SubBytesIns_Inst_Sbox_11_L14}), .c ({new_AGEMA_signal_7306, SubBytesIns_Inst_Sbox_11_L28}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L29_U1 ( .a ({new_AGEMA_signal_7093, SubBytesIns_Inst_Sbox_11_L11}), .b ({new_AGEMA_signal_6911, SubBytesIns_Inst_Sbox_11_L17}), .c ({new_AGEMA_signal_7307, SubBytesIns_Inst_Sbox_11_L29}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_S0_U1 ( .a ({new_AGEMA_signal_7089, SubBytesIns_Inst_Sbox_11_L6}), .b ({new_AGEMA_signal_7302, SubBytesIns_Inst_Sbox_11_L24}), .c ({new_AGEMA_signal_7462, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_S1_U1 ( .a ({new_AGEMA_signal_7299, SubBytesIns_Inst_Sbox_11_L16}), .b ({new_AGEMA_signal_7304, SubBytesIns_Inst_Sbox_11_L26}), .c ({new_AGEMA_signal_7463, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_S2_U1 ( .a ({new_AGEMA_signal_7094, SubBytesIns_Inst_Sbox_11_L19}), .b ({new_AGEMA_signal_7306, SubBytesIns_Inst_Sbox_11_L28}), .c ({new_AGEMA_signal_7464, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_S3_U1 ( .a ({new_AGEMA_signal_7089, SubBytesIns_Inst_Sbox_11_L6}), .b ({new_AGEMA_signal_7301, SubBytesIns_Inst_Sbox_11_L21}), .c ({new_AGEMA_signal_7465, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_S4_U1 ( .a ({new_AGEMA_signal_7300, SubBytesIns_Inst_Sbox_11_L20}), .b ({new_AGEMA_signal_7095, SubBytesIns_Inst_Sbox_11_L22}), .c ({new_AGEMA_signal_7466, MixColumnsInput[91]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_S5_U1 ( .a ({new_AGEMA_signal_7303, SubBytesIns_Inst_Sbox_11_L25}), .b ({new_AGEMA_signal_7307, SubBytesIns_Inst_Sbox_11_L29}), .c ({new_AGEMA_signal_7467, MixColumnsInput[90]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_S6_U1 ( .a ({new_AGEMA_signal_7298, SubBytesIns_Inst_Sbox_11_L13}), .b ({new_AGEMA_signal_7305, SubBytesIns_Inst_Sbox_11_L27}), .c ({new_AGEMA_signal_7468, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_S7_U1 ( .a ({new_AGEMA_signal_7089, SubBytesIns_Inst_Sbox_11_L6}), .b ({new_AGEMA_signal_7096, SubBytesIns_Inst_Sbox_11_L23}), .c ({new_AGEMA_signal_7308, MixColumnsInput[88]}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M46_U1 ( .a ({new_AGEMA_signal_6468, SubBytesIns_Inst_Sbox_12_M44}), .b ({new_AGEMA_signal_12898, new_AGEMA_signal_12895}), .clk (clk), .r ({Fresh[1073], Fresh[1072]}), .c ({new_AGEMA_signal_6706, SubBytesIns_Inst_Sbox_12_M46}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M47_U1 ( .a ({new_AGEMA_signal_6260, SubBytesIns_Inst_Sbox_12_M40}), .b ({new_AGEMA_signal_12904, new_AGEMA_signal_12901}), .clk (clk), .r ({Fresh[1075], Fresh[1074]}), .c ({new_AGEMA_signal_6469, SubBytesIns_Inst_Sbox_12_M47}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M48_U1 ( .a ({new_AGEMA_signal_6259, SubBytesIns_Inst_Sbox_12_M39}), .b ({new_AGEMA_signal_12910, new_AGEMA_signal_12907}), .clk (clk), .r ({Fresh[1077], Fresh[1076]}), .c ({new_AGEMA_signal_6470, SubBytesIns_Inst_Sbox_12_M48}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M49_U1 ( .a ({new_AGEMA_signal_6467, SubBytesIns_Inst_Sbox_12_M43}), .b ({new_AGEMA_signal_12916, new_AGEMA_signal_12913}), .clk (clk), .r ({Fresh[1079], Fresh[1078]}), .c ({new_AGEMA_signal_6707, SubBytesIns_Inst_Sbox_12_M49}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M50_U1 ( .a ({new_AGEMA_signal_6258, SubBytesIns_Inst_Sbox_12_M38}), .b ({new_AGEMA_signal_12922, new_AGEMA_signal_12919}), .clk (clk), .r ({Fresh[1081], Fresh[1080]}), .c ({new_AGEMA_signal_6471, SubBytesIns_Inst_Sbox_12_M50}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M51_U1 ( .a ({new_AGEMA_signal_6257, SubBytesIns_Inst_Sbox_12_M37}), .b ({new_AGEMA_signal_12928, new_AGEMA_signal_12925}), .clk (clk), .r ({Fresh[1083], Fresh[1082]}), .c ({new_AGEMA_signal_6472, SubBytesIns_Inst_Sbox_12_M51}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M52_U1 ( .a ({new_AGEMA_signal_6466, SubBytesIns_Inst_Sbox_12_M42}), .b ({new_AGEMA_signal_12934, new_AGEMA_signal_12931}), .clk (clk), .r ({Fresh[1085], Fresh[1084]}), .c ({new_AGEMA_signal_6708, SubBytesIns_Inst_Sbox_12_M52}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M53_U1 ( .a ({new_AGEMA_signal_6705, SubBytesIns_Inst_Sbox_12_M45}), .b ({new_AGEMA_signal_12940, new_AGEMA_signal_12937}), .clk (clk), .r ({Fresh[1087], Fresh[1086]}), .c ({new_AGEMA_signal_6913, SubBytesIns_Inst_Sbox_12_M53}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M54_U1 ( .a ({new_AGEMA_signal_6465, SubBytesIns_Inst_Sbox_12_M41}), .b ({new_AGEMA_signal_12946, new_AGEMA_signal_12943}), .clk (clk), .r ({Fresh[1089], Fresh[1088]}), .c ({new_AGEMA_signal_6709, SubBytesIns_Inst_Sbox_12_M54}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M55_U1 ( .a ({new_AGEMA_signal_6468, SubBytesIns_Inst_Sbox_12_M44}), .b ({new_AGEMA_signal_12952, new_AGEMA_signal_12949}), .clk (clk), .r ({Fresh[1091], Fresh[1090]}), .c ({new_AGEMA_signal_6710, SubBytesIns_Inst_Sbox_12_M55}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M56_U1 ( .a ({new_AGEMA_signal_6260, SubBytesIns_Inst_Sbox_12_M40}), .b ({new_AGEMA_signal_12958, new_AGEMA_signal_12955}), .clk (clk), .r ({Fresh[1093], Fresh[1092]}), .c ({new_AGEMA_signal_6473, SubBytesIns_Inst_Sbox_12_M56}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M57_U1 ( .a ({new_AGEMA_signal_6259, SubBytesIns_Inst_Sbox_12_M39}), .b ({new_AGEMA_signal_12964, new_AGEMA_signal_12961}), .clk (clk), .r ({Fresh[1095], Fresh[1094]}), .c ({new_AGEMA_signal_6474, SubBytesIns_Inst_Sbox_12_M57}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M58_U1 ( .a ({new_AGEMA_signal_6467, SubBytesIns_Inst_Sbox_12_M43}), .b ({new_AGEMA_signal_12970, new_AGEMA_signal_12967}), .clk (clk), .r ({Fresh[1097], Fresh[1096]}), .c ({new_AGEMA_signal_6711, SubBytesIns_Inst_Sbox_12_M58}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M59_U1 ( .a ({new_AGEMA_signal_6258, SubBytesIns_Inst_Sbox_12_M38}), .b ({new_AGEMA_signal_12976, new_AGEMA_signal_12973}), .clk (clk), .r ({Fresh[1099], Fresh[1098]}), .c ({new_AGEMA_signal_6475, SubBytesIns_Inst_Sbox_12_M59}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M60_U1 ( .a ({new_AGEMA_signal_6257, SubBytesIns_Inst_Sbox_12_M37}), .b ({new_AGEMA_signal_12982, new_AGEMA_signal_12979}), .clk (clk), .r ({Fresh[1101], Fresh[1100]}), .c ({new_AGEMA_signal_6476, SubBytesIns_Inst_Sbox_12_M60}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M61_U1 ( .a ({new_AGEMA_signal_6466, SubBytesIns_Inst_Sbox_12_M42}), .b ({new_AGEMA_signal_12988, new_AGEMA_signal_12985}), .clk (clk), .r ({Fresh[1103], Fresh[1102]}), .c ({new_AGEMA_signal_6712, SubBytesIns_Inst_Sbox_12_M61}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M62_U1 ( .a ({new_AGEMA_signal_6705, SubBytesIns_Inst_Sbox_12_M45}), .b ({new_AGEMA_signal_12994, new_AGEMA_signal_12991}), .clk (clk), .r ({Fresh[1105], Fresh[1104]}), .c ({new_AGEMA_signal_6914, SubBytesIns_Inst_Sbox_12_M62}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M63_U1 ( .a ({new_AGEMA_signal_6465, SubBytesIns_Inst_Sbox_12_M41}), .b ({new_AGEMA_signal_13000, new_AGEMA_signal_12997}), .clk (clk), .r ({Fresh[1107], Fresh[1106]}), .c ({new_AGEMA_signal_6713, SubBytesIns_Inst_Sbox_12_M63}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L0_U1 ( .a ({new_AGEMA_signal_6712, SubBytesIns_Inst_Sbox_12_M61}), .b ({new_AGEMA_signal_6914, SubBytesIns_Inst_Sbox_12_M62}), .c ({new_AGEMA_signal_7097, SubBytesIns_Inst_Sbox_12_L0}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L1_U1 ( .a ({new_AGEMA_signal_6471, SubBytesIns_Inst_Sbox_12_M50}), .b ({new_AGEMA_signal_6473, SubBytesIns_Inst_Sbox_12_M56}), .c ({new_AGEMA_signal_6714, SubBytesIns_Inst_Sbox_12_L1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L2_U1 ( .a ({new_AGEMA_signal_6706, SubBytesIns_Inst_Sbox_12_M46}), .b ({new_AGEMA_signal_6470, SubBytesIns_Inst_Sbox_12_M48}), .c ({new_AGEMA_signal_6915, SubBytesIns_Inst_Sbox_12_L2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L3_U1 ( .a ({new_AGEMA_signal_6469, SubBytesIns_Inst_Sbox_12_M47}), .b ({new_AGEMA_signal_6710, SubBytesIns_Inst_Sbox_12_M55}), .c ({new_AGEMA_signal_6916, SubBytesIns_Inst_Sbox_12_L3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L4_U1 ( .a ({new_AGEMA_signal_6709, SubBytesIns_Inst_Sbox_12_M54}), .b ({new_AGEMA_signal_6711, SubBytesIns_Inst_Sbox_12_M58}), .c ({new_AGEMA_signal_6917, SubBytesIns_Inst_Sbox_12_L4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L5_U1 ( .a ({new_AGEMA_signal_6707, SubBytesIns_Inst_Sbox_12_M49}), .b ({new_AGEMA_signal_6712, SubBytesIns_Inst_Sbox_12_M61}), .c ({new_AGEMA_signal_6918, SubBytesIns_Inst_Sbox_12_L5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L6_U1 ( .a ({new_AGEMA_signal_6914, SubBytesIns_Inst_Sbox_12_M62}), .b ({new_AGEMA_signal_6918, SubBytesIns_Inst_Sbox_12_L5}), .c ({new_AGEMA_signal_7098, SubBytesIns_Inst_Sbox_12_L6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L7_U1 ( .a ({new_AGEMA_signal_6706, SubBytesIns_Inst_Sbox_12_M46}), .b ({new_AGEMA_signal_6916, SubBytesIns_Inst_Sbox_12_L3}), .c ({new_AGEMA_signal_7099, SubBytesIns_Inst_Sbox_12_L7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L8_U1 ( .a ({new_AGEMA_signal_6472, SubBytesIns_Inst_Sbox_12_M51}), .b ({new_AGEMA_signal_6475, SubBytesIns_Inst_Sbox_12_M59}), .c ({new_AGEMA_signal_6715, SubBytesIns_Inst_Sbox_12_L8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L9_U1 ( .a ({new_AGEMA_signal_6708, SubBytesIns_Inst_Sbox_12_M52}), .b ({new_AGEMA_signal_6913, SubBytesIns_Inst_Sbox_12_M53}), .c ({new_AGEMA_signal_7100, SubBytesIns_Inst_Sbox_12_L9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L10_U1 ( .a ({new_AGEMA_signal_6913, SubBytesIns_Inst_Sbox_12_M53}), .b ({new_AGEMA_signal_6917, SubBytesIns_Inst_Sbox_12_L4}), .c ({new_AGEMA_signal_7101, SubBytesIns_Inst_Sbox_12_L10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L11_U1 ( .a ({new_AGEMA_signal_6476, SubBytesIns_Inst_Sbox_12_M60}), .b ({new_AGEMA_signal_6915, SubBytesIns_Inst_Sbox_12_L2}), .c ({new_AGEMA_signal_7102, SubBytesIns_Inst_Sbox_12_L11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L12_U1 ( .a ({new_AGEMA_signal_6470, SubBytesIns_Inst_Sbox_12_M48}), .b ({new_AGEMA_signal_6472, SubBytesIns_Inst_Sbox_12_M51}), .c ({new_AGEMA_signal_6716, SubBytesIns_Inst_Sbox_12_L12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L13_U1 ( .a ({new_AGEMA_signal_6471, SubBytesIns_Inst_Sbox_12_M50}), .b ({new_AGEMA_signal_7097, SubBytesIns_Inst_Sbox_12_L0}), .c ({new_AGEMA_signal_7309, SubBytesIns_Inst_Sbox_12_L13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L14_U1 ( .a ({new_AGEMA_signal_6708, SubBytesIns_Inst_Sbox_12_M52}), .b ({new_AGEMA_signal_6712, SubBytesIns_Inst_Sbox_12_M61}), .c ({new_AGEMA_signal_6919, SubBytesIns_Inst_Sbox_12_L14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L15_U1 ( .a ({new_AGEMA_signal_6710, SubBytesIns_Inst_Sbox_12_M55}), .b ({new_AGEMA_signal_6714, SubBytesIns_Inst_Sbox_12_L1}), .c ({new_AGEMA_signal_6920, SubBytesIns_Inst_Sbox_12_L15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L16_U1 ( .a ({new_AGEMA_signal_6473, SubBytesIns_Inst_Sbox_12_M56}), .b ({new_AGEMA_signal_7097, SubBytesIns_Inst_Sbox_12_L0}), .c ({new_AGEMA_signal_7310, SubBytesIns_Inst_Sbox_12_L16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L17_U1 ( .a ({new_AGEMA_signal_6474, SubBytesIns_Inst_Sbox_12_M57}), .b ({new_AGEMA_signal_6714, SubBytesIns_Inst_Sbox_12_L1}), .c ({new_AGEMA_signal_6921, SubBytesIns_Inst_Sbox_12_L17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L18_U1 ( .a ({new_AGEMA_signal_6711, SubBytesIns_Inst_Sbox_12_M58}), .b ({new_AGEMA_signal_6715, SubBytesIns_Inst_Sbox_12_L8}), .c ({new_AGEMA_signal_6922, SubBytesIns_Inst_Sbox_12_L18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L19_U1 ( .a ({new_AGEMA_signal_6713, SubBytesIns_Inst_Sbox_12_M63}), .b ({new_AGEMA_signal_6917, SubBytesIns_Inst_Sbox_12_L4}), .c ({new_AGEMA_signal_7103, SubBytesIns_Inst_Sbox_12_L19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L20_U1 ( .a ({new_AGEMA_signal_7097, SubBytesIns_Inst_Sbox_12_L0}), .b ({new_AGEMA_signal_6714, SubBytesIns_Inst_Sbox_12_L1}), .c ({new_AGEMA_signal_7311, SubBytesIns_Inst_Sbox_12_L20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L21_U1 ( .a ({new_AGEMA_signal_6714, SubBytesIns_Inst_Sbox_12_L1}), .b ({new_AGEMA_signal_7099, SubBytesIns_Inst_Sbox_12_L7}), .c ({new_AGEMA_signal_7312, SubBytesIns_Inst_Sbox_12_L21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L22_U1 ( .a ({new_AGEMA_signal_6916, SubBytesIns_Inst_Sbox_12_L3}), .b ({new_AGEMA_signal_6716, SubBytesIns_Inst_Sbox_12_L12}), .c ({new_AGEMA_signal_7104, SubBytesIns_Inst_Sbox_12_L22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L23_U1 ( .a ({new_AGEMA_signal_6922, SubBytesIns_Inst_Sbox_12_L18}), .b ({new_AGEMA_signal_6915, SubBytesIns_Inst_Sbox_12_L2}), .c ({new_AGEMA_signal_7105, SubBytesIns_Inst_Sbox_12_L23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L24_U1 ( .a ({new_AGEMA_signal_6920, SubBytesIns_Inst_Sbox_12_L15}), .b ({new_AGEMA_signal_7100, SubBytesIns_Inst_Sbox_12_L9}), .c ({new_AGEMA_signal_7313, SubBytesIns_Inst_Sbox_12_L24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L25_U1 ( .a ({new_AGEMA_signal_7098, SubBytesIns_Inst_Sbox_12_L6}), .b ({new_AGEMA_signal_7101, SubBytesIns_Inst_Sbox_12_L10}), .c ({new_AGEMA_signal_7314, SubBytesIns_Inst_Sbox_12_L25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L26_U1 ( .a ({new_AGEMA_signal_7099, SubBytesIns_Inst_Sbox_12_L7}), .b ({new_AGEMA_signal_7100, SubBytesIns_Inst_Sbox_12_L9}), .c ({new_AGEMA_signal_7315, SubBytesIns_Inst_Sbox_12_L26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L27_U1 ( .a ({new_AGEMA_signal_6715, SubBytesIns_Inst_Sbox_12_L8}), .b ({new_AGEMA_signal_7101, SubBytesIns_Inst_Sbox_12_L10}), .c ({new_AGEMA_signal_7316, SubBytesIns_Inst_Sbox_12_L27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L28_U1 ( .a ({new_AGEMA_signal_7102, SubBytesIns_Inst_Sbox_12_L11}), .b ({new_AGEMA_signal_6919, SubBytesIns_Inst_Sbox_12_L14}), .c ({new_AGEMA_signal_7317, SubBytesIns_Inst_Sbox_12_L28}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L29_U1 ( .a ({new_AGEMA_signal_7102, SubBytesIns_Inst_Sbox_12_L11}), .b ({new_AGEMA_signal_6921, SubBytesIns_Inst_Sbox_12_L17}), .c ({new_AGEMA_signal_7318, SubBytesIns_Inst_Sbox_12_L29}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_S0_U1 ( .a ({new_AGEMA_signal_7098, SubBytesIns_Inst_Sbox_12_L6}), .b ({new_AGEMA_signal_7313, SubBytesIns_Inst_Sbox_12_L24}), .c ({new_AGEMA_signal_7469, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_S1_U1 ( .a ({new_AGEMA_signal_7310, SubBytesIns_Inst_Sbox_12_L16}), .b ({new_AGEMA_signal_7315, SubBytesIns_Inst_Sbox_12_L26}), .c ({new_AGEMA_signal_7470, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_S2_U1 ( .a ({new_AGEMA_signal_7103, SubBytesIns_Inst_Sbox_12_L19}), .b ({new_AGEMA_signal_7317, SubBytesIns_Inst_Sbox_12_L28}), .c ({new_AGEMA_signal_7471, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_S3_U1 ( .a ({new_AGEMA_signal_7098, SubBytesIns_Inst_Sbox_12_L6}), .b ({new_AGEMA_signal_7312, SubBytesIns_Inst_Sbox_12_L21}), .c ({new_AGEMA_signal_7472, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_S4_U1 ( .a ({new_AGEMA_signal_7311, SubBytesIns_Inst_Sbox_12_L20}), .b ({new_AGEMA_signal_7104, SubBytesIns_Inst_Sbox_12_L22}), .c ({new_AGEMA_signal_7473, MixColumnsInput[67]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_S5_U1 ( .a ({new_AGEMA_signal_7314, SubBytesIns_Inst_Sbox_12_L25}), .b ({new_AGEMA_signal_7318, SubBytesIns_Inst_Sbox_12_L29}), .c ({new_AGEMA_signal_7474, MixColumnsInput[66]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_S6_U1 ( .a ({new_AGEMA_signal_7309, SubBytesIns_Inst_Sbox_12_L13}), .b ({new_AGEMA_signal_7316, SubBytesIns_Inst_Sbox_12_L27}), .c ({new_AGEMA_signal_7475, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_S7_U1 ( .a ({new_AGEMA_signal_7098, SubBytesIns_Inst_Sbox_12_L6}), .b ({new_AGEMA_signal_7105, SubBytesIns_Inst_Sbox_12_L23}), .c ({new_AGEMA_signal_7319, MixColumnsInput[64]}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M46_U1 ( .a ({new_AGEMA_signal_6480, SubBytesIns_Inst_Sbox_13_M44}), .b ({new_AGEMA_signal_13006, new_AGEMA_signal_13003}), .clk (clk), .r ({Fresh[1109], Fresh[1108]}), .c ({new_AGEMA_signal_6718, SubBytesIns_Inst_Sbox_13_M46}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M47_U1 ( .a ({new_AGEMA_signal_6264, SubBytesIns_Inst_Sbox_13_M40}), .b ({new_AGEMA_signal_13012, new_AGEMA_signal_13009}), .clk (clk), .r ({Fresh[1111], Fresh[1110]}), .c ({new_AGEMA_signal_6481, SubBytesIns_Inst_Sbox_13_M47}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M48_U1 ( .a ({new_AGEMA_signal_6263, SubBytesIns_Inst_Sbox_13_M39}), .b ({new_AGEMA_signal_13018, new_AGEMA_signal_13015}), .clk (clk), .r ({Fresh[1113], Fresh[1112]}), .c ({new_AGEMA_signal_6482, SubBytesIns_Inst_Sbox_13_M48}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M49_U1 ( .a ({new_AGEMA_signal_6479, SubBytesIns_Inst_Sbox_13_M43}), .b ({new_AGEMA_signal_13024, new_AGEMA_signal_13021}), .clk (clk), .r ({Fresh[1115], Fresh[1114]}), .c ({new_AGEMA_signal_6719, SubBytesIns_Inst_Sbox_13_M49}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M50_U1 ( .a ({new_AGEMA_signal_6262, SubBytesIns_Inst_Sbox_13_M38}), .b ({new_AGEMA_signal_13030, new_AGEMA_signal_13027}), .clk (clk), .r ({Fresh[1117], Fresh[1116]}), .c ({new_AGEMA_signal_6483, SubBytesIns_Inst_Sbox_13_M50}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M51_U1 ( .a ({new_AGEMA_signal_6261, SubBytesIns_Inst_Sbox_13_M37}), .b ({new_AGEMA_signal_13036, new_AGEMA_signal_13033}), .clk (clk), .r ({Fresh[1119], Fresh[1118]}), .c ({new_AGEMA_signal_6484, SubBytesIns_Inst_Sbox_13_M51}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M52_U1 ( .a ({new_AGEMA_signal_6478, SubBytesIns_Inst_Sbox_13_M42}), .b ({new_AGEMA_signal_13042, new_AGEMA_signal_13039}), .clk (clk), .r ({Fresh[1121], Fresh[1120]}), .c ({new_AGEMA_signal_6720, SubBytesIns_Inst_Sbox_13_M52}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M53_U1 ( .a ({new_AGEMA_signal_6717, SubBytesIns_Inst_Sbox_13_M45}), .b ({new_AGEMA_signal_13048, new_AGEMA_signal_13045}), .clk (clk), .r ({Fresh[1123], Fresh[1122]}), .c ({new_AGEMA_signal_6923, SubBytesIns_Inst_Sbox_13_M53}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M54_U1 ( .a ({new_AGEMA_signal_6477, SubBytesIns_Inst_Sbox_13_M41}), .b ({new_AGEMA_signal_13054, new_AGEMA_signal_13051}), .clk (clk), .r ({Fresh[1125], Fresh[1124]}), .c ({new_AGEMA_signal_6721, SubBytesIns_Inst_Sbox_13_M54}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M55_U1 ( .a ({new_AGEMA_signal_6480, SubBytesIns_Inst_Sbox_13_M44}), .b ({new_AGEMA_signal_13060, new_AGEMA_signal_13057}), .clk (clk), .r ({Fresh[1127], Fresh[1126]}), .c ({new_AGEMA_signal_6722, SubBytesIns_Inst_Sbox_13_M55}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M56_U1 ( .a ({new_AGEMA_signal_6264, SubBytesIns_Inst_Sbox_13_M40}), .b ({new_AGEMA_signal_13066, new_AGEMA_signal_13063}), .clk (clk), .r ({Fresh[1129], Fresh[1128]}), .c ({new_AGEMA_signal_6485, SubBytesIns_Inst_Sbox_13_M56}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M57_U1 ( .a ({new_AGEMA_signal_6263, SubBytesIns_Inst_Sbox_13_M39}), .b ({new_AGEMA_signal_13072, new_AGEMA_signal_13069}), .clk (clk), .r ({Fresh[1131], Fresh[1130]}), .c ({new_AGEMA_signal_6486, SubBytesIns_Inst_Sbox_13_M57}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M58_U1 ( .a ({new_AGEMA_signal_6479, SubBytesIns_Inst_Sbox_13_M43}), .b ({new_AGEMA_signal_13078, new_AGEMA_signal_13075}), .clk (clk), .r ({Fresh[1133], Fresh[1132]}), .c ({new_AGEMA_signal_6723, SubBytesIns_Inst_Sbox_13_M58}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M59_U1 ( .a ({new_AGEMA_signal_6262, SubBytesIns_Inst_Sbox_13_M38}), .b ({new_AGEMA_signal_13084, new_AGEMA_signal_13081}), .clk (clk), .r ({Fresh[1135], Fresh[1134]}), .c ({new_AGEMA_signal_6487, SubBytesIns_Inst_Sbox_13_M59}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M60_U1 ( .a ({new_AGEMA_signal_6261, SubBytesIns_Inst_Sbox_13_M37}), .b ({new_AGEMA_signal_13090, new_AGEMA_signal_13087}), .clk (clk), .r ({Fresh[1137], Fresh[1136]}), .c ({new_AGEMA_signal_6488, SubBytesIns_Inst_Sbox_13_M60}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M61_U1 ( .a ({new_AGEMA_signal_6478, SubBytesIns_Inst_Sbox_13_M42}), .b ({new_AGEMA_signal_13096, new_AGEMA_signal_13093}), .clk (clk), .r ({Fresh[1139], Fresh[1138]}), .c ({new_AGEMA_signal_6724, SubBytesIns_Inst_Sbox_13_M61}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M62_U1 ( .a ({new_AGEMA_signal_6717, SubBytesIns_Inst_Sbox_13_M45}), .b ({new_AGEMA_signal_13102, new_AGEMA_signal_13099}), .clk (clk), .r ({Fresh[1141], Fresh[1140]}), .c ({new_AGEMA_signal_6924, SubBytesIns_Inst_Sbox_13_M62}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M63_U1 ( .a ({new_AGEMA_signal_6477, SubBytesIns_Inst_Sbox_13_M41}), .b ({new_AGEMA_signal_13108, new_AGEMA_signal_13105}), .clk (clk), .r ({Fresh[1143], Fresh[1142]}), .c ({new_AGEMA_signal_6725, SubBytesIns_Inst_Sbox_13_M63}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L0_U1 ( .a ({new_AGEMA_signal_6724, SubBytesIns_Inst_Sbox_13_M61}), .b ({new_AGEMA_signal_6924, SubBytesIns_Inst_Sbox_13_M62}), .c ({new_AGEMA_signal_7106, SubBytesIns_Inst_Sbox_13_L0}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L1_U1 ( .a ({new_AGEMA_signal_6483, SubBytesIns_Inst_Sbox_13_M50}), .b ({new_AGEMA_signal_6485, SubBytesIns_Inst_Sbox_13_M56}), .c ({new_AGEMA_signal_6726, SubBytesIns_Inst_Sbox_13_L1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L2_U1 ( .a ({new_AGEMA_signal_6718, SubBytesIns_Inst_Sbox_13_M46}), .b ({new_AGEMA_signal_6482, SubBytesIns_Inst_Sbox_13_M48}), .c ({new_AGEMA_signal_6925, SubBytesIns_Inst_Sbox_13_L2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L3_U1 ( .a ({new_AGEMA_signal_6481, SubBytesIns_Inst_Sbox_13_M47}), .b ({new_AGEMA_signal_6722, SubBytesIns_Inst_Sbox_13_M55}), .c ({new_AGEMA_signal_6926, SubBytesIns_Inst_Sbox_13_L3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L4_U1 ( .a ({new_AGEMA_signal_6721, SubBytesIns_Inst_Sbox_13_M54}), .b ({new_AGEMA_signal_6723, SubBytesIns_Inst_Sbox_13_M58}), .c ({new_AGEMA_signal_6927, SubBytesIns_Inst_Sbox_13_L4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L5_U1 ( .a ({new_AGEMA_signal_6719, SubBytesIns_Inst_Sbox_13_M49}), .b ({new_AGEMA_signal_6724, SubBytesIns_Inst_Sbox_13_M61}), .c ({new_AGEMA_signal_6928, SubBytesIns_Inst_Sbox_13_L5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L6_U1 ( .a ({new_AGEMA_signal_6924, SubBytesIns_Inst_Sbox_13_M62}), .b ({new_AGEMA_signal_6928, SubBytesIns_Inst_Sbox_13_L5}), .c ({new_AGEMA_signal_7107, SubBytesIns_Inst_Sbox_13_L6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L7_U1 ( .a ({new_AGEMA_signal_6718, SubBytesIns_Inst_Sbox_13_M46}), .b ({new_AGEMA_signal_6926, SubBytesIns_Inst_Sbox_13_L3}), .c ({new_AGEMA_signal_7108, SubBytesIns_Inst_Sbox_13_L7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L8_U1 ( .a ({new_AGEMA_signal_6484, SubBytesIns_Inst_Sbox_13_M51}), .b ({new_AGEMA_signal_6487, SubBytesIns_Inst_Sbox_13_M59}), .c ({new_AGEMA_signal_6727, SubBytesIns_Inst_Sbox_13_L8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L9_U1 ( .a ({new_AGEMA_signal_6720, SubBytesIns_Inst_Sbox_13_M52}), .b ({new_AGEMA_signal_6923, SubBytesIns_Inst_Sbox_13_M53}), .c ({new_AGEMA_signal_7109, SubBytesIns_Inst_Sbox_13_L9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L10_U1 ( .a ({new_AGEMA_signal_6923, SubBytesIns_Inst_Sbox_13_M53}), .b ({new_AGEMA_signal_6927, SubBytesIns_Inst_Sbox_13_L4}), .c ({new_AGEMA_signal_7110, SubBytesIns_Inst_Sbox_13_L10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L11_U1 ( .a ({new_AGEMA_signal_6488, SubBytesIns_Inst_Sbox_13_M60}), .b ({new_AGEMA_signal_6925, SubBytesIns_Inst_Sbox_13_L2}), .c ({new_AGEMA_signal_7111, SubBytesIns_Inst_Sbox_13_L11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L12_U1 ( .a ({new_AGEMA_signal_6482, SubBytesIns_Inst_Sbox_13_M48}), .b ({new_AGEMA_signal_6484, SubBytesIns_Inst_Sbox_13_M51}), .c ({new_AGEMA_signal_6728, SubBytesIns_Inst_Sbox_13_L12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L13_U1 ( .a ({new_AGEMA_signal_6483, SubBytesIns_Inst_Sbox_13_M50}), .b ({new_AGEMA_signal_7106, SubBytesIns_Inst_Sbox_13_L0}), .c ({new_AGEMA_signal_7320, SubBytesIns_Inst_Sbox_13_L13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L14_U1 ( .a ({new_AGEMA_signal_6720, SubBytesIns_Inst_Sbox_13_M52}), .b ({new_AGEMA_signal_6724, SubBytesIns_Inst_Sbox_13_M61}), .c ({new_AGEMA_signal_6929, SubBytesIns_Inst_Sbox_13_L14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L15_U1 ( .a ({new_AGEMA_signal_6722, SubBytesIns_Inst_Sbox_13_M55}), .b ({new_AGEMA_signal_6726, SubBytesIns_Inst_Sbox_13_L1}), .c ({new_AGEMA_signal_6930, SubBytesIns_Inst_Sbox_13_L15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L16_U1 ( .a ({new_AGEMA_signal_6485, SubBytesIns_Inst_Sbox_13_M56}), .b ({new_AGEMA_signal_7106, SubBytesIns_Inst_Sbox_13_L0}), .c ({new_AGEMA_signal_7321, SubBytesIns_Inst_Sbox_13_L16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L17_U1 ( .a ({new_AGEMA_signal_6486, SubBytesIns_Inst_Sbox_13_M57}), .b ({new_AGEMA_signal_6726, SubBytesIns_Inst_Sbox_13_L1}), .c ({new_AGEMA_signal_6931, SubBytesIns_Inst_Sbox_13_L17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L18_U1 ( .a ({new_AGEMA_signal_6723, SubBytesIns_Inst_Sbox_13_M58}), .b ({new_AGEMA_signal_6727, SubBytesIns_Inst_Sbox_13_L8}), .c ({new_AGEMA_signal_6932, SubBytesIns_Inst_Sbox_13_L18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L19_U1 ( .a ({new_AGEMA_signal_6725, SubBytesIns_Inst_Sbox_13_M63}), .b ({new_AGEMA_signal_6927, SubBytesIns_Inst_Sbox_13_L4}), .c ({new_AGEMA_signal_7112, SubBytesIns_Inst_Sbox_13_L19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L20_U1 ( .a ({new_AGEMA_signal_7106, SubBytesIns_Inst_Sbox_13_L0}), .b ({new_AGEMA_signal_6726, SubBytesIns_Inst_Sbox_13_L1}), .c ({new_AGEMA_signal_7322, SubBytesIns_Inst_Sbox_13_L20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L21_U1 ( .a ({new_AGEMA_signal_6726, SubBytesIns_Inst_Sbox_13_L1}), .b ({new_AGEMA_signal_7108, SubBytesIns_Inst_Sbox_13_L7}), .c ({new_AGEMA_signal_7323, SubBytesIns_Inst_Sbox_13_L21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L22_U1 ( .a ({new_AGEMA_signal_6926, SubBytesIns_Inst_Sbox_13_L3}), .b ({new_AGEMA_signal_6728, SubBytesIns_Inst_Sbox_13_L12}), .c ({new_AGEMA_signal_7113, SubBytesIns_Inst_Sbox_13_L22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L23_U1 ( .a ({new_AGEMA_signal_6932, SubBytesIns_Inst_Sbox_13_L18}), .b ({new_AGEMA_signal_6925, SubBytesIns_Inst_Sbox_13_L2}), .c ({new_AGEMA_signal_7114, SubBytesIns_Inst_Sbox_13_L23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L24_U1 ( .a ({new_AGEMA_signal_6930, SubBytesIns_Inst_Sbox_13_L15}), .b ({new_AGEMA_signal_7109, SubBytesIns_Inst_Sbox_13_L9}), .c ({new_AGEMA_signal_7324, SubBytesIns_Inst_Sbox_13_L24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L25_U1 ( .a ({new_AGEMA_signal_7107, SubBytesIns_Inst_Sbox_13_L6}), .b ({new_AGEMA_signal_7110, SubBytesIns_Inst_Sbox_13_L10}), .c ({new_AGEMA_signal_7325, SubBytesIns_Inst_Sbox_13_L25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L26_U1 ( .a ({new_AGEMA_signal_7108, SubBytesIns_Inst_Sbox_13_L7}), .b ({new_AGEMA_signal_7109, SubBytesIns_Inst_Sbox_13_L9}), .c ({new_AGEMA_signal_7326, SubBytesIns_Inst_Sbox_13_L26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L27_U1 ( .a ({new_AGEMA_signal_6727, SubBytesIns_Inst_Sbox_13_L8}), .b ({new_AGEMA_signal_7110, SubBytesIns_Inst_Sbox_13_L10}), .c ({new_AGEMA_signal_7327, SubBytesIns_Inst_Sbox_13_L27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L28_U1 ( .a ({new_AGEMA_signal_7111, SubBytesIns_Inst_Sbox_13_L11}), .b ({new_AGEMA_signal_6929, SubBytesIns_Inst_Sbox_13_L14}), .c ({new_AGEMA_signal_7328, SubBytesIns_Inst_Sbox_13_L28}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L29_U1 ( .a ({new_AGEMA_signal_7111, SubBytesIns_Inst_Sbox_13_L11}), .b ({new_AGEMA_signal_6931, SubBytesIns_Inst_Sbox_13_L17}), .c ({new_AGEMA_signal_7329, SubBytesIns_Inst_Sbox_13_L29}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_S0_U1 ( .a ({new_AGEMA_signal_7107, SubBytesIns_Inst_Sbox_13_L6}), .b ({new_AGEMA_signal_7324, SubBytesIns_Inst_Sbox_13_L24}), .c ({new_AGEMA_signal_7476, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_S1_U1 ( .a ({new_AGEMA_signal_7321, SubBytesIns_Inst_Sbox_13_L16}), .b ({new_AGEMA_signal_7326, SubBytesIns_Inst_Sbox_13_L26}), .c ({new_AGEMA_signal_7477, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_S2_U1 ( .a ({new_AGEMA_signal_7112, SubBytesIns_Inst_Sbox_13_L19}), .b ({new_AGEMA_signal_7328, SubBytesIns_Inst_Sbox_13_L28}), .c ({new_AGEMA_signal_7478, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_S3_U1 ( .a ({new_AGEMA_signal_7107, SubBytesIns_Inst_Sbox_13_L6}), .b ({new_AGEMA_signal_7323, SubBytesIns_Inst_Sbox_13_L21}), .c ({new_AGEMA_signal_7479, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_S4_U1 ( .a ({new_AGEMA_signal_7322, SubBytesIns_Inst_Sbox_13_L20}), .b ({new_AGEMA_signal_7113, SubBytesIns_Inst_Sbox_13_L22}), .c ({new_AGEMA_signal_7480, MixColumnsInput[43]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_S5_U1 ( .a ({new_AGEMA_signal_7325, SubBytesIns_Inst_Sbox_13_L25}), .b ({new_AGEMA_signal_7329, SubBytesIns_Inst_Sbox_13_L29}), .c ({new_AGEMA_signal_7481, MixColumnsInput[42]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_S6_U1 ( .a ({new_AGEMA_signal_7320, SubBytesIns_Inst_Sbox_13_L13}), .b ({new_AGEMA_signal_7327, SubBytesIns_Inst_Sbox_13_L27}), .c ({new_AGEMA_signal_7482, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_S7_U1 ( .a ({new_AGEMA_signal_7107, SubBytesIns_Inst_Sbox_13_L6}), .b ({new_AGEMA_signal_7114, SubBytesIns_Inst_Sbox_13_L23}), .c ({new_AGEMA_signal_7330, MixColumnsInput[40]}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M46_U1 ( .a ({new_AGEMA_signal_6492, SubBytesIns_Inst_Sbox_14_M44}), .b ({new_AGEMA_signal_13114, new_AGEMA_signal_13111}), .clk (clk), .r ({Fresh[1145], Fresh[1144]}), .c ({new_AGEMA_signal_6730, SubBytesIns_Inst_Sbox_14_M46}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M47_U1 ( .a ({new_AGEMA_signal_6268, SubBytesIns_Inst_Sbox_14_M40}), .b ({new_AGEMA_signal_13120, new_AGEMA_signal_13117}), .clk (clk), .r ({Fresh[1147], Fresh[1146]}), .c ({new_AGEMA_signal_6493, SubBytesIns_Inst_Sbox_14_M47}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M48_U1 ( .a ({new_AGEMA_signal_6267, SubBytesIns_Inst_Sbox_14_M39}), .b ({new_AGEMA_signal_13126, new_AGEMA_signal_13123}), .clk (clk), .r ({Fresh[1149], Fresh[1148]}), .c ({new_AGEMA_signal_6494, SubBytesIns_Inst_Sbox_14_M48}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M49_U1 ( .a ({new_AGEMA_signal_6491, SubBytesIns_Inst_Sbox_14_M43}), .b ({new_AGEMA_signal_13132, new_AGEMA_signal_13129}), .clk (clk), .r ({Fresh[1151], Fresh[1150]}), .c ({new_AGEMA_signal_6731, SubBytesIns_Inst_Sbox_14_M49}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M50_U1 ( .a ({new_AGEMA_signal_6266, SubBytesIns_Inst_Sbox_14_M38}), .b ({new_AGEMA_signal_13138, new_AGEMA_signal_13135}), .clk (clk), .r ({Fresh[1153], Fresh[1152]}), .c ({new_AGEMA_signal_6495, SubBytesIns_Inst_Sbox_14_M50}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M51_U1 ( .a ({new_AGEMA_signal_6265, SubBytesIns_Inst_Sbox_14_M37}), .b ({new_AGEMA_signal_13144, new_AGEMA_signal_13141}), .clk (clk), .r ({Fresh[1155], Fresh[1154]}), .c ({new_AGEMA_signal_6496, SubBytesIns_Inst_Sbox_14_M51}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M52_U1 ( .a ({new_AGEMA_signal_6490, SubBytesIns_Inst_Sbox_14_M42}), .b ({new_AGEMA_signal_13150, new_AGEMA_signal_13147}), .clk (clk), .r ({Fresh[1157], Fresh[1156]}), .c ({new_AGEMA_signal_6732, SubBytesIns_Inst_Sbox_14_M52}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M53_U1 ( .a ({new_AGEMA_signal_6729, SubBytesIns_Inst_Sbox_14_M45}), .b ({new_AGEMA_signal_13156, new_AGEMA_signal_13153}), .clk (clk), .r ({Fresh[1159], Fresh[1158]}), .c ({new_AGEMA_signal_6933, SubBytesIns_Inst_Sbox_14_M53}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M54_U1 ( .a ({new_AGEMA_signal_6489, SubBytesIns_Inst_Sbox_14_M41}), .b ({new_AGEMA_signal_13162, new_AGEMA_signal_13159}), .clk (clk), .r ({Fresh[1161], Fresh[1160]}), .c ({new_AGEMA_signal_6733, SubBytesIns_Inst_Sbox_14_M54}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M55_U1 ( .a ({new_AGEMA_signal_6492, SubBytesIns_Inst_Sbox_14_M44}), .b ({new_AGEMA_signal_13168, new_AGEMA_signal_13165}), .clk (clk), .r ({Fresh[1163], Fresh[1162]}), .c ({new_AGEMA_signal_6734, SubBytesIns_Inst_Sbox_14_M55}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M56_U1 ( .a ({new_AGEMA_signal_6268, SubBytesIns_Inst_Sbox_14_M40}), .b ({new_AGEMA_signal_13174, new_AGEMA_signal_13171}), .clk (clk), .r ({Fresh[1165], Fresh[1164]}), .c ({new_AGEMA_signal_6497, SubBytesIns_Inst_Sbox_14_M56}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M57_U1 ( .a ({new_AGEMA_signal_6267, SubBytesIns_Inst_Sbox_14_M39}), .b ({new_AGEMA_signal_13180, new_AGEMA_signal_13177}), .clk (clk), .r ({Fresh[1167], Fresh[1166]}), .c ({new_AGEMA_signal_6498, SubBytesIns_Inst_Sbox_14_M57}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M58_U1 ( .a ({new_AGEMA_signal_6491, SubBytesIns_Inst_Sbox_14_M43}), .b ({new_AGEMA_signal_13186, new_AGEMA_signal_13183}), .clk (clk), .r ({Fresh[1169], Fresh[1168]}), .c ({new_AGEMA_signal_6735, SubBytesIns_Inst_Sbox_14_M58}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M59_U1 ( .a ({new_AGEMA_signal_6266, SubBytesIns_Inst_Sbox_14_M38}), .b ({new_AGEMA_signal_13192, new_AGEMA_signal_13189}), .clk (clk), .r ({Fresh[1171], Fresh[1170]}), .c ({new_AGEMA_signal_6499, SubBytesIns_Inst_Sbox_14_M59}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M60_U1 ( .a ({new_AGEMA_signal_6265, SubBytesIns_Inst_Sbox_14_M37}), .b ({new_AGEMA_signal_13198, new_AGEMA_signal_13195}), .clk (clk), .r ({Fresh[1173], Fresh[1172]}), .c ({new_AGEMA_signal_6500, SubBytesIns_Inst_Sbox_14_M60}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M61_U1 ( .a ({new_AGEMA_signal_6490, SubBytesIns_Inst_Sbox_14_M42}), .b ({new_AGEMA_signal_13204, new_AGEMA_signal_13201}), .clk (clk), .r ({Fresh[1175], Fresh[1174]}), .c ({new_AGEMA_signal_6736, SubBytesIns_Inst_Sbox_14_M61}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M62_U1 ( .a ({new_AGEMA_signal_6729, SubBytesIns_Inst_Sbox_14_M45}), .b ({new_AGEMA_signal_13210, new_AGEMA_signal_13207}), .clk (clk), .r ({Fresh[1177], Fresh[1176]}), .c ({new_AGEMA_signal_6934, SubBytesIns_Inst_Sbox_14_M62}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M63_U1 ( .a ({new_AGEMA_signal_6489, SubBytesIns_Inst_Sbox_14_M41}), .b ({new_AGEMA_signal_13216, new_AGEMA_signal_13213}), .clk (clk), .r ({Fresh[1179], Fresh[1178]}), .c ({new_AGEMA_signal_6737, SubBytesIns_Inst_Sbox_14_M63}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L0_U1 ( .a ({new_AGEMA_signal_6736, SubBytesIns_Inst_Sbox_14_M61}), .b ({new_AGEMA_signal_6934, SubBytesIns_Inst_Sbox_14_M62}), .c ({new_AGEMA_signal_7115, SubBytesIns_Inst_Sbox_14_L0}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L1_U1 ( .a ({new_AGEMA_signal_6495, SubBytesIns_Inst_Sbox_14_M50}), .b ({new_AGEMA_signal_6497, SubBytesIns_Inst_Sbox_14_M56}), .c ({new_AGEMA_signal_6738, SubBytesIns_Inst_Sbox_14_L1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L2_U1 ( .a ({new_AGEMA_signal_6730, SubBytesIns_Inst_Sbox_14_M46}), .b ({new_AGEMA_signal_6494, SubBytesIns_Inst_Sbox_14_M48}), .c ({new_AGEMA_signal_6935, SubBytesIns_Inst_Sbox_14_L2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L3_U1 ( .a ({new_AGEMA_signal_6493, SubBytesIns_Inst_Sbox_14_M47}), .b ({new_AGEMA_signal_6734, SubBytesIns_Inst_Sbox_14_M55}), .c ({new_AGEMA_signal_6936, SubBytesIns_Inst_Sbox_14_L3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L4_U1 ( .a ({new_AGEMA_signal_6733, SubBytesIns_Inst_Sbox_14_M54}), .b ({new_AGEMA_signal_6735, SubBytesIns_Inst_Sbox_14_M58}), .c ({new_AGEMA_signal_6937, SubBytesIns_Inst_Sbox_14_L4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L5_U1 ( .a ({new_AGEMA_signal_6731, SubBytesIns_Inst_Sbox_14_M49}), .b ({new_AGEMA_signal_6736, SubBytesIns_Inst_Sbox_14_M61}), .c ({new_AGEMA_signal_6938, SubBytesIns_Inst_Sbox_14_L5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L6_U1 ( .a ({new_AGEMA_signal_6934, SubBytesIns_Inst_Sbox_14_M62}), .b ({new_AGEMA_signal_6938, SubBytesIns_Inst_Sbox_14_L5}), .c ({new_AGEMA_signal_7116, SubBytesIns_Inst_Sbox_14_L6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L7_U1 ( .a ({new_AGEMA_signal_6730, SubBytesIns_Inst_Sbox_14_M46}), .b ({new_AGEMA_signal_6936, SubBytesIns_Inst_Sbox_14_L3}), .c ({new_AGEMA_signal_7117, SubBytesIns_Inst_Sbox_14_L7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L8_U1 ( .a ({new_AGEMA_signal_6496, SubBytesIns_Inst_Sbox_14_M51}), .b ({new_AGEMA_signal_6499, SubBytesIns_Inst_Sbox_14_M59}), .c ({new_AGEMA_signal_6739, SubBytesIns_Inst_Sbox_14_L8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L9_U1 ( .a ({new_AGEMA_signal_6732, SubBytesIns_Inst_Sbox_14_M52}), .b ({new_AGEMA_signal_6933, SubBytesIns_Inst_Sbox_14_M53}), .c ({new_AGEMA_signal_7118, SubBytesIns_Inst_Sbox_14_L9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L10_U1 ( .a ({new_AGEMA_signal_6933, SubBytesIns_Inst_Sbox_14_M53}), .b ({new_AGEMA_signal_6937, SubBytesIns_Inst_Sbox_14_L4}), .c ({new_AGEMA_signal_7119, SubBytesIns_Inst_Sbox_14_L10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L11_U1 ( .a ({new_AGEMA_signal_6500, SubBytesIns_Inst_Sbox_14_M60}), .b ({new_AGEMA_signal_6935, SubBytesIns_Inst_Sbox_14_L2}), .c ({new_AGEMA_signal_7120, SubBytesIns_Inst_Sbox_14_L11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L12_U1 ( .a ({new_AGEMA_signal_6494, SubBytesIns_Inst_Sbox_14_M48}), .b ({new_AGEMA_signal_6496, SubBytesIns_Inst_Sbox_14_M51}), .c ({new_AGEMA_signal_6740, SubBytesIns_Inst_Sbox_14_L12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L13_U1 ( .a ({new_AGEMA_signal_6495, SubBytesIns_Inst_Sbox_14_M50}), .b ({new_AGEMA_signal_7115, SubBytesIns_Inst_Sbox_14_L0}), .c ({new_AGEMA_signal_7331, SubBytesIns_Inst_Sbox_14_L13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L14_U1 ( .a ({new_AGEMA_signal_6732, SubBytesIns_Inst_Sbox_14_M52}), .b ({new_AGEMA_signal_6736, SubBytesIns_Inst_Sbox_14_M61}), .c ({new_AGEMA_signal_6939, SubBytesIns_Inst_Sbox_14_L14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L15_U1 ( .a ({new_AGEMA_signal_6734, SubBytesIns_Inst_Sbox_14_M55}), .b ({new_AGEMA_signal_6738, SubBytesIns_Inst_Sbox_14_L1}), .c ({new_AGEMA_signal_6940, SubBytesIns_Inst_Sbox_14_L15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L16_U1 ( .a ({new_AGEMA_signal_6497, SubBytesIns_Inst_Sbox_14_M56}), .b ({new_AGEMA_signal_7115, SubBytesIns_Inst_Sbox_14_L0}), .c ({new_AGEMA_signal_7332, SubBytesIns_Inst_Sbox_14_L16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L17_U1 ( .a ({new_AGEMA_signal_6498, SubBytesIns_Inst_Sbox_14_M57}), .b ({new_AGEMA_signal_6738, SubBytesIns_Inst_Sbox_14_L1}), .c ({new_AGEMA_signal_6941, SubBytesIns_Inst_Sbox_14_L17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L18_U1 ( .a ({new_AGEMA_signal_6735, SubBytesIns_Inst_Sbox_14_M58}), .b ({new_AGEMA_signal_6739, SubBytesIns_Inst_Sbox_14_L8}), .c ({new_AGEMA_signal_6942, SubBytesIns_Inst_Sbox_14_L18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L19_U1 ( .a ({new_AGEMA_signal_6737, SubBytesIns_Inst_Sbox_14_M63}), .b ({new_AGEMA_signal_6937, SubBytesIns_Inst_Sbox_14_L4}), .c ({new_AGEMA_signal_7121, SubBytesIns_Inst_Sbox_14_L19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L20_U1 ( .a ({new_AGEMA_signal_7115, SubBytesIns_Inst_Sbox_14_L0}), .b ({new_AGEMA_signal_6738, SubBytesIns_Inst_Sbox_14_L1}), .c ({new_AGEMA_signal_7333, SubBytesIns_Inst_Sbox_14_L20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L21_U1 ( .a ({new_AGEMA_signal_6738, SubBytesIns_Inst_Sbox_14_L1}), .b ({new_AGEMA_signal_7117, SubBytesIns_Inst_Sbox_14_L7}), .c ({new_AGEMA_signal_7334, SubBytesIns_Inst_Sbox_14_L21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L22_U1 ( .a ({new_AGEMA_signal_6936, SubBytesIns_Inst_Sbox_14_L3}), .b ({new_AGEMA_signal_6740, SubBytesIns_Inst_Sbox_14_L12}), .c ({new_AGEMA_signal_7122, SubBytesIns_Inst_Sbox_14_L22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L23_U1 ( .a ({new_AGEMA_signal_6942, SubBytesIns_Inst_Sbox_14_L18}), .b ({new_AGEMA_signal_6935, SubBytesIns_Inst_Sbox_14_L2}), .c ({new_AGEMA_signal_7123, SubBytesIns_Inst_Sbox_14_L23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L24_U1 ( .a ({new_AGEMA_signal_6940, SubBytesIns_Inst_Sbox_14_L15}), .b ({new_AGEMA_signal_7118, SubBytesIns_Inst_Sbox_14_L9}), .c ({new_AGEMA_signal_7335, SubBytesIns_Inst_Sbox_14_L24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L25_U1 ( .a ({new_AGEMA_signal_7116, SubBytesIns_Inst_Sbox_14_L6}), .b ({new_AGEMA_signal_7119, SubBytesIns_Inst_Sbox_14_L10}), .c ({new_AGEMA_signal_7336, SubBytesIns_Inst_Sbox_14_L25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L26_U1 ( .a ({new_AGEMA_signal_7117, SubBytesIns_Inst_Sbox_14_L7}), .b ({new_AGEMA_signal_7118, SubBytesIns_Inst_Sbox_14_L9}), .c ({new_AGEMA_signal_7337, SubBytesIns_Inst_Sbox_14_L26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L27_U1 ( .a ({new_AGEMA_signal_6739, SubBytesIns_Inst_Sbox_14_L8}), .b ({new_AGEMA_signal_7119, SubBytesIns_Inst_Sbox_14_L10}), .c ({new_AGEMA_signal_7338, SubBytesIns_Inst_Sbox_14_L27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L28_U1 ( .a ({new_AGEMA_signal_7120, SubBytesIns_Inst_Sbox_14_L11}), .b ({new_AGEMA_signal_6939, SubBytesIns_Inst_Sbox_14_L14}), .c ({new_AGEMA_signal_7339, SubBytesIns_Inst_Sbox_14_L28}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L29_U1 ( .a ({new_AGEMA_signal_7120, SubBytesIns_Inst_Sbox_14_L11}), .b ({new_AGEMA_signal_6941, SubBytesIns_Inst_Sbox_14_L17}), .c ({new_AGEMA_signal_7340, SubBytesIns_Inst_Sbox_14_L29}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_S0_U1 ( .a ({new_AGEMA_signal_7116, SubBytesIns_Inst_Sbox_14_L6}), .b ({new_AGEMA_signal_7335, SubBytesIns_Inst_Sbox_14_L24}), .c ({new_AGEMA_signal_7483, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_S1_U1 ( .a ({new_AGEMA_signal_7332, SubBytesIns_Inst_Sbox_14_L16}), .b ({new_AGEMA_signal_7337, SubBytesIns_Inst_Sbox_14_L26}), .c ({new_AGEMA_signal_7484, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_S2_U1 ( .a ({new_AGEMA_signal_7121, SubBytesIns_Inst_Sbox_14_L19}), .b ({new_AGEMA_signal_7339, SubBytesIns_Inst_Sbox_14_L28}), .c ({new_AGEMA_signal_7485, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_S3_U1 ( .a ({new_AGEMA_signal_7116, SubBytesIns_Inst_Sbox_14_L6}), .b ({new_AGEMA_signal_7334, SubBytesIns_Inst_Sbox_14_L21}), .c ({new_AGEMA_signal_7486, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_S4_U1 ( .a ({new_AGEMA_signal_7333, SubBytesIns_Inst_Sbox_14_L20}), .b ({new_AGEMA_signal_7122, SubBytesIns_Inst_Sbox_14_L22}), .c ({new_AGEMA_signal_7487, MixColumnsInput[19]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_S5_U1 ( .a ({new_AGEMA_signal_7336, SubBytesIns_Inst_Sbox_14_L25}), .b ({new_AGEMA_signal_7340, SubBytesIns_Inst_Sbox_14_L29}), .c ({new_AGEMA_signal_7488, MixColumnsInput[18]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_S6_U1 ( .a ({new_AGEMA_signal_7331, SubBytesIns_Inst_Sbox_14_L13}), .b ({new_AGEMA_signal_7338, SubBytesIns_Inst_Sbox_14_L27}), .c ({new_AGEMA_signal_7489, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_S7_U1 ( .a ({new_AGEMA_signal_7116, SubBytesIns_Inst_Sbox_14_L6}), .b ({new_AGEMA_signal_7123, SubBytesIns_Inst_Sbox_14_L23}), .c ({new_AGEMA_signal_7341, MixColumnsInput[16]}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M46_U1 ( .a ({new_AGEMA_signal_6504, SubBytesIns_Inst_Sbox_15_M44}), .b ({new_AGEMA_signal_13222, new_AGEMA_signal_13219}), .clk (clk), .r ({Fresh[1181], Fresh[1180]}), .c ({new_AGEMA_signal_6742, SubBytesIns_Inst_Sbox_15_M46}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M47_U1 ( .a ({new_AGEMA_signal_6272, SubBytesIns_Inst_Sbox_15_M40}), .b ({new_AGEMA_signal_13228, new_AGEMA_signal_13225}), .clk (clk), .r ({Fresh[1183], Fresh[1182]}), .c ({new_AGEMA_signal_6505, SubBytesIns_Inst_Sbox_15_M47}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M48_U1 ( .a ({new_AGEMA_signal_6271, SubBytesIns_Inst_Sbox_15_M39}), .b ({new_AGEMA_signal_13234, new_AGEMA_signal_13231}), .clk (clk), .r ({Fresh[1185], Fresh[1184]}), .c ({new_AGEMA_signal_6506, SubBytesIns_Inst_Sbox_15_M48}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M49_U1 ( .a ({new_AGEMA_signal_6503, SubBytesIns_Inst_Sbox_15_M43}), .b ({new_AGEMA_signal_13240, new_AGEMA_signal_13237}), .clk (clk), .r ({Fresh[1187], Fresh[1186]}), .c ({new_AGEMA_signal_6743, SubBytesIns_Inst_Sbox_15_M49}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M50_U1 ( .a ({new_AGEMA_signal_6270, SubBytesIns_Inst_Sbox_15_M38}), .b ({new_AGEMA_signal_13246, new_AGEMA_signal_13243}), .clk (clk), .r ({Fresh[1189], Fresh[1188]}), .c ({new_AGEMA_signal_6507, SubBytesIns_Inst_Sbox_15_M50}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M51_U1 ( .a ({new_AGEMA_signal_6269, SubBytesIns_Inst_Sbox_15_M37}), .b ({new_AGEMA_signal_13252, new_AGEMA_signal_13249}), .clk (clk), .r ({Fresh[1191], Fresh[1190]}), .c ({new_AGEMA_signal_6508, SubBytesIns_Inst_Sbox_15_M51}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M52_U1 ( .a ({new_AGEMA_signal_6502, SubBytesIns_Inst_Sbox_15_M42}), .b ({new_AGEMA_signal_13258, new_AGEMA_signal_13255}), .clk (clk), .r ({Fresh[1193], Fresh[1192]}), .c ({new_AGEMA_signal_6744, SubBytesIns_Inst_Sbox_15_M52}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M53_U1 ( .a ({new_AGEMA_signal_6741, SubBytesIns_Inst_Sbox_15_M45}), .b ({new_AGEMA_signal_13264, new_AGEMA_signal_13261}), .clk (clk), .r ({Fresh[1195], Fresh[1194]}), .c ({new_AGEMA_signal_6943, SubBytesIns_Inst_Sbox_15_M53}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M54_U1 ( .a ({new_AGEMA_signal_6501, SubBytesIns_Inst_Sbox_15_M41}), .b ({new_AGEMA_signal_13270, new_AGEMA_signal_13267}), .clk (clk), .r ({Fresh[1197], Fresh[1196]}), .c ({new_AGEMA_signal_6745, SubBytesIns_Inst_Sbox_15_M54}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M55_U1 ( .a ({new_AGEMA_signal_6504, SubBytesIns_Inst_Sbox_15_M44}), .b ({new_AGEMA_signal_13276, new_AGEMA_signal_13273}), .clk (clk), .r ({Fresh[1199], Fresh[1198]}), .c ({new_AGEMA_signal_6746, SubBytesIns_Inst_Sbox_15_M55}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M56_U1 ( .a ({new_AGEMA_signal_6272, SubBytesIns_Inst_Sbox_15_M40}), .b ({new_AGEMA_signal_13282, new_AGEMA_signal_13279}), .clk (clk), .r ({Fresh[1201], Fresh[1200]}), .c ({new_AGEMA_signal_6509, SubBytesIns_Inst_Sbox_15_M56}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M57_U1 ( .a ({new_AGEMA_signal_6271, SubBytesIns_Inst_Sbox_15_M39}), .b ({new_AGEMA_signal_13288, new_AGEMA_signal_13285}), .clk (clk), .r ({Fresh[1203], Fresh[1202]}), .c ({new_AGEMA_signal_6510, SubBytesIns_Inst_Sbox_15_M57}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M58_U1 ( .a ({new_AGEMA_signal_6503, SubBytesIns_Inst_Sbox_15_M43}), .b ({new_AGEMA_signal_13294, new_AGEMA_signal_13291}), .clk (clk), .r ({Fresh[1205], Fresh[1204]}), .c ({new_AGEMA_signal_6747, SubBytesIns_Inst_Sbox_15_M58}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M59_U1 ( .a ({new_AGEMA_signal_6270, SubBytesIns_Inst_Sbox_15_M38}), .b ({new_AGEMA_signal_13300, new_AGEMA_signal_13297}), .clk (clk), .r ({Fresh[1207], Fresh[1206]}), .c ({new_AGEMA_signal_6511, SubBytesIns_Inst_Sbox_15_M59}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M60_U1 ( .a ({new_AGEMA_signal_6269, SubBytesIns_Inst_Sbox_15_M37}), .b ({new_AGEMA_signal_13306, new_AGEMA_signal_13303}), .clk (clk), .r ({Fresh[1209], Fresh[1208]}), .c ({new_AGEMA_signal_6512, SubBytesIns_Inst_Sbox_15_M60}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M61_U1 ( .a ({new_AGEMA_signal_6502, SubBytesIns_Inst_Sbox_15_M42}), .b ({new_AGEMA_signal_13312, new_AGEMA_signal_13309}), .clk (clk), .r ({Fresh[1211], Fresh[1210]}), .c ({new_AGEMA_signal_6748, SubBytesIns_Inst_Sbox_15_M61}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M62_U1 ( .a ({new_AGEMA_signal_6741, SubBytesIns_Inst_Sbox_15_M45}), .b ({new_AGEMA_signal_13318, new_AGEMA_signal_13315}), .clk (clk), .r ({Fresh[1213], Fresh[1212]}), .c ({new_AGEMA_signal_6944, SubBytesIns_Inst_Sbox_15_M62}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M63_U1 ( .a ({new_AGEMA_signal_6501, SubBytesIns_Inst_Sbox_15_M41}), .b ({new_AGEMA_signal_13324, new_AGEMA_signal_13321}), .clk (clk), .r ({Fresh[1215], Fresh[1214]}), .c ({new_AGEMA_signal_6749, SubBytesIns_Inst_Sbox_15_M63}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L0_U1 ( .a ({new_AGEMA_signal_6748, SubBytesIns_Inst_Sbox_15_M61}), .b ({new_AGEMA_signal_6944, SubBytesIns_Inst_Sbox_15_M62}), .c ({new_AGEMA_signal_7124, SubBytesIns_Inst_Sbox_15_L0}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L1_U1 ( .a ({new_AGEMA_signal_6507, SubBytesIns_Inst_Sbox_15_M50}), .b ({new_AGEMA_signal_6509, SubBytesIns_Inst_Sbox_15_M56}), .c ({new_AGEMA_signal_6750, SubBytesIns_Inst_Sbox_15_L1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L2_U1 ( .a ({new_AGEMA_signal_6742, SubBytesIns_Inst_Sbox_15_M46}), .b ({new_AGEMA_signal_6506, SubBytesIns_Inst_Sbox_15_M48}), .c ({new_AGEMA_signal_6945, SubBytesIns_Inst_Sbox_15_L2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L3_U1 ( .a ({new_AGEMA_signal_6505, SubBytesIns_Inst_Sbox_15_M47}), .b ({new_AGEMA_signal_6746, SubBytesIns_Inst_Sbox_15_M55}), .c ({new_AGEMA_signal_6946, SubBytesIns_Inst_Sbox_15_L3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L4_U1 ( .a ({new_AGEMA_signal_6745, SubBytesIns_Inst_Sbox_15_M54}), .b ({new_AGEMA_signal_6747, SubBytesIns_Inst_Sbox_15_M58}), .c ({new_AGEMA_signal_6947, SubBytesIns_Inst_Sbox_15_L4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L5_U1 ( .a ({new_AGEMA_signal_6743, SubBytesIns_Inst_Sbox_15_M49}), .b ({new_AGEMA_signal_6748, SubBytesIns_Inst_Sbox_15_M61}), .c ({new_AGEMA_signal_6948, SubBytesIns_Inst_Sbox_15_L5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L6_U1 ( .a ({new_AGEMA_signal_6944, SubBytesIns_Inst_Sbox_15_M62}), .b ({new_AGEMA_signal_6948, SubBytesIns_Inst_Sbox_15_L5}), .c ({new_AGEMA_signal_7125, SubBytesIns_Inst_Sbox_15_L6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L7_U1 ( .a ({new_AGEMA_signal_6742, SubBytesIns_Inst_Sbox_15_M46}), .b ({new_AGEMA_signal_6946, SubBytesIns_Inst_Sbox_15_L3}), .c ({new_AGEMA_signal_7126, SubBytesIns_Inst_Sbox_15_L7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L8_U1 ( .a ({new_AGEMA_signal_6508, SubBytesIns_Inst_Sbox_15_M51}), .b ({new_AGEMA_signal_6511, SubBytesIns_Inst_Sbox_15_M59}), .c ({new_AGEMA_signal_6751, SubBytesIns_Inst_Sbox_15_L8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L9_U1 ( .a ({new_AGEMA_signal_6744, SubBytesIns_Inst_Sbox_15_M52}), .b ({new_AGEMA_signal_6943, SubBytesIns_Inst_Sbox_15_M53}), .c ({new_AGEMA_signal_7127, SubBytesIns_Inst_Sbox_15_L9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L10_U1 ( .a ({new_AGEMA_signal_6943, SubBytesIns_Inst_Sbox_15_M53}), .b ({new_AGEMA_signal_6947, SubBytesIns_Inst_Sbox_15_L4}), .c ({new_AGEMA_signal_7128, SubBytesIns_Inst_Sbox_15_L10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L11_U1 ( .a ({new_AGEMA_signal_6512, SubBytesIns_Inst_Sbox_15_M60}), .b ({new_AGEMA_signal_6945, SubBytesIns_Inst_Sbox_15_L2}), .c ({new_AGEMA_signal_7129, SubBytesIns_Inst_Sbox_15_L11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L12_U1 ( .a ({new_AGEMA_signal_6506, SubBytesIns_Inst_Sbox_15_M48}), .b ({new_AGEMA_signal_6508, SubBytesIns_Inst_Sbox_15_M51}), .c ({new_AGEMA_signal_6752, SubBytesIns_Inst_Sbox_15_L12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L13_U1 ( .a ({new_AGEMA_signal_6507, SubBytesIns_Inst_Sbox_15_M50}), .b ({new_AGEMA_signal_7124, SubBytesIns_Inst_Sbox_15_L0}), .c ({new_AGEMA_signal_7342, SubBytesIns_Inst_Sbox_15_L13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L14_U1 ( .a ({new_AGEMA_signal_6744, SubBytesIns_Inst_Sbox_15_M52}), .b ({new_AGEMA_signal_6748, SubBytesIns_Inst_Sbox_15_M61}), .c ({new_AGEMA_signal_6949, SubBytesIns_Inst_Sbox_15_L14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L15_U1 ( .a ({new_AGEMA_signal_6746, SubBytesIns_Inst_Sbox_15_M55}), .b ({new_AGEMA_signal_6750, SubBytesIns_Inst_Sbox_15_L1}), .c ({new_AGEMA_signal_6950, SubBytesIns_Inst_Sbox_15_L15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L16_U1 ( .a ({new_AGEMA_signal_6509, SubBytesIns_Inst_Sbox_15_M56}), .b ({new_AGEMA_signal_7124, SubBytesIns_Inst_Sbox_15_L0}), .c ({new_AGEMA_signal_7343, SubBytesIns_Inst_Sbox_15_L16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L17_U1 ( .a ({new_AGEMA_signal_6510, SubBytesIns_Inst_Sbox_15_M57}), .b ({new_AGEMA_signal_6750, SubBytesIns_Inst_Sbox_15_L1}), .c ({new_AGEMA_signal_6951, SubBytesIns_Inst_Sbox_15_L17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L18_U1 ( .a ({new_AGEMA_signal_6747, SubBytesIns_Inst_Sbox_15_M58}), .b ({new_AGEMA_signal_6751, SubBytesIns_Inst_Sbox_15_L8}), .c ({new_AGEMA_signal_6952, SubBytesIns_Inst_Sbox_15_L18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L19_U1 ( .a ({new_AGEMA_signal_6749, SubBytesIns_Inst_Sbox_15_M63}), .b ({new_AGEMA_signal_6947, SubBytesIns_Inst_Sbox_15_L4}), .c ({new_AGEMA_signal_7130, SubBytesIns_Inst_Sbox_15_L19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L20_U1 ( .a ({new_AGEMA_signal_7124, SubBytesIns_Inst_Sbox_15_L0}), .b ({new_AGEMA_signal_6750, SubBytesIns_Inst_Sbox_15_L1}), .c ({new_AGEMA_signal_7344, SubBytesIns_Inst_Sbox_15_L20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L21_U1 ( .a ({new_AGEMA_signal_6750, SubBytesIns_Inst_Sbox_15_L1}), .b ({new_AGEMA_signal_7126, SubBytesIns_Inst_Sbox_15_L7}), .c ({new_AGEMA_signal_7345, SubBytesIns_Inst_Sbox_15_L21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L22_U1 ( .a ({new_AGEMA_signal_6946, SubBytesIns_Inst_Sbox_15_L3}), .b ({new_AGEMA_signal_6752, SubBytesIns_Inst_Sbox_15_L12}), .c ({new_AGEMA_signal_7131, SubBytesIns_Inst_Sbox_15_L22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L23_U1 ( .a ({new_AGEMA_signal_6952, SubBytesIns_Inst_Sbox_15_L18}), .b ({new_AGEMA_signal_6945, SubBytesIns_Inst_Sbox_15_L2}), .c ({new_AGEMA_signal_7132, SubBytesIns_Inst_Sbox_15_L23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L24_U1 ( .a ({new_AGEMA_signal_6950, SubBytesIns_Inst_Sbox_15_L15}), .b ({new_AGEMA_signal_7127, SubBytesIns_Inst_Sbox_15_L9}), .c ({new_AGEMA_signal_7346, SubBytesIns_Inst_Sbox_15_L24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L25_U1 ( .a ({new_AGEMA_signal_7125, SubBytesIns_Inst_Sbox_15_L6}), .b ({new_AGEMA_signal_7128, SubBytesIns_Inst_Sbox_15_L10}), .c ({new_AGEMA_signal_7347, SubBytesIns_Inst_Sbox_15_L25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L26_U1 ( .a ({new_AGEMA_signal_7126, SubBytesIns_Inst_Sbox_15_L7}), .b ({new_AGEMA_signal_7127, SubBytesIns_Inst_Sbox_15_L9}), .c ({new_AGEMA_signal_7348, SubBytesIns_Inst_Sbox_15_L26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L27_U1 ( .a ({new_AGEMA_signal_6751, SubBytesIns_Inst_Sbox_15_L8}), .b ({new_AGEMA_signal_7128, SubBytesIns_Inst_Sbox_15_L10}), .c ({new_AGEMA_signal_7349, SubBytesIns_Inst_Sbox_15_L27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L28_U1 ( .a ({new_AGEMA_signal_7129, SubBytesIns_Inst_Sbox_15_L11}), .b ({new_AGEMA_signal_6949, SubBytesIns_Inst_Sbox_15_L14}), .c ({new_AGEMA_signal_7350, SubBytesIns_Inst_Sbox_15_L28}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L29_U1 ( .a ({new_AGEMA_signal_7129, SubBytesIns_Inst_Sbox_15_L11}), .b ({new_AGEMA_signal_6951, SubBytesIns_Inst_Sbox_15_L17}), .c ({new_AGEMA_signal_7351, SubBytesIns_Inst_Sbox_15_L29}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_S0_U1 ( .a ({new_AGEMA_signal_7125, SubBytesIns_Inst_Sbox_15_L6}), .b ({new_AGEMA_signal_7346, SubBytesIns_Inst_Sbox_15_L24}), .c ({new_AGEMA_signal_7490, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_S1_U1 ( .a ({new_AGEMA_signal_7343, SubBytesIns_Inst_Sbox_15_L16}), .b ({new_AGEMA_signal_7348, SubBytesIns_Inst_Sbox_15_L26}), .c ({new_AGEMA_signal_7491, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_S2_U1 ( .a ({new_AGEMA_signal_7130, SubBytesIns_Inst_Sbox_15_L19}), .b ({new_AGEMA_signal_7350, SubBytesIns_Inst_Sbox_15_L28}), .c ({new_AGEMA_signal_7492, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_S3_U1 ( .a ({new_AGEMA_signal_7125, SubBytesIns_Inst_Sbox_15_L6}), .b ({new_AGEMA_signal_7345, SubBytesIns_Inst_Sbox_15_L21}), .c ({new_AGEMA_signal_7493, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_S4_U1 ( .a ({new_AGEMA_signal_7344, SubBytesIns_Inst_Sbox_15_L20}), .b ({new_AGEMA_signal_7131, SubBytesIns_Inst_Sbox_15_L22}), .c ({new_AGEMA_signal_7494, MixColumnsInput[123]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_S5_U1 ( .a ({new_AGEMA_signal_7347, SubBytesIns_Inst_Sbox_15_L25}), .b ({new_AGEMA_signal_7351, SubBytesIns_Inst_Sbox_15_L29}), .c ({new_AGEMA_signal_7495, MixColumnsInput[122]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_S6_U1 ( .a ({new_AGEMA_signal_7342, SubBytesIns_Inst_Sbox_15_L13}), .b ({new_AGEMA_signal_7349, SubBytesIns_Inst_Sbox_15_L27}), .c ({new_AGEMA_signal_7496, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_S7_U1 ( .a ({new_AGEMA_signal_7125, SubBytesIns_Inst_Sbox_15_L6}), .b ({new_AGEMA_signal_7132, SubBytesIns_Inst_Sbox_15_L23}), .c ({new_AGEMA_signal_7352, MixColumnsInput[120]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U96 ( .a ({new_AGEMA_signal_7969, MixColumnsIns_MixOneColumnInst_0_n64}), .b ({new_AGEMA_signal_7461, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]}), .c ({new_AGEMA_signal_8270, MixColumnsOutput[105]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U95 ( .a ({new_AGEMA_signal_7766, MixColumnsIns_MixOneColumnInst_0_n63}), .b ({new_AGEMA_signal_7762, MixColumnsIns_MixOneColumnInst_0_n62}), .c ({new_AGEMA_signal_7969, MixColumnsIns_MixOneColumnInst_0_n64}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U94 ( .a ({new_AGEMA_signal_7745, MixColumnsIns_MixOneColumnInst_0_n61}), .b ({new_AGEMA_signal_7544, MixColumnsIns_MixOneColumnInst_0_n60}), .c ({new_AGEMA_signal_7970, MixColumnsOutput[104]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U93 ( .a ({new_AGEMA_signal_7554, MixColumnsIns_MixOneColumnInst_0_n59}), .b ({new_AGEMA_signal_7297, MixColumnsInput[112]}), .c ({new_AGEMA_signal_7745, MixColumnsIns_MixOneColumnInst_0_n61}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U92 ( .a ({new_AGEMA_signal_7746, MixColumnsIns_MixOneColumnInst_0_n58}), .b ({new_AGEMA_signal_7535, MixColumnsIns_MixOneColumnInst_0_n57}), .c ({new_AGEMA_signal_7971, MixColumnsOutput[103]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U91 ( .a ({new_AGEMA_signal_7546, MixColumnsIns_MixOneColumnInst_0_n56}), .b ({new_AGEMA_signal_7420, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .c ({new_AGEMA_signal_7746, MixColumnsIns_MixOneColumnInst_0_n58}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U90 ( .a ({new_AGEMA_signal_7747, MixColumnsIns_MixOneColumnInst_0_n55}), .b ({new_AGEMA_signal_7536, MixColumnsIns_MixOneColumnInst_0_n54}), .c ({new_AGEMA_signal_7972, MixColumnsOutput[102]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U89 ( .a ({new_AGEMA_signal_7548, MixColumnsIns_MixOneColumnInst_0_n53}), .b ({new_AGEMA_signal_7421, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]}), .c ({new_AGEMA_signal_7747, MixColumnsIns_MixOneColumnInst_0_n55}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U88 ( .a ({new_AGEMA_signal_7748, MixColumnsIns_MixOneColumnInst_0_n52}), .b ({new_AGEMA_signal_7537, MixColumnsIns_MixOneColumnInst_0_n51}), .c ({new_AGEMA_signal_7973, MixColumnsOutput[101]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U87 ( .a ({new_AGEMA_signal_7550, MixColumnsIns_MixOneColumnInst_0_n50}), .b ({new_AGEMA_signal_7422, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]}), .c ({new_AGEMA_signal_7748, MixColumnsIns_MixOneColumnInst_0_n52}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U86 ( .a ({new_AGEMA_signal_7974, MixColumnsIns_MixOneColumnInst_0_n49}), .b ({new_AGEMA_signal_7753, MixColumnsIns_MixOneColumnInst_0_n48}), .c ({new_AGEMA_signal_8271, MixColumnsOutput[100]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U85 ( .a ({new_AGEMA_signal_7772, MixColumnsIns_MixOneColumnInst_0_n47}), .b ({new_AGEMA_signal_7423, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]}), .c ({new_AGEMA_signal_7974, MixColumnsIns_MixOneColumnInst_0_n49}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U84 ( .a ({new_AGEMA_signal_7975, MixColumnsIns_MixOneColumnInst_0_n46}), .b ({new_AGEMA_signal_7754, MixColumnsIns_MixOneColumnInst_0_n45}), .c ({new_AGEMA_signal_8272, MixColumnsOutput[99]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U83 ( .a ({new_AGEMA_signal_7774, MixColumnsIns_MixOneColumnInst_0_n44}), .b ({new_AGEMA_signal_7424, MixColumnsInput[107]}), .c ({new_AGEMA_signal_7975, MixColumnsIns_MixOneColumnInst_0_n46}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U82 ( .a ({new_AGEMA_signal_7749, MixColumnsIns_MixOneColumnInst_0_n43}), .b ({new_AGEMA_signal_7535, MixColumnsIns_MixOneColumnInst_0_n57}), .c ({new_AGEMA_signal_7976, MixColumnsOutput[127]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U81 ( .a ({new_AGEMA_signal_7455, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .b ({new_AGEMA_signal_7491, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]}), .c ({new_AGEMA_signal_7535, MixColumnsIns_MixOneColumnInst_0_n57}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U80 ( .a ({new_AGEMA_signal_7385, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_7539, MixColumnsIns_MixOneColumnInst_0_n42}), .c ({new_AGEMA_signal_7749, MixColumnsIns_MixOneColumnInst_0_n43}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U79 ( .a ({new_AGEMA_signal_7750, MixColumnsIns_MixOneColumnInst_0_n41}), .b ({new_AGEMA_signal_7536, MixColumnsIns_MixOneColumnInst_0_n54}), .c ({new_AGEMA_signal_7977, MixColumnsOutput[126]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U78 ( .a ({new_AGEMA_signal_7456, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]}), .b ({new_AGEMA_signal_7492, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]}), .c ({new_AGEMA_signal_7536, MixColumnsIns_MixOneColumnInst_0_n54}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U77 ( .a ({new_AGEMA_signal_7386, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]}), .b ({new_AGEMA_signal_7540, MixColumnsIns_MixOneColumnInst_0_n40}), .c ({new_AGEMA_signal_7750, MixColumnsIns_MixOneColumnInst_0_n41}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U76 ( .a ({new_AGEMA_signal_7751, MixColumnsIns_MixOneColumnInst_0_n39}), .b ({new_AGEMA_signal_7538, MixColumnsIns_MixOneColumnInst_0_n38}), .c ({new_AGEMA_signal_7978, MixColumnsOutput[98]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U75 ( .a ({new_AGEMA_signal_7552, MixColumnsIns_MixOneColumnInst_0_n37}), .b ({new_AGEMA_signal_7425, MixColumnsInput[106]}), .c ({new_AGEMA_signal_7751, MixColumnsIns_MixOneColumnInst_0_n39}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U74 ( .a ({new_AGEMA_signal_7752, MixColumnsIns_MixOneColumnInst_0_n36}), .b ({new_AGEMA_signal_7537, MixColumnsIns_MixOneColumnInst_0_n51}), .c ({new_AGEMA_signal_7979, MixColumnsOutput[125]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U73 ( .a ({new_AGEMA_signal_7457, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]}), .b ({new_AGEMA_signal_7493, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]}), .c ({new_AGEMA_signal_7537, MixColumnsIns_MixOneColumnInst_0_n51}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U72 ( .a ({new_AGEMA_signal_7387, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]}), .b ({new_AGEMA_signal_7541, MixColumnsIns_MixOneColumnInst_0_n35}), .c ({new_AGEMA_signal_7752, MixColumnsIns_MixOneColumnInst_0_n36}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U71 ( .a ({new_AGEMA_signal_7980, MixColumnsIns_MixOneColumnInst_0_n34}), .b ({new_AGEMA_signal_7753, MixColumnsIns_MixOneColumnInst_0_n48}), .c ({new_AGEMA_signal_8273, MixColumnsOutput[124]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U70 ( .a ({new_AGEMA_signal_7458, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]}), .b ({new_AGEMA_signal_7555, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[28]}), .c ({new_AGEMA_signal_7753, MixColumnsIns_MixOneColumnInst_0_n48}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U69 ( .a ({new_AGEMA_signal_7388, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]}), .b ({new_AGEMA_signal_7760, MixColumnsIns_MixOneColumnInst_0_n33}), .c ({new_AGEMA_signal_7980, MixColumnsIns_MixOneColumnInst_0_n34}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U68 ( .a ({new_AGEMA_signal_7981, MixColumnsIns_MixOneColumnInst_0_n32}), .b ({new_AGEMA_signal_7754, MixColumnsIns_MixOneColumnInst_0_n45}), .c ({new_AGEMA_signal_8274, MixColumnsOutput[123]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U67 ( .a ({new_AGEMA_signal_7459, MixColumnsInput[115]}), .b ({new_AGEMA_signal_7556, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[27]}), .c ({new_AGEMA_signal_7754, MixColumnsIns_MixOneColumnInst_0_n45}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U66 ( .a ({new_AGEMA_signal_7389, MixColumnsInput[99]}), .b ({new_AGEMA_signal_7763, MixColumnsIns_MixOneColumnInst_0_n31}), .c ({new_AGEMA_signal_7981, MixColumnsIns_MixOneColumnInst_0_n32}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U65 ( .a ({new_AGEMA_signal_7755, MixColumnsIns_MixOneColumnInst_0_n30}), .b ({new_AGEMA_signal_7538, MixColumnsIns_MixOneColumnInst_0_n38}), .c ({new_AGEMA_signal_7982, MixColumnsOutput[122]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U64 ( .a ({new_AGEMA_signal_7460, MixColumnsInput[114]}), .b ({new_AGEMA_signal_7496, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]}), .c ({new_AGEMA_signal_7538, MixColumnsIns_MixOneColumnInst_0_n38}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U63 ( .a ({new_AGEMA_signal_7390, MixColumnsInput[98]}), .b ({new_AGEMA_signal_7542, MixColumnsIns_MixOneColumnInst_0_n29}), .c ({new_AGEMA_signal_7755, MixColumnsIns_MixOneColumnInst_0_n30}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U62 ( .a ({new_AGEMA_signal_7983, MixColumnsIns_MixOneColumnInst_0_n28}), .b ({new_AGEMA_signal_7761, MixColumnsIns_MixOneColumnInst_0_n27}), .c ({new_AGEMA_signal_8275, MixColumnsOutput[121]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U61 ( .a ({new_AGEMA_signal_7391, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]}), .b ({new_AGEMA_signal_7765, MixColumnsIns_MixOneColumnInst_0_n26}), .c ({new_AGEMA_signal_7983, MixColumnsIns_MixOneColumnInst_0_n28}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U60 ( .a ({new_AGEMA_signal_7756, MixColumnsIns_MixOneColumnInst_0_n25}), .b ({new_AGEMA_signal_7543, MixColumnsIns_MixOneColumnInst_0_n24}), .c ({new_AGEMA_signal_7984, MixColumnsOutput[120]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U59 ( .a ({new_AGEMA_signal_7553, MixColumnsIns_MixOneColumnInst_0_n23}), .b ({new_AGEMA_signal_7187, MixColumnsInput[96]}), .c ({new_AGEMA_signal_7756, MixColumnsIns_MixOneColumnInst_0_n25}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U58 ( .a ({new_AGEMA_signal_7757, MixColumnsIns_MixOneColumnInst_0_n22}), .b ({new_AGEMA_signal_7539, MixColumnsIns_MixOneColumnInst_0_n42}), .c ({new_AGEMA_signal_7985, MixColumnsOutput[119]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U57 ( .a ({new_AGEMA_signal_7420, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .b ({new_AGEMA_signal_7456, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]}), .c ({new_AGEMA_signal_7539, MixColumnsIns_MixOneColumnInst_0_n42}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U56 ( .a ({new_AGEMA_signal_7490, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .b ({new_AGEMA_signal_7545, MixColumnsIns_MixOneColumnInst_0_n21}), .c ({new_AGEMA_signal_7757, MixColumnsIns_MixOneColumnInst_0_n22}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U55 ( .a ({new_AGEMA_signal_7758, MixColumnsIns_MixOneColumnInst_0_n20}), .b ({new_AGEMA_signal_7540, MixColumnsIns_MixOneColumnInst_0_n40}), .c ({new_AGEMA_signal_7986, MixColumnsOutput[118]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U54 ( .a ({new_AGEMA_signal_7421, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]}), .b ({new_AGEMA_signal_7457, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]}), .c ({new_AGEMA_signal_7540, MixColumnsIns_MixOneColumnInst_0_n40}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U53 ( .a ({new_AGEMA_signal_7491, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]}), .b ({new_AGEMA_signal_7547, MixColumnsIns_MixOneColumnInst_0_n19}), .c ({new_AGEMA_signal_7758, MixColumnsIns_MixOneColumnInst_0_n20}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U52 ( .a ({new_AGEMA_signal_7759, MixColumnsIns_MixOneColumnInst_0_n18}), .b ({new_AGEMA_signal_7541, MixColumnsIns_MixOneColumnInst_0_n35}), .c ({new_AGEMA_signal_7987, MixColumnsOutput[117]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U51 ( .a ({new_AGEMA_signal_7422, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]}), .b ({new_AGEMA_signal_7458, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]}), .c ({new_AGEMA_signal_7541, MixColumnsIns_MixOneColumnInst_0_n35}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U50 ( .a ({new_AGEMA_signal_7492, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]}), .b ({new_AGEMA_signal_7549, MixColumnsIns_MixOneColumnInst_0_n17}), .c ({new_AGEMA_signal_7759, MixColumnsIns_MixOneColumnInst_0_n18}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U49 ( .a ({new_AGEMA_signal_7988, MixColumnsIns_MixOneColumnInst_0_n16}), .b ({new_AGEMA_signal_7760, MixColumnsIns_MixOneColumnInst_0_n33}), .c ({new_AGEMA_signal_8276, MixColumnsOutput[116]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U48 ( .a ({new_AGEMA_signal_7423, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]}), .b ({new_AGEMA_signal_7558, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[20]}), .c ({new_AGEMA_signal_7760, MixColumnsIns_MixOneColumnInst_0_n33}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U47 ( .a ({new_AGEMA_signal_7493, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]}), .b ({new_AGEMA_signal_7771, MixColumnsIns_MixOneColumnInst_0_n15}), .c ({new_AGEMA_signal_7988, MixColumnsIns_MixOneColumnInst_0_n16}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U46 ( .a ({new_AGEMA_signal_7989, MixColumnsIns_MixOneColumnInst_0_n14}), .b ({new_AGEMA_signal_7761, MixColumnsIns_MixOneColumnInst_0_n27}), .c ({new_AGEMA_signal_8277, MixColumnsOutput[97]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U45 ( .a ({new_AGEMA_signal_7461, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]}), .b ({new_AGEMA_signal_7557, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[25]}), .c ({new_AGEMA_signal_7761, MixColumnsIns_MixOneColumnInst_0_n27}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U44 ( .a ({new_AGEMA_signal_7426, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]}), .b ({new_AGEMA_signal_7762, MixColumnsIns_MixOneColumnInst_0_n62}), .c ({new_AGEMA_signal_7989, MixColumnsIns_MixOneColumnInst_0_n14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U43 ( .a ({new_AGEMA_signal_7496, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]}), .b ({new_AGEMA_signal_7566, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[1]}), .c ({new_AGEMA_signal_7762, MixColumnsIns_MixOneColumnInst_0_n62}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U42 ( .a ({new_AGEMA_signal_7990, MixColumnsIns_MixOneColumnInst_0_n13}), .b ({new_AGEMA_signal_7763, MixColumnsIns_MixOneColumnInst_0_n31}), .c ({new_AGEMA_signal_8278, MixColumnsOutput[115]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U41 ( .a ({new_AGEMA_signal_7424, MixColumnsInput[107]}), .b ({new_AGEMA_signal_7559, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[19]}), .c ({new_AGEMA_signal_7763, MixColumnsIns_MixOneColumnInst_0_n31}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U40 ( .a ({new_AGEMA_signal_7494, MixColumnsInput[123]}), .b ({new_AGEMA_signal_7773, MixColumnsIns_MixOneColumnInst_0_n12}), .c ({new_AGEMA_signal_7990, MixColumnsIns_MixOneColumnInst_0_n13}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U39 ( .a ({new_AGEMA_signal_7764, MixColumnsIns_MixOneColumnInst_0_n11}), .b ({new_AGEMA_signal_7542, MixColumnsIns_MixOneColumnInst_0_n29}), .c ({new_AGEMA_signal_7991, MixColumnsOutput[114]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U38 ( .a ({new_AGEMA_signal_7425, MixColumnsInput[106]}), .b ({new_AGEMA_signal_7461, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]}), .c ({new_AGEMA_signal_7542, MixColumnsIns_MixOneColumnInst_0_n29}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U37 ( .a ({new_AGEMA_signal_7495, MixColumnsInput[122]}), .b ({new_AGEMA_signal_7551, MixColumnsIns_MixOneColumnInst_0_n10}), .c ({new_AGEMA_signal_7764, MixColumnsIns_MixOneColumnInst_0_n11}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U36 ( .a ({new_AGEMA_signal_7992, MixColumnsIns_MixOneColumnInst_0_n9}), .b ({new_AGEMA_signal_7765, MixColumnsIns_MixOneColumnInst_0_n26}), .c ({new_AGEMA_signal_8279, MixColumnsOutput[113]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U35 ( .a ({new_AGEMA_signal_7560, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[17]}), .b ({new_AGEMA_signal_7426, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]}), .c ({new_AGEMA_signal_7765, MixColumnsIns_MixOneColumnInst_0_n26}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U34 ( .a ({new_AGEMA_signal_7766, MixColumnsIns_MixOneColumnInst_0_n63}), .b ({new_AGEMA_signal_7496, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]}), .c ({new_AGEMA_signal_7992, MixColumnsIns_MixOneColumnInst_0_n9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U33 ( .a ({new_AGEMA_signal_7563, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[9]}), .b ({new_AGEMA_signal_7391, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]}), .c ({new_AGEMA_signal_7766, MixColumnsIns_MixOneColumnInst_0_n63}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U32 ( .a ({new_AGEMA_signal_7767, MixColumnsIns_MixOneColumnInst_0_n8}), .b ({new_AGEMA_signal_7543, MixColumnsIns_MixOneColumnInst_0_n24}), .c ({new_AGEMA_signal_7993, MixColumnsOutput[112]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U31 ( .a ({new_AGEMA_signal_7242, MixColumnsInput[104]}), .b ({new_AGEMA_signal_7455, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .c ({new_AGEMA_signal_7543, MixColumnsIns_MixOneColumnInst_0_n24}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U30 ( .a ({new_AGEMA_signal_7352, MixColumnsInput[120]}), .b ({new_AGEMA_signal_7544, MixColumnsIns_MixOneColumnInst_0_n60}), .c ({new_AGEMA_signal_7767, MixColumnsIns_MixOneColumnInst_0_n8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U29 ( .a ({new_AGEMA_signal_7420, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .b ({new_AGEMA_signal_7187, MixColumnsInput[96]}), .c ({new_AGEMA_signal_7544, MixColumnsIns_MixOneColumnInst_0_n60}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U28 ( .a ({new_AGEMA_signal_7768, MixColumnsIns_MixOneColumnInst_0_n7}), .b ({new_AGEMA_signal_7545, MixColumnsIns_MixOneColumnInst_0_n21}), .c ({new_AGEMA_signal_7994, MixColumnsOutput[111]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U27 ( .a ({new_AGEMA_signal_7385, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_7421, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]}), .c ({new_AGEMA_signal_7545, MixColumnsIns_MixOneColumnInst_0_n21}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U26 ( .a ({new_AGEMA_signal_7546, MixColumnsIns_MixOneColumnInst_0_n56}), .b ({new_AGEMA_signal_7455, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .c ({new_AGEMA_signal_7768, MixColumnsIns_MixOneColumnInst_0_n7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U25 ( .a ({new_AGEMA_signal_7386, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]}), .b ({new_AGEMA_signal_7490, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .c ({new_AGEMA_signal_7546, MixColumnsIns_MixOneColumnInst_0_n56}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U24 ( .a ({new_AGEMA_signal_7769, MixColumnsIns_MixOneColumnInst_0_n6}), .b ({new_AGEMA_signal_7547, MixColumnsIns_MixOneColumnInst_0_n19}), .c ({new_AGEMA_signal_7995, MixColumnsOutput[110]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U23 ( .a ({new_AGEMA_signal_7386, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]}), .b ({new_AGEMA_signal_7422, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]}), .c ({new_AGEMA_signal_7547, MixColumnsIns_MixOneColumnInst_0_n19}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U22 ( .a ({new_AGEMA_signal_7548, MixColumnsIns_MixOneColumnInst_0_n53}), .b ({new_AGEMA_signal_7456, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]}), .c ({new_AGEMA_signal_7769, MixColumnsIns_MixOneColumnInst_0_n6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U21 ( .a ({new_AGEMA_signal_7387, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]}), .b ({new_AGEMA_signal_7491, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]}), .c ({new_AGEMA_signal_7548, MixColumnsIns_MixOneColumnInst_0_n53}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U20 ( .a ({new_AGEMA_signal_7770, MixColumnsIns_MixOneColumnInst_0_n5}), .b ({new_AGEMA_signal_7549, MixColumnsIns_MixOneColumnInst_0_n17}), .c ({new_AGEMA_signal_7996, MixColumnsOutput[109]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U19 ( .a ({new_AGEMA_signal_7387, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]}), .b ({new_AGEMA_signal_7423, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]}), .c ({new_AGEMA_signal_7549, MixColumnsIns_MixOneColumnInst_0_n17}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U18 ( .a ({new_AGEMA_signal_7550, MixColumnsIns_MixOneColumnInst_0_n50}), .b ({new_AGEMA_signal_7457, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]}), .c ({new_AGEMA_signal_7770, MixColumnsIns_MixOneColumnInst_0_n5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U17 ( .a ({new_AGEMA_signal_7388, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]}), .b ({new_AGEMA_signal_7492, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]}), .c ({new_AGEMA_signal_7550, MixColumnsIns_MixOneColumnInst_0_n50}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U16 ( .a ({new_AGEMA_signal_7997, MixColumnsIns_MixOneColumnInst_0_n4}), .b ({new_AGEMA_signal_7771, MixColumnsIns_MixOneColumnInst_0_n15}), .c ({new_AGEMA_signal_8280, MixColumnsOutput[108]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U15 ( .a ({new_AGEMA_signal_7388, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]}), .b ({new_AGEMA_signal_7561, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[12]}), .c ({new_AGEMA_signal_7771, MixColumnsIns_MixOneColumnInst_0_n15}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U14 ( .a ({new_AGEMA_signal_7772, MixColumnsIns_MixOneColumnInst_0_n47}), .b ({new_AGEMA_signal_7458, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]}), .c ({new_AGEMA_signal_7997, MixColumnsIns_MixOneColumnInst_0_n4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U13 ( .a ({new_AGEMA_signal_7564, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[4]}), .b ({new_AGEMA_signal_7493, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]}), .c ({new_AGEMA_signal_7772, MixColumnsIns_MixOneColumnInst_0_n47}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U12 ( .a ({new_AGEMA_signal_7998, MixColumnsIns_MixOneColumnInst_0_n3}), .b ({new_AGEMA_signal_7773, MixColumnsIns_MixOneColumnInst_0_n12}), .c ({new_AGEMA_signal_8281, MixColumnsOutput[107]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U11 ( .a ({new_AGEMA_signal_7389, MixColumnsInput[99]}), .b ({new_AGEMA_signal_7562, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[11]}), .c ({new_AGEMA_signal_7773, MixColumnsIns_MixOneColumnInst_0_n12}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U10 ( .a ({new_AGEMA_signal_7774, MixColumnsIns_MixOneColumnInst_0_n44}), .b ({new_AGEMA_signal_7459, MixColumnsInput[115]}), .c ({new_AGEMA_signal_7998, MixColumnsIns_MixOneColumnInst_0_n3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U9 ( .a ({new_AGEMA_signal_7565, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[3]}), .b ({new_AGEMA_signal_7494, MixColumnsInput[123]}), .c ({new_AGEMA_signal_7774, MixColumnsIns_MixOneColumnInst_0_n44}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U8 ( .a ({new_AGEMA_signal_7775, MixColumnsIns_MixOneColumnInst_0_n2}), .b ({new_AGEMA_signal_7551, MixColumnsIns_MixOneColumnInst_0_n10}), .c ({new_AGEMA_signal_7999, MixColumnsOutput[106]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U7 ( .a ({new_AGEMA_signal_7390, MixColumnsInput[98]}), .b ({new_AGEMA_signal_7426, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]}), .c ({new_AGEMA_signal_7551, MixColumnsIns_MixOneColumnInst_0_n10}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U6 ( .a ({new_AGEMA_signal_7552, MixColumnsIns_MixOneColumnInst_0_n37}), .b ({new_AGEMA_signal_7460, MixColumnsInput[114]}), .c ({new_AGEMA_signal_7775, MixColumnsIns_MixOneColumnInst_0_n2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U5 ( .a ({new_AGEMA_signal_7391, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]}), .b ({new_AGEMA_signal_7495, MixColumnsInput[122]}), .c ({new_AGEMA_signal_7552, MixColumnsIns_MixOneColumnInst_0_n37}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U4 ( .a ({new_AGEMA_signal_7776, MixColumnsIns_MixOneColumnInst_0_n1}), .b ({new_AGEMA_signal_7242, MixColumnsInput[104]}), .c ({new_AGEMA_signal_8000, MixColumnsOutput[96]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U3 ( .a ({new_AGEMA_signal_7554, MixColumnsIns_MixOneColumnInst_0_n59}), .b ({new_AGEMA_signal_7553, MixColumnsIns_MixOneColumnInst_0_n23}), .c ({new_AGEMA_signal_7776, MixColumnsIns_MixOneColumnInst_0_n1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U2 ( .a ({new_AGEMA_signal_7297, MixColumnsInput[112]}), .b ({new_AGEMA_signal_7490, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .c ({new_AGEMA_signal_7553, MixColumnsIns_MixOneColumnInst_0_n23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U1 ( .a ({new_AGEMA_signal_7385, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_7352, MixColumnsInput[120]}), .c ({new_AGEMA_signal_7554, MixColumnsIns_MixOneColumnInst_0_n59}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_0_U3 ( .a ({new_AGEMA_signal_7490, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .b ({new_AGEMA_signal_7494, MixColumnsInput[123]}), .c ({new_AGEMA_signal_7555, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[28]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_0_U2 ( .a ({new_AGEMA_signal_7490, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .b ({new_AGEMA_signal_7495, MixColumnsInput[122]}), .c ({new_AGEMA_signal_7556, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[27]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_0_U1 ( .a ({new_AGEMA_signal_7490, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .b ({new_AGEMA_signal_7352, MixColumnsInput[120]}), .c ({new_AGEMA_signal_7557, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[25]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_1_U3 ( .a ({new_AGEMA_signal_7455, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .b ({new_AGEMA_signal_7459, MixColumnsInput[115]}), .c ({new_AGEMA_signal_7558, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[20]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_1_U2 ( .a ({new_AGEMA_signal_7455, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .b ({new_AGEMA_signal_7460, MixColumnsInput[114]}), .c ({new_AGEMA_signal_7559, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[19]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_1_U1 ( .a ({new_AGEMA_signal_7455, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .b ({new_AGEMA_signal_7297, MixColumnsInput[112]}), .c ({new_AGEMA_signal_7560, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[17]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_2_U3 ( .a ({new_AGEMA_signal_7420, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .b ({new_AGEMA_signal_7424, MixColumnsInput[107]}), .c ({new_AGEMA_signal_7561, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[12]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_2_U2 ( .a ({new_AGEMA_signal_7420, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .b ({new_AGEMA_signal_7425, MixColumnsInput[106]}), .c ({new_AGEMA_signal_7562, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[11]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_2_U1 ( .a ({new_AGEMA_signal_7420, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .b ({new_AGEMA_signal_7242, MixColumnsInput[104]}), .c ({new_AGEMA_signal_7563, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[9]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_3_U3 ( .a ({new_AGEMA_signal_7385, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_7389, MixColumnsInput[99]}), .c ({new_AGEMA_signal_7564, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[4]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_3_U2 ( .a ({new_AGEMA_signal_7385, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_7390, MixColumnsInput[98]}), .c ({new_AGEMA_signal_7565, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[3]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_3_U1 ( .a ({new_AGEMA_signal_7385, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_7187, MixColumnsInput[96]}), .c ({new_AGEMA_signal_7566, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[1]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U96 ( .a ({new_AGEMA_signal_8001, MixColumnsIns_MixOneColumnInst_1_n64}), .b ({new_AGEMA_signal_7433, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]}), .c ({new_AGEMA_signal_8282, MixColumnsOutput[73]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U95 ( .a ({new_AGEMA_signal_7798, MixColumnsIns_MixOneColumnInst_1_n63}), .b ({new_AGEMA_signal_7794, MixColumnsIns_MixOneColumnInst_1_n62}), .c ({new_AGEMA_signal_8001, MixColumnsIns_MixOneColumnInst_1_n64}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U94 ( .a ({new_AGEMA_signal_7777, MixColumnsIns_MixOneColumnInst_1_n61}), .b ({new_AGEMA_signal_7576, MixColumnsIns_MixOneColumnInst_1_n60}), .c ({new_AGEMA_signal_8002, MixColumnsOutput[72]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U93 ( .a ({new_AGEMA_signal_7586, MixColumnsIns_MixOneColumnInst_1_n59}), .b ({new_AGEMA_signal_7253, MixColumnsInput[80]}), .c ({new_AGEMA_signal_7777, MixColumnsIns_MixOneColumnInst_1_n61}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U92 ( .a ({new_AGEMA_signal_7778, MixColumnsIns_MixOneColumnInst_1_n58}), .b ({new_AGEMA_signal_7567, MixColumnsIns_MixOneColumnInst_1_n57}), .c ({new_AGEMA_signal_8003, MixColumnsOutput[71]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U91 ( .a ({new_AGEMA_signal_7578, MixColumnsIns_MixOneColumnInst_1_n56}), .b ({new_AGEMA_signal_7392, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .c ({new_AGEMA_signal_7778, MixColumnsIns_MixOneColumnInst_1_n58}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U90 ( .a ({new_AGEMA_signal_7779, MixColumnsIns_MixOneColumnInst_1_n55}), .b ({new_AGEMA_signal_7568, MixColumnsIns_MixOneColumnInst_1_n54}), .c ({new_AGEMA_signal_8004, MixColumnsOutput[70]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U89 ( .a ({new_AGEMA_signal_7580, MixColumnsIns_MixOneColumnInst_1_n53}), .b ({new_AGEMA_signal_7393, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]}), .c ({new_AGEMA_signal_7779, MixColumnsIns_MixOneColumnInst_1_n55}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U88 ( .a ({new_AGEMA_signal_7780, MixColumnsIns_MixOneColumnInst_1_n52}), .b ({new_AGEMA_signal_7569, MixColumnsIns_MixOneColumnInst_1_n51}), .c ({new_AGEMA_signal_8005, MixColumnsOutput[69]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U87 ( .a ({new_AGEMA_signal_7582, MixColumnsIns_MixOneColumnInst_1_n50}), .b ({new_AGEMA_signal_7394, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]}), .c ({new_AGEMA_signal_7780, MixColumnsIns_MixOneColumnInst_1_n52}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U86 ( .a ({new_AGEMA_signal_8006, MixColumnsIns_MixOneColumnInst_1_n49}), .b ({new_AGEMA_signal_7785, MixColumnsIns_MixOneColumnInst_1_n48}), .c ({new_AGEMA_signal_8283, MixColumnsOutput[68]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U85 ( .a ({new_AGEMA_signal_7804, MixColumnsIns_MixOneColumnInst_1_n47}), .b ({new_AGEMA_signal_7395, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]}), .c ({new_AGEMA_signal_8006, MixColumnsIns_MixOneColumnInst_1_n49}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U84 ( .a ({new_AGEMA_signal_8007, MixColumnsIns_MixOneColumnInst_1_n46}), .b ({new_AGEMA_signal_7786, MixColumnsIns_MixOneColumnInst_1_n45}), .c ({new_AGEMA_signal_8284, MixColumnsOutput[67]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U83 ( .a ({new_AGEMA_signal_7806, MixColumnsIns_MixOneColumnInst_1_n44}), .b ({new_AGEMA_signal_7396, MixColumnsInput[75]}), .c ({new_AGEMA_signal_8007, MixColumnsIns_MixOneColumnInst_1_n46}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U82 ( .a ({new_AGEMA_signal_7781, MixColumnsIns_MixOneColumnInst_1_n43}), .b ({new_AGEMA_signal_7567, MixColumnsIns_MixOneColumnInst_1_n57}), .c ({new_AGEMA_signal_8008, MixColumnsOutput[95]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U81 ( .a ({new_AGEMA_signal_7427, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .b ({new_AGEMA_signal_7463, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]}), .c ({new_AGEMA_signal_7567, MixColumnsIns_MixOneColumnInst_1_n57}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U80 ( .a ({new_AGEMA_signal_7469, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_7571, MixColumnsIns_MixOneColumnInst_1_n42}), .c ({new_AGEMA_signal_7781, MixColumnsIns_MixOneColumnInst_1_n43}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U79 ( .a ({new_AGEMA_signal_7782, MixColumnsIns_MixOneColumnInst_1_n41}), .b ({new_AGEMA_signal_7568, MixColumnsIns_MixOneColumnInst_1_n54}), .c ({new_AGEMA_signal_8009, MixColumnsOutput[94]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U78 ( .a ({new_AGEMA_signal_7428, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]}), .b ({new_AGEMA_signal_7464, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]}), .c ({new_AGEMA_signal_7568, MixColumnsIns_MixOneColumnInst_1_n54}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U77 ( .a ({new_AGEMA_signal_7470, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]}), .b ({new_AGEMA_signal_7572, MixColumnsIns_MixOneColumnInst_1_n40}), .c ({new_AGEMA_signal_7782, MixColumnsIns_MixOneColumnInst_1_n41}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U76 ( .a ({new_AGEMA_signal_7783, MixColumnsIns_MixOneColumnInst_1_n39}), .b ({new_AGEMA_signal_7570, MixColumnsIns_MixOneColumnInst_1_n38}), .c ({new_AGEMA_signal_8010, MixColumnsOutput[66]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U75 ( .a ({new_AGEMA_signal_7584, MixColumnsIns_MixOneColumnInst_1_n37}), .b ({new_AGEMA_signal_7397, MixColumnsInput[74]}), .c ({new_AGEMA_signal_7783, MixColumnsIns_MixOneColumnInst_1_n39}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U74 ( .a ({new_AGEMA_signal_7784, MixColumnsIns_MixOneColumnInst_1_n36}), .b ({new_AGEMA_signal_7569, MixColumnsIns_MixOneColumnInst_1_n51}), .c ({new_AGEMA_signal_8011, MixColumnsOutput[93]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U73 ( .a ({new_AGEMA_signal_7429, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]}), .b ({new_AGEMA_signal_7465, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]}), .c ({new_AGEMA_signal_7569, MixColumnsIns_MixOneColumnInst_1_n51}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U72 ( .a ({new_AGEMA_signal_7471, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]}), .b ({new_AGEMA_signal_7573, MixColumnsIns_MixOneColumnInst_1_n35}), .c ({new_AGEMA_signal_7784, MixColumnsIns_MixOneColumnInst_1_n36}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U71 ( .a ({new_AGEMA_signal_8012, MixColumnsIns_MixOneColumnInst_1_n34}), .b ({new_AGEMA_signal_7785, MixColumnsIns_MixOneColumnInst_1_n48}), .c ({new_AGEMA_signal_8285, MixColumnsOutput[92]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U70 ( .a ({new_AGEMA_signal_7430, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]}), .b ({new_AGEMA_signal_7587, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[28]}), .c ({new_AGEMA_signal_7785, MixColumnsIns_MixOneColumnInst_1_n48}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U69 ( .a ({new_AGEMA_signal_7472, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]}), .b ({new_AGEMA_signal_7792, MixColumnsIns_MixOneColumnInst_1_n33}), .c ({new_AGEMA_signal_8012, MixColumnsIns_MixOneColumnInst_1_n34}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U68 ( .a ({new_AGEMA_signal_8013, MixColumnsIns_MixOneColumnInst_1_n32}), .b ({new_AGEMA_signal_7786, MixColumnsIns_MixOneColumnInst_1_n45}), .c ({new_AGEMA_signal_8286, MixColumnsOutput[91]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U67 ( .a ({new_AGEMA_signal_7431, MixColumnsInput[83]}), .b ({new_AGEMA_signal_7588, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[27]}), .c ({new_AGEMA_signal_7786, MixColumnsIns_MixOneColumnInst_1_n45}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U66 ( .a ({new_AGEMA_signal_7473, MixColumnsInput[67]}), .b ({new_AGEMA_signal_7795, MixColumnsIns_MixOneColumnInst_1_n31}), .c ({new_AGEMA_signal_8013, MixColumnsIns_MixOneColumnInst_1_n32}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U65 ( .a ({new_AGEMA_signal_7787, MixColumnsIns_MixOneColumnInst_1_n30}), .b ({new_AGEMA_signal_7570, MixColumnsIns_MixOneColumnInst_1_n38}), .c ({new_AGEMA_signal_8014, MixColumnsOutput[90]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U64 ( .a ({new_AGEMA_signal_7432, MixColumnsInput[82]}), .b ({new_AGEMA_signal_7468, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]}), .c ({new_AGEMA_signal_7570, MixColumnsIns_MixOneColumnInst_1_n38}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U63 ( .a ({new_AGEMA_signal_7474, MixColumnsInput[66]}), .b ({new_AGEMA_signal_7574, MixColumnsIns_MixOneColumnInst_1_n29}), .c ({new_AGEMA_signal_7787, MixColumnsIns_MixOneColumnInst_1_n30}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U62 ( .a ({new_AGEMA_signal_8015, MixColumnsIns_MixOneColumnInst_1_n28}), .b ({new_AGEMA_signal_7793, MixColumnsIns_MixOneColumnInst_1_n27}), .c ({new_AGEMA_signal_8287, MixColumnsOutput[89]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U61 ( .a ({new_AGEMA_signal_7475, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]}), .b ({new_AGEMA_signal_7797, MixColumnsIns_MixOneColumnInst_1_n26}), .c ({new_AGEMA_signal_8015, MixColumnsIns_MixOneColumnInst_1_n28}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U60 ( .a ({new_AGEMA_signal_7788, MixColumnsIns_MixOneColumnInst_1_n25}), .b ({new_AGEMA_signal_7575, MixColumnsIns_MixOneColumnInst_1_n24}), .c ({new_AGEMA_signal_8016, MixColumnsOutput[88]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U59 ( .a ({new_AGEMA_signal_7585, MixColumnsIns_MixOneColumnInst_1_n23}), .b ({new_AGEMA_signal_7319, MixColumnsInput[64]}), .c ({new_AGEMA_signal_7788, MixColumnsIns_MixOneColumnInst_1_n25}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U58 ( .a ({new_AGEMA_signal_7789, MixColumnsIns_MixOneColumnInst_1_n22}), .b ({new_AGEMA_signal_7571, MixColumnsIns_MixOneColumnInst_1_n42}), .c ({new_AGEMA_signal_8017, MixColumnsOutput[87]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U57 ( .a ({new_AGEMA_signal_7392, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .b ({new_AGEMA_signal_7428, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]}), .c ({new_AGEMA_signal_7571, MixColumnsIns_MixOneColumnInst_1_n42}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U56 ( .a ({new_AGEMA_signal_7462, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .b ({new_AGEMA_signal_7577, MixColumnsIns_MixOneColumnInst_1_n21}), .c ({new_AGEMA_signal_7789, MixColumnsIns_MixOneColumnInst_1_n22}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U55 ( .a ({new_AGEMA_signal_7790, MixColumnsIns_MixOneColumnInst_1_n20}), .b ({new_AGEMA_signal_7572, MixColumnsIns_MixOneColumnInst_1_n40}), .c ({new_AGEMA_signal_8018, MixColumnsOutput[86]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U54 ( .a ({new_AGEMA_signal_7393, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]}), .b ({new_AGEMA_signal_7429, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]}), .c ({new_AGEMA_signal_7572, MixColumnsIns_MixOneColumnInst_1_n40}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U53 ( .a ({new_AGEMA_signal_7463, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]}), .b ({new_AGEMA_signal_7579, MixColumnsIns_MixOneColumnInst_1_n19}), .c ({new_AGEMA_signal_7790, MixColumnsIns_MixOneColumnInst_1_n20}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U52 ( .a ({new_AGEMA_signal_7791, MixColumnsIns_MixOneColumnInst_1_n18}), .b ({new_AGEMA_signal_7573, MixColumnsIns_MixOneColumnInst_1_n35}), .c ({new_AGEMA_signal_8019, MixColumnsOutput[85]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U51 ( .a ({new_AGEMA_signal_7394, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]}), .b ({new_AGEMA_signal_7430, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]}), .c ({new_AGEMA_signal_7573, MixColumnsIns_MixOneColumnInst_1_n35}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U50 ( .a ({new_AGEMA_signal_7464, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]}), .b ({new_AGEMA_signal_7581, MixColumnsIns_MixOneColumnInst_1_n17}), .c ({new_AGEMA_signal_7791, MixColumnsIns_MixOneColumnInst_1_n18}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U49 ( .a ({new_AGEMA_signal_8020, MixColumnsIns_MixOneColumnInst_1_n16}), .b ({new_AGEMA_signal_7792, MixColumnsIns_MixOneColumnInst_1_n33}), .c ({new_AGEMA_signal_8288, MixColumnsOutput[84]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U48 ( .a ({new_AGEMA_signal_7395, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]}), .b ({new_AGEMA_signal_7590, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[20]}), .c ({new_AGEMA_signal_7792, MixColumnsIns_MixOneColumnInst_1_n33}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U47 ( .a ({new_AGEMA_signal_7465, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]}), .b ({new_AGEMA_signal_7803, MixColumnsIns_MixOneColumnInst_1_n15}), .c ({new_AGEMA_signal_8020, MixColumnsIns_MixOneColumnInst_1_n16}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U46 ( .a ({new_AGEMA_signal_8021, MixColumnsIns_MixOneColumnInst_1_n14}), .b ({new_AGEMA_signal_7793, MixColumnsIns_MixOneColumnInst_1_n27}), .c ({new_AGEMA_signal_8289, MixColumnsOutput[65]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U45 ( .a ({new_AGEMA_signal_7433, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]}), .b ({new_AGEMA_signal_7589, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[25]}), .c ({new_AGEMA_signal_7793, MixColumnsIns_MixOneColumnInst_1_n27}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U44 ( .a ({new_AGEMA_signal_7398, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]}), .b ({new_AGEMA_signal_7794, MixColumnsIns_MixOneColumnInst_1_n62}), .c ({new_AGEMA_signal_8021, MixColumnsIns_MixOneColumnInst_1_n14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U43 ( .a ({new_AGEMA_signal_7468, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]}), .b ({new_AGEMA_signal_7598, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[1]}), .c ({new_AGEMA_signal_7794, MixColumnsIns_MixOneColumnInst_1_n62}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U42 ( .a ({new_AGEMA_signal_8022, MixColumnsIns_MixOneColumnInst_1_n13}), .b ({new_AGEMA_signal_7795, MixColumnsIns_MixOneColumnInst_1_n31}), .c ({new_AGEMA_signal_8290, MixColumnsOutput[83]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U41 ( .a ({new_AGEMA_signal_7396, MixColumnsInput[75]}), .b ({new_AGEMA_signal_7591, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[19]}), .c ({new_AGEMA_signal_7795, MixColumnsIns_MixOneColumnInst_1_n31}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U40 ( .a ({new_AGEMA_signal_7466, MixColumnsInput[91]}), .b ({new_AGEMA_signal_7805, MixColumnsIns_MixOneColumnInst_1_n12}), .c ({new_AGEMA_signal_8022, MixColumnsIns_MixOneColumnInst_1_n13}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U39 ( .a ({new_AGEMA_signal_7796, MixColumnsIns_MixOneColumnInst_1_n11}), .b ({new_AGEMA_signal_7574, MixColumnsIns_MixOneColumnInst_1_n29}), .c ({new_AGEMA_signal_8023, MixColumnsOutput[82]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U38 ( .a ({new_AGEMA_signal_7397, MixColumnsInput[74]}), .b ({new_AGEMA_signal_7433, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]}), .c ({new_AGEMA_signal_7574, MixColumnsIns_MixOneColumnInst_1_n29}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U37 ( .a ({new_AGEMA_signal_7467, MixColumnsInput[90]}), .b ({new_AGEMA_signal_7583, MixColumnsIns_MixOneColumnInst_1_n10}), .c ({new_AGEMA_signal_7796, MixColumnsIns_MixOneColumnInst_1_n11}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U36 ( .a ({new_AGEMA_signal_8024, MixColumnsIns_MixOneColumnInst_1_n9}), .b ({new_AGEMA_signal_7797, MixColumnsIns_MixOneColumnInst_1_n26}), .c ({new_AGEMA_signal_8291, MixColumnsOutput[81]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U35 ( .a ({new_AGEMA_signal_7592, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[17]}), .b ({new_AGEMA_signal_7398, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]}), .c ({new_AGEMA_signal_7797, MixColumnsIns_MixOneColumnInst_1_n26}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U34 ( .a ({new_AGEMA_signal_7798, MixColumnsIns_MixOneColumnInst_1_n63}), .b ({new_AGEMA_signal_7468, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]}), .c ({new_AGEMA_signal_8024, MixColumnsIns_MixOneColumnInst_1_n9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U33 ( .a ({new_AGEMA_signal_7595, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[9]}), .b ({new_AGEMA_signal_7475, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]}), .c ({new_AGEMA_signal_7798, MixColumnsIns_MixOneColumnInst_1_n63}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U32 ( .a ({new_AGEMA_signal_7799, MixColumnsIns_MixOneColumnInst_1_n8}), .b ({new_AGEMA_signal_7575, MixColumnsIns_MixOneColumnInst_1_n24}), .c ({new_AGEMA_signal_8025, MixColumnsOutput[80]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U31 ( .a ({new_AGEMA_signal_7198, MixColumnsInput[72]}), .b ({new_AGEMA_signal_7427, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .c ({new_AGEMA_signal_7575, MixColumnsIns_MixOneColumnInst_1_n24}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U30 ( .a ({new_AGEMA_signal_7308, MixColumnsInput[88]}), .b ({new_AGEMA_signal_7576, MixColumnsIns_MixOneColumnInst_1_n60}), .c ({new_AGEMA_signal_7799, MixColumnsIns_MixOneColumnInst_1_n8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U29 ( .a ({new_AGEMA_signal_7392, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .b ({new_AGEMA_signal_7319, MixColumnsInput[64]}), .c ({new_AGEMA_signal_7576, MixColumnsIns_MixOneColumnInst_1_n60}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U28 ( .a ({new_AGEMA_signal_7800, MixColumnsIns_MixOneColumnInst_1_n7}), .b ({new_AGEMA_signal_7577, MixColumnsIns_MixOneColumnInst_1_n21}), .c ({new_AGEMA_signal_8026, MixColumnsOutput[79]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U27 ( .a ({new_AGEMA_signal_7469, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_7393, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]}), .c ({new_AGEMA_signal_7577, MixColumnsIns_MixOneColumnInst_1_n21}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U26 ( .a ({new_AGEMA_signal_7578, MixColumnsIns_MixOneColumnInst_1_n56}), .b ({new_AGEMA_signal_7427, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .c ({new_AGEMA_signal_7800, MixColumnsIns_MixOneColumnInst_1_n7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U25 ( .a ({new_AGEMA_signal_7470, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]}), .b ({new_AGEMA_signal_7462, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .c ({new_AGEMA_signal_7578, MixColumnsIns_MixOneColumnInst_1_n56}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U24 ( .a ({new_AGEMA_signal_7801, MixColumnsIns_MixOneColumnInst_1_n6}), .b ({new_AGEMA_signal_7579, MixColumnsIns_MixOneColumnInst_1_n19}), .c ({new_AGEMA_signal_8027, MixColumnsOutput[78]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U23 ( .a ({new_AGEMA_signal_7470, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]}), .b ({new_AGEMA_signal_7394, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]}), .c ({new_AGEMA_signal_7579, MixColumnsIns_MixOneColumnInst_1_n19}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U22 ( .a ({new_AGEMA_signal_7580, MixColumnsIns_MixOneColumnInst_1_n53}), .b ({new_AGEMA_signal_7428, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]}), .c ({new_AGEMA_signal_7801, MixColumnsIns_MixOneColumnInst_1_n6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U21 ( .a ({new_AGEMA_signal_7471, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]}), .b ({new_AGEMA_signal_7463, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]}), .c ({new_AGEMA_signal_7580, MixColumnsIns_MixOneColumnInst_1_n53}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U20 ( .a ({new_AGEMA_signal_7802, MixColumnsIns_MixOneColumnInst_1_n5}), .b ({new_AGEMA_signal_7581, MixColumnsIns_MixOneColumnInst_1_n17}), .c ({new_AGEMA_signal_8028, MixColumnsOutput[77]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U19 ( .a ({new_AGEMA_signal_7471, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]}), .b ({new_AGEMA_signal_7395, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]}), .c ({new_AGEMA_signal_7581, MixColumnsIns_MixOneColumnInst_1_n17}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U18 ( .a ({new_AGEMA_signal_7582, MixColumnsIns_MixOneColumnInst_1_n50}), .b ({new_AGEMA_signal_7429, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]}), .c ({new_AGEMA_signal_7802, MixColumnsIns_MixOneColumnInst_1_n5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U17 ( .a ({new_AGEMA_signal_7472, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]}), .b ({new_AGEMA_signal_7464, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]}), .c ({new_AGEMA_signal_7582, MixColumnsIns_MixOneColumnInst_1_n50}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U16 ( .a ({new_AGEMA_signal_8029, MixColumnsIns_MixOneColumnInst_1_n4}), .b ({new_AGEMA_signal_7803, MixColumnsIns_MixOneColumnInst_1_n15}), .c ({new_AGEMA_signal_8292, MixColumnsOutput[76]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U15 ( .a ({new_AGEMA_signal_7472, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]}), .b ({new_AGEMA_signal_7593, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[12]}), .c ({new_AGEMA_signal_7803, MixColumnsIns_MixOneColumnInst_1_n15}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U14 ( .a ({new_AGEMA_signal_7804, MixColumnsIns_MixOneColumnInst_1_n47}), .b ({new_AGEMA_signal_7430, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]}), .c ({new_AGEMA_signal_8029, MixColumnsIns_MixOneColumnInst_1_n4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U13 ( .a ({new_AGEMA_signal_7596, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[4]}), .b ({new_AGEMA_signal_7465, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]}), .c ({new_AGEMA_signal_7804, MixColumnsIns_MixOneColumnInst_1_n47}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U12 ( .a ({new_AGEMA_signal_8030, MixColumnsIns_MixOneColumnInst_1_n3}), .b ({new_AGEMA_signal_7805, MixColumnsIns_MixOneColumnInst_1_n12}), .c ({new_AGEMA_signal_8293, MixColumnsOutput[75]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U11 ( .a ({new_AGEMA_signal_7473, MixColumnsInput[67]}), .b ({new_AGEMA_signal_7594, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[11]}), .c ({new_AGEMA_signal_7805, MixColumnsIns_MixOneColumnInst_1_n12}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U10 ( .a ({new_AGEMA_signal_7806, MixColumnsIns_MixOneColumnInst_1_n44}), .b ({new_AGEMA_signal_7431, MixColumnsInput[83]}), .c ({new_AGEMA_signal_8030, MixColumnsIns_MixOneColumnInst_1_n3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U9 ( .a ({new_AGEMA_signal_7597, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[3]}), .b ({new_AGEMA_signal_7466, MixColumnsInput[91]}), .c ({new_AGEMA_signal_7806, MixColumnsIns_MixOneColumnInst_1_n44}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U8 ( .a ({new_AGEMA_signal_7807, MixColumnsIns_MixOneColumnInst_1_n2}), .b ({new_AGEMA_signal_7583, MixColumnsIns_MixOneColumnInst_1_n10}), .c ({new_AGEMA_signal_8031, MixColumnsOutput[74]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U7 ( .a ({new_AGEMA_signal_7474, MixColumnsInput[66]}), .b ({new_AGEMA_signal_7398, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]}), .c ({new_AGEMA_signal_7583, MixColumnsIns_MixOneColumnInst_1_n10}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U6 ( .a ({new_AGEMA_signal_7584, MixColumnsIns_MixOneColumnInst_1_n37}), .b ({new_AGEMA_signal_7432, MixColumnsInput[82]}), .c ({new_AGEMA_signal_7807, MixColumnsIns_MixOneColumnInst_1_n2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U5 ( .a ({new_AGEMA_signal_7475, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]}), .b ({new_AGEMA_signal_7467, MixColumnsInput[90]}), .c ({new_AGEMA_signal_7584, MixColumnsIns_MixOneColumnInst_1_n37}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U4 ( .a ({new_AGEMA_signal_7808, MixColumnsIns_MixOneColumnInst_1_n1}), .b ({new_AGEMA_signal_7198, MixColumnsInput[72]}), .c ({new_AGEMA_signal_8032, MixColumnsOutput[64]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U3 ( .a ({new_AGEMA_signal_7586, MixColumnsIns_MixOneColumnInst_1_n59}), .b ({new_AGEMA_signal_7585, MixColumnsIns_MixOneColumnInst_1_n23}), .c ({new_AGEMA_signal_7808, MixColumnsIns_MixOneColumnInst_1_n1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U2 ( .a ({new_AGEMA_signal_7253, MixColumnsInput[80]}), .b ({new_AGEMA_signal_7462, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .c ({new_AGEMA_signal_7585, MixColumnsIns_MixOneColumnInst_1_n23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U1 ( .a ({new_AGEMA_signal_7469, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_7308, MixColumnsInput[88]}), .c ({new_AGEMA_signal_7586, MixColumnsIns_MixOneColumnInst_1_n59}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_0_U3 ( .a ({new_AGEMA_signal_7462, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .b ({new_AGEMA_signal_7466, MixColumnsInput[91]}), .c ({new_AGEMA_signal_7587, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[28]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_0_U2 ( .a ({new_AGEMA_signal_7462, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .b ({new_AGEMA_signal_7467, MixColumnsInput[90]}), .c ({new_AGEMA_signal_7588, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[27]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_0_U1 ( .a ({new_AGEMA_signal_7462, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .b ({new_AGEMA_signal_7308, MixColumnsInput[88]}), .c ({new_AGEMA_signal_7589, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[25]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_1_U3 ( .a ({new_AGEMA_signal_7427, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .b ({new_AGEMA_signal_7431, MixColumnsInput[83]}), .c ({new_AGEMA_signal_7590, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[20]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_1_U2 ( .a ({new_AGEMA_signal_7427, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .b ({new_AGEMA_signal_7432, MixColumnsInput[82]}), .c ({new_AGEMA_signal_7591, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[19]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_1_U1 ( .a ({new_AGEMA_signal_7427, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .b ({new_AGEMA_signal_7253, MixColumnsInput[80]}), .c ({new_AGEMA_signal_7592, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[17]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_2_U3 ( .a ({new_AGEMA_signal_7392, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .b ({new_AGEMA_signal_7396, MixColumnsInput[75]}), .c ({new_AGEMA_signal_7593, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[12]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_2_U2 ( .a ({new_AGEMA_signal_7392, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .b ({new_AGEMA_signal_7397, MixColumnsInput[74]}), .c ({new_AGEMA_signal_7594, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[11]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_2_U1 ( .a ({new_AGEMA_signal_7392, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .b ({new_AGEMA_signal_7198, MixColumnsInput[72]}), .c ({new_AGEMA_signal_7595, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[9]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_3_U3 ( .a ({new_AGEMA_signal_7469, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_7473, MixColumnsInput[67]}), .c ({new_AGEMA_signal_7596, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[4]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_3_U2 ( .a ({new_AGEMA_signal_7469, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_7474, MixColumnsInput[66]}), .c ({new_AGEMA_signal_7597, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[3]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_3_U1 ( .a ({new_AGEMA_signal_7469, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_7319, MixColumnsInput[64]}), .c ({new_AGEMA_signal_7598, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[1]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U96 ( .a ({new_AGEMA_signal_8033, MixColumnsIns_MixOneColumnInst_2_n64}), .b ({new_AGEMA_signal_7405, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]}), .c ({new_AGEMA_signal_8294, MixColumnsOutput[41]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U95 ( .a ({new_AGEMA_signal_7830, MixColumnsIns_MixOneColumnInst_2_n63}), .b ({new_AGEMA_signal_7826, MixColumnsIns_MixOneColumnInst_2_n62}), .c ({new_AGEMA_signal_8033, MixColumnsIns_MixOneColumnInst_2_n64}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U94 ( .a ({new_AGEMA_signal_7809, MixColumnsIns_MixOneColumnInst_2_n61}), .b ({new_AGEMA_signal_7608, MixColumnsIns_MixOneColumnInst_2_n60}), .c ({new_AGEMA_signal_8034, MixColumnsOutput[40]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U93 ( .a ({new_AGEMA_signal_7618, MixColumnsIns_MixOneColumnInst_2_n59}), .b ({new_AGEMA_signal_7209, MixColumnsInput[48]}), .c ({new_AGEMA_signal_7809, MixColumnsIns_MixOneColumnInst_2_n61}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U92 ( .a ({new_AGEMA_signal_7810, MixColumnsIns_MixOneColumnInst_2_n58}), .b ({new_AGEMA_signal_7599, MixColumnsIns_MixOneColumnInst_2_n57}), .c ({new_AGEMA_signal_8035, MixColumnsOutput[39]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U91 ( .a ({new_AGEMA_signal_7610, MixColumnsIns_MixOneColumnInst_2_n56}), .b ({new_AGEMA_signal_7476, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .c ({new_AGEMA_signal_7810, MixColumnsIns_MixOneColumnInst_2_n58}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U90 ( .a ({new_AGEMA_signal_7811, MixColumnsIns_MixOneColumnInst_2_n55}), .b ({new_AGEMA_signal_7600, MixColumnsIns_MixOneColumnInst_2_n54}), .c ({new_AGEMA_signal_8036, MixColumnsOutput[38]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U89 ( .a ({new_AGEMA_signal_7612, MixColumnsIns_MixOneColumnInst_2_n53}), .b ({new_AGEMA_signal_7477, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]}), .c ({new_AGEMA_signal_7811, MixColumnsIns_MixOneColumnInst_2_n55}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U88 ( .a ({new_AGEMA_signal_7812, MixColumnsIns_MixOneColumnInst_2_n52}), .b ({new_AGEMA_signal_7601, MixColumnsIns_MixOneColumnInst_2_n51}), .c ({new_AGEMA_signal_8037, MixColumnsOutput[37]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U87 ( .a ({new_AGEMA_signal_7614, MixColumnsIns_MixOneColumnInst_2_n50}), .b ({new_AGEMA_signal_7478, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]}), .c ({new_AGEMA_signal_7812, MixColumnsIns_MixOneColumnInst_2_n52}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U86 ( .a ({new_AGEMA_signal_8038, MixColumnsIns_MixOneColumnInst_2_n49}), .b ({new_AGEMA_signal_7817, MixColumnsIns_MixOneColumnInst_2_n48}), .c ({new_AGEMA_signal_8295, MixColumnsOutput[36]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U85 ( .a ({new_AGEMA_signal_7836, MixColumnsIns_MixOneColumnInst_2_n47}), .b ({new_AGEMA_signal_7479, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]}), .c ({new_AGEMA_signal_8038, MixColumnsIns_MixOneColumnInst_2_n49}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U84 ( .a ({new_AGEMA_signal_8039, MixColumnsIns_MixOneColumnInst_2_n46}), .b ({new_AGEMA_signal_7818, MixColumnsIns_MixOneColumnInst_2_n45}), .c ({new_AGEMA_signal_8296, MixColumnsOutput[35]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U83 ( .a ({new_AGEMA_signal_7838, MixColumnsIns_MixOneColumnInst_2_n44}), .b ({new_AGEMA_signal_7480, MixColumnsInput[43]}), .c ({new_AGEMA_signal_8039, MixColumnsIns_MixOneColumnInst_2_n46}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U82 ( .a ({new_AGEMA_signal_7813, MixColumnsIns_MixOneColumnInst_2_n43}), .b ({new_AGEMA_signal_7599, MixColumnsIns_MixOneColumnInst_2_n57}), .c ({new_AGEMA_signal_8040, MixColumnsOutput[63]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U81 ( .a ({new_AGEMA_signal_7399, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .b ({new_AGEMA_signal_7435, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]}), .c ({new_AGEMA_signal_7599, MixColumnsIns_MixOneColumnInst_2_n57}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U80 ( .a ({new_AGEMA_signal_7441, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_7603, MixColumnsIns_MixOneColumnInst_2_n42}), .c ({new_AGEMA_signal_7813, MixColumnsIns_MixOneColumnInst_2_n43}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U79 ( .a ({new_AGEMA_signal_7814, MixColumnsIns_MixOneColumnInst_2_n41}), .b ({new_AGEMA_signal_7600, MixColumnsIns_MixOneColumnInst_2_n54}), .c ({new_AGEMA_signal_8041, MixColumnsOutput[62]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U78 ( .a ({new_AGEMA_signal_7400, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]}), .b ({new_AGEMA_signal_7436, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]}), .c ({new_AGEMA_signal_7600, MixColumnsIns_MixOneColumnInst_2_n54}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U77 ( .a ({new_AGEMA_signal_7442, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]}), .b ({new_AGEMA_signal_7604, MixColumnsIns_MixOneColumnInst_2_n40}), .c ({new_AGEMA_signal_7814, MixColumnsIns_MixOneColumnInst_2_n41}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U76 ( .a ({new_AGEMA_signal_7815, MixColumnsIns_MixOneColumnInst_2_n39}), .b ({new_AGEMA_signal_7602, MixColumnsIns_MixOneColumnInst_2_n38}), .c ({new_AGEMA_signal_8042, MixColumnsOutput[34]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U75 ( .a ({new_AGEMA_signal_7616, MixColumnsIns_MixOneColumnInst_2_n37}), .b ({new_AGEMA_signal_7481, MixColumnsInput[42]}), .c ({new_AGEMA_signal_7815, MixColumnsIns_MixOneColumnInst_2_n39}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U74 ( .a ({new_AGEMA_signal_7816, MixColumnsIns_MixOneColumnInst_2_n36}), .b ({new_AGEMA_signal_7601, MixColumnsIns_MixOneColumnInst_2_n51}), .c ({new_AGEMA_signal_8043, MixColumnsOutput[61]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U73 ( .a ({new_AGEMA_signal_7401, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]}), .b ({new_AGEMA_signal_7437, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]}), .c ({new_AGEMA_signal_7601, MixColumnsIns_MixOneColumnInst_2_n51}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U72 ( .a ({new_AGEMA_signal_7443, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]}), .b ({new_AGEMA_signal_7605, MixColumnsIns_MixOneColumnInst_2_n35}), .c ({new_AGEMA_signal_7816, MixColumnsIns_MixOneColumnInst_2_n36}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U71 ( .a ({new_AGEMA_signal_8044, MixColumnsIns_MixOneColumnInst_2_n34}), .b ({new_AGEMA_signal_7817, MixColumnsIns_MixOneColumnInst_2_n48}), .c ({new_AGEMA_signal_8297, MixColumnsOutput[60]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U70 ( .a ({new_AGEMA_signal_7402, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]}), .b ({new_AGEMA_signal_7619, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[28]}), .c ({new_AGEMA_signal_7817, MixColumnsIns_MixOneColumnInst_2_n48}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U69 ( .a ({new_AGEMA_signal_7444, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]}), .b ({new_AGEMA_signal_7824, MixColumnsIns_MixOneColumnInst_2_n33}), .c ({new_AGEMA_signal_8044, MixColumnsIns_MixOneColumnInst_2_n34}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U68 ( .a ({new_AGEMA_signal_8045, MixColumnsIns_MixOneColumnInst_2_n32}), .b ({new_AGEMA_signal_7818, MixColumnsIns_MixOneColumnInst_2_n45}), .c ({new_AGEMA_signal_8298, MixColumnsOutput[59]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U67 ( .a ({new_AGEMA_signal_7403, MixColumnsInput[51]}), .b ({new_AGEMA_signal_7620, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[27]}), .c ({new_AGEMA_signal_7818, MixColumnsIns_MixOneColumnInst_2_n45}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U66 ( .a ({new_AGEMA_signal_7445, MixColumnsInput[35]}), .b ({new_AGEMA_signal_7827, MixColumnsIns_MixOneColumnInst_2_n31}), .c ({new_AGEMA_signal_8045, MixColumnsIns_MixOneColumnInst_2_n32}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U65 ( .a ({new_AGEMA_signal_7819, MixColumnsIns_MixOneColumnInst_2_n30}), .b ({new_AGEMA_signal_7602, MixColumnsIns_MixOneColumnInst_2_n38}), .c ({new_AGEMA_signal_8046, MixColumnsOutput[58]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U64 ( .a ({new_AGEMA_signal_7404, MixColumnsInput[50]}), .b ({new_AGEMA_signal_7440, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]}), .c ({new_AGEMA_signal_7602, MixColumnsIns_MixOneColumnInst_2_n38}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U63 ( .a ({new_AGEMA_signal_7446, MixColumnsInput[34]}), .b ({new_AGEMA_signal_7606, MixColumnsIns_MixOneColumnInst_2_n29}), .c ({new_AGEMA_signal_7819, MixColumnsIns_MixOneColumnInst_2_n30}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U62 ( .a ({new_AGEMA_signal_8047, MixColumnsIns_MixOneColumnInst_2_n28}), .b ({new_AGEMA_signal_7825, MixColumnsIns_MixOneColumnInst_2_n27}), .c ({new_AGEMA_signal_8299, MixColumnsOutput[57]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U61 ( .a ({new_AGEMA_signal_7447, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]}), .b ({new_AGEMA_signal_7829, MixColumnsIns_MixOneColumnInst_2_n26}), .c ({new_AGEMA_signal_8047, MixColumnsIns_MixOneColumnInst_2_n28}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U60 ( .a ({new_AGEMA_signal_7820, MixColumnsIns_MixOneColumnInst_2_n25}), .b ({new_AGEMA_signal_7607, MixColumnsIns_MixOneColumnInst_2_n24}), .c ({new_AGEMA_signal_8048, MixColumnsOutput[56]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U59 ( .a ({new_AGEMA_signal_7617, MixColumnsIns_MixOneColumnInst_2_n23}), .b ({new_AGEMA_signal_7275, MixColumnsInput[32]}), .c ({new_AGEMA_signal_7820, MixColumnsIns_MixOneColumnInst_2_n25}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U58 ( .a ({new_AGEMA_signal_7821, MixColumnsIns_MixOneColumnInst_2_n22}), .b ({new_AGEMA_signal_7603, MixColumnsIns_MixOneColumnInst_2_n42}), .c ({new_AGEMA_signal_8049, MixColumnsOutput[55]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U57 ( .a ({new_AGEMA_signal_7476, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .b ({new_AGEMA_signal_7400, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]}), .c ({new_AGEMA_signal_7603, MixColumnsIns_MixOneColumnInst_2_n42}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U56 ( .a ({new_AGEMA_signal_7434, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .b ({new_AGEMA_signal_7609, MixColumnsIns_MixOneColumnInst_2_n21}), .c ({new_AGEMA_signal_7821, MixColumnsIns_MixOneColumnInst_2_n22}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U55 ( .a ({new_AGEMA_signal_7822, MixColumnsIns_MixOneColumnInst_2_n20}), .b ({new_AGEMA_signal_7604, MixColumnsIns_MixOneColumnInst_2_n40}), .c ({new_AGEMA_signal_8050, MixColumnsOutput[54]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U54 ( .a ({new_AGEMA_signal_7477, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]}), .b ({new_AGEMA_signal_7401, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]}), .c ({new_AGEMA_signal_7604, MixColumnsIns_MixOneColumnInst_2_n40}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U53 ( .a ({new_AGEMA_signal_7435, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]}), .b ({new_AGEMA_signal_7611, MixColumnsIns_MixOneColumnInst_2_n19}), .c ({new_AGEMA_signal_7822, MixColumnsIns_MixOneColumnInst_2_n20}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U52 ( .a ({new_AGEMA_signal_7823, MixColumnsIns_MixOneColumnInst_2_n18}), .b ({new_AGEMA_signal_7605, MixColumnsIns_MixOneColumnInst_2_n35}), .c ({new_AGEMA_signal_8051, MixColumnsOutput[53]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U51 ( .a ({new_AGEMA_signal_7478, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]}), .b ({new_AGEMA_signal_7402, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]}), .c ({new_AGEMA_signal_7605, MixColumnsIns_MixOneColumnInst_2_n35}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U50 ( .a ({new_AGEMA_signal_7436, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]}), .b ({new_AGEMA_signal_7613, MixColumnsIns_MixOneColumnInst_2_n17}), .c ({new_AGEMA_signal_7823, MixColumnsIns_MixOneColumnInst_2_n18}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U49 ( .a ({new_AGEMA_signal_8052, MixColumnsIns_MixOneColumnInst_2_n16}), .b ({new_AGEMA_signal_7824, MixColumnsIns_MixOneColumnInst_2_n33}), .c ({new_AGEMA_signal_8300, MixColumnsOutput[52]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U48 ( .a ({new_AGEMA_signal_7479, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]}), .b ({new_AGEMA_signal_7622, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[20]}), .c ({new_AGEMA_signal_7824, MixColumnsIns_MixOneColumnInst_2_n33}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U47 ( .a ({new_AGEMA_signal_7437, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]}), .b ({new_AGEMA_signal_7835, MixColumnsIns_MixOneColumnInst_2_n15}), .c ({new_AGEMA_signal_8052, MixColumnsIns_MixOneColumnInst_2_n16}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U46 ( .a ({new_AGEMA_signal_8053, MixColumnsIns_MixOneColumnInst_2_n14}), .b ({new_AGEMA_signal_7825, MixColumnsIns_MixOneColumnInst_2_n27}), .c ({new_AGEMA_signal_8301, MixColumnsOutput[33]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U45 ( .a ({new_AGEMA_signal_7405, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]}), .b ({new_AGEMA_signal_7621, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[25]}), .c ({new_AGEMA_signal_7825, MixColumnsIns_MixOneColumnInst_2_n27}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U44 ( .a ({new_AGEMA_signal_7482, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]}), .b ({new_AGEMA_signal_7826, MixColumnsIns_MixOneColumnInst_2_n62}), .c ({new_AGEMA_signal_8053, MixColumnsIns_MixOneColumnInst_2_n14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U43 ( .a ({new_AGEMA_signal_7440, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]}), .b ({new_AGEMA_signal_7630, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[1]}), .c ({new_AGEMA_signal_7826, MixColumnsIns_MixOneColumnInst_2_n62}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U42 ( .a ({new_AGEMA_signal_8054, MixColumnsIns_MixOneColumnInst_2_n13}), .b ({new_AGEMA_signal_7827, MixColumnsIns_MixOneColumnInst_2_n31}), .c ({new_AGEMA_signal_8302, MixColumnsOutput[51]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U41 ( .a ({new_AGEMA_signal_7480, MixColumnsInput[43]}), .b ({new_AGEMA_signal_7623, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[19]}), .c ({new_AGEMA_signal_7827, MixColumnsIns_MixOneColumnInst_2_n31}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U40 ( .a ({new_AGEMA_signal_7438, MixColumnsInput[59]}), .b ({new_AGEMA_signal_7837, MixColumnsIns_MixOneColumnInst_2_n12}), .c ({new_AGEMA_signal_8054, MixColumnsIns_MixOneColumnInst_2_n13}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U39 ( .a ({new_AGEMA_signal_7828, MixColumnsIns_MixOneColumnInst_2_n11}), .b ({new_AGEMA_signal_7606, MixColumnsIns_MixOneColumnInst_2_n29}), .c ({new_AGEMA_signal_8055, MixColumnsOutput[50]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U38 ( .a ({new_AGEMA_signal_7481, MixColumnsInput[42]}), .b ({new_AGEMA_signal_7405, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]}), .c ({new_AGEMA_signal_7606, MixColumnsIns_MixOneColumnInst_2_n29}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U37 ( .a ({new_AGEMA_signal_7439, MixColumnsInput[58]}), .b ({new_AGEMA_signal_7615, MixColumnsIns_MixOneColumnInst_2_n10}), .c ({new_AGEMA_signal_7828, MixColumnsIns_MixOneColumnInst_2_n11}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U36 ( .a ({new_AGEMA_signal_8056, MixColumnsIns_MixOneColumnInst_2_n9}), .b ({new_AGEMA_signal_7829, MixColumnsIns_MixOneColumnInst_2_n26}), .c ({new_AGEMA_signal_8303, MixColumnsOutput[49]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U35 ( .a ({new_AGEMA_signal_7624, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[17]}), .b ({new_AGEMA_signal_7482, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]}), .c ({new_AGEMA_signal_7829, MixColumnsIns_MixOneColumnInst_2_n26}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U34 ( .a ({new_AGEMA_signal_7830, MixColumnsIns_MixOneColumnInst_2_n63}), .b ({new_AGEMA_signal_7440, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]}), .c ({new_AGEMA_signal_8056, MixColumnsIns_MixOneColumnInst_2_n9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U33 ( .a ({new_AGEMA_signal_7627, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[9]}), .b ({new_AGEMA_signal_7447, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]}), .c ({new_AGEMA_signal_7830, MixColumnsIns_MixOneColumnInst_2_n63}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U32 ( .a ({new_AGEMA_signal_7831, MixColumnsIns_MixOneColumnInst_2_n8}), .b ({new_AGEMA_signal_7607, MixColumnsIns_MixOneColumnInst_2_n24}), .c ({new_AGEMA_signal_8057, MixColumnsOutput[48]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U31 ( .a ({new_AGEMA_signal_7330, MixColumnsInput[40]}), .b ({new_AGEMA_signal_7399, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .c ({new_AGEMA_signal_7607, MixColumnsIns_MixOneColumnInst_2_n24}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U30 ( .a ({new_AGEMA_signal_7264, MixColumnsInput[56]}), .b ({new_AGEMA_signal_7608, MixColumnsIns_MixOneColumnInst_2_n60}), .c ({new_AGEMA_signal_7831, MixColumnsIns_MixOneColumnInst_2_n8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U29 ( .a ({new_AGEMA_signal_7476, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .b ({new_AGEMA_signal_7275, MixColumnsInput[32]}), .c ({new_AGEMA_signal_7608, MixColumnsIns_MixOneColumnInst_2_n60}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U28 ( .a ({new_AGEMA_signal_7832, MixColumnsIns_MixOneColumnInst_2_n7}), .b ({new_AGEMA_signal_7609, MixColumnsIns_MixOneColumnInst_2_n21}), .c ({new_AGEMA_signal_8058, MixColumnsOutput[47]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U27 ( .a ({new_AGEMA_signal_7441, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_7477, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]}), .c ({new_AGEMA_signal_7609, MixColumnsIns_MixOneColumnInst_2_n21}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U26 ( .a ({new_AGEMA_signal_7610, MixColumnsIns_MixOneColumnInst_2_n56}), .b ({new_AGEMA_signal_7399, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .c ({new_AGEMA_signal_7832, MixColumnsIns_MixOneColumnInst_2_n7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U25 ( .a ({new_AGEMA_signal_7442, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]}), .b ({new_AGEMA_signal_7434, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .c ({new_AGEMA_signal_7610, MixColumnsIns_MixOneColumnInst_2_n56}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U24 ( .a ({new_AGEMA_signal_7833, MixColumnsIns_MixOneColumnInst_2_n6}), .b ({new_AGEMA_signal_7611, MixColumnsIns_MixOneColumnInst_2_n19}), .c ({new_AGEMA_signal_8059, MixColumnsOutput[46]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U23 ( .a ({new_AGEMA_signal_7442, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]}), .b ({new_AGEMA_signal_7478, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]}), .c ({new_AGEMA_signal_7611, MixColumnsIns_MixOneColumnInst_2_n19}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U22 ( .a ({new_AGEMA_signal_7612, MixColumnsIns_MixOneColumnInst_2_n53}), .b ({new_AGEMA_signal_7400, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]}), .c ({new_AGEMA_signal_7833, MixColumnsIns_MixOneColumnInst_2_n6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U21 ( .a ({new_AGEMA_signal_7443, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]}), .b ({new_AGEMA_signal_7435, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]}), .c ({new_AGEMA_signal_7612, MixColumnsIns_MixOneColumnInst_2_n53}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U20 ( .a ({new_AGEMA_signal_7834, MixColumnsIns_MixOneColumnInst_2_n5}), .b ({new_AGEMA_signal_7613, MixColumnsIns_MixOneColumnInst_2_n17}), .c ({new_AGEMA_signal_8060, MixColumnsOutput[45]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U19 ( .a ({new_AGEMA_signal_7443, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]}), .b ({new_AGEMA_signal_7479, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]}), .c ({new_AGEMA_signal_7613, MixColumnsIns_MixOneColumnInst_2_n17}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U18 ( .a ({new_AGEMA_signal_7614, MixColumnsIns_MixOneColumnInst_2_n50}), .b ({new_AGEMA_signal_7401, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]}), .c ({new_AGEMA_signal_7834, MixColumnsIns_MixOneColumnInst_2_n5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U17 ( .a ({new_AGEMA_signal_7444, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]}), .b ({new_AGEMA_signal_7436, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]}), .c ({new_AGEMA_signal_7614, MixColumnsIns_MixOneColumnInst_2_n50}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U16 ( .a ({new_AGEMA_signal_8061, MixColumnsIns_MixOneColumnInst_2_n4}), .b ({new_AGEMA_signal_7835, MixColumnsIns_MixOneColumnInst_2_n15}), .c ({new_AGEMA_signal_8304, MixColumnsOutput[44]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U15 ( .a ({new_AGEMA_signal_7444, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]}), .b ({new_AGEMA_signal_7625, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[12]}), .c ({new_AGEMA_signal_7835, MixColumnsIns_MixOneColumnInst_2_n15}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U14 ( .a ({new_AGEMA_signal_7836, MixColumnsIns_MixOneColumnInst_2_n47}), .b ({new_AGEMA_signal_7402, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]}), .c ({new_AGEMA_signal_8061, MixColumnsIns_MixOneColumnInst_2_n4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U13 ( .a ({new_AGEMA_signal_7628, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[4]}), .b ({new_AGEMA_signal_7437, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]}), .c ({new_AGEMA_signal_7836, MixColumnsIns_MixOneColumnInst_2_n47}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U12 ( .a ({new_AGEMA_signal_8062, MixColumnsIns_MixOneColumnInst_2_n3}), .b ({new_AGEMA_signal_7837, MixColumnsIns_MixOneColumnInst_2_n12}), .c ({new_AGEMA_signal_8305, MixColumnsOutput[43]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U11 ( .a ({new_AGEMA_signal_7445, MixColumnsInput[35]}), .b ({new_AGEMA_signal_7626, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[11]}), .c ({new_AGEMA_signal_7837, MixColumnsIns_MixOneColumnInst_2_n12}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U10 ( .a ({new_AGEMA_signal_7838, MixColumnsIns_MixOneColumnInst_2_n44}), .b ({new_AGEMA_signal_7403, MixColumnsInput[51]}), .c ({new_AGEMA_signal_8062, MixColumnsIns_MixOneColumnInst_2_n3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U9 ( .a ({new_AGEMA_signal_7629, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[3]}), .b ({new_AGEMA_signal_7438, MixColumnsInput[59]}), .c ({new_AGEMA_signal_7838, MixColumnsIns_MixOneColumnInst_2_n44}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U8 ( .a ({new_AGEMA_signal_7839, MixColumnsIns_MixOneColumnInst_2_n2}), .b ({new_AGEMA_signal_7615, MixColumnsIns_MixOneColumnInst_2_n10}), .c ({new_AGEMA_signal_8063, MixColumnsOutput[42]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U7 ( .a ({new_AGEMA_signal_7446, MixColumnsInput[34]}), .b ({new_AGEMA_signal_7482, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]}), .c ({new_AGEMA_signal_7615, MixColumnsIns_MixOneColumnInst_2_n10}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U6 ( .a ({new_AGEMA_signal_7616, MixColumnsIns_MixOneColumnInst_2_n37}), .b ({new_AGEMA_signal_7404, MixColumnsInput[50]}), .c ({new_AGEMA_signal_7839, MixColumnsIns_MixOneColumnInst_2_n2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U5 ( .a ({new_AGEMA_signal_7447, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]}), .b ({new_AGEMA_signal_7439, MixColumnsInput[58]}), .c ({new_AGEMA_signal_7616, MixColumnsIns_MixOneColumnInst_2_n37}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U4 ( .a ({new_AGEMA_signal_7840, MixColumnsIns_MixOneColumnInst_2_n1}), .b ({new_AGEMA_signal_7330, MixColumnsInput[40]}), .c ({new_AGEMA_signal_8064, MixColumnsOutput[32]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U3 ( .a ({new_AGEMA_signal_7618, MixColumnsIns_MixOneColumnInst_2_n59}), .b ({new_AGEMA_signal_7617, MixColumnsIns_MixOneColumnInst_2_n23}), .c ({new_AGEMA_signal_7840, MixColumnsIns_MixOneColumnInst_2_n1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U2 ( .a ({new_AGEMA_signal_7209, MixColumnsInput[48]}), .b ({new_AGEMA_signal_7434, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .c ({new_AGEMA_signal_7617, MixColumnsIns_MixOneColumnInst_2_n23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U1 ( .a ({new_AGEMA_signal_7441, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_7264, MixColumnsInput[56]}), .c ({new_AGEMA_signal_7618, MixColumnsIns_MixOneColumnInst_2_n59}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_0_U3 ( .a ({new_AGEMA_signal_7434, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .b ({new_AGEMA_signal_7438, MixColumnsInput[59]}), .c ({new_AGEMA_signal_7619, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[28]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_0_U2 ( .a ({new_AGEMA_signal_7434, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .b ({new_AGEMA_signal_7439, MixColumnsInput[58]}), .c ({new_AGEMA_signal_7620, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[27]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_0_U1 ( .a ({new_AGEMA_signal_7434, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .b ({new_AGEMA_signal_7264, MixColumnsInput[56]}), .c ({new_AGEMA_signal_7621, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[25]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_1_U3 ( .a ({new_AGEMA_signal_7399, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .b ({new_AGEMA_signal_7403, MixColumnsInput[51]}), .c ({new_AGEMA_signal_7622, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[20]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_1_U2 ( .a ({new_AGEMA_signal_7399, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .b ({new_AGEMA_signal_7404, MixColumnsInput[50]}), .c ({new_AGEMA_signal_7623, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[19]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_1_U1 ( .a ({new_AGEMA_signal_7399, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .b ({new_AGEMA_signal_7209, MixColumnsInput[48]}), .c ({new_AGEMA_signal_7624, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[17]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_2_U3 ( .a ({new_AGEMA_signal_7476, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .b ({new_AGEMA_signal_7480, MixColumnsInput[43]}), .c ({new_AGEMA_signal_7625, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[12]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_2_U2 ( .a ({new_AGEMA_signal_7476, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .b ({new_AGEMA_signal_7481, MixColumnsInput[42]}), .c ({new_AGEMA_signal_7626, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[11]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_2_U1 ( .a ({new_AGEMA_signal_7476, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .b ({new_AGEMA_signal_7330, MixColumnsInput[40]}), .c ({new_AGEMA_signal_7627, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[9]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_3_U3 ( .a ({new_AGEMA_signal_7441, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_7445, MixColumnsInput[35]}), .c ({new_AGEMA_signal_7628, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[4]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_3_U2 ( .a ({new_AGEMA_signal_7441, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_7446, MixColumnsInput[34]}), .c ({new_AGEMA_signal_7629, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[3]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_3_U1 ( .a ({new_AGEMA_signal_7441, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_7275, MixColumnsInput[32]}), .c ({new_AGEMA_signal_7630, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[1]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U96 ( .a ({new_AGEMA_signal_8065, MixColumnsIns_MixOneColumnInst_3_n64}), .b ({new_AGEMA_signal_7489, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]}), .c ({new_AGEMA_signal_8306, MixColumnsOutput[9]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U95 ( .a ({new_AGEMA_signal_7862, MixColumnsIns_MixOneColumnInst_3_n63}), .b ({new_AGEMA_signal_7858, MixColumnsIns_MixOneColumnInst_3_n62}), .c ({new_AGEMA_signal_8065, MixColumnsIns_MixOneColumnInst_3_n64}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U94 ( .a ({new_AGEMA_signal_7841, MixColumnsIns_MixOneColumnInst_3_n61}), .b ({new_AGEMA_signal_7640, MixColumnsIns_MixOneColumnInst_3_n60}), .c ({new_AGEMA_signal_8066, MixColumnsOutput[8]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U93 ( .a ({new_AGEMA_signal_7650, MixColumnsIns_MixOneColumnInst_3_n59}), .b ({new_AGEMA_signal_7341, MixColumnsInput[16]}), .c ({new_AGEMA_signal_7841, MixColumnsIns_MixOneColumnInst_3_n61}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U92 ( .a ({new_AGEMA_signal_7842, MixColumnsIns_MixOneColumnInst_3_n58}), .b ({new_AGEMA_signal_7631, MixColumnsIns_MixOneColumnInst_3_n57}), .c ({new_AGEMA_signal_8067, MixColumnsOutput[7]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U91 ( .a ({new_AGEMA_signal_7642, MixColumnsIns_MixOneColumnInst_3_n56}), .b ({new_AGEMA_signal_7448, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .c ({new_AGEMA_signal_7842, MixColumnsIns_MixOneColumnInst_3_n58}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U90 ( .a ({new_AGEMA_signal_7843, MixColumnsIns_MixOneColumnInst_3_n55}), .b ({new_AGEMA_signal_7632, MixColumnsIns_MixOneColumnInst_3_n54}), .c ({new_AGEMA_signal_8068, MixColumnsOutput[6]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U89 ( .a ({new_AGEMA_signal_7644, MixColumnsIns_MixOneColumnInst_3_n53}), .b ({new_AGEMA_signal_7449, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]}), .c ({new_AGEMA_signal_7843, MixColumnsIns_MixOneColumnInst_3_n55}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U88 ( .a ({new_AGEMA_signal_7844, MixColumnsIns_MixOneColumnInst_3_n52}), .b ({new_AGEMA_signal_7633, MixColumnsIns_MixOneColumnInst_3_n51}), .c ({new_AGEMA_signal_8069, MixColumnsOutput[5]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U87 ( .a ({new_AGEMA_signal_7646, MixColumnsIns_MixOneColumnInst_3_n50}), .b ({new_AGEMA_signal_7450, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]}), .c ({new_AGEMA_signal_7844, MixColumnsIns_MixOneColumnInst_3_n52}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U86 ( .a ({new_AGEMA_signal_8070, MixColumnsIns_MixOneColumnInst_3_n49}), .b ({new_AGEMA_signal_7849, MixColumnsIns_MixOneColumnInst_3_n48}), .c ({new_AGEMA_signal_8307, MixColumnsOutput[4]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U85 ( .a ({new_AGEMA_signal_7868, MixColumnsIns_MixOneColumnInst_3_n47}), .b ({new_AGEMA_signal_7451, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]}), .c ({new_AGEMA_signal_8070, MixColumnsIns_MixOneColumnInst_3_n49}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U84 ( .a ({new_AGEMA_signal_8071, MixColumnsIns_MixOneColumnInst_3_n46}), .b ({new_AGEMA_signal_7850, MixColumnsIns_MixOneColumnInst_3_n45}), .c ({new_AGEMA_signal_8308, MixColumnsOutput[3]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U83 ( .a ({new_AGEMA_signal_7870, MixColumnsIns_MixOneColumnInst_3_n44}), .b ({new_AGEMA_signal_7452, MixColumnsInput[11]}), .c ({new_AGEMA_signal_8071, MixColumnsIns_MixOneColumnInst_3_n46}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U82 ( .a ({new_AGEMA_signal_7845, MixColumnsIns_MixOneColumnInst_3_n43}), .b ({new_AGEMA_signal_7631, MixColumnsIns_MixOneColumnInst_3_n57}), .c ({new_AGEMA_signal_8072, MixColumnsOutput[31]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U81 ( .a ({new_AGEMA_signal_7483, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .b ({new_AGEMA_signal_7407, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]}), .c ({new_AGEMA_signal_7631, MixColumnsIns_MixOneColumnInst_3_n57}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U80 ( .a ({new_AGEMA_signal_7413, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_7635, MixColumnsIns_MixOneColumnInst_3_n42}), .c ({new_AGEMA_signal_7845, MixColumnsIns_MixOneColumnInst_3_n43}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U79 ( .a ({new_AGEMA_signal_7846, MixColumnsIns_MixOneColumnInst_3_n41}), .b ({new_AGEMA_signal_7632, MixColumnsIns_MixOneColumnInst_3_n54}), .c ({new_AGEMA_signal_8073, MixColumnsOutput[30]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U78 ( .a ({new_AGEMA_signal_7484, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]}), .b ({new_AGEMA_signal_7408, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]}), .c ({new_AGEMA_signal_7632, MixColumnsIns_MixOneColumnInst_3_n54}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U77 ( .a ({new_AGEMA_signal_7414, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]}), .b ({new_AGEMA_signal_7636, MixColumnsIns_MixOneColumnInst_3_n40}), .c ({new_AGEMA_signal_7846, MixColumnsIns_MixOneColumnInst_3_n41}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U76 ( .a ({new_AGEMA_signal_7847, MixColumnsIns_MixOneColumnInst_3_n39}), .b ({new_AGEMA_signal_7634, MixColumnsIns_MixOneColumnInst_3_n38}), .c ({new_AGEMA_signal_8074, MixColumnsOutput[2]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U75 ( .a ({new_AGEMA_signal_7648, MixColumnsIns_MixOneColumnInst_3_n37}), .b ({new_AGEMA_signal_7453, MixColumnsInput[10]}), .c ({new_AGEMA_signal_7847, MixColumnsIns_MixOneColumnInst_3_n39}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U74 ( .a ({new_AGEMA_signal_7848, MixColumnsIns_MixOneColumnInst_3_n36}), .b ({new_AGEMA_signal_7633, MixColumnsIns_MixOneColumnInst_3_n51}), .c ({new_AGEMA_signal_8075, MixColumnsOutput[29]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U73 ( .a ({new_AGEMA_signal_7485, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]}), .b ({new_AGEMA_signal_7409, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]}), .c ({new_AGEMA_signal_7633, MixColumnsIns_MixOneColumnInst_3_n51}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U72 ( .a ({new_AGEMA_signal_7415, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]}), .b ({new_AGEMA_signal_7637, MixColumnsIns_MixOneColumnInst_3_n35}), .c ({new_AGEMA_signal_7848, MixColumnsIns_MixOneColumnInst_3_n36}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U71 ( .a ({new_AGEMA_signal_8076, MixColumnsIns_MixOneColumnInst_3_n34}), .b ({new_AGEMA_signal_7849, MixColumnsIns_MixOneColumnInst_3_n48}), .c ({new_AGEMA_signal_8309, MixColumnsOutput[28]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U70 ( .a ({new_AGEMA_signal_7486, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]}), .b ({new_AGEMA_signal_7651, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[28]}), .c ({new_AGEMA_signal_7849, MixColumnsIns_MixOneColumnInst_3_n48}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U69 ( .a ({new_AGEMA_signal_7416, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]}), .b ({new_AGEMA_signal_7856, MixColumnsIns_MixOneColumnInst_3_n33}), .c ({new_AGEMA_signal_8076, MixColumnsIns_MixOneColumnInst_3_n34}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U68 ( .a ({new_AGEMA_signal_8077, MixColumnsIns_MixOneColumnInst_3_n32}), .b ({new_AGEMA_signal_7850, MixColumnsIns_MixOneColumnInst_3_n45}), .c ({new_AGEMA_signal_8310, MixColumnsOutput[27]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U67 ( .a ({new_AGEMA_signal_7487, MixColumnsInput[19]}), .b ({new_AGEMA_signal_7652, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[27]}), .c ({new_AGEMA_signal_7850, MixColumnsIns_MixOneColumnInst_3_n45}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U66 ( .a ({new_AGEMA_signal_7417, MixColumnsInput[3]}), .b ({new_AGEMA_signal_7859, MixColumnsIns_MixOneColumnInst_3_n31}), .c ({new_AGEMA_signal_8077, MixColumnsIns_MixOneColumnInst_3_n32}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U65 ( .a ({new_AGEMA_signal_7851, MixColumnsIns_MixOneColumnInst_3_n30}), .b ({new_AGEMA_signal_7634, MixColumnsIns_MixOneColumnInst_3_n38}), .c ({new_AGEMA_signal_8078, MixColumnsOutput[26]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U64 ( .a ({new_AGEMA_signal_7488, MixColumnsInput[18]}), .b ({new_AGEMA_signal_7412, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]}), .c ({new_AGEMA_signal_7634, MixColumnsIns_MixOneColumnInst_3_n38}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U63 ( .a ({new_AGEMA_signal_7418, MixColumnsInput[2]}), .b ({new_AGEMA_signal_7638, MixColumnsIns_MixOneColumnInst_3_n29}), .c ({new_AGEMA_signal_7851, MixColumnsIns_MixOneColumnInst_3_n30}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U62 ( .a ({new_AGEMA_signal_8079, MixColumnsIns_MixOneColumnInst_3_n28}), .b ({new_AGEMA_signal_7857, MixColumnsIns_MixOneColumnInst_3_n27}), .c ({new_AGEMA_signal_8311, MixColumnsOutput[25]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U61 ( .a ({new_AGEMA_signal_7419, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]}), .b ({new_AGEMA_signal_7861, MixColumnsIns_MixOneColumnInst_3_n26}), .c ({new_AGEMA_signal_8079, MixColumnsIns_MixOneColumnInst_3_n28}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U60 ( .a ({new_AGEMA_signal_7852, MixColumnsIns_MixOneColumnInst_3_n25}), .b ({new_AGEMA_signal_7639, MixColumnsIns_MixOneColumnInst_3_n24}), .c ({new_AGEMA_signal_8080, MixColumnsOutput[24]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U59 ( .a ({new_AGEMA_signal_7649, MixColumnsIns_MixOneColumnInst_3_n23}), .b ({new_AGEMA_signal_7231, MixColumnsInput[0]}), .c ({new_AGEMA_signal_7852, MixColumnsIns_MixOneColumnInst_3_n25}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U58 ( .a ({new_AGEMA_signal_7853, MixColumnsIns_MixOneColumnInst_3_n22}), .b ({new_AGEMA_signal_7635, MixColumnsIns_MixOneColumnInst_3_n42}), .c ({new_AGEMA_signal_8081, MixColumnsOutput[23]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U57 ( .a ({new_AGEMA_signal_7448, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .b ({new_AGEMA_signal_7484, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]}), .c ({new_AGEMA_signal_7635, MixColumnsIns_MixOneColumnInst_3_n42}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U56 ( .a ({new_AGEMA_signal_7406, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .b ({new_AGEMA_signal_7641, MixColumnsIns_MixOneColumnInst_3_n21}), .c ({new_AGEMA_signal_7853, MixColumnsIns_MixOneColumnInst_3_n22}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U55 ( .a ({new_AGEMA_signal_7854, MixColumnsIns_MixOneColumnInst_3_n20}), .b ({new_AGEMA_signal_7636, MixColumnsIns_MixOneColumnInst_3_n40}), .c ({new_AGEMA_signal_8082, MixColumnsOutput[22]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U54 ( .a ({new_AGEMA_signal_7449, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]}), .b ({new_AGEMA_signal_7485, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]}), .c ({new_AGEMA_signal_7636, MixColumnsIns_MixOneColumnInst_3_n40}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U53 ( .a ({new_AGEMA_signal_7407, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]}), .b ({new_AGEMA_signal_7643, MixColumnsIns_MixOneColumnInst_3_n19}), .c ({new_AGEMA_signal_7854, MixColumnsIns_MixOneColumnInst_3_n20}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U52 ( .a ({new_AGEMA_signal_7855, MixColumnsIns_MixOneColumnInst_3_n18}), .b ({new_AGEMA_signal_7637, MixColumnsIns_MixOneColumnInst_3_n35}), .c ({new_AGEMA_signal_8083, MixColumnsOutput[21]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U51 ( .a ({new_AGEMA_signal_7450, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]}), .b ({new_AGEMA_signal_7486, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]}), .c ({new_AGEMA_signal_7637, MixColumnsIns_MixOneColumnInst_3_n35}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U50 ( .a ({new_AGEMA_signal_7408, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]}), .b ({new_AGEMA_signal_7645, MixColumnsIns_MixOneColumnInst_3_n17}), .c ({new_AGEMA_signal_7855, MixColumnsIns_MixOneColumnInst_3_n18}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U49 ( .a ({new_AGEMA_signal_8084, MixColumnsIns_MixOneColumnInst_3_n16}), .b ({new_AGEMA_signal_7856, MixColumnsIns_MixOneColumnInst_3_n33}), .c ({new_AGEMA_signal_8312, MixColumnsOutput[20]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U48 ( .a ({new_AGEMA_signal_7451, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]}), .b ({new_AGEMA_signal_7654, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[20]}), .c ({new_AGEMA_signal_7856, MixColumnsIns_MixOneColumnInst_3_n33}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U47 ( .a ({new_AGEMA_signal_7409, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]}), .b ({new_AGEMA_signal_7867, MixColumnsIns_MixOneColumnInst_3_n15}), .c ({new_AGEMA_signal_8084, MixColumnsIns_MixOneColumnInst_3_n16}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U46 ( .a ({new_AGEMA_signal_8085, MixColumnsIns_MixOneColumnInst_3_n14}), .b ({new_AGEMA_signal_7857, MixColumnsIns_MixOneColumnInst_3_n27}), .c ({new_AGEMA_signal_8313, MixColumnsOutput[1]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U45 ( .a ({new_AGEMA_signal_7489, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]}), .b ({new_AGEMA_signal_7653, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[25]}), .c ({new_AGEMA_signal_7857, MixColumnsIns_MixOneColumnInst_3_n27}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U44 ( .a ({new_AGEMA_signal_7454, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]}), .b ({new_AGEMA_signal_7858, MixColumnsIns_MixOneColumnInst_3_n62}), .c ({new_AGEMA_signal_8085, MixColumnsIns_MixOneColumnInst_3_n14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U43 ( .a ({new_AGEMA_signal_7412, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]}), .b ({new_AGEMA_signal_7662, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[1]}), .c ({new_AGEMA_signal_7858, MixColumnsIns_MixOneColumnInst_3_n62}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U42 ( .a ({new_AGEMA_signal_8086, MixColumnsIns_MixOneColumnInst_3_n13}), .b ({new_AGEMA_signal_7859, MixColumnsIns_MixOneColumnInst_3_n31}), .c ({new_AGEMA_signal_8314, MixColumnsOutput[19]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U41 ( .a ({new_AGEMA_signal_7452, MixColumnsInput[11]}), .b ({new_AGEMA_signal_7655, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[19]}), .c ({new_AGEMA_signal_7859, MixColumnsIns_MixOneColumnInst_3_n31}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U40 ( .a ({new_AGEMA_signal_7410, MixColumnsInput[27]}), .b ({new_AGEMA_signal_7869, MixColumnsIns_MixOneColumnInst_3_n12}), .c ({new_AGEMA_signal_8086, MixColumnsIns_MixOneColumnInst_3_n13}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U39 ( .a ({new_AGEMA_signal_7860, MixColumnsIns_MixOneColumnInst_3_n11}), .b ({new_AGEMA_signal_7638, MixColumnsIns_MixOneColumnInst_3_n29}), .c ({new_AGEMA_signal_8087, MixColumnsOutput[18]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U38 ( .a ({new_AGEMA_signal_7453, MixColumnsInput[10]}), .b ({new_AGEMA_signal_7489, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]}), .c ({new_AGEMA_signal_7638, MixColumnsIns_MixOneColumnInst_3_n29}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U37 ( .a ({new_AGEMA_signal_7411, MixColumnsInput[26]}), .b ({new_AGEMA_signal_7647, MixColumnsIns_MixOneColumnInst_3_n10}), .c ({new_AGEMA_signal_7860, MixColumnsIns_MixOneColumnInst_3_n11}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U36 ( .a ({new_AGEMA_signal_8088, MixColumnsIns_MixOneColumnInst_3_n9}), .b ({new_AGEMA_signal_7861, MixColumnsIns_MixOneColumnInst_3_n26}), .c ({new_AGEMA_signal_8315, MixColumnsOutput[17]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U35 ( .a ({new_AGEMA_signal_7656, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[17]}), .b ({new_AGEMA_signal_7454, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]}), .c ({new_AGEMA_signal_7861, MixColumnsIns_MixOneColumnInst_3_n26}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U34 ( .a ({new_AGEMA_signal_7862, MixColumnsIns_MixOneColumnInst_3_n63}), .b ({new_AGEMA_signal_7412, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]}), .c ({new_AGEMA_signal_8088, MixColumnsIns_MixOneColumnInst_3_n9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U33 ( .a ({new_AGEMA_signal_7659, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[9]}), .b ({new_AGEMA_signal_7419, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]}), .c ({new_AGEMA_signal_7862, MixColumnsIns_MixOneColumnInst_3_n63}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U32 ( .a ({new_AGEMA_signal_7863, MixColumnsIns_MixOneColumnInst_3_n8}), .b ({new_AGEMA_signal_7639, MixColumnsIns_MixOneColumnInst_3_n24}), .c ({new_AGEMA_signal_8089, MixColumnsOutput[16]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U31 ( .a ({new_AGEMA_signal_7286, MixColumnsInput[8]}), .b ({new_AGEMA_signal_7483, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .c ({new_AGEMA_signal_7639, MixColumnsIns_MixOneColumnInst_3_n24}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U30 ( .a ({new_AGEMA_signal_7220, MixColumnsInput[24]}), .b ({new_AGEMA_signal_7640, MixColumnsIns_MixOneColumnInst_3_n60}), .c ({new_AGEMA_signal_7863, MixColumnsIns_MixOneColumnInst_3_n8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U29 ( .a ({new_AGEMA_signal_7448, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .b ({new_AGEMA_signal_7231, MixColumnsInput[0]}), .c ({new_AGEMA_signal_7640, MixColumnsIns_MixOneColumnInst_3_n60}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U28 ( .a ({new_AGEMA_signal_7864, MixColumnsIns_MixOneColumnInst_3_n7}), .b ({new_AGEMA_signal_7641, MixColumnsIns_MixOneColumnInst_3_n21}), .c ({new_AGEMA_signal_8090, MixColumnsOutput[15]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U27 ( .a ({new_AGEMA_signal_7413, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_7449, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]}), .c ({new_AGEMA_signal_7641, MixColumnsIns_MixOneColumnInst_3_n21}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U26 ( .a ({new_AGEMA_signal_7642, MixColumnsIns_MixOneColumnInst_3_n56}), .b ({new_AGEMA_signal_7483, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .c ({new_AGEMA_signal_7864, MixColumnsIns_MixOneColumnInst_3_n7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U25 ( .a ({new_AGEMA_signal_7414, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]}), .b ({new_AGEMA_signal_7406, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .c ({new_AGEMA_signal_7642, MixColumnsIns_MixOneColumnInst_3_n56}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U24 ( .a ({new_AGEMA_signal_7865, MixColumnsIns_MixOneColumnInst_3_n6}), .b ({new_AGEMA_signal_7643, MixColumnsIns_MixOneColumnInst_3_n19}), .c ({new_AGEMA_signal_8091, MixColumnsOutput[14]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U23 ( .a ({new_AGEMA_signal_7414, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]}), .b ({new_AGEMA_signal_7450, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]}), .c ({new_AGEMA_signal_7643, MixColumnsIns_MixOneColumnInst_3_n19}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U22 ( .a ({new_AGEMA_signal_7644, MixColumnsIns_MixOneColumnInst_3_n53}), .b ({new_AGEMA_signal_7484, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]}), .c ({new_AGEMA_signal_7865, MixColumnsIns_MixOneColumnInst_3_n6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U21 ( .a ({new_AGEMA_signal_7415, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]}), .b ({new_AGEMA_signal_7407, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]}), .c ({new_AGEMA_signal_7644, MixColumnsIns_MixOneColumnInst_3_n53}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U20 ( .a ({new_AGEMA_signal_7866, MixColumnsIns_MixOneColumnInst_3_n5}), .b ({new_AGEMA_signal_7645, MixColumnsIns_MixOneColumnInst_3_n17}), .c ({new_AGEMA_signal_8092, MixColumnsOutput[13]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U19 ( .a ({new_AGEMA_signal_7415, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]}), .b ({new_AGEMA_signal_7451, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]}), .c ({new_AGEMA_signal_7645, MixColumnsIns_MixOneColumnInst_3_n17}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U18 ( .a ({new_AGEMA_signal_7646, MixColumnsIns_MixOneColumnInst_3_n50}), .b ({new_AGEMA_signal_7485, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]}), .c ({new_AGEMA_signal_7866, MixColumnsIns_MixOneColumnInst_3_n5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U17 ( .a ({new_AGEMA_signal_7416, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]}), .b ({new_AGEMA_signal_7408, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]}), .c ({new_AGEMA_signal_7646, MixColumnsIns_MixOneColumnInst_3_n50}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U16 ( .a ({new_AGEMA_signal_8093, MixColumnsIns_MixOneColumnInst_3_n4}), .b ({new_AGEMA_signal_7867, MixColumnsIns_MixOneColumnInst_3_n15}), .c ({new_AGEMA_signal_8316, MixColumnsOutput[12]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U15 ( .a ({new_AGEMA_signal_7416, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]}), .b ({new_AGEMA_signal_7657, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[12]}), .c ({new_AGEMA_signal_7867, MixColumnsIns_MixOneColumnInst_3_n15}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U14 ( .a ({new_AGEMA_signal_7868, MixColumnsIns_MixOneColumnInst_3_n47}), .b ({new_AGEMA_signal_7486, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]}), .c ({new_AGEMA_signal_8093, MixColumnsIns_MixOneColumnInst_3_n4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U13 ( .a ({new_AGEMA_signal_7660, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[4]}), .b ({new_AGEMA_signal_7409, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]}), .c ({new_AGEMA_signal_7868, MixColumnsIns_MixOneColumnInst_3_n47}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U12 ( .a ({new_AGEMA_signal_8094, MixColumnsIns_MixOneColumnInst_3_n3}), .b ({new_AGEMA_signal_7869, MixColumnsIns_MixOneColumnInst_3_n12}), .c ({new_AGEMA_signal_8317, MixColumnsOutput[11]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U11 ( .a ({new_AGEMA_signal_7417, MixColumnsInput[3]}), .b ({new_AGEMA_signal_7658, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[11]}), .c ({new_AGEMA_signal_7869, MixColumnsIns_MixOneColumnInst_3_n12}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U10 ( .a ({new_AGEMA_signal_7870, MixColumnsIns_MixOneColumnInst_3_n44}), .b ({new_AGEMA_signal_7487, MixColumnsInput[19]}), .c ({new_AGEMA_signal_8094, MixColumnsIns_MixOneColumnInst_3_n3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U9 ( .a ({new_AGEMA_signal_7661, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[3]}), .b ({new_AGEMA_signal_7410, MixColumnsInput[27]}), .c ({new_AGEMA_signal_7870, MixColumnsIns_MixOneColumnInst_3_n44}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U8 ( .a ({new_AGEMA_signal_7871, MixColumnsIns_MixOneColumnInst_3_n2}), .b ({new_AGEMA_signal_7647, MixColumnsIns_MixOneColumnInst_3_n10}), .c ({new_AGEMA_signal_8095, MixColumnsOutput[10]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U7 ( .a ({new_AGEMA_signal_7418, MixColumnsInput[2]}), .b ({new_AGEMA_signal_7454, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]}), .c ({new_AGEMA_signal_7647, MixColumnsIns_MixOneColumnInst_3_n10}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U6 ( .a ({new_AGEMA_signal_7648, MixColumnsIns_MixOneColumnInst_3_n37}), .b ({new_AGEMA_signal_7488, MixColumnsInput[18]}), .c ({new_AGEMA_signal_7871, MixColumnsIns_MixOneColumnInst_3_n2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U5 ( .a ({new_AGEMA_signal_7419, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]}), .b ({new_AGEMA_signal_7411, MixColumnsInput[26]}), .c ({new_AGEMA_signal_7648, MixColumnsIns_MixOneColumnInst_3_n37}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U4 ( .a ({new_AGEMA_signal_7872, MixColumnsIns_MixOneColumnInst_3_n1}), .b ({new_AGEMA_signal_7286, MixColumnsInput[8]}), .c ({new_AGEMA_signal_8096, MixColumnsOutput[0]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U3 ( .a ({new_AGEMA_signal_7650, MixColumnsIns_MixOneColumnInst_3_n59}), .b ({new_AGEMA_signal_7649, MixColumnsIns_MixOneColumnInst_3_n23}), .c ({new_AGEMA_signal_7872, MixColumnsIns_MixOneColumnInst_3_n1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U2 ( .a ({new_AGEMA_signal_7341, MixColumnsInput[16]}), .b ({new_AGEMA_signal_7406, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .c ({new_AGEMA_signal_7649, MixColumnsIns_MixOneColumnInst_3_n23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U1 ( .a ({new_AGEMA_signal_7413, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_7220, MixColumnsInput[24]}), .c ({new_AGEMA_signal_7650, MixColumnsIns_MixOneColumnInst_3_n59}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_0_U3 ( .a ({new_AGEMA_signal_7406, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .b ({new_AGEMA_signal_7410, MixColumnsInput[27]}), .c ({new_AGEMA_signal_7651, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[28]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_0_U2 ( .a ({new_AGEMA_signal_7406, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .b ({new_AGEMA_signal_7411, MixColumnsInput[26]}), .c ({new_AGEMA_signal_7652, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[27]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_0_U1 ( .a ({new_AGEMA_signal_7406, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .b ({new_AGEMA_signal_7220, MixColumnsInput[24]}), .c ({new_AGEMA_signal_7653, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[25]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_1_U3 ( .a ({new_AGEMA_signal_7483, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .b ({new_AGEMA_signal_7487, MixColumnsInput[19]}), .c ({new_AGEMA_signal_7654, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[20]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_1_U2 ( .a ({new_AGEMA_signal_7483, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .b ({new_AGEMA_signal_7488, MixColumnsInput[18]}), .c ({new_AGEMA_signal_7655, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[19]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_1_U1 ( .a ({new_AGEMA_signal_7483, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .b ({new_AGEMA_signal_7341, MixColumnsInput[16]}), .c ({new_AGEMA_signal_7656, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[17]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_2_U3 ( .a ({new_AGEMA_signal_7448, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .b ({new_AGEMA_signal_7452, MixColumnsInput[11]}), .c ({new_AGEMA_signal_7657, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[12]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_2_U2 ( .a ({new_AGEMA_signal_7448, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .b ({new_AGEMA_signal_7453, MixColumnsInput[10]}), .c ({new_AGEMA_signal_7658, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[11]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_2_U1 ( .a ({new_AGEMA_signal_7448, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .b ({new_AGEMA_signal_7286, MixColumnsInput[8]}), .c ({new_AGEMA_signal_7659, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[9]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_3_U3 ( .a ({new_AGEMA_signal_7413, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_7417, MixColumnsInput[3]}), .c ({new_AGEMA_signal_7660, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[4]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_3_U2 ( .a ({new_AGEMA_signal_7413, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_7418, MixColumnsInput[2]}), .c ({new_AGEMA_signal_7661, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[3]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_3_U1 ( .a ({new_AGEMA_signal_7413, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_7231, MixColumnsInput[0]}), .c ({new_AGEMA_signal_7662, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_0_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7968, KeyExpansionOutput[0]}), .a ({new_AGEMA_signal_13332, new_AGEMA_signal_13328}), .c ({new_AGEMA_signal_8098, KeyReg_Inst_ff_SDE_0_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_1_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8180, KeyExpansionOutput[1]}), .a ({new_AGEMA_signal_13340, new_AGEMA_signal_13336}), .c ({new_AGEMA_signal_8319, KeyReg_Inst_ff_SDE_1_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_2_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8169, KeyExpansionOutput[2]}), .a ({new_AGEMA_signal_13348, new_AGEMA_signal_13344}), .c ({new_AGEMA_signal_8321, KeyReg_Inst_ff_SDE_2_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_3_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8166, KeyExpansionOutput[3]}), .a ({new_AGEMA_signal_13356, new_AGEMA_signal_13352}), .c ({new_AGEMA_signal_8323, KeyReg_Inst_ff_SDE_3_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_4_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8165, KeyExpansionOutput[4]}), .a ({new_AGEMA_signal_13364, new_AGEMA_signal_13360}), .c ({new_AGEMA_signal_8325, KeyReg_Inst_ff_SDE_4_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_5_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8164, KeyExpansionOutput[5]}), .a ({new_AGEMA_signal_13372, new_AGEMA_signal_13368}), .c ({new_AGEMA_signal_8327, KeyReg_Inst_ff_SDE_5_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_6_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8163, KeyExpansionOutput[6]}), .a ({new_AGEMA_signal_13380, new_AGEMA_signal_13376}), .c ({new_AGEMA_signal_8329, KeyReg_Inst_ff_SDE_6_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_7_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8162, KeyExpansionOutput[7]}), .a ({new_AGEMA_signal_13388, new_AGEMA_signal_13384}), .c ({new_AGEMA_signal_8331, KeyReg_Inst_ff_SDE_7_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_8_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7937, KeyExpansionOutput[8]}), .a ({new_AGEMA_signal_13396, new_AGEMA_signal_13392}), .c ({new_AGEMA_signal_8100, KeyReg_Inst_ff_SDE_8_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_9_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8161, KeyExpansionOutput[9]}), .a ({new_AGEMA_signal_13404, new_AGEMA_signal_13400}), .c ({new_AGEMA_signal_8333, KeyReg_Inst_ff_SDE_9_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_10_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8189, KeyExpansionOutput[10]}), .a ({new_AGEMA_signal_13412, new_AGEMA_signal_13408}), .c ({new_AGEMA_signal_8335, KeyReg_Inst_ff_SDE_10_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_11_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8188, KeyExpansionOutput[11]}), .a ({new_AGEMA_signal_13420, new_AGEMA_signal_13416}), .c ({new_AGEMA_signal_8337, KeyReg_Inst_ff_SDE_11_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_12_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8187, KeyExpansionOutput[12]}), .a ({new_AGEMA_signal_13428, new_AGEMA_signal_13424}), .c ({new_AGEMA_signal_8339, KeyReg_Inst_ff_SDE_12_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_13_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8186, KeyExpansionOutput[13]}), .a ({new_AGEMA_signal_13436, new_AGEMA_signal_13432}), .c ({new_AGEMA_signal_8341, KeyReg_Inst_ff_SDE_13_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_14_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8185, KeyExpansionOutput[14]}), .a ({new_AGEMA_signal_13444, new_AGEMA_signal_13440}), .c ({new_AGEMA_signal_8343, KeyReg_Inst_ff_SDE_14_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_15_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8184, KeyExpansionOutput[15]}), .a ({new_AGEMA_signal_13452, new_AGEMA_signal_13448}), .c ({new_AGEMA_signal_8345, KeyReg_Inst_ff_SDE_15_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_16_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7961, KeyExpansionOutput[16]}), .a ({new_AGEMA_signal_13460, new_AGEMA_signal_13456}), .c ({new_AGEMA_signal_8102, KeyReg_Inst_ff_SDE_16_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_17_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8183, KeyExpansionOutput[17]}), .a ({new_AGEMA_signal_13468, new_AGEMA_signal_13464}), .c ({new_AGEMA_signal_8347, KeyReg_Inst_ff_SDE_17_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_18_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8182, KeyExpansionOutput[18]}), .a ({new_AGEMA_signal_13476, new_AGEMA_signal_13472}), .c ({new_AGEMA_signal_8349, KeyReg_Inst_ff_SDE_18_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_19_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8181, KeyExpansionOutput[19]}), .a ({new_AGEMA_signal_13484, new_AGEMA_signal_13480}), .c ({new_AGEMA_signal_8351, KeyReg_Inst_ff_SDE_19_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_20_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8179, KeyExpansionOutput[20]}), .a ({new_AGEMA_signal_13492, new_AGEMA_signal_13488}), .c ({new_AGEMA_signal_8353, KeyReg_Inst_ff_SDE_20_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_21_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8178, KeyExpansionOutput[21]}), .a ({new_AGEMA_signal_13500, new_AGEMA_signal_13496}), .c ({new_AGEMA_signal_8355, KeyReg_Inst_ff_SDE_21_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_22_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8177, KeyExpansionOutput[22]}), .a ({new_AGEMA_signal_13508, new_AGEMA_signal_13504}), .c ({new_AGEMA_signal_8357, KeyReg_Inst_ff_SDE_22_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_23_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8176, KeyExpansionOutput[23]}), .a ({new_AGEMA_signal_13516, new_AGEMA_signal_13512}), .c ({new_AGEMA_signal_8359, KeyReg_Inst_ff_SDE_23_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_24_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8175, KeyExpansionOutput[24]}), .a ({new_AGEMA_signal_13524, new_AGEMA_signal_13520}), .c ({new_AGEMA_signal_8361, KeyReg_Inst_ff_SDE_24_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_25_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8382, KeyExpansionOutput[25]}), .a ({new_AGEMA_signal_13532, new_AGEMA_signal_13528}), .c ({new_AGEMA_signal_8592, KeyReg_Inst_ff_SDE_25_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_26_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8381, KeyExpansionOutput[26]}), .a ({new_AGEMA_signal_13540, new_AGEMA_signal_13536}), .c ({new_AGEMA_signal_8594, KeyReg_Inst_ff_SDE_26_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_27_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8380, KeyExpansionOutput[27]}), .a ({new_AGEMA_signal_13548, new_AGEMA_signal_13544}), .c ({new_AGEMA_signal_8596, KeyReg_Inst_ff_SDE_27_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_28_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8379, KeyExpansionOutput[28]}), .a ({new_AGEMA_signal_13556, new_AGEMA_signal_13552}), .c ({new_AGEMA_signal_8598, KeyReg_Inst_ff_SDE_28_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_29_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8378, KeyExpansionOutput[29]}), .a ({new_AGEMA_signal_13564, new_AGEMA_signal_13560}), .c ({new_AGEMA_signal_8600, KeyReg_Inst_ff_SDE_29_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_30_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8377, KeyExpansionOutput[30]}), .a ({new_AGEMA_signal_13572, new_AGEMA_signal_13568}), .c ({new_AGEMA_signal_8602, KeyReg_Inst_ff_SDE_30_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_31_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8376, KeyExpansionOutput[31]}), .a ({new_AGEMA_signal_13580, new_AGEMA_signal_13576}), .c ({new_AGEMA_signal_8604, KeyReg_Inst_ff_SDE_31_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_32_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7744, KeyExpansionOutput[32]}), .a ({new_AGEMA_signal_13588, new_AGEMA_signal_13584}), .c ({new_AGEMA_signal_7874, KeyReg_Inst_ff_SDE_32_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_33_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7957, KeyExpansionOutput[33]}), .a ({new_AGEMA_signal_13596, new_AGEMA_signal_13592}), .c ({new_AGEMA_signal_8104, KeyReg_Inst_ff_SDE_33_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_34_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7946, KeyExpansionOutput[34]}), .a ({new_AGEMA_signal_13604, new_AGEMA_signal_13600}), .c ({new_AGEMA_signal_8106, KeyReg_Inst_ff_SDE_34_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_35_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7943, KeyExpansionOutput[35]}), .a ({new_AGEMA_signal_13612, new_AGEMA_signal_13608}), .c ({new_AGEMA_signal_8108, KeyReg_Inst_ff_SDE_35_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_36_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7942, KeyExpansionOutput[36]}), .a ({new_AGEMA_signal_13620, new_AGEMA_signal_13616}), .c ({new_AGEMA_signal_8110, KeyReg_Inst_ff_SDE_36_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_37_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7941, KeyExpansionOutput[37]}), .a ({new_AGEMA_signal_13628, new_AGEMA_signal_13624}), .c ({new_AGEMA_signal_8112, KeyReg_Inst_ff_SDE_37_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_38_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7940, KeyExpansionOutput[38]}), .a ({new_AGEMA_signal_13636, new_AGEMA_signal_13632}), .c ({new_AGEMA_signal_8114, KeyReg_Inst_ff_SDE_38_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_39_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7939, KeyExpansionOutput[39]}), .a ({new_AGEMA_signal_13644, new_AGEMA_signal_13640}), .c ({new_AGEMA_signal_8116, KeyReg_Inst_ff_SDE_39_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_40_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7714, KeyExpansionOutput[40]}), .a ({new_AGEMA_signal_13652, new_AGEMA_signal_13648}), .c ({new_AGEMA_signal_7876, KeyReg_Inst_ff_SDE_40_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_41_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7938, KeyExpansionOutput[41]}), .a ({new_AGEMA_signal_13660, new_AGEMA_signal_13656}), .c ({new_AGEMA_signal_8118, KeyReg_Inst_ff_SDE_41_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_42_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7967, KeyExpansionOutput[42]}), .a ({new_AGEMA_signal_13668, new_AGEMA_signal_13664}), .c ({new_AGEMA_signal_8120, KeyReg_Inst_ff_SDE_42_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_43_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7966, KeyExpansionOutput[43]}), .a ({new_AGEMA_signal_13676, new_AGEMA_signal_13672}), .c ({new_AGEMA_signal_8122, KeyReg_Inst_ff_SDE_43_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_44_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7965, KeyExpansionOutput[44]}), .a ({new_AGEMA_signal_13684, new_AGEMA_signal_13680}), .c ({new_AGEMA_signal_8124, KeyReg_Inst_ff_SDE_44_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_45_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7964, KeyExpansionOutput[45]}), .a ({new_AGEMA_signal_13692, new_AGEMA_signal_13688}), .c ({new_AGEMA_signal_8126, KeyReg_Inst_ff_SDE_45_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_46_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7963, KeyExpansionOutput[46]}), .a ({new_AGEMA_signal_13700, new_AGEMA_signal_13696}), .c ({new_AGEMA_signal_8128, KeyReg_Inst_ff_SDE_46_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_47_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7962, KeyExpansionOutput[47]}), .a ({new_AGEMA_signal_13708, new_AGEMA_signal_13704}), .c ({new_AGEMA_signal_8130, KeyReg_Inst_ff_SDE_47_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_48_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7730, KeyExpansionOutput[48]}), .a ({new_AGEMA_signal_13716, new_AGEMA_signal_13712}), .c ({new_AGEMA_signal_7878, KeyReg_Inst_ff_SDE_48_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_49_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7960, KeyExpansionOutput[49]}), .a ({new_AGEMA_signal_13724, new_AGEMA_signal_13720}), .c ({new_AGEMA_signal_8132, KeyReg_Inst_ff_SDE_49_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_50_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7959, KeyExpansionOutput[50]}), .a ({new_AGEMA_signal_13732, new_AGEMA_signal_13728}), .c ({new_AGEMA_signal_8134, KeyReg_Inst_ff_SDE_50_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_51_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7958, KeyExpansionOutput[51]}), .a ({new_AGEMA_signal_13740, new_AGEMA_signal_13736}), .c ({new_AGEMA_signal_8136, KeyReg_Inst_ff_SDE_51_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_52_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7956, KeyExpansionOutput[52]}), .a ({new_AGEMA_signal_13748, new_AGEMA_signal_13744}), .c ({new_AGEMA_signal_8138, KeyReg_Inst_ff_SDE_52_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_53_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7955, KeyExpansionOutput[53]}), .a ({new_AGEMA_signal_13756, new_AGEMA_signal_13752}), .c ({new_AGEMA_signal_8140, KeyReg_Inst_ff_SDE_53_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_54_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7954, KeyExpansionOutput[54]}), .a ({new_AGEMA_signal_13764, new_AGEMA_signal_13760}), .c ({new_AGEMA_signal_8142, KeyReg_Inst_ff_SDE_54_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_55_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7953, KeyExpansionOutput[55]}), .a ({new_AGEMA_signal_13772, new_AGEMA_signal_13768}), .c ({new_AGEMA_signal_8144, KeyReg_Inst_ff_SDE_55_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_56_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7952, KeyExpansionOutput[56]}), .a ({new_AGEMA_signal_13780, new_AGEMA_signal_13776}), .c ({new_AGEMA_signal_8146, KeyReg_Inst_ff_SDE_56_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_57_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8174, KeyExpansionOutput[57]}), .a ({new_AGEMA_signal_13788, new_AGEMA_signal_13784}), .c ({new_AGEMA_signal_8363, KeyReg_Inst_ff_SDE_57_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_58_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8173, KeyExpansionOutput[58]}), .a ({new_AGEMA_signal_13796, new_AGEMA_signal_13792}), .c ({new_AGEMA_signal_8365, KeyReg_Inst_ff_SDE_58_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_59_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8172, KeyExpansionOutput[59]}), .a ({new_AGEMA_signal_13804, new_AGEMA_signal_13800}), .c ({new_AGEMA_signal_8367, KeyReg_Inst_ff_SDE_59_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_60_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8171, KeyExpansionOutput[60]}), .a ({new_AGEMA_signal_13812, new_AGEMA_signal_13808}), .c ({new_AGEMA_signal_8369, KeyReg_Inst_ff_SDE_60_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_61_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8170, KeyExpansionOutput[61]}), .a ({new_AGEMA_signal_13820, new_AGEMA_signal_13816}), .c ({new_AGEMA_signal_8371, KeyReg_Inst_ff_SDE_61_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_62_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8168, KeyExpansionOutput[62]}), .a ({new_AGEMA_signal_13828, new_AGEMA_signal_13824}), .c ({new_AGEMA_signal_8373, KeyReg_Inst_ff_SDE_62_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_63_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_8167, KeyExpansionOutput[63]}), .a ({new_AGEMA_signal_13836, new_AGEMA_signal_13832}), .c ({new_AGEMA_signal_8375, KeyReg_Inst_ff_SDE_63_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_64_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7527, KeyExpansionOutput[64]}), .a ({new_AGEMA_signal_13844, new_AGEMA_signal_13840}), .c ({new_AGEMA_signal_7664, KeyReg_Inst_ff_SDE_64_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_65_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7726, KeyExpansionOutput[65]}), .a ({new_AGEMA_signal_13852, new_AGEMA_signal_13848}), .c ({new_AGEMA_signal_7880, KeyReg_Inst_ff_SDE_65_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_66_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7720, KeyExpansionOutput[66]}), .a ({new_AGEMA_signal_13860, new_AGEMA_signal_13856}), .c ({new_AGEMA_signal_7882, KeyReg_Inst_ff_SDE_66_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_67_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7719, KeyExpansionOutput[67]}), .a ({new_AGEMA_signal_13868, new_AGEMA_signal_13864}), .c ({new_AGEMA_signal_7884, KeyReg_Inst_ff_SDE_67_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_68_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7718, KeyExpansionOutput[68]}), .a ({new_AGEMA_signal_13876, new_AGEMA_signal_13872}), .c ({new_AGEMA_signal_7886, KeyReg_Inst_ff_SDE_68_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_69_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7717, KeyExpansionOutput[69]}), .a ({new_AGEMA_signal_13884, new_AGEMA_signal_13880}), .c ({new_AGEMA_signal_7888, KeyReg_Inst_ff_SDE_69_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_70_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7716, KeyExpansionOutput[70]}), .a ({new_AGEMA_signal_13892, new_AGEMA_signal_13888}), .c ({new_AGEMA_signal_7890, KeyReg_Inst_ff_SDE_70_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_71_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7715, KeyExpansionOutput[71]}), .a ({new_AGEMA_signal_13900, new_AGEMA_signal_13896}), .c ({new_AGEMA_signal_7892, KeyReg_Inst_ff_SDE_71_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_72_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7503, KeyExpansionOutput[72]}), .a ({new_AGEMA_signal_13908, new_AGEMA_signal_13904}), .c ({new_AGEMA_signal_7666, KeyReg_Inst_ff_SDE_72_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_73_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7713, KeyExpansionOutput[73]}), .a ({new_AGEMA_signal_13916, new_AGEMA_signal_13912}), .c ({new_AGEMA_signal_7894, KeyReg_Inst_ff_SDE_73_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_74_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7743, KeyExpansionOutput[74]}), .a ({new_AGEMA_signal_13924, new_AGEMA_signal_13920}), .c ({new_AGEMA_signal_7896, KeyReg_Inst_ff_SDE_74_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_75_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7742, KeyExpansionOutput[75]}), .a ({new_AGEMA_signal_13932, new_AGEMA_signal_13928}), .c ({new_AGEMA_signal_7898, KeyReg_Inst_ff_SDE_75_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_76_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7734, KeyExpansionOutput[76]}), .a ({new_AGEMA_signal_13940, new_AGEMA_signal_13936}), .c ({new_AGEMA_signal_7900, KeyReg_Inst_ff_SDE_76_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_77_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7733, KeyExpansionOutput[77]}), .a ({new_AGEMA_signal_13948, new_AGEMA_signal_13944}), .c ({new_AGEMA_signal_7902, KeyReg_Inst_ff_SDE_77_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_78_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7732, KeyExpansionOutput[78]}), .a ({new_AGEMA_signal_13956, new_AGEMA_signal_13952}), .c ({new_AGEMA_signal_7904, KeyReg_Inst_ff_SDE_78_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_79_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7731, KeyExpansionOutput[79]}), .a ({new_AGEMA_signal_13964, new_AGEMA_signal_13960}), .c ({new_AGEMA_signal_7906, KeyReg_Inst_ff_SDE_79_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_80_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7507, KeyExpansionOutput[80]}), .a ({new_AGEMA_signal_13972, new_AGEMA_signal_13968}), .c ({new_AGEMA_signal_7668, KeyReg_Inst_ff_SDE_80_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_81_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7729, KeyExpansionOutput[81]}), .a ({new_AGEMA_signal_13980, new_AGEMA_signal_13976}), .c ({new_AGEMA_signal_7908, KeyReg_Inst_ff_SDE_81_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_82_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7728, KeyExpansionOutput[82]}), .a ({new_AGEMA_signal_13988, new_AGEMA_signal_13984}), .c ({new_AGEMA_signal_7910, KeyReg_Inst_ff_SDE_82_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_83_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7727, KeyExpansionOutput[83]}), .a ({new_AGEMA_signal_13996, new_AGEMA_signal_13992}), .c ({new_AGEMA_signal_7912, KeyReg_Inst_ff_SDE_83_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_84_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7725, KeyExpansionOutput[84]}), .a ({new_AGEMA_signal_14004, new_AGEMA_signal_14000}), .c ({new_AGEMA_signal_7914, KeyReg_Inst_ff_SDE_84_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_85_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7724, KeyExpansionOutput[85]}), .a ({new_AGEMA_signal_14012, new_AGEMA_signal_14008}), .c ({new_AGEMA_signal_7916, KeyReg_Inst_ff_SDE_85_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_86_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7723, KeyExpansionOutput[86]}), .a ({new_AGEMA_signal_14020, new_AGEMA_signal_14016}), .c ({new_AGEMA_signal_7918, KeyReg_Inst_ff_SDE_86_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_87_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7722, KeyExpansionOutput[87]}), .a ({new_AGEMA_signal_14028, new_AGEMA_signal_14024}), .c ({new_AGEMA_signal_7920, KeyReg_Inst_ff_SDE_87_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_88_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7721, KeyExpansionOutput[88]}), .a ({new_AGEMA_signal_14036, new_AGEMA_signal_14032}), .c ({new_AGEMA_signal_7922, KeyReg_Inst_ff_SDE_88_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_89_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7951, KeyExpansionOutput[89]}), .a ({new_AGEMA_signal_14044, new_AGEMA_signal_14040}), .c ({new_AGEMA_signal_8148, KeyReg_Inst_ff_SDE_89_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_90_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7950, KeyExpansionOutput[90]}), .a ({new_AGEMA_signal_14052, new_AGEMA_signal_14048}), .c ({new_AGEMA_signal_8150, KeyReg_Inst_ff_SDE_90_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_91_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7949, KeyExpansionOutput[91]}), .a ({new_AGEMA_signal_14060, new_AGEMA_signal_14056}), .c ({new_AGEMA_signal_8152, KeyReg_Inst_ff_SDE_91_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_92_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7948, KeyExpansionOutput[92]}), .a ({new_AGEMA_signal_14068, new_AGEMA_signal_14064}), .c ({new_AGEMA_signal_8154, KeyReg_Inst_ff_SDE_92_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_93_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7947, KeyExpansionOutput[93]}), .a ({new_AGEMA_signal_14076, new_AGEMA_signal_14072}), .c ({new_AGEMA_signal_8156, KeyReg_Inst_ff_SDE_93_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_94_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7945, KeyExpansionOutput[94]}), .a ({new_AGEMA_signal_14084, new_AGEMA_signal_14080}), .c ({new_AGEMA_signal_8158, KeyReg_Inst_ff_SDE_94_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_95_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7944, KeyExpansionOutput[95]}), .a ({new_AGEMA_signal_14092, new_AGEMA_signal_14088}), .c ({new_AGEMA_signal_8160, KeyReg_Inst_ff_SDE_95_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_96_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7355, KeyExpansionOutput[96]}), .a ({new_AGEMA_signal_14100, new_AGEMA_signal_14096}), .c ({new_AGEMA_signal_7498, KeyReg_Inst_ff_SDE_96_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_97_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7506, KeyExpansionOutput[97]}), .a ({new_AGEMA_signal_14108, new_AGEMA_signal_14104}), .c ({new_AGEMA_signal_7670, KeyReg_Inst_ff_SDE_97_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_98_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7505, KeyExpansionOutput[98]}), .a ({new_AGEMA_signal_14116, new_AGEMA_signal_14112}), .c ({new_AGEMA_signal_7672, KeyReg_Inst_ff_SDE_98_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_99_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7504, KeyExpansionOutput[99]}), .a ({new_AGEMA_signal_14124, new_AGEMA_signal_14120}), .c ({new_AGEMA_signal_7674, KeyReg_Inst_ff_SDE_99_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_100_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7526, KeyExpansionOutput[100]}), .a ({new_AGEMA_signal_14132, new_AGEMA_signal_14128}), .c ({new_AGEMA_signal_7676, KeyReg_Inst_ff_SDE_100_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_101_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7525, KeyExpansionOutput[101]}), .a ({new_AGEMA_signal_14140, new_AGEMA_signal_14136}), .c ({new_AGEMA_signal_7678, KeyReg_Inst_ff_SDE_101_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_102_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7524, KeyExpansionOutput[102]}), .a ({new_AGEMA_signal_14148, new_AGEMA_signal_14144}), .c ({new_AGEMA_signal_7680, KeyReg_Inst_ff_SDE_102_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_103_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7523, KeyExpansionOutput[103]}), .a ({new_AGEMA_signal_14156, new_AGEMA_signal_14152}), .c ({new_AGEMA_signal_7682, KeyReg_Inst_ff_SDE_103_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_104_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7354, KeyExpansionOutput[104]}), .a ({new_AGEMA_signal_14164, new_AGEMA_signal_14160}), .c ({new_AGEMA_signal_7500, KeyReg_Inst_ff_SDE_104_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_105_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7522, KeyExpansionOutput[105]}), .a ({new_AGEMA_signal_14172, new_AGEMA_signal_14168}), .c ({new_AGEMA_signal_7684, KeyReg_Inst_ff_SDE_105_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_106_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7521, KeyExpansionOutput[106]}), .a ({new_AGEMA_signal_14180, new_AGEMA_signal_14176}), .c ({new_AGEMA_signal_7686, KeyReg_Inst_ff_SDE_106_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_107_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7520, KeyExpansionOutput[107]}), .a ({new_AGEMA_signal_14188, new_AGEMA_signal_14184}), .c ({new_AGEMA_signal_7688, KeyReg_Inst_ff_SDE_107_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_108_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7519, KeyExpansionOutput[108]}), .a ({new_AGEMA_signal_14196, new_AGEMA_signal_14192}), .c ({new_AGEMA_signal_7690, KeyReg_Inst_ff_SDE_108_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_109_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7518, KeyExpansionOutput[109]}), .a ({new_AGEMA_signal_14204, new_AGEMA_signal_14200}), .c ({new_AGEMA_signal_7692, KeyReg_Inst_ff_SDE_109_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_110_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7517, KeyExpansionOutput[110]}), .a ({new_AGEMA_signal_14212, new_AGEMA_signal_14208}), .c ({new_AGEMA_signal_7694, KeyReg_Inst_ff_SDE_110_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_111_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7516, KeyExpansionOutput[111]}), .a ({new_AGEMA_signal_14220, new_AGEMA_signal_14216}), .c ({new_AGEMA_signal_7696, KeyReg_Inst_ff_SDE_111_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_112_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7353, KeyExpansionOutput[112]}), .a ({new_AGEMA_signal_14228, new_AGEMA_signal_14224}), .c ({new_AGEMA_signal_7502, KeyReg_Inst_ff_SDE_112_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_113_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7515, KeyExpansionOutput[113]}), .a ({new_AGEMA_signal_14236, new_AGEMA_signal_14232}), .c ({new_AGEMA_signal_7698, KeyReg_Inst_ff_SDE_113_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_114_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7514, KeyExpansionOutput[114]}), .a ({new_AGEMA_signal_14244, new_AGEMA_signal_14240}), .c ({new_AGEMA_signal_7700, KeyReg_Inst_ff_SDE_114_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_115_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7513, KeyExpansionOutput[115]}), .a ({new_AGEMA_signal_14252, new_AGEMA_signal_14248}), .c ({new_AGEMA_signal_7702, KeyReg_Inst_ff_SDE_115_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_116_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7512, KeyExpansionOutput[116]}), .a ({new_AGEMA_signal_14260, new_AGEMA_signal_14256}), .c ({new_AGEMA_signal_7704, KeyReg_Inst_ff_SDE_116_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_117_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7511, KeyExpansionOutput[117]}), .a ({new_AGEMA_signal_14268, new_AGEMA_signal_14264}), .c ({new_AGEMA_signal_7706, KeyReg_Inst_ff_SDE_117_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_118_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7510, KeyExpansionOutput[118]}), .a ({new_AGEMA_signal_14276, new_AGEMA_signal_14272}), .c ({new_AGEMA_signal_7708, KeyReg_Inst_ff_SDE_118_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_119_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7509, KeyExpansionOutput[119]}), .a ({new_AGEMA_signal_14284, new_AGEMA_signal_14280}), .c ({new_AGEMA_signal_7710, KeyReg_Inst_ff_SDE_119_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_120_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7508, KeyExpansionOutput[120]}), .a ({new_AGEMA_signal_14292, new_AGEMA_signal_14288}), .c ({new_AGEMA_signal_7712, KeyReg_Inst_ff_SDE_120_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_121_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7741, KeyExpansionOutput[121]}), .a ({new_AGEMA_signal_14300, new_AGEMA_signal_14296}), .c ({new_AGEMA_signal_7924, KeyReg_Inst_ff_SDE_121_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_122_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7740, KeyExpansionOutput[122]}), .a ({new_AGEMA_signal_14308, new_AGEMA_signal_14304}), .c ({new_AGEMA_signal_7926, KeyReg_Inst_ff_SDE_122_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_123_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7739, KeyExpansionOutput[123]}), .a ({new_AGEMA_signal_14316, new_AGEMA_signal_14312}), .c ({new_AGEMA_signal_7928, KeyReg_Inst_ff_SDE_123_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_124_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7738, KeyExpansionOutput[124]}), .a ({new_AGEMA_signal_14324, new_AGEMA_signal_14320}), .c ({new_AGEMA_signal_7930, KeyReg_Inst_ff_SDE_124_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_125_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7737, KeyExpansionOutput[125]}), .a ({new_AGEMA_signal_14332, new_AGEMA_signal_14328}), .c ({new_AGEMA_signal_7932, KeyReg_Inst_ff_SDE_125_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_126_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7736, KeyExpansionOutput[126]}), .a ({new_AGEMA_signal_14340, new_AGEMA_signal_14336}), .c ({new_AGEMA_signal_7934, KeyReg_Inst_ff_SDE_126_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_127_MUX_inst_U1 ( .s (new_AGEMA_signal_10572), .b ({new_AGEMA_signal_7735, KeyExpansionOutput[127]}), .a ({new_AGEMA_signal_14348, new_AGEMA_signal_14344}), .c ({new_AGEMA_signal_7936, KeyReg_Inst_ff_SDE_127_next_state}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U128 ( .a ({new_AGEMA_signal_14356, new_AGEMA_signal_14352}), .b ({new_AGEMA_signal_7938, KeyExpansionOutput[41]}), .c ({new_AGEMA_signal_8161, KeyExpansionOutput[9]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U127 ( .a ({new_AGEMA_signal_14364, new_AGEMA_signal_14360}), .b ({new_AGEMA_signal_7714, KeyExpansionOutput[40]}), .c ({new_AGEMA_signal_7937, KeyExpansionOutput[8]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U126 ( .a ({new_AGEMA_signal_14372, new_AGEMA_signal_14368}), .b ({new_AGEMA_signal_7939, KeyExpansionOutput[39]}), .c ({new_AGEMA_signal_8162, KeyExpansionOutput[7]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U125 ( .a ({new_AGEMA_signal_14380, new_AGEMA_signal_14376}), .b ({new_AGEMA_signal_7940, KeyExpansionOutput[38]}), .c ({new_AGEMA_signal_8163, KeyExpansionOutput[6]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U124 ( .a ({new_AGEMA_signal_14388, new_AGEMA_signal_14384}), .b ({new_AGEMA_signal_7941, KeyExpansionOutput[37]}), .c ({new_AGEMA_signal_8164, KeyExpansionOutput[5]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U123 ( .a ({new_AGEMA_signal_14396, new_AGEMA_signal_14392}), .b ({new_AGEMA_signal_7942, KeyExpansionOutput[36]}), .c ({new_AGEMA_signal_8165, KeyExpansionOutput[4]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U122 ( .a ({new_AGEMA_signal_14404, new_AGEMA_signal_14400}), .b ({new_AGEMA_signal_7713, KeyExpansionOutput[73]}), .c ({new_AGEMA_signal_7938, KeyExpansionOutput[41]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U121 ( .a ({new_AGEMA_signal_14412, new_AGEMA_signal_14408}), .b ({new_AGEMA_signal_7522, KeyExpansionOutput[105]}), .c ({new_AGEMA_signal_7713, KeyExpansionOutput[73]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U120 ( .a ({new_AGEMA_signal_14420, new_AGEMA_signal_14416}), .b ({new_AGEMA_signal_7503, KeyExpansionOutput[72]}), .c ({new_AGEMA_signal_7714, KeyExpansionOutput[40]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U119 ( .a ({new_AGEMA_signal_14428, new_AGEMA_signal_14424}), .b ({new_AGEMA_signal_7354, KeyExpansionOutput[104]}), .c ({new_AGEMA_signal_7503, KeyExpansionOutput[72]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U118 ( .a ({new_AGEMA_signal_14436, new_AGEMA_signal_14432}), .b ({new_AGEMA_signal_7943, KeyExpansionOutput[35]}), .c ({new_AGEMA_signal_8166, KeyExpansionOutput[3]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U117 ( .a ({new_AGEMA_signal_14444, new_AGEMA_signal_14440}), .b ({new_AGEMA_signal_7715, KeyExpansionOutput[71]}), .c ({new_AGEMA_signal_7939, KeyExpansionOutput[39]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U116 ( .a ({new_AGEMA_signal_14452, new_AGEMA_signal_14448}), .b ({new_AGEMA_signal_7523, KeyExpansionOutput[103]}), .c ({new_AGEMA_signal_7715, KeyExpansionOutput[71]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U115 ( .a ({new_AGEMA_signal_14460, new_AGEMA_signal_14456}), .b ({new_AGEMA_signal_7716, KeyExpansionOutput[70]}), .c ({new_AGEMA_signal_7940, KeyExpansionOutput[38]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U114 ( .a ({new_AGEMA_signal_14468, new_AGEMA_signal_14464}), .b ({new_AGEMA_signal_7524, KeyExpansionOutput[102]}), .c ({new_AGEMA_signal_7716, KeyExpansionOutput[70]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U113 ( .a ({new_AGEMA_signal_14476, new_AGEMA_signal_14472}), .b ({new_AGEMA_signal_7717, KeyExpansionOutput[69]}), .c ({new_AGEMA_signal_7941, KeyExpansionOutput[37]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U112 ( .a ({new_AGEMA_signal_14484, new_AGEMA_signal_14480}), .b ({new_AGEMA_signal_7525, KeyExpansionOutput[101]}), .c ({new_AGEMA_signal_7717, KeyExpansionOutput[69]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U111 ( .a ({new_AGEMA_signal_14492, new_AGEMA_signal_14488}), .b ({new_AGEMA_signal_7718, KeyExpansionOutput[68]}), .c ({new_AGEMA_signal_7942, KeyExpansionOutput[36]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U110 ( .a ({new_AGEMA_signal_14500, new_AGEMA_signal_14496}), .b ({new_AGEMA_signal_7526, KeyExpansionOutput[100]}), .c ({new_AGEMA_signal_7718, KeyExpansionOutput[68]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U109 ( .a ({new_AGEMA_signal_14508, new_AGEMA_signal_14504}), .b ({new_AGEMA_signal_7719, KeyExpansionOutput[67]}), .c ({new_AGEMA_signal_7943, KeyExpansionOutput[35]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U108 ( .a ({new_AGEMA_signal_14516, new_AGEMA_signal_14512}), .b ({new_AGEMA_signal_7504, KeyExpansionOutput[99]}), .c ({new_AGEMA_signal_7719, KeyExpansionOutput[67]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U107 ( .a ({new_AGEMA_signal_14524, new_AGEMA_signal_14520}), .b ({new_AGEMA_signal_7382, KeyExpansionIns_tmp[3]}), .c ({new_AGEMA_signal_7504, KeyExpansionOutput[99]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U106 ( .a ({new_AGEMA_signal_14532, new_AGEMA_signal_14528}), .b ({new_AGEMA_signal_8167, KeyExpansionOutput[63]}), .c ({new_AGEMA_signal_8376, KeyExpansionOutput[31]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U105 ( .a ({new_AGEMA_signal_14540, new_AGEMA_signal_14536}), .b ({new_AGEMA_signal_7944, KeyExpansionOutput[95]}), .c ({new_AGEMA_signal_8167, KeyExpansionOutput[63]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U104 ( .a ({new_AGEMA_signal_14548, new_AGEMA_signal_14544}), .b ({new_AGEMA_signal_7735, KeyExpansionOutput[127]}), .c ({new_AGEMA_signal_7944, KeyExpansionOutput[95]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U103 ( .a ({new_AGEMA_signal_14556, new_AGEMA_signal_14552}), .b ({new_AGEMA_signal_8168, KeyExpansionOutput[62]}), .c ({new_AGEMA_signal_8377, KeyExpansionOutput[30]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U102 ( .a ({new_AGEMA_signal_14564, new_AGEMA_signal_14560}), .b ({new_AGEMA_signal_7945, KeyExpansionOutput[94]}), .c ({new_AGEMA_signal_8168, KeyExpansionOutput[62]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U101 ( .a ({new_AGEMA_signal_14572, new_AGEMA_signal_14568}), .b ({new_AGEMA_signal_7736, KeyExpansionOutput[126]}), .c ({new_AGEMA_signal_7945, KeyExpansionOutput[94]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U100 ( .a ({new_AGEMA_signal_14580, new_AGEMA_signal_14576}), .b ({new_AGEMA_signal_7946, KeyExpansionOutput[34]}), .c ({new_AGEMA_signal_8169, KeyExpansionOutput[2]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U99 ( .a ({new_AGEMA_signal_14588, new_AGEMA_signal_14584}), .b ({new_AGEMA_signal_7720, KeyExpansionOutput[66]}), .c ({new_AGEMA_signal_7946, KeyExpansionOutput[34]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U98 ( .a ({new_AGEMA_signal_14596, new_AGEMA_signal_14592}), .b ({new_AGEMA_signal_7505, KeyExpansionOutput[98]}), .c ({new_AGEMA_signal_7720, KeyExpansionOutput[66]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U97 ( .a ({new_AGEMA_signal_14604, new_AGEMA_signal_14600}), .b ({new_AGEMA_signal_7383, KeyExpansionIns_tmp[2]}), .c ({new_AGEMA_signal_7505, KeyExpansionOutput[98]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U96 ( .a ({new_AGEMA_signal_14612, new_AGEMA_signal_14608}), .b ({new_AGEMA_signal_8170, KeyExpansionOutput[61]}), .c ({new_AGEMA_signal_8378, KeyExpansionOutput[29]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U95 ( .a ({new_AGEMA_signal_14620, new_AGEMA_signal_14616}), .b ({new_AGEMA_signal_7947, KeyExpansionOutput[93]}), .c ({new_AGEMA_signal_8170, KeyExpansionOutput[61]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U94 ( .a ({new_AGEMA_signal_14628, new_AGEMA_signal_14624}), .b ({new_AGEMA_signal_7737, KeyExpansionOutput[125]}), .c ({new_AGEMA_signal_7947, KeyExpansionOutput[93]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U93 ( .a ({new_AGEMA_signal_14636, new_AGEMA_signal_14632}), .b ({new_AGEMA_signal_8171, KeyExpansionOutput[60]}), .c ({new_AGEMA_signal_8379, KeyExpansionOutput[28]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U92 ( .a ({new_AGEMA_signal_14644, new_AGEMA_signal_14640}), .b ({new_AGEMA_signal_7948, KeyExpansionOutput[92]}), .c ({new_AGEMA_signal_8171, KeyExpansionOutput[60]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U91 ( .a ({new_AGEMA_signal_14652, new_AGEMA_signal_14648}), .b ({new_AGEMA_signal_7738, KeyExpansionOutput[124]}), .c ({new_AGEMA_signal_7948, KeyExpansionOutput[92]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U90 ( .a ({new_AGEMA_signal_14660, new_AGEMA_signal_14656}), .b ({new_AGEMA_signal_8172, KeyExpansionOutput[59]}), .c ({new_AGEMA_signal_8380, KeyExpansionOutput[27]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U89 ( .a ({new_AGEMA_signal_14668, new_AGEMA_signal_14664}), .b ({new_AGEMA_signal_7949, KeyExpansionOutput[91]}), .c ({new_AGEMA_signal_8172, KeyExpansionOutput[59]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U88 ( .a ({new_AGEMA_signal_14676, new_AGEMA_signal_14672}), .b ({new_AGEMA_signal_7739, KeyExpansionOutput[123]}), .c ({new_AGEMA_signal_7949, KeyExpansionOutput[91]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U87 ( .a ({new_AGEMA_signal_14684, new_AGEMA_signal_14680}), .b ({new_AGEMA_signal_8173, KeyExpansionOutput[58]}), .c ({new_AGEMA_signal_8381, KeyExpansionOutput[26]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U86 ( .a ({new_AGEMA_signal_14692, new_AGEMA_signal_14688}), .b ({new_AGEMA_signal_7950, KeyExpansionOutput[90]}), .c ({new_AGEMA_signal_8173, KeyExpansionOutput[58]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U85 ( .a ({new_AGEMA_signal_14700, new_AGEMA_signal_14696}), .b ({new_AGEMA_signal_7740, KeyExpansionOutput[122]}), .c ({new_AGEMA_signal_7950, KeyExpansionOutput[90]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U84 ( .a ({new_AGEMA_signal_14708, new_AGEMA_signal_14704}), .b ({new_AGEMA_signal_8174, KeyExpansionOutput[57]}), .c ({new_AGEMA_signal_8382, KeyExpansionOutput[25]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U83 ( .a ({new_AGEMA_signal_14716, new_AGEMA_signal_14712}), .b ({new_AGEMA_signal_7951, KeyExpansionOutput[89]}), .c ({new_AGEMA_signal_8174, KeyExpansionOutput[57]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U82 ( .a ({new_AGEMA_signal_14724, new_AGEMA_signal_14720}), .b ({new_AGEMA_signal_7741, KeyExpansionOutput[121]}), .c ({new_AGEMA_signal_7951, KeyExpansionOutput[89]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U81 ( .a ({new_AGEMA_signal_14732, new_AGEMA_signal_14728}), .b ({new_AGEMA_signal_7952, KeyExpansionOutput[56]}), .c ({new_AGEMA_signal_8175, KeyExpansionOutput[24]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U80 ( .a ({new_AGEMA_signal_14740, new_AGEMA_signal_14736}), .b ({new_AGEMA_signal_7721, KeyExpansionOutput[88]}), .c ({new_AGEMA_signal_7952, KeyExpansionOutput[56]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U79 ( .a ({new_AGEMA_signal_14748, new_AGEMA_signal_14744}), .b ({new_AGEMA_signal_7508, KeyExpansionOutput[120]}), .c ({new_AGEMA_signal_7721, KeyExpansionOutput[88]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U78 ( .a ({new_AGEMA_signal_14756, new_AGEMA_signal_14752}), .b ({new_AGEMA_signal_7953, KeyExpansionOutput[55]}), .c ({new_AGEMA_signal_8176, KeyExpansionOutput[23]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U77 ( .a ({new_AGEMA_signal_14764, new_AGEMA_signal_14760}), .b ({new_AGEMA_signal_7722, KeyExpansionOutput[87]}), .c ({new_AGEMA_signal_7953, KeyExpansionOutput[55]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U76 ( .a ({new_AGEMA_signal_14772, new_AGEMA_signal_14768}), .b ({new_AGEMA_signal_7509, KeyExpansionOutput[119]}), .c ({new_AGEMA_signal_7722, KeyExpansionOutput[87]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U75 ( .a ({new_AGEMA_signal_14780, new_AGEMA_signal_14776}), .b ({new_AGEMA_signal_7954, KeyExpansionOutput[54]}), .c ({new_AGEMA_signal_8177, KeyExpansionOutput[22]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U74 ( .a ({new_AGEMA_signal_14788, new_AGEMA_signal_14784}), .b ({new_AGEMA_signal_7723, KeyExpansionOutput[86]}), .c ({new_AGEMA_signal_7954, KeyExpansionOutput[54]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U73 ( .a ({new_AGEMA_signal_14796, new_AGEMA_signal_14792}), .b ({new_AGEMA_signal_7510, KeyExpansionOutput[118]}), .c ({new_AGEMA_signal_7723, KeyExpansionOutput[86]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U72 ( .a ({new_AGEMA_signal_14804, new_AGEMA_signal_14800}), .b ({new_AGEMA_signal_7955, KeyExpansionOutput[53]}), .c ({new_AGEMA_signal_8178, KeyExpansionOutput[21]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U71 ( .a ({new_AGEMA_signal_14812, new_AGEMA_signal_14808}), .b ({new_AGEMA_signal_7724, KeyExpansionOutput[85]}), .c ({new_AGEMA_signal_7955, KeyExpansionOutput[53]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U70 ( .a ({new_AGEMA_signal_14820, new_AGEMA_signal_14816}), .b ({new_AGEMA_signal_7511, KeyExpansionOutput[117]}), .c ({new_AGEMA_signal_7724, KeyExpansionOutput[85]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U69 ( .a ({new_AGEMA_signal_14828, new_AGEMA_signal_14824}), .b ({new_AGEMA_signal_7956, KeyExpansionOutput[52]}), .c ({new_AGEMA_signal_8179, KeyExpansionOutput[20]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U68 ( .a ({new_AGEMA_signal_14836, new_AGEMA_signal_14832}), .b ({new_AGEMA_signal_7725, KeyExpansionOutput[84]}), .c ({new_AGEMA_signal_7956, KeyExpansionOutput[52]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U67 ( .a ({new_AGEMA_signal_14844, new_AGEMA_signal_14840}), .b ({new_AGEMA_signal_7512, KeyExpansionOutput[116]}), .c ({new_AGEMA_signal_7725, KeyExpansionOutput[84]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U66 ( .a ({new_AGEMA_signal_14852, new_AGEMA_signal_14848}), .b ({new_AGEMA_signal_7957, KeyExpansionOutput[33]}), .c ({new_AGEMA_signal_8180, KeyExpansionOutput[1]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U65 ( .a ({new_AGEMA_signal_14860, new_AGEMA_signal_14856}), .b ({new_AGEMA_signal_7726, KeyExpansionOutput[65]}), .c ({new_AGEMA_signal_7957, KeyExpansionOutput[33]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U64 ( .a ({new_AGEMA_signal_14868, new_AGEMA_signal_14864}), .b ({new_AGEMA_signal_7506, KeyExpansionOutput[97]}), .c ({new_AGEMA_signal_7726, KeyExpansionOutput[65]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U63 ( .a ({new_AGEMA_signal_14876, new_AGEMA_signal_14872}), .b ({new_AGEMA_signal_7384, KeyExpansionIns_tmp[1]}), .c ({new_AGEMA_signal_7506, KeyExpansionOutput[97]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U62 ( .a ({new_AGEMA_signal_14884, new_AGEMA_signal_14880}), .b ({new_AGEMA_signal_7958, KeyExpansionOutput[51]}), .c ({new_AGEMA_signal_8181, KeyExpansionOutput[19]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U61 ( .a ({new_AGEMA_signal_14892, new_AGEMA_signal_14888}), .b ({new_AGEMA_signal_7727, KeyExpansionOutput[83]}), .c ({new_AGEMA_signal_7958, KeyExpansionOutput[51]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U60 ( .a ({new_AGEMA_signal_14900, new_AGEMA_signal_14896}), .b ({new_AGEMA_signal_7513, KeyExpansionOutput[115]}), .c ({new_AGEMA_signal_7727, KeyExpansionOutput[83]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U59 ( .a ({new_AGEMA_signal_14908, new_AGEMA_signal_14904}), .b ({new_AGEMA_signal_7959, KeyExpansionOutput[50]}), .c ({new_AGEMA_signal_8182, KeyExpansionOutput[18]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U58 ( .a ({new_AGEMA_signal_14916, new_AGEMA_signal_14912}), .b ({new_AGEMA_signal_7728, KeyExpansionOutput[82]}), .c ({new_AGEMA_signal_7959, KeyExpansionOutput[50]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U57 ( .a ({new_AGEMA_signal_14924, new_AGEMA_signal_14920}), .b ({new_AGEMA_signal_7514, KeyExpansionOutput[114]}), .c ({new_AGEMA_signal_7728, KeyExpansionOutput[82]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U56 ( .a ({new_AGEMA_signal_14932, new_AGEMA_signal_14928}), .b ({new_AGEMA_signal_7960, KeyExpansionOutput[49]}), .c ({new_AGEMA_signal_8183, KeyExpansionOutput[17]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U55 ( .a ({new_AGEMA_signal_14940, new_AGEMA_signal_14936}), .b ({new_AGEMA_signal_7729, KeyExpansionOutput[81]}), .c ({new_AGEMA_signal_7960, KeyExpansionOutput[49]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U54 ( .a ({new_AGEMA_signal_14948, new_AGEMA_signal_14944}), .b ({new_AGEMA_signal_7515, KeyExpansionOutput[113]}), .c ({new_AGEMA_signal_7729, KeyExpansionOutput[81]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U53 ( .a ({new_AGEMA_signal_14956, new_AGEMA_signal_14952}), .b ({new_AGEMA_signal_7730, KeyExpansionOutput[48]}), .c ({new_AGEMA_signal_7961, KeyExpansionOutput[16]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U52 ( .a ({new_AGEMA_signal_14964, new_AGEMA_signal_14960}), .b ({new_AGEMA_signal_7507, KeyExpansionOutput[80]}), .c ({new_AGEMA_signal_7730, KeyExpansionOutput[48]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U51 ( .a ({new_AGEMA_signal_14972, new_AGEMA_signal_14968}), .b ({new_AGEMA_signal_7353, KeyExpansionOutput[112]}), .c ({new_AGEMA_signal_7507, KeyExpansionOutput[80]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U50 ( .a ({new_AGEMA_signal_14980, new_AGEMA_signal_14976}), .b ({new_AGEMA_signal_7962, KeyExpansionOutput[47]}), .c ({new_AGEMA_signal_8184, KeyExpansionOutput[15]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U49 ( .a ({new_AGEMA_signal_14988, new_AGEMA_signal_14984}), .b ({new_AGEMA_signal_7731, KeyExpansionOutput[79]}), .c ({new_AGEMA_signal_7962, KeyExpansionOutput[47]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U48 ( .a ({new_AGEMA_signal_14996, new_AGEMA_signal_14992}), .b ({new_AGEMA_signal_7516, KeyExpansionOutput[111]}), .c ({new_AGEMA_signal_7731, KeyExpansionOutput[79]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U47 ( .a ({new_AGEMA_signal_15004, new_AGEMA_signal_15000}), .b ({new_AGEMA_signal_7963, KeyExpansionOutput[46]}), .c ({new_AGEMA_signal_8185, KeyExpansionOutput[14]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U46 ( .a ({new_AGEMA_signal_15012, new_AGEMA_signal_15008}), .b ({new_AGEMA_signal_7732, KeyExpansionOutput[78]}), .c ({new_AGEMA_signal_7963, KeyExpansionOutput[46]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U45 ( .a ({new_AGEMA_signal_15020, new_AGEMA_signal_15016}), .b ({new_AGEMA_signal_7517, KeyExpansionOutput[110]}), .c ({new_AGEMA_signal_7732, KeyExpansionOutput[78]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U44 ( .a ({new_AGEMA_signal_15028, new_AGEMA_signal_15024}), .b ({new_AGEMA_signal_7964, KeyExpansionOutput[45]}), .c ({new_AGEMA_signal_8186, KeyExpansionOutput[13]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U43 ( .a ({new_AGEMA_signal_15036, new_AGEMA_signal_15032}), .b ({new_AGEMA_signal_7733, KeyExpansionOutput[77]}), .c ({new_AGEMA_signal_7964, KeyExpansionOutput[45]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U42 ( .a ({new_AGEMA_signal_15044, new_AGEMA_signal_15040}), .b ({new_AGEMA_signal_7518, KeyExpansionOutput[109]}), .c ({new_AGEMA_signal_7733, KeyExpansionOutput[77]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U41 ( .a ({new_AGEMA_signal_15052, new_AGEMA_signal_15048}), .b ({new_AGEMA_signal_7965, KeyExpansionOutput[44]}), .c ({new_AGEMA_signal_8187, KeyExpansionOutput[12]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U40 ( .a ({new_AGEMA_signal_15060, new_AGEMA_signal_15056}), .b ({new_AGEMA_signal_7734, KeyExpansionOutput[76]}), .c ({new_AGEMA_signal_7965, KeyExpansionOutput[44]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U39 ( .a ({new_AGEMA_signal_15068, new_AGEMA_signal_15064}), .b ({new_AGEMA_signal_7519, KeyExpansionOutput[108]}), .c ({new_AGEMA_signal_7734, KeyExpansionOutput[76]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U38 ( .a ({new_AGEMA_signal_15076, new_AGEMA_signal_15072}), .b ({new_AGEMA_signal_7528, KeyExpansionIns_tmp[31]}), .c ({new_AGEMA_signal_7735, KeyExpansionOutput[127]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U37 ( .a ({new_AGEMA_signal_15084, new_AGEMA_signal_15080}), .b ({new_AGEMA_signal_7529, KeyExpansionIns_tmp[30]}), .c ({new_AGEMA_signal_7736, KeyExpansionOutput[126]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U36 ( .a ({new_AGEMA_signal_15092, new_AGEMA_signal_15088}), .b ({new_AGEMA_signal_7530, KeyExpansionIns_tmp[29]}), .c ({new_AGEMA_signal_7737, KeyExpansionOutput[125]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U35 ( .a ({new_AGEMA_signal_15100, new_AGEMA_signal_15096}), .b ({new_AGEMA_signal_7531, KeyExpansionIns_tmp[28]}), .c ({new_AGEMA_signal_7738, KeyExpansionOutput[124]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U34 ( .a ({new_AGEMA_signal_15108, new_AGEMA_signal_15104}), .b ({new_AGEMA_signal_7532, KeyExpansionIns_tmp[27]}), .c ({new_AGEMA_signal_7739, KeyExpansionOutput[123]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U33 ( .a ({new_AGEMA_signal_15116, new_AGEMA_signal_15112}), .b ({new_AGEMA_signal_7533, KeyExpansionIns_tmp[26]}), .c ({new_AGEMA_signal_7740, KeyExpansionOutput[122]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U32 ( .a ({new_AGEMA_signal_15124, new_AGEMA_signal_15120}), .b ({new_AGEMA_signal_7534, KeyExpansionIns_tmp[25]}), .c ({new_AGEMA_signal_7741, KeyExpansionOutput[121]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U31 ( .a ({new_AGEMA_signal_15132, new_AGEMA_signal_15128}), .b ({new_AGEMA_signal_7356, KeyExpansionIns_tmp[24]}), .c ({new_AGEMA_signal_7508, KeyExpansionOutput[120]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U30 ( .a ({new_AGEMA_signal_15140, new_AGEMA_signal_15136}), .b ({new_AGEMA_signal_7966, KeyExpansionOutput[43]}), .c ({new_AGEMA_signal_8188, KeyExpansionOutput[11]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U29 ( .a ({new_AGEMA_signal_15148, new_AGEMA_signal_15144}), .b ({new_AGEMA_signal_7742, KeyExpansionOutput[75]}), .c ({new_AGEMA_signal_7966, KeyExpansionOutput[43]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U28 ( .a ({new_AGEMA_signal_15156, new_AGEMA_signal_15152}), .b ({new_AGEMA_signal_7520, KeyExpansionOutput[107]}), .c ({new_AGEMA_signal_7742, KeyExpansionOutput[75]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U27 ( .a ({new_AGEMA_signal_15164, new_AGEMA_signal_15160}), .b ({new_AGEMA_signal_7364, KeyExpansionIns_tmp[23]}), .c ({new_AGEMA_signal_7509, KeyExpansionOutput[119]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U26 ( .a ({new_AGEMA_signal_15172, new_AGEMA_signal_15168}), .b ({new_AGEMA_signal_7365, KeyExpansionIns_tmp[22]}), .c ({new_AGEMA_signal_7510, KeyExpansionOutput[118]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U25 ( .a ({new_AGEMA_signal_15180, new_AGEMA_signal_15176}), .b ({new_AGEMA_signal_7366, KeyExpansionIns_tmp[21]}), .c ({new_AGEMA_signal_7511, KeyExpansionOutput[117]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U24 ( .a ({new_AGEMA_signal_15188, new_AGEMA_signal_15184}), .b ({new_AGEMA_signal_7367, KeyExpansionIns_tmp[20]}), .c ({new_AGEMA_signal_7512, KeyExpansionOutput[116]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U23 ( .a ({new_AGEMA_signal_15196, new_AGEMA_signal_15192}), .b ({new_AGEMA_signal_7368, KeyExpansionIns_tmp[19]}), .c ({new_AGEMA_signal_7513, KeyExpansionOutput[115]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U22 ( .a ({new_AGEMA_signal_15204, new_AGEMA_signal_15200}), .b ({new_AGEMA_signal_7369, KeyExpansionIns_tmp[18]}), .c ({new_AGEMA_signal_7514, KeyExpansionOutput[114]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U21 ( .a ({new_AGEMA_signal_15212, new_AGEMA_signal_15208}), .b ({new_AGEMA_signal_7370, KeyExpansionIns_tmp[17]}), .c ({new_AGEMA_signal_7515, KeyExpansionOutput[113]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U20 ( .a ({new_AGEMA_signal_15220, new_AGEMA_signal_15216}), .b ({new_AGEMA_signal_7154, KeyExpansionIns_tmp[16]}), .c ({new_AGEMA_signal_7353, KeyExpansionOutput[112]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U19 ( .a ({new_AGEMA_signal_15228, new_AGEMA_signal_15224}), .b ({new_AGEMA_signal_7371, KeyExpansionIns_tmp[15]}), .c ({new_AGEMA_signal_7516, KeyExpansionOutput[111]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U18 ( .a ({new_AGEMA_signal_15236, new_AGEMA_signal_15232}), .b ({new_AGEMA_signal_7372, KeyExpansionIns_tmp[14]}), .c ({new_AGEMA_signal_7517, KeyExpansionOutput[110]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U17 ( .a ({new_AGEMA_signal_15244, new_AGEMA_signal_15240}), .b ({new_AGEMA_signal_7967, KeyExpansionOutput[42]}), .c ({new_AGEMA_signal_8189, KeyExpansionOutput[10]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U16 ( .a ({new_AGEMA_signal_15252, new_AGEMA_signal_15248}), .b ({new_AGEMA_signal_7743, KeyExpansionOutput[74]}), .c ({new_AGEMA_signal_7967, KeyExpansionOutput[42]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U15 ( .a ({new_AGEMA_signal_15260, new_AGEMA_signal_15256}), .b ({new_AGEMA_signal_7521, KeyExpansionOutput[106]}), .c ({new_AGEMA_signal_7743, KeyExpansionOutput[74]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U14 ( .a ({new_AGEMA_signal_15268, new_AGEMA_signal_15264}), .b ({new_AGEMA_signal_7373, KeyExpansionIns_tmp[13]}), .c ({new_AGEMA_signal_7518, KeyExpansionOutput[109]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U13 ( .a ({new_AGEMA_signal_15276, new_AGEMA_signal_15272}), .b ({new_AGEMA_signal_7374, KeyExpansionIns_tmp[12]}), .c ({new_AGEMA_signal_7519, KeyExpansionOutput[108]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U12 ( .a ({new_AGEMA_signal_15284, new_AGEMA_signal_15280}), .b ({new_AGEMA_signal_7375, KeyExpansionIns_tmp[11]}), .c ({new_AGEMA_signal_7520, KeyExpansionOutput[107]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U11 ( .a ({new_AGEMA_signal_15292, new_AGEMA_signal_15288}), .b ({new_AGEMA_signal_7376, KeyExpansionIns_tmp[10]}), .c ({new_AGEMA_signal_7521, KeyExpansionOutput[106]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U10 ( .a ({new_AGEMA_signal_15300, new_AGEMA_signal_15296}), .b ({new_AGEMA_signal_7377, KeyExpansionIns_tmp[9]}), .c ({new_AGEMA_signal_7522, KeyExpansionOutput[105]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U9 ( .a ({new_AGEMA_signal_15308, new_AGEMA_signal_15304}), .b ({new_AGEMA_signal_7165, KeyExpansionIns_tmp[8]}), .c ({new_AGEMA_signal_7354, KeyExpansionOutput[104]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U8 ( .a ({new_AGEMA_signal_15316, new_AGEMA_signal_15312}), .b ({new_AGEMA_signal_7378, KeyExpansionIns_tmp[7]}), .c ({new_AGEMA_signal_7523, KeyExpansionOutput[103]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U7 ( .a ({new_AGEMA_signal_15324, new_AGEMA_signal_15320}), .b ({new_AGEMA_signal_7379, KeyExpansionIns_tmp[6]}), .c ({new_AGEMA_signal_7524, KeyExpansionOutput[102]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U6 ( .a ({new_AGEMA_signal_15332, new_AGEMA_signal_15328}), .b ({new_AGEMA_signal_7380, KeyExpansionIns_tmp[5]}), .c ({new_AGEMA_signal_7525, KeyExpansionOutput[101]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U5 ( .a ({new_AGEMA_signal_15340, new_AGEMA_signal_15336}), .b ({new_AGEMA_signal_7381, KeyExpansionIns_tmp[4]}), .c ({new_AGEMA_signal_7526, KeyExpansionOutput[100]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U4 ( .a ({new_AGEMA_signal_15348, new_AGEMA_signal_15344}), .b ({new_AGEMA_signal_7744, KeyExpansionOutput[32]}), .c ({new_AGEMA_signal_7968, KeyExpansionOutput[0]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U3 ( .a ({new_AGEMA_signal_15356, new_AGEMA_signal_15352}), .b ({new_AGEMA_signal_7527, KeyExpansionOutput[64]}), .c ({new_AGEMA_signal_7744, KeyExpansionOutput[32]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U2 ( .a ({new_AGEMA_signal_15364, new_AGEMA_signal_15360}), .b ({new_AGEMA_signal_7355, KeyExpansionOutput[96]}), .c ({new_AGEMA_signal_7527, KeyExpansionOutput[64]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U1 ( .a ({new_AGEMA_signal_15372, new_AGEMA_signal_15368}), .b ({new_AGEMA_signal_7176, KeyExpansionIns_tmp[0]}), .c ({new_AGEMA_signal_7355, KeyExpansionOutput[96]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U8 ( .a ({new_AGEMA_signal_7357, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__7_}), .b ({1'b0, new_AGEMA_signal_15376}), .c ({new_AGEMA_signal_7528, KeyExpansionIns_tmp[31]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U7 ( .a ({new_AGEMA_signal_7358, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__6_}), .b ({1'b0, new_AGEMA_signal_15380}), .c ({new_AGEMA_signal_7529, KeyExpansionIns_tmp[30]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U6 ( .a ({new_AGEMA_signal_7359, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__5_}), .b ({1'b0, new_AGEMA_signal_15384}), .c ({new_AGEMA_signal_7530, KeyExpansionIns_tmp[29]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U5 ( .a ({new_AGEMA_signal_7360, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__4_}), .b ({1'b0, new_AGEMA_signal_15388}), .c ({new_AGEMA_signal_7531, KeyExpansionIns_tmp[28]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U4 ( .a ({new_AGEMA_signal_7361, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__3_}), .b ({1'b0, new_AGEMA_signal_15392}), .c ({new_AGEMA_signal_7532, KeyExpansionIns_tmp[27]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U3 ( .a ({new_AGEMA_signal_7362, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__2_}), .b ({1'b0, new_AGEMA_signal_15396}), .c ({new_AGEMA_signal_7533, KeyExpansionIns_tmp[26]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U2 ( .a ({new_AGEMA_signal_7363, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__1_}), .b ({1'b0, new_AGEMA_signal_15400}), .c ({new_AGEMA_signal_7534, KeyExpansionIns_tmp[25]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U1 ( .a ({new_AGEMA_signal_7143, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__0_}), .b ({1'b0, new_AGEMA_signal_15404}), .c ({new_AGEMA_signal_7356, KeyExpansionIns_tmp[24]}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M46_U1 ( .a ({new_AGEMA_signal_6276, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_15410, new_AGEMA_signal_15407}), .clk (clk), .r ({Fresh[1217], Fresh[1216]}), .c ({new_AGEMA_signal_6514, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M47_U1 ( .a ({new_AGEMA_signal_6196, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_15416, new_AGEMA_signal_15413}), .clk (clk), .r ({Fresh[1219], Fresh[1218]}), .c ({new_AGEMA_signal_6277, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M47}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M48_U1 ( .a ({new_AGEMA_signal_6195, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_14955, new_AGEMA_signal_14951}), .clk (clk), .r ({Fresh[1221], Fresh[1220]}), .c ({new_AGEMA_signal_6278, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M49_U1 ( .a ({new_AGEMA_signal_6275, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_15422, new_AGEMA_signal_15419}), .clk (clk), .r ({Fresh[1223], Fresh[1222]}), .c ({new_AGEMA_signal_6515, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M49}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M50_U1 ( .a ({new_AGEMA_signal_6194, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_15428, new_AGEMA_signal_15425}), .clk (clk), .r ({Fresh[1225], Fresh[1224]}), .c ({new_AGEMA_signal_6279, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M51_U1 ( .a ({new_AGEMA_signal_6193, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_15434, new_AGEMA_signal_15431}), .clk (clk), .r ({Fresh[1227], Fresh[1226]}), .c ({new_AGEMA_signal_6280, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M52_U1 ( .a ({new_AGEMA_signal_6274, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_15440, new_AGEMA_signal_15437}), .clk (clk), .r ({Fresh[1229], Fresh[1228]}), .c ({new_AGEMA_signal_6516, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M53_U1 ( .a ({new_AGEMA_signal_6513, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_15446, new_AGEMA_signal_15443}), .clk (clk), .r ({Fresh[1231], Fresh[1230]}), .c ({new_AGEMA_signal_6753, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M54_U1 ( .a ({new_AGEMA_signal_6273, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_15452, new_AGEMA_signal_15449}), .clk (clk), .r ({Fresh[1233], Fresh[1232]}), .c ({new_AGEMA_signal_6517, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M54}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M55_U1 ( .a ({new_AGEMA_signal_6276, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_15458, new_AGEMA_signal_15455}), .clk (clk), .r ({Fresh[1235], Fresh[1234]}), .c ({new_AGEMA_signal_6518, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M56_U1 ( .a ({new_AGEMA_signal_6196, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_15464, new_AGEMA_signal_15461}), .clk (clk), .r ({Fresh[1237], Fresh[1236]}), .c ({new_AGEMA_signal_6281, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M57_U1 ( .a ({new_AGEMA_signal_6195, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_15470, new_AGEMA_signal_15467}), .clk (clk), .r ({Fresh[1239], Fresh[1238]}), .c ({new_AGEMA_signal_6282, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M57}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M58_U1 ( .a ({new_AGEMA_signal_6275, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_15476, new_AGEMA_signal_15473}), .clk (clk), .r ({Fresh[1241], Fresh[1240]}), .c ({new_AGEMA_signal_6519, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M59_U1 ( .a ({new_AGEMA_signal_6194, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_15482, new_AGEMA_signal_15479}), .clk (clk), .r ({Fresh[1243], Fresh[1242]}), .c ({new_AGEMA_signal_6283, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M59}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M60_U1 ( .a ({new_AGEMA_signal_6193, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_15488, new_AGEMA_signal_15485}), .clk (clk), .r ({Fresh[1245], Fresh[1244]}), .c ({new_AGEMA_signal_6284, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M60}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M61_U1 ( .a ({new_AGEMA_signal_6274, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_15494, new_AGEMA_signal_15491}), .clk (clk), .r ({Fresh[1247], Fresh[1246]}), .c ({new_AGEMA_signal_6520, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M62_U1 ( .a ({new_AGEMA_signal_6513, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_15500, new_AGEMA_signal_15497}), .clk (clk), .r ({Fresh[1249], Fresh[1248]}), .c ({new_AGEMA_signal_6754, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M63_U1 ( .a ({new_AGEMA_signal_6273, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_15506, new_AGEMA_signal_15503}), .clk (clk), .r ({Fresh[1251], Fresh[1250]}), .c ({new_AGEMA_signal_6521, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M63}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L0_U1 ( .a ({new_AGEMA_signal_6520, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61}), .b ({new_AGEMA_signal_6754, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62}), .c ({new_AGEMA_signal_6953, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L1_U1 ( .a ({new_AGEMA_signal_6279, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_6281, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56}), .c ({new_AGEMA_signal_6522, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L2_U1 ( .a ({new_AGEMA_signal_6514, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_6278, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48}), .c ({new_AGEMA_signal_6755, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L3_U1 ( .a ({new_AGEMA_signal_6277, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M47}), .b ({new_AGEMA_signal_6518, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55}), .c ({new_AGEMA_signal_6756, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L4_U1 ( .a ({new_AGEMA_signal_6517, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M54}), .b ({new_AGEMA_signal_6519, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58}), .c ({new_AGEMA_signal_6757, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L5_U1 ( .a ({new_AGEMA_signal_6515, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M49}), .b ({new_AGEMA_signal_6520, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_6758, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L6_U1 ( .a ({new_AGEMA_signal_6754, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62}), .b ({new_AGEMA_signal_6758, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L5}), .c ({new_AGEMA_signal_6954, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L7_U1 ( .a ({new_AGEMA_signal_6514, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_6756, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3}), .c ({new_AGEMA_signal_6955, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L8_U1 ( .a ({new_AGEMA_signal_6280, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51}), .b ({new_AGEMA_signal_6283, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M59}), .c ({new_AGEMA_signal_6523, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L9_U1 ( .a ({new_AGEMA_signal_6516, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_6753, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53}), .c ({new_AGEMA_signal_6956, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L10_U1 ( .a ({new_AGEMA_signal_6753, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53}), .b ({new_AGEMA_signal_6757, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_6957, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L11_U1 ( .a ({new_AGEMA_signal_6284, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M60}), .b ({new_AGEMA_signal_6755, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_6958, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L12_U1 ( .a ({new_AGEMA_signal_6278, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48}), .b ({new_AGEMA_signal_6280, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51}), .c ({new_AGEMA_signal_6524, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L13_U1 ( .a ({new_AGEMA_signal_6279, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_6953, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_7133, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L14_U1 ( .a ({new_AGEMA_signal_6516, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_6520, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_6759, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L15_U1 ( .a ({new_AGEMA_signal_6518, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55}), .b ({new_AGEMA_signal_6522, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_6760, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L16_U1 ( .a ({new_AGEMA_signal_6281, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56}), .b ({new_AGEMA_signal_6953, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_7134, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L17_U1 ( .a ({new_AGEMA_signal_6282, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M57}), .b ({new_AGEMA_signal_6522, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_6761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L18_U1 ( .a ({new_AGEMA_signal_6519, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58}), .b ({new_AGEMA_signal_6523, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8}), .c ({new_AGEMA_signal_6762, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L19_U1 ( .a ({new_AGEMA_signal_6521, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M63}), .b ({new_AGEMA_signal_6757, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_6959, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L20_U1 ( .a ({new_AGEMA_signal_6953, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0}), .b ({new_AGEMA_signal_6522, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_7135, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L21_U1 ( .a ({new_AGEMA_signal_6522, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1}), .b ({new_AGEMA_signal_6955, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7}), .c ({new_AGEMA_signal_7136, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L22_U1 ( .a ({new_AGEMA_signal_6756, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3}), .b ({new_AGEMA_signal_6524, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L12}), .c ({new_AGEMA_signal_6960, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L23_U1 ( .a ({new_AGEMA_signal_6762, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L18}), .b ({new_AGEMA_signal_6755, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_6961, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L24_U1 ( .a ({new_AGEMA_signal_6760, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L15}), .b ({new_AGEMA_signal_6956, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_7137, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L25_U1 ( .a ({new_AGEMA_signal_6954, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_6957, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_7138, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L26_U1 ( .a ({new_AGEMA_signal_6955, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7}), .b ({new_AGEMA_signal_6956, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_7139, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L27_U1 ( .a ({new_AGEMA_signal_6523, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8}), .b ({new_AGEMA_signal_6957, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_7140, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L28_U1 ( .a ({new_AGEMA_signal_6958, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_6759, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L14}), .c ({new_AGEMA_signal_7141, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L28}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L29_U1 ( .a ({new_AGEMA_signal_6958, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_6761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L17}), .c ({new_AGEMA_signal_7142, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L29}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S0_U1 ( .a ({new_AGEMA_signal_6954, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_7137, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L24}), .c ({new_AGEMA_signal_7357, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__7_}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S1_U1 ( .a ({new_AGEMA_signal_7134, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L16}), .b ({new_AGEMA_signal_7139, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L26}), .c ({new_AGEMA_signal_7358, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__6_}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S2_U1 ( .a ({new_AGEMA_signal_6959, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L19}), .b ({new_AGEMA_signal_7141, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L28}), .c ({new_AGEMA_signal_7359, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__5_}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S3_U1 ( .a ({new_AGEMA_signal_6954, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_7136, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L21}), .c ({new_AGEMA_signal_7360, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__4_}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S4_U1 ( .a ({new_AGEMA_signal_7135, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L20}), .b ({new_AGEMA_signal_6960, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L22}), .c ({new_AGEMA_signal_7361, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__3_}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S5_U1 ( .a ({new_AGEMA_signal_7138, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L25}), .b ({new_AGEMA_signal_7142, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L29}), .c ({new_AGEMA_signal_7362, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__2_}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S6_U1 ( .a ({new_AGEMA_signal_7133, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L13}), .b ({new_AGEMA_signal_7140, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L27}), .c ({new_AGEMA_signal_7363, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__1_}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S7_U1 ( .a ({new_AGEMA_signal_6954, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_6961, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L23}), .c ({new_AGEMA_signal_7143, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__0_}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M46_U1 ( .a ({new_AGEMA_signal_6288, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_15512, new_AGEMA_signal_15509}), .clk (clk), .r ({Fresh[1253], Fresh[1252]}), .c ({new_AGEMA_signal_6526, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M47_U1 ( .a ({new_AGEMA_signal_6200, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_15518, new_AGEMA_signal_15515}), .clk (clk), .r ({Fresh[1255], Fresh[1254]}), .c ({new_AGEMA_signal_6289, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M47}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M48_U1 ( .a ({new_AGEMA_signal_6199, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_14363, new_AGEMA_signal_14359}), .clk (clk), .r ({Fresh[1257], Fresh[1256]}), .c ({new_AGEMA_signal_6290, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M49_U1 ( .a ({new_AGEMA_signal_6287, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_15524, new_AGEMA_signal_15521}), .clk (clk), .r ({Fresh[1259], Fresh[1258]}), .c ({new_AGEMA_signal_6527, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M49}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M50_U1 ( .a ({new_AGEMA_signal_6198, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_15530, new_AGEMA_signal_15527}), .clk (clk), .r ({Fresh[1261], Fresh[1260]}), .c ({new_AGEMA_signal_6291, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M51_U1 ( .a ({new_AGEMA_signal_6197, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_15536, new_AGEMA_signal_15533}), .clk (clk), .r ({Fresh[1263], Fresh[1262]}), .c ({new_AGEMA_signal_6292, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M52_U1 ( .a ({new_AGEMA_signal_6286, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_15542, new_AGEMA_signal_15539}), .clk (clk), .r ({Fresh[1265], Fresh[1264]}), .c ({new_AGEMA_signal_6528, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M53_U1 ( .a ({new_AGEMA_signal_6525, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_15548, new_AGEMA_signal_15545}), .clk (clk), .r ({Fresh[1267], Fresh[1266]}), .c ({new_AGEMA_signal_6763, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M54_U1 ( .a ({new_AGEMA_signal_6285, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_15554, new_AGEMA_signal_15551}), .clk (clk), .r ({Fresh[1269], Fresh[1268]}), .c ({new_AGEMA_signal_6529, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M54}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M55_U1 ( .a ({new_AGEMA_signal_6288, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_15560, new_AGEMA_signal_15557}), .clk (clk), .r ({Fresh[1271], Fresh[1270]}), .c ({new_AGEMA_signal_6530, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M56_U1 ( .a ({new_AGEMA_signal_6200, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_15566, new_AGEMA_signal_15563}), .clk (clk), .r ({Fresh[1273], Fresh[1272]}), .c ({new_AGEMA_signal_6293, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M57_U1 ( .a ({new_AGEMA_signal_6199, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_15572, new_AGEMA_signal_15569}), .clk (clk), .r ({Fresh[1275], Fresh[1274]}), .c ({new_AGEMA_signal_6294, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M57}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M58_U1 ( .a ({new_AGEMA_signal_6287, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_15578, new_AGEMA_signal_15575}), .clk (clk), .r ({Fresh[1277], Fresh[1276]}), .c ({new_AGEMA_signal_6531, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M59_U1 ( .a ({new_AGEMA_signal_6198, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_15584, new_AGEMA_signal_15581}), .clk (clk), .r ({Fresh[1279], Fresh[1278]}), .c ({new_AGEMA_signal_6295, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M59}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M60_U1 ( .a ({new_AGEMA_signal_6197, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_15590, new_AGEMA_signal_15587}), .clk (clk), .r ({Fresh[1281], Fresh[1280]}), .c ({new_AGEMA_signal_6296, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M60}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M61_U1 ( .a ({new_AGEMA_signal_6286, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_15596, new_AGEMA_signal_15593}), .clk (clk), .r ({Fresh[1283], Fresh[1282]}), .c ({new_AGEMA_signal_6532, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M62_U1 ( .a ({new_AGEMA_signal_6525, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_15602, new_AGEMA_signal_15599}), .clk (clk), .r ({Fresh[1285], Fresh[1284]}), .c ({new_AGEMA_signal_6764, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M63_U1 ( .a ({new_AGEMA_signal_6285, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_15608, new_AGEMA_signal_15605}), .clk (clk), .r ({Fresh[1287], Fresh[1286]}), .c ({new_AGEMA_signal_6533, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M63}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L0_U1 ( .a ({new_AGEMA_signal_6532, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61}), .b ({new_AGEMA_signal_6764, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62}), .c ({new_AGEMA_signal_6962, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L1_U1 ( .a ({new_AGEMA_signal_6291, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_6293, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56}), .c ({new_AGEMA_signal_6534, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L2_U1 ( .a ({new_AGEMA_signal_6526, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_6290, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48}), .c ({new_AGEMA_signal_6765, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L3_U1 ( .a ({new_AGEMA_signal_6289, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M47}), .b ({new_AGEMA_signal_6530, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55}), .c ({new_AGEMA_signal_6766, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L4_U1 ( .a ({new_AGEMA_signal_6529, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M54}), .b ({new_AGEMA_signal_6531, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58}), .c ({new_AGEMA_signal_6767, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L5_U1 ( .a ({new_AGEMA_signal_6527, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M49}), .b ({new_AGEMA_signal_6532, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_6768, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L6_U1 ( .a ({new_AGEMA_signal_6764, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62}), .b ({new_AGEMA_signal_6768, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L5}), .c ({new_AGEMA_signal_6963, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L7_U1 ( .a ({new_AGEMA_signal_6526, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_6766, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3}), .c ({new_AGEMA_signal_6964, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L8_U1 ( .a ({new_AGEMA_signal_6292, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51}), .b ({new_AGEMA_signal_6295, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M59}), .c ({new_AGEMA_signal_6535, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L9_U1 ( .a ({new_AGEMA_signal_6528, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_6763, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53}), .c ({new_AGEMA_signal_6965, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L10_U1 ( .a ({new_AGEMA_signal_6763, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53}), .b ({new_AGEMA_signal_6767, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_6966, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L11_U1 ( .a ({new_AGEMA_signal_6296, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M60}), .b ({new_AGEMA_signal_6765, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_6967, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L12_U1 ( .a ({new_AGEMA_signal_6290, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48}), .b ({new_AGEMA_signal_6292, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51}), .c ({new_AGEMA_signal_6536, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L13_U1 ( .a ({new_AGEMA_signal_6291, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_6962, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_7144, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L14_U1 ( .a ({new_AGEMA_signal_6528, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_6532, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_6769, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L15_U1 ( .a ({new_AGEMA_signal_6530, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55}), .b ({new_AGEMA_signal_6534, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_6770, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L16_U1 ( .a ({new_AGEMA_signal_6293, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56}), .b ({new_AGEMA_signal_6962, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_7145, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L17_U1 ( .a ({new_AGEMA_signal_6294, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M57}), .b ({new_AGEMA_signal_6534, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_6771, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L18_U1 ( .a ({new_AGEMA_signal_6531, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58}), .b ({new_AGEMA_signal_6535, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8}), .c ({new_AGEMA_signal_6772, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L19_U1 ( .a ({new_AGEMA_signal_6533, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M63}), .b ({new_AGEMA_signal_6767, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_6968, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L20_U1 ( .a ({new_AGEMA_signal_6962, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0}), .b ({new_AGEMA_signal_6534, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_7146, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L21_U1 ( .a ({new_AGEMA_signal_6534, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1}), .b ({new_AGEMA_signal_6964, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7}), .c ({new_AGEMA_signal_7147, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L22_U1 ( .a ({new_AGEMA_signal_6766, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3}), .b ({new_AGEMA_signal_6536, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L12}), .c ({new_AGEMA_signal_6969, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L23_U1 ( .a ({new_AGEMA_signal_6772, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L18}), .b ({new_AGEMA_signal_6765, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_6970, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L24_U1 ( .a ({new_AGEMA_signal_6770, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L15}), .b ({new_AGEMA_signal_6965, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_7148, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L25_U1 ( .a ({new_AGEMA_signal_6963, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_6966, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_7149, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L26_U1 ( .a ({new_AGEMA_signal_6964, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7}), .b ({new_AGEMA_signal_6965, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_7150, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L27_U1 ( .a ({new_AGEMA_signal_6535, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8}), .b ({new_AGEMA_signal_6966, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_7151, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L28_U1 ( .a ({new_AGEMA_signal_6967, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_6769, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L14}), .c ({new_AGEMA_signal_7152, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L28}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L29_U1 ( .a ({new_AGEMA_signal_6967, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_6771, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L17}), .c ({new_AGEMA_signal_7153, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L29}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S0_U1 ( .a ({new_AGEMA_signal_6963, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_7148, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L24}), .c ({new_AGEMA_signal_7364, KeyExpansionIns_tmp[23]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S1_U1 ( .a ({new_AGEMA_signal_7145, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L16}), .b ({new_AGEMA_signal_7150, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L26}), .c ({new_AGEMA_signal_7365, KeyExpansionIns_tmp[22]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S2_U1 ( .a ({new_AGEMA_signal_6968, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L19}), .b ({new_AGEMA_signal_7152, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L28}), .c ({new_AGEMA_signal_7366, KeyExpansionIns_tmp[21]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S3_U1 ( .a ({new_AGEMA_signal_6963, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_7147, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L21}), .c ({new_AGEMA_signal_7367, KeyExpansionIns_tmp[20]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S4_U1 ( .a ({new_AGEMA_signal_7146, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L20}), .b ({new_AGEMA_signal_6969, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L22}), .c ({new_AGEMA_signal_7368, KeyExpansionIns_tmp[19]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S5_U1 ( .a ({new_AGEMA_signal_7149, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L25}), .b ({new_AGEMA_signal_7153, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L29}), .c ({new_AGEMA_signal_7369, KeyExpansionIns_tmp[18]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S6_U1 ( .a ({new_AGEMA_signal_7144, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L13}), .b ({new_AGEMA_signal_7151, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L27}), .c ({new_AGEMA_signal_7370, KeyExpansionIns_tmp[17]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S7_U1 ( .a ({new_AGEMA_signal_6963, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_6970, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L23}), .c ({new_AGEMA_signal_7154, KeyExpansionIns_tmp[16]}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M46_U1 ( .a ({new_AGEMA_signal_6300, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_15614, new_AGEMA_signal_15611}), .clk (clk), .r ({Fresh[1289], Fresh[1288]}), .c ({new_AGEMA_signal_6538, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M47_U1 ( .a ({new_AGEMA_signal_6204, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_15620, new_AGEMA_signal_15617}), .clk (clk), .r ({Fresh[1291], Fresh[1290]}), .c ({new_AGEMA_signal_6301, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M47}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M48_U1 ( .a ({new_AGEMA_signal_6203, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_15347, new_AGEMA_signal_15343}), .clk (clk), .r ({Fresh[1293], Fresh[1292]}), .c ({new_AGEMA_signal_6302, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M49_U1 ( .a ({new_AGEMA_signal_6299, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_15626, new_AGEMA_signal_15623}), .clk (clk), .r ({Fresh[1295], Fresh[1294]}), .c ({new_AGEMA_signal_6539, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M49}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M50_U1 ( .a ({new_AGEMA_signal_6202, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_15632, new_AGEMA_signal_15629}), .clk (clk), .r ({Fresh[1297], Fresh[1296]}), .c ({new_AGEMA_signal_6303, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M51_U1 ( .a ({new_AGEMA_signal_6201, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_15638, new_AGEMA_signal_15635}), .clk (clk), .r ({Fresh[1299], Fresh[1298]}), .c ({new_AGEMA_signal_6304, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M52_U1 ( .a ({new_AGEMA_signal_6298, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_15644, new_AGEMA_signal_15641}), .clk (clk), .r ({Fresh[1301], Fresh[1300]}), .c ({new_AGEMA_signal_6540, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M53_U1 ( .a ({new_AGEMA_signal_6537, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_15650, new_AGEMA_signal_15647}), .clk (clk), .r ({Fresh[1303], Fresh[1302]}), .c ({new_AGEMA_signal_6773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M54_U1 ( .a ({new_AGEMA_signal_6297, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_15656, new_AGEMA_signal_15653}), .clk (clk), .r ({Fresh[1305], Fresh[1304]}), .c ({new_AGEMA_signal_6541, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M54}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M55_U1 ( .a ({new_AGEMA_signal_6300, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_15662, new_AGEMA_signal_15659}), .clk (clk), .r ({Fresh[1307], Fresh[1306]}), .c ({new_AGEMA_signal_6542, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M56_U1 ( .a ({new_AGEMA_signal_6204, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_15668, new_AGEMA_signal_15665}), .clk (clk), .r ({Fresh[1309], Fresh[1308]}), .c ({new_AGEMA_signal_6305, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M57_U1 ( .a ({new_AGEMA_signal_6203, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_15674, new_AGEMA_signal_15671}), .clk (clk), .r ({Fresh[1311], Fresh[1310]}), .c ({new_AGEMA_signal_6306, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M57}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M58_U1 ( .a ({new_AGEMA_signal_6299, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_15680, new_AGEMA_signal_15677}), .clk (clk), .r ({Fresh[1313], Fresh[1312]}), .c ({new_AGEMA_signal_6543, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M59_U1 ( .a ({new_AGEMA_signal_6202, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_15686, new_AGEMA_signal_15683}), .clk (clk), .r ({Fresh[1315], Fresh[1314]}), .c ({new_AGEMA_signal_6307, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M59}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M60_U1 ( .a ({new_AGEMA_signal_6201, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_15692, new_AGEMA_signal_15689}), .clk (clk), .r ({Fresh[1317], Fresh[1316]}), .c ({new_AGEMA_signal_6308, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M60}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M61_U1 ( .a ({new_AGEMA_signal_6298, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_15698, new_AGEMA_signal_15695}), .clk (clk), .r ({Fresh[1319], Fresh[1318]}), .c ({new_AGEMA_signal_6544, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M62_U1 ( .a ({new_AGEMA_signal_6537, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_15704, new_AGEMA_signal_15701}), .clk (clk), .r ({Fresh[1321], Fresh[1320]}), .c ({new_AGEMA_signal_6774, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M63_U1 ( .a ({new_AGEMA_signal_6297, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_15710, new_AGEMA_signal_15707}), .clk (clk), .r ({Fresh[1323], Fresh[1322]}), .c ({new_AGEMA_signal_6545, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M63}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L0_U1 ( .a ({new_AGEMA_signal_6544, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61}), .b ({new_AGEMA_signal_6774, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62}), .c ({new_AGEMA_signal_6971, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L1_U1 ( .a ({new_AGEMA_signal_6303, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_6305, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56}), .c ({new_AGEMA_signal_6546, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L2_U1 ( .a ({new_AGEMA_signal_6538, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_6302, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48}), .c ({new_AGEMA_signal_6775, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L3_U1 ( .a ({new_AGEMA_signal_6301, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M47}), .b ({new_AGEMA_signal_6542, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55}), .c ({new_AGEMA_signal_6776, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L4_U1 ( .a ({new_AGEMA_signal_6541, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M54}), .b ({new_AGEMA_signal_6543, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58}), .c ({new_AGEMA_signal_6777, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L5_U1 ( .a ({new_AGEMA_signal_6539, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M49}), .b ({new_AGEMA_signal_6544, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_6778, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L6_U1 ( .a ({new_AGEMA_signal_6774, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62}), .b ({new_AGEMA_signal_6778, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L5}), .c ({new_AGEMA_signal_6972, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L7_U1 ( .a ({new_AGEMA_signal_6538, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_6776, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3}), .c ({new_AGEMA_signal_6973, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L8_U1 ( .a ({new_AGEMA_signal_6304, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51}), .b ({new_AGEMA_signal_6307, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M59}), .c ({new_AGEMA_signal_6547, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L9_U1 ( .a ({new_AGEMA_signal_6540, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_6773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53}), .c ({new_AGEMA_signal_6974, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L10_U1 ( .a ({new_AGEMA_signal_6773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53}), .b ({new_AGEMA_signal_6777, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_6975, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L11_U1 ( .a ({new_AGEMA_signal_6308, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M60}), .b ({new_AGEMA_signal_6775, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_6976, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L12_U1 ( .a ({new_AGEMA_signal_6302, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48}), .b ({new_AGEMA_signal_6304, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51}), .c ({new_AGEMA_signal_6548, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L13_U1 ( .a ({new_AGEMA_signal_6303, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_6971, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_7155, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L14_U1 ( .a ({new_AGEMA_signal_6540, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_6544, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_6779, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L15_U1 ( .a ({new_AGEMA_signal_6542, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55}), .b ({new_AGEMA_signal_6546, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_6780, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L16_U1 ( .a ({new_AGEMA_signal_6305, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56}), .b ({new_AGEMA_signal_6971, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_7156, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L17_U1 ( .a ({new_AGEMA_signal_6306, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M57}), .b ({new_AGEMA_signal_6546, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_6781, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L18_U1 ( .a ({new_AGEMA_signal_6543, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58}), .b ({new_AGEMA_signal_6547, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8}), .c ({new_AGEMA_signal_6782, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L19_U1 ( .a ({new_AGEMA_signal_6545, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M63}), .b ({new_AGEMA_signal_6777, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_6977, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L20_U1 ( .a ({new_AGEMA_signal_6971, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0}), .b ({new_AGEMA_signal_6546, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_7157, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L21_U1 ( .a ({new_AGEMA_signal_6546, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1}), .b ({new_AGEMA_signal_6973, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7}), .c ({new_AGEMA_signal_7158, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L22_U1 ( .a ({new_AGEMA_signal_6776, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3}), .b ({new_AGEMA_signal_6548, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L12}), .c ({new_AGEMA_signal_6978, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L23_U1 ( .a ({new_AGEMA_signal_6782, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L18}), .b ({new_AGEMA_signal_6775, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_6979, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L24_U1 ( .a ({new_AGEMA_signal_6780, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L15}), .b ({new_AGEMA_signal_6974, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_7159, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L25_U1 ( .a ({new_AGEMA_signal_6972, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_6975, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_7160, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L26_U1 ( .a ({new_AGEMA_signal_6973, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7}), .b ({new_AGEMA_signal_6974, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_7161, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L27_U1 ( .a ({new_AGEMA_signal_6547, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8}), .b ({new_AGEMA_signal_6975, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_7162, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L28_U1 ( .a ({new_AGEMA_signal_6976, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_6779, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L14}), .c ({new_AGEMA_signal_7163, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L28}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L29_U1 ( .a ({new_AGEMA_signal_6976, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_6781, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L17}), .c ({new_AGEMA_signal_7164, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L29}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S0_U1 ( .a ({new_AGEMA_signal_6972, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_7159, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L24}), .c ({new_AGEMA_signal_7371, KeyExpansionIns_tmp[15]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S1_U1 ( .a ({new_AGEMA_signal_7156, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L16}), .b ({new_AGEMA_signal_7161, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L26}), .c ({new_AGEMA_signal_7372, KeyExpansionIns_tmp[14]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S2_U1 ( .a ({new_AGEMA_signal_6977, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L19}), .b ({new_AGEMA_signal_7163, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L28}), .c ({new_AGEMA_signal_7373, KeyExpansionIns_tmp[13]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S3_U1 ( .a ({new_AGEMA_signal_6972, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_7158, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L21}), .c ({new_AGEMA_signal_7374, KeyExpansionIns_tmp[12]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S4_U1 ( .a ({new_AGEMA_signal_7157, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L20}), .b ({new_AGEMA_signal_6978, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L22}), .c ({new_AGEMA_signal_7375, KeyExpansionIns_tmp[11]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S5_U1 ( .a ({new_AGEMA_signal_7160, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L25}), .b ({new_AGEMA_signal_7164, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L29}), .c ({new_AGEMA_signal_7376, KeyExpansionIns_tmp[10]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S6_U1 ( .a ({new_AGEMA_signal_7155, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L13}), .b ({new_AGEMA_signal_7162, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L27}), .c ({new_AGEMA_signal_7377, KeyExpansionIns_tmp[9]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S7_U1 ( .a ({new_AGEMA_signal_6972, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_6979, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L23}), .c ({new_AGEMA_signal_7165, KeyExpansionIns_tmp[8]}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M46_U1 ( .a ({new_AGEMA_signal_6312, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_15716, new_AGEMA_signal_15713}), .clk (clk), .r ({Fresh[1325], Fresh[1324]}), .c ({new_AGEMA_signal_6550, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M47_U1 ( .a ({new_AGEMA_signal_6208, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_15722, new_AGEMA_signal_15719}), .clk (clk), .r ({Fresh[1327], Fresh[1326]}), .c ({new_AGEMA_signal_6313, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M47}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M48_U1 ( .a ({new_AGEMA_signal_6207, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_14731, new_AGEMA_signal_14727}), .clk (clk), .r ({Fresh[1329], Fresh[1328]}), .c ({new_AGEMA_signal_6314, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M49_U1 ( .a ({new_AGEMA_signal_6311, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_15728, new_AGEMA_signal_15725}), .clk (clk), .r ({Fresh[1331], Fresh[1330]}), .c ({new_AGEMA_signal_6551, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M49}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M50_U1 ( .a ({new_AGEMA_signal_6206, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_15734, new_AGEMA_signal_15731}), .clk (clk), .r ({Fresh[1333], Fresh[1332]}), .c ({new_AGEMA_signal_6315, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M51_U1 ( .a ({new_AGEMA_signal_6205, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_15740, new_AGEMA_signal_15737}), .clk (clk), .r ({Fresh[1335], Fresh[1334]}), .c ({new_AGEMA_signal_6316, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M52_U1 ( .a ({new_AGEMA_signal_6310, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_15746, new_AGEMA_signal_15743}), .clk (clk), .r ({Fresh[1337], Fresh[1336]}), .c ({new_AGEMA_signal_6552, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M53_U1 ( .a ({new_AGEMA_signal_6549, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_15752, new_AGEMA_signal_15749}), .clk (clk), .r ({Fresh[1339], Fresh[1338]}), .c ({new_AGEMA_signal_6783, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M54_U1 ( .a ({new_AGEMA_signal_6309, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_15758, new_AGEMA_signal_15755}), .clk (clk), .r ({Fresh[1341], Fresh[1340]}), .c ({new_AGEMA_signal_6553, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M54}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M55_U1 ( .a ({new_AGEMA_signal_6312, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_15764, new_AGEMA_signal_15761}), .clk (clk), .r ({Fresh[1343], Fresh[1342]}), .c ({new_AGEMA_signal_6554, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M56_U1 ( .a ({new_AGEMA_signal_6208, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_15770, new_AGEMA_signal_15767}), .clk (clk), .r ({Fresh[1345], Fresh[1344]}), .c ({new_AGEMA_signal_6317, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M57_U1 ( .a ({new_AGEMA_signal_6207, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_15776, new_AGEMA_signal_15773}), .clk (clk), .r ({Fresh[1347], Fresh[1346]}), .c ({new_AGEMA_signal_6318, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M57}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M58_U1 ( .a ({new_AGEMA_signal_6311, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_15782, new_AGEMA_signal_15779}), .clk (clk), .r ({Fresh[1349], Fresh[1348]}), .c ({new_AGEMA_signal_6555, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M59_U1 ( .a ({new_AGEMA_signal_6206, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_15788, new_AGEMA_signal_15785}), .clk (clk), .r ({Fresh[1351], Fresh[1350]}), .c ({new_AGEMA_signal_6319, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M59}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M60_U1 ( .a ({new_AGEMA_signal_6205, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_15794, new_AGEMA_signal_15791}), .clk (clk), .r ({Fresh[1353], Fresh[1352]}), .c ({new_AGEMA_signal_6320, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M60}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M61_U1 ( .a ({new_AGEMA_signal_6310, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_15800, new_AGEMA_signal_15797}), .clk (clk), .r ({Fresh[1355], Fresh[1354]}), .c ({new_AGEMA_signal_6556, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M62_U1 ( .a ({new_AGEMA_signal_6549, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_15806, new_AGEMA_signal_15803}), .clk (clk), .r ({Fresh[1357], Fresh[1356]}), .c ({new_AGEMA_signal_6784, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M63_U1 ( .a ({new_AGEMA_signal_6309, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_15812, new_AGEMA_signal_15809}), .clk (clk), .r ({Fresh[1359], Fresh[1358]}), .c ({new_AGEMA_signal_6557, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M63}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L0_U1 ( .a ({new_AGEMA_signal_6556, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61}), .b ({new_AGEMA_signal_6784, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62}), .c ({new_AGEMA_signal_6980, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L1_U1 ( .a ({new_AGEMA_signal_6315, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_6317, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56}), .c ({new_AGEMA_signal_6558, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L2_U1 ( .a ({new_AGEMA_signal_6550, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_6314, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48}), .c ({new_AGEMA_signal_6785, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L3_U1 ( .a ({new_AGEMA_signal_6313, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M47}), .b ({new_AGEMA_signal_6554, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55}), .c ({new_AGEMA_signal_6786, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L4_U1 ( .a ({new_AGEMA_signal_6553, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M54}), .b ({new_AGEMA_signal_6555, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58}), .c ({new_AGEMA_signal_6787, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L5_U1 ( .a ({new_AGEMA_signal_6551, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M49}), .b ({new_AGEMA_signal_6556, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_6788, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L6_U1 ( .a ({new_AGEMA_signal_6784, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62}), .b ({new_AGEMA_signal_6788, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L5}), .c ({new_AGEMA_signal_6981, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L7_U1 ( .a ({new_AGEMA_signal_6550, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_6786, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3}), .c ({new_AGEMA_signal_6982, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L8_U1 ( .a ({new_AGEMA_signal_6316, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51}), .b ({new_AGEMA_signal_6319, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M59}), .c ({new_AGEMA_signal_6559, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L9_U1 ( .a ({new_AGEMA_signal_6552, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_6783, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53}), .c ({new_AGEMA_signal_6983, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L10_U1 ( .a ({new_AGEMA_signal_6783, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53}), .b ({new_AGEMA_signal_6787, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_6984, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L11_U1 ( .a ({new_AGEMA_signal_6320, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M60}), .b ({new_AGEMA_signal_6785, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_6985, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L12_U1 ( .a ({new_AGEMA_signal_6314, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48}), .b ({new_AGEMA_signal_6316, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51}), .c ({new_AGEMA_signal_6560, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L13_U1 ( .a ({new_AGEMA_signal_6315, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_6980, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_7166, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L14_U1 ( .a ({new_AGEMA_signal_6552, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_6556, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_6789, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L15_U1 ( .a ({new_AGEMA_signal_6554, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55}), .b ({new_AGEMA_signal_6558, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_6790, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L16_U1 ( .a ({new_AGEMA_signal_6317, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56}), .b ({new_AGEMA_signal_6980, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_7167, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L17_U1 ( .a ({new_AGEMA_signal_6318, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M57}), .b ({new_AGEMA_signal_6558, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_6791, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L18_U1 ( .a ({new_AGEMA_signal_6555, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58}), .b ({new_AGEMA_signal_6559, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8}), .c ({new_AGEMA_signal_6792, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L19_U1 ( .a ({new_AGEMA_signal_6557, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M63}), .b ({new_AGEMA_signal_6787, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_6986, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L20_U1 ( .a ({new_AGEMA_signal_6980, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0}), .b ({new_AGEMA_signal_6558, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_7168, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L21_U1 ( .a ({new_AGEMA_signal_6558, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1}), .b ({new_AGEMA_signal_6982, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7}), .c ({new_AGEMA_signal_7169, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L22_U1 ( .a ({new_AGEMA_signal_6786, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3}), .b ({new_AGEMA_signal_6560, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L12}), .c ({new_AGEMA_signal_6987, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L23_U1 ( .a ({new_AGEMA_signal_6792, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L18}), .b ({new_AGEMA_signal_6785, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_6988, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L24_U1 ( .a ({new_AGEMA_signal_6790, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L15}), .b ({new_AGEMA_signal_6983, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_7170, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L25_U1 ( .a ({new_AGEMA_signal_6981, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_6984, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_7171, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L26_U1 ( .a ({new_AGEMA_signal_6982, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7}), .b ({new_AGEMA_signal_6983, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_7172, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L27_U1 ( .a ({new_AGEMA_signal_6559, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8}), .b ({new_AGEMA_signal_6984, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_7173, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L28_U1 ( .a ({new_AGEMA_signal_6985, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_6789, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L14}), .c ({new_AGEMA_signal_7174, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L28}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L29_U1 ( .a ({new_AGEMA_signal_6985, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_6791, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L17}), .c ({new_AGEMA_signal_7175, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L29}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S0_U1 ( .a ({new_AGEMA_signal_6981, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_7170, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L24}), .c ({new_AGEMA_signal_7378, KeyExpansionIns_tmp[7]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S1_U1 ( .a ({new_AGEMA_signal_7167, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L16}), .b ({new_AGEMA_signal_7172, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L26}), .c ({new_AGEMA_signal_7379, KeyExpansionIns_tmp[6]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S2_U1 ( .a ({new_AGEMA_signal_6986, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L19}), .b ({new_AGEMA_signal_7174, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L28}), .c ({new_AGEMA_signal_7380, KeyExpansionIns_tmp[5]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S3_U1 ( .a ({new_AGEMA_signal_6981, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_7169, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L21}), .c ({new_AGEMA_signal_7381, KeyExpansionIns_tmp[4]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S4_U1 ( .a ({new_AGEMA_signal_7168, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L20}), .b ({new_AGEMA_signal_6987, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L22}), .c ({new_AGEMA_signal_7382, KeyExpansionIns_tmp[3]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S5_U1 ( .a ({new_AGEMA_signal_7171, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L25}), .b ({new_AGEMA_signal_7175, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L29}), .c ({new_AGEMA_signal_7383, KeyExpansionIns_tmp[2]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S6_U1 ( .a ({new_AGEMA_signal_7166, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L13}), .b ({new_AGEMA_signal_7173, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L27}), .c ({new_AGEMA_signal_7384, KeyExpansionIns_tmp[1]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S7_U1 ( .a ({new_AGEMA_signal_6981, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_6988, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L23}), .c ({new_AGEMA_signal_7176, KeyExpansionIns_tmp[0]}) ) ;
    buf_clk new_AGEMA_reg_buffer_4692 ( .C (clk), .D (new_AGEMA_signal_10543), .Q (new_AGEMA_signal_10544) ) ;
    buf_clk new_AGEMA_reg_buffer_4696 ( .C (clk), .D (new_AGEMA_signal_10547), .Q (new_AGEMA_signal_10548) ) ;
    buf_clk new_AGEMA_reg_buffer_4700 ( .C (clk), .D (new_AGEMA_signal_10551), .Q (new_AGEMA_signal_10552) ) ;
    buf_clk new_AGEMA_reg_buffer_4704 ( .C (clk), .D (new_AGEMA_signal_10555), .Q (new_AGEMA_signal_10556) ) ;
    buf_clk new_AGEMA_reg_buffer_4708 ( .C (clk), .D (new_AGEMA_signal_10559), .Q (new_AGEMA_signal_10560) ) ;
    buf_clk new_AGEMA_reg_buffer_4712 ( .C (clk), .D (new_AGEMA_signal_10563), .Q (new_AGEMA_signal_10564) ) ;
    buf_clk new_AGEMA_reg_buffer_4716 ( .C (clk), .D (new_AGEMA_signal_10567), .Q (new_AGEMA_signal_10568) ) ;
    buf_clk new_AGEMA_reg_buffer_4720 ( .C (clk), .D (new_AGEMA_signal_10571), .Q (new_AGEMA_signal_10572) ) ;
    buf_clk new_AGEMA_reg_buffer_4724 ( .C (clk), .D (new_AGEMA_signal_10575), .Q (new_AGEMA_signal_10576) ) ;
    buf_clk new_AGEMA_reg_buffer_4728 ( .C (clk), .D (new_AGEMA_signal_10579), .Q (new_AGEMA_signal_10580) ) ;
    buf_clk new_AGEMA_reg_buffer_4732 ( .C (clk), .D (new_AGEMA_signal_10583), .Q (new_AGEMA_signal_10584) ) ;
    buf_clk new_AGEMA_reg_buffer_4736 ( .C (clk), .D (new_AGEMA_signal_10587), .Q (new_AGEMA_signal_10588) ) ;
    buf_clk new_AGEMA_reg_buffer_4740 ( .C (clk), .D (new_AGEMA_signal_10591), .Q (new_AGEMA_signal_10592) ) ;
    buf_clk new_AGEMA_reg_buffer_4744 ( .C (clk), .D (new_AGEMA_signal_10595), .Q (new_AGEMA_signal_10596) ) ;
    buf_clk new_AGEMA_reg_buffer_4748 ( .C (clk), .D (new_AGEMA_signal_10599), .Q (new_AGEMA_signal_10600) ) ;
    buf_clk new_AGEMA_reg_buffer_4752 ( .C (clk), .D (new_AGEMA_signal_10603), .Q (new_AGEMA_signal_10604) ) ;
    buf_clk new_AGEMA_reg_buffer_4756 ( .C (clk), .D (new_AGEMA_signal_10607), .Q (new_AGEMA_signal_10608) ) ;
    buf_clk new_AGEMA_reg_buffer_4760 ( .C (clk), .D (new_AGEMA_signal_10611), .Q (new_AGEMA_signal_10612) ) ;
    buf_clk new_AGEMA_reg_buffer_4764 ( .C (clk), .D (new_AGEMA_signal_10615), .Q (new_AGEMA_signal_10616) ) ;
    buf_clk new_AGEMA_reg_buffer_4768 ( .C (clk), .D (new_AGEMA_signal_10619), .Q (new_AGEMA_signal_10620) ) ;
    buf_clk new_AGEMA_reg_buffer_4772 ( .C (clk), .D (new_AGEMA_signal_10623), .Q (new_AGEMA_signal_10624) ) ;
    buf_clk new_AGEMA_reg_buffer_4776 ( .C (clk), .D (new_AGEMA_signal_10627), .Q (new_AGEMA_signal_10628) ) ;
    buf_clk new_AGEMA_reg_buffer_4780 ( .C (clk), .D (new_AGEMA_signal_10631), .Q (new_AGEMA_signal_10632) ) ;
    buf_clk new_AGEMA_reg_buffer_4784 ( .C (clk), .D (new_AGEMA_signal_10635), .Q (new_AGEMA_signal_10636) ) ;
    buf_clk new_AGEMA_reg_buffer_4788 ( .C (clk), .D (new_AGEMA_signal_10639), .Q (new_AGEMA_signal_10640) ) ;
    buf_clk new_AGEMA_reg_buffer_4792 ( .C (clk), .D (new_AGEMA_signal_10643), .Q (new_AGEMA_signal_10644) ) ;
    buf_clk new_AGEMA_reg_buffer_4796 ( .C (clk), .D (new_AGEMA_signal_10647), .Q (new_AGEMA_signal_10648) ) ;
    buf_clk new_AGEMA_reg_buffer_4800 ( .C (clk), .D (new_AGEMA_signal_10651), .Q (new_AGEMA_signal_10652) ) ;
    buf_clk new_AGEMA_reg_buffer_4804 ( .C (clk), .D (new_AGEMA_signal_10655), .Q (new_AGEMA_signal_10656) ) ;
    buf_clk new_AGEMA_reg_buffer_4808 ( .C (clk), .D (new_AGEMA_signal_10659), .Q (new_AGEMA_signal_10660) ) ;
    buf_clk new_AGEMA_reg_buffer_4812 ( .C (clk), .D (new_AGEMA_signal_10663), .Q (new_AGEMA_signal_10664) ) ;
    buf_clk new_AGEMA_reg_buffer_4816 ( .C (clk), .D (new_AGEMA_signal_10667), .Q (new_AGEMA_signal_10668) ) ;
    buf_clk new_AGEMA_reg_buffer_4820 ( .C (clk), .D (new_AGEMA_signal_10671), .Q (new_AGEMA_signal_10672) ) ;
    buf_clk new_AGEMA_reg_buffer_4824 ( .C (clk), .D (new_AGEMA_signal_10675), .Q (new_AGEMA_signal_10676) ) ;
    buf_clk new_AGEMA_reg_buffer_4828 ( .C (clk), .D (new_AGEMA_signal_10679), .Q (new_AGEMA_signal_10680) ) ;
    buf_clk new_AGEMA_reg_buffer_4832 ( .C (clk), .D (new_AGEMA_signal_10683), .Q (new_AGEMA_signal_10684) ) ;
    buf_clk new_AGEMA_reg_buffer_4836 ( .C (clk), .D (new_AGEMA_signal_10687), .Q (new_AGEMA_signal_10688) ) ;
    buf_clk new_AGEMA_reg_buffer_4840 ( .C (clk), .D (new_AGEMA_signal_10691), .Q (new_AGEMA_signal_10692) ) ;
    buf_clk new_AGEMA_reg_buffer_4844 ( .C (clk), .D (new_AGEMA_signal_10695), .Q (new_AGEMA_signal_10696) ) ;
    buf_clk new_AGEMA_reg_buffer_4848 ( .C (clk), .D (new_AGEMA_signal_10699), .Q (new_AGEMA_signal_10700) ) ;
    buf_clk new_AGEMA_reg_buffer_4852 ( .C (clk), .D (new_AGEMA_signal_10703), .Q (new_AGEMA_signal_10704) ) ;
    buf_clk new_AGEMA_reg_buffer_4856 ( .C (clk), .D (new_AGEMA_signal_10707), .Q (new_AGEMA_signal_10708) ) ;
    buf_clk new_AGEMA_reg_buffer_4860 ( .C (clk), .D (new_AGEMA_signal_10711), .Q (new_AGEMA_signal_10712) ) ;
    buf_clk new_AGEMA_reg_buffer_4864 ( .C (clk), .D (new_AGEMA_signal_10715), .Q (new_AGEMA_signal_10716) ) ;
    buf_clk new_AGEMA_reg_buffer_4868 ( .C (clk), .D (new_AGEMA_signal_10719), .Q (new_AGEMA_signal_10720) ) ;
    buf_clk new_AGEMA_reg_buffer_4872 ( .C (clk), .D (new_AGEMA_signal_10723), .Q (new_AGEMA_signal_10724) ) ;
    buf_clk new_AGEMA_reg_buffer_4876 ( .C (clk), .D (new_AGEMA_signal_10727), .Q (new_AGEMA_signal_10728) ) ;
    buf_clk new_AGEMA_reg_buffer_4880 ( .C (clk), .D (new_AGEMA_signal_10731), .Q (new_AGEMA_signal_10732) ) ;
    buf_clk new_AGEMA_reg_buffer_4884 ( .C (clk), .D (new_AGEMA_signal_10735), .Q (new_AGEMA_signal_10736) ) ;
    buf_clk new_AGEMA_reg_buffer_4888 ( .C (clk), .D (new_AGEMA_signal_10739), .Q (new_AGEMA_signal_10740) ) ;
    buf_clk new_AGEMA_reg_buffer_4892 ( .C (clk), .D (new_AGEMA_signal_10743), .Q (new_AGEMA_signal_10744) ) ;
    buf_clk new_AGEMA_reg_buffer_4896 ( .C (clk), .D (new_AGEMA_signal_10747), .Q (new_AGEMA_signal_10748) ) ;
    buf_clk new_AGEMA_reg_buffer_4900 ( .C (clk), .D (new_AGEMA_signal_10751), .Q (new_AGEMA_signal_10752) ) ;
    buf_clk new_AGEMA_reg_buffer_4904 ( .C (clk), .D (new_AGEMA_signal_10755), .Q (new_AGEMA_signal_10756) ) ;
    buf_clk new_AGEMA_reg_buffer_4908 ( .C (clk), .D (new_AGEMA_signal_10759), .Q (new_AGEMA_signal_10760) ) ;
    buf_clk new_AGEMA_reg_buffer_4912 ( .C (clk), .D (new_AGEMA_signal_10763), .Q (new_AGEMA_signal_10764) ) ;
    buf_clk new_AGEMA_reg_buffer_4916 ( .C (clk), .D (new_AGEMA_signal_10767), .Q (new_AGEMA_signal_10768) ) ;
    buf_clk new_AGEMA_reg_buffer_4920 ( .C (clk), .D (new_AGEMA_signal_10771), .Q (new_AGEMA_signal_10772) ) ;
    buf_clk new_AGEMA_reg_buffer_4924 ( .C (clk), .D (new_AGEMA_signal_10775), .Q (new_AGEMA_signal_10776) ) ;
    buf_clk new_AGEMA_reg_buffer_4928 ( .C (clk), .D (new_AGEMA_signal_10779), .Q (new_AGEMA_signal_10780) ) ;
    buf_clk new_AGEMA_reg_buffer_4932 ( .C (clk), .D (new_AGEMA_signal_10783), .Q (new_AGEMA_signal_10784) ) ;
    buf_clk new_AGEMA_reg_buffer_4936 ( .C (clk), .D (new_AGEMA_signal_10787), .Q (new_AGEMA_signal_10788) ) ;
    buf_clk new_AGEMA_reg_buffer_4940 ( .C (clk), .D (new_AGEMA_signal_10791), .Q (new_AGEMA_signal_10792) ) ;
    buf_clk new_AGEMA_reg_buffer_4944 ( .C (clk), .D (new_AGEMA_signal_10795), .Q (new_AGEMA_signal_10796) ) ;
    buf_clk new_AGEMA_reg_buffer_4948 ( .C (clk), .D (new_AGEMA_signal_10799), .Q (new_AGEMA_signal_10800) ) ;
    buf_clk new_AGEMA_reg_buffer_4952 ( .C (clk), .D (new_AGEMA_signal_10803), .Q (new_AGEMA_signal_10804) ) ;
    buf_clk new_AGEMA_reg_buffer_4956 ( .C (clk), .D (new_AGEMA_signal_10807), .Q (new_AGEMA_signal_10808) ) ;
    buf_clk new_AGEMA_reg_buffer_4960 ( .C (clk), .D (new_AGEMA_signal_10811), .Q (new_AGEMA_signal_10812) ) ;
    buf_clk new_AGEMA_reg_buffer_4964 ( .C (clk), .D (new_AGEMA_signal_10815), .Q (new_AGEMA_signal_10816) ) ;
    buf_clk new_AGEMA_reg_buffer_4968 ( .C (clk), .D (new_AGEMA_signal_10819), .Q (new_AGEMA_signal_10820) ) ;
    buf_clk new_AGEMA_reg_buffer_4972 ( .C (clk), .D (new_AGEMA_signal_10823), .Q (new_AGEMA_signal_10824) ) ;
    buf_clk new_AGEMA_reg_buffer_4976 ( .C (clk), .D (new_AGEMA_signal_10827), .Q (new_AGEMA_signal_10828) ) ;
    buf_clk new_AGEMA_reg_buffer_4980 ( .C (clk), .D (new_AGEMA_signal_10831), .Q (new_AGEMA_signal_10832) ) ;
    buf_clk new_AGEMA_reg_buffer_4984 ( .C (clk), .D (new_AGEMA_signal_10835), .Q (new_AGEMA_signal_10836) ) ;
    buf_clk new_AGEMA_reg_buffer_4988 ( .C (clk), .D (new_AGEMA_signal_10839), .Q (new_AGEMA_signal_10840) ) ;
    buf_clk new_AGEMA_reg_buffer_4992 ( .C (clk), .D (new_AGEMA_signal_10843), .Q (new_AGEMA_signal_10844) ) ;
    buf_clk new_AGEMA_reg_buffer_4996 ( .C (clk), .D (new_AGEMA_signal_10847), .Q (new_AGEMA_signal_10848) ) ;
    buf_clk new_AGEMA_reg_buffer_5000 ( .C (clk), .D (new_AGEMA_signal_10851), .Q (new_AGEMA_signal_10852) ) ;
    buf_clk new_AGEMA_reg_buffer_5004 ( .C (clk), .D (new_AGEMA_signal_10855), .Q (new_AGEMA_signal_10856) ) ;
    buf_clk new_AGEMA_reg_buffer_5008 ( .C (clk), .D (new_AGEMA_signal_10859), .Q (new_AGEMA_signal_10860) ) ;
    buf_clk new_AGEMA_reg_buffer_5012 ( .C (clk), .D (new_AGEMA_signal_10863), .Q (new_AGEMA_signal_10864) ) ;
    buf_clk new_AGEMA_reg_buffer_5016 ( .C (clk), .D (new_AGEMA_signal_10867), .Q (new_AGEMA_signal_10868) ) ;
    buf_clk new_AGEMA_reg_buffer_5020 ( .C (clk), .D (new_AGEMA_signal_10871), .Q (new_AGEMA_signal_10872) ) ;
    buf_clk new_AGEMA_reg_buffer_5024 ( .C (clk), .D (new_AGEMA_signal_10875), .Q (new_AGEMA_signal_10876) ) ;
    buf_clk new_AGEMA_reg_buffer_5028 ( .C (clk), .D (new_AGEMA_signal_10879), .Q (new_AGEMA_signal_10880) ) ;
    buf_clk new_AGEMA_reg_buffer_5032 ( .C (clk), .D (new_AGEMA_signal_10883), .Q (new_AGEMA_signal_10884) ) ;
    buf_clk new_AGEMA_reg_buffer_5036 ( .C (clk), .D (new_AGEMA_signal_10887), .Q (new_AGEMA_signal_10888) ) ;
    buf_clk new_AGEMA_reg_buffer_5040 ( .C (clk), .D (new_AGEMA_signal_10891), .Q (new_AGEMA_signal_10892) ) ;
    buf_clk new_AGEMA_reg_buffer_5044 ( .C (clk), .D (new_AGEMA_signal_10895), .Q (new_AGEMA_signal_10896) ) ;
    buf_clk new_AGEMA_reg_buffer_5048 ( .C (clk), .D (new_AGEMA_signal_10899), .Q (new_AGEMA_signal_10900) ) ;
    buf_clk new_AGEMA_reg_buffer_5052 ( .C (clk), .D (new_AGEMA_signal_10903), .Q (new_AGEMA_signal_10904) ) ;
    buf_clk new_AGEMA_reg_buffer_5056 ( .C (clk), .D (new_AGEMA_signal_10907), .Q (new_AGEMA_signal_10908) ) ;
    buf_clk new_AGEMA_reg_buffer_5060 ( .C (clk), .D (new_AGEMA_signal_10911), .Q (new_AGEMA_signal_10912) ) ;
    buf_clk new_AGEMA_reg_buffer_5064 ( .C (clk), .D (new_AGEMA_signal_10915), .Q (new_AGEMA_signal_10916) ) ;
    buf_clk new_AGEMA_reg_buffer_5068 ( .C (clk), .D (new_AGEMA_signal_10919), .Q (new_AGEMA_signal_10920) ) ;
    buf_clk new_AGEMA_reg_buffer_5072 ( .C (clk), .D (new_AGEMA_signal_10923), .Q (new_AGEMA_signal_10924) ) ;
    buf_clk new_AGEMA_reg_buffer_5076 ( .C (clk), .D (new_AGEMA_signal_10927), .Q (new_AGEMA_signal_10928) ) ;
    buf_clk new_AGEMA_reg_buffer_5080 ( .C (clk), .D (new_AGEMA_signal_10931), .Q (new_AGEMA_signal_10932) ) ;
    buf_clk new_AGEMA_reg_buffer_5084 ( .C (clk), .D (new_AGEMA_signal_10935), .Q (new_AGEMA_signal_10936) ) ;
    buf_clk new_AGEMA_reg_buffer_5088 ( .C (clk), .D (new_AGEMA_signal_10939), .Q (new_AGEMA_signal_10940) ) ;
    buf_clk new_AGEMA_reg_buffer_5092 ( .C (clk), .D (new_AGEMA_signal_10943), .Q (new_AGEMA_signal_10944) ) ;
    buf_clk new_AGEMA_reg_buffer_5096 ( .C (clk), .D (new_AGEMA_signal_10947), .Q (new_AGEMA_signal_10948) ) ;
    buf_clk new_AGEMA_reg_buffer_5100 ( .C (clk), .D (new_AGEMA_signal_10951), .Q (new_AGEMA_signal_10952) ) ;
    buf_clk new_AGEMA_reg_buffer_5104 ( .C (clk), .D (new_AGEMA_signal_10955), .Q (new_AGEMA_signal_10956) ) ;
    buf_clk new_AGEMA_reg_buffer_5108 ( .C (clk), .D (new_AGEMA_signal_10959), .Q (new_AGEMA_signal_10960) ) ;
    buf_clk new_AGEMA_reg_buffer_5112 ( .C (clk), .D (new_AGEMA_signal_10963), .Q (new_AGEMA_signal_10964) ) ;
    buf_clk new_AGEMA_reg_buffer_5116 ( .C (clk), .D (new_AGEMA_signal_10967), .Q (new_AGEMA_signal_10968) ) ;
    buf_clk new_AGEMA_reg_buffer_5120 ( .C (clk), .D (new_AGEMA_signal_10971), .Q (new_AGEMA_signal_10972) ) ;
    buf_clk new_AGEMA_reg_buffer_5124 ( .C (clk), .D (new_AGEMA_signal_10975), .Q (new_AGEMA_signal_10976) ) ;
    buf_clk new_AGEMA_reg_buffer_5128 ( .C (clk), .D (new_AGEMA_signal_10979), .Q (new_AGEMA_signal_10980) ) ;
    buf_clk new_AGEMA_reg_buffer_5132 ( .C (clk), .D (new_AGEMA_signal_10983), .Q (new_AGEMA_signal_10984) ) ;
    buf_clk new_AGEMA_reg_buffer_5136 ( .C (clk), .D (new_AGEMA_signal_10987), .Q (new_AGEMA_signal_10988) ) ;
    buf_clk new_AGEMA_reg_buffer_5140 ( .C (clk), .D (new_AGEMA_signal_10991), .Q (new_AGEMA_signal_10992) ) ;
    buf_clk new_AGEMA_reg_buffer_5144 ( .C (clk), .D (new_AGEMA_signal_10995), .Q (new_AGEMA_signal_10996) ) ;
    buf_clk new_AGEMA_reg_buffer_5148 ( .C (clk), .D (new_AGEMA_signal_10999), .Q (new_AGEMA_signal_11000) ) ;
    buf_clk new_AGEMA_reg_buffer_5152 ( .C (clk), .D (new_AGEMA_signal_11003), .Q (new_AGEMA_signal_11004) ) ;
    buf_clk new_AGEMA_reg_buffer_5156 ( .C (clk), .D (new_AGEMA_signal_11007), .Q (new_AGEMA_signal_11008) ) ;
    buf_clk new_AGEMA_reg_buffer_5160 ( .C (clk), .D (new_AGEMA_signal_11011), .Q (new_AGEMA_signal_11012) ) ;
    buf_clk new_AGEMA_reg_buffer_5164 ( .C (clk), .D (new_AGEMA_signal_11015), .Q (new_AGEMA_signal_11016) ) ;
    buf_clk new_AGEMA_reg_buffer_5168 ( .C (clk), .D (new_AGEMA_signal_11019), .Q (new_AGEMA_signal_11020) ) ;
    buf_clk new_AGEMA_reg_buffer_5172 ( .C (clk), .D (new_AGEMA_signal_11023), .Q (new_AGEMA_signal_11024) ) ;
    buf_clk new_AGEMA_reg_buffer_5176 ( .C (clk), .D (new_AGEMA_signal_11027), .Q (new_AGEMA_signal_11028) ) ;
    buf_clk new_AGEMA_reg_buffer_5180 ( .C (clk), .D (new_AGEMA_signal_11031), .Q (new_AGEMA_signal_11032) ) ;
    buf_clk new_AGEMA_reg_buffer_5184 ( .C (clk), .D (new_AGEMA_signal_11035), .Q (new_AGEMA_signal_11036) ) ;
    buf_clk new_AGEMA_reg_buffer_5188 ( .C (clk), .D (new_AGEMA_signal_11039), .Q (new_AGEMA_signal_11040) ) ;
    buf_clk new_AGEMA_reg_buffer_5192 ( .C (clk), .D (new_AGEMA_signal_11043), .Q (new_AGEMA_signal_11044) ) ;
    buf_clk new_AGEMA_reg_buffer_5196 ( .C (clk), .D (new_AGEMA_signal_11047), .Q (new_AGEMA_signal_11048) ) ;
    buf_clk new_AGEMA_reg_buffer_5200 ( .C (clk), .D (new_AGEMA_signal_11051), .Q (new_AGEMA_signal_11052) ) ;
    buf_clk new_AGEMA_reg_buffer_5204 ( .C (clk), .D (new_AGEMA_signal_11055), .Q (new_AGEMA_signal_11056) ) ;
    buf_clk new_AGEMA_reg_buffer_5208 ( .C (clk), .D (new_AGEMA_signal_11059), .Q (new_AGEMA_signal_11060) ) ;
    buf_clk new_AGEMA_reg_buffer_5212 ( .C (clk), .D (new_AGEMA_signal_11063), .Q (new_AGEMA_signal_11064) ) ;
    buf_clk new_AGEMA_reg_buffer_5216 ( .C (clk), .D (new_AGEMA_signal_11067), .Q (new_AGEMA_signal_11068) ) ;
    buf_clk new_AGEMA_reg_buffer_5220 ( .C (clk), .D (new_AGEMA_signal_11071), .Q (new_AGEMA_signal_11072) ) ;
    buf_clk new_AGEMA_reg_buffer_5224 ( .C (clk), .D (new_AGEMA_signal_11075), .Q (new_AGEMA_signal_11076) ) ;
    buf_clk new_AGEMA_reg_buffer_5228 ( .C (clk), .D (new_AGEMA_signal_11079), .Q (new_AGEMA_signal_11080) ) ;
    buf_clk new_AGEMA_reg_buffer_5232 ( .C (clk), .D (new_AGEMA_signal_11083), .Q (new_AGEMA_signal_11084) ) ;
    buf_clk new_AGEMA_reg_buffer_5236 ( .C (clk), .D (new_AGEMA_signal_11087), .Q (new_AGEMA_signal_11088) ) ;
    buf_clk new_AGEMA_reg_buffer_5240 ( .C (clk), .D (new_AGEMA_signal_11091), .Q (new_AGEMA_signal_11092) ) ;
    buf_clk new_AGEMA_reg_buffer_5244 ( .C (clk), .D (new_AGEMA_signal_11095), .Q (new_AGEMA_signal_11096) ) ;
    buf_clk new_AGEMA_reg_buffer_5248 ( .C (clk), .D (new_AGEMA_signal_11099), .Q (new_AGEMA_signal_11100) ) ;
    buf_clk new_AGEMA_reg_buffer_5252 ( .C (clk), .D (new_AGEMA_signal_11103), .Q (new_AGEMA_signal_11104) ) ;
    buf_clk new_AGEMA_reg_buffer_5256 ( .C (clk), .D (new_AGEMA_signal_11107), .Q (new_AGEMA_signal_11108) ) ;
    buf_clk new_AGEMA_reg_buffer_5260 ( .C (clk), .D (new_AGEMA_signal_11111), .Q (new_AGEMA_signal_11112) ) ;
    buf_clk new_AGEMA_reg_buffer_5264 ( .C (clk), .D (new_AGEMA_signal_11115), .Q (new_AGEMA_signal_11116) ) ;
    buf_clk new_AGEMA_reg_buffer_5268 ( .C (clk), .D (new_AGEMA_signal_11119), .Q (new_AGEMA_signal_11120) ) ;
    buf_clk new_AGEMA_reg_buffer_5272 ( .C (clk), .D (new_AGEMA_signal_11123), .Q (new_AGEMA_signal_11124) ) ;
    buf_clk new_AGEMA_reg_buffer_5276 ( .C (clk), .D (new_AGEMA_signal_11127), .Q (new_AGEMA_signal_11128) ) ;
    buf_clk new_AGEMA_reg_buffer_5280 ( .C (clk), .D (new_AGEMA_signal_11131), .Q (new_AGEMA_signal_11132) ) ;
    buf_clk new_AGEMA_reg_buffer_5284 ( .C (clk), .D (new_AGEMA_signal_11135), .Q (new_AGEMA_signal_11136) ) ;
    buf_clk new_AGEMA_reg_buffer_5288 ( .C (clk), .D (new_AGEMA_signal_11139), .Q (new_AGEMA_signal_11140) ) ;
    buf_clk new_AGEMA_reg_buffer_5292 ( .C (clk), .D (new_AGEMA_signal_11143), .Q (new_AGEMA_signal_11144) ) ;
    buf_clk new_AGEMA_reg_buffer_5296 ( .C (clk), .D (new_AGEMA_signal_11147), .Q (new_AGEMA_signal_11148) ) ;
    buf_clk new_AGEMA_reg_buffer_5300 ( .C (clk), .D (new_AGEMA_signal_11151), .Q (new_AGEMA_signal_11152) ) ;
    buf_clk new_AGEMA_reg_buffer_5304 ( .C (clk), .D (new_AGEMA_signal_11155), .Q (new_AGEMA_signal_11156) ) ;
    buf_clk new_AGEMA_reg_buffer_5308 ( .C (clk), .D (new_AGEMA_signal_11159), .Q (new_AGEMA_signal_11160) ) ;
    buf_clk new_AGEMA_reg_buffer_5312 ( .C (clk), .D (new_AGEMA_signal_11163), .Q (new_AGEMA_signal_11164) ) ;
    buf_clk new_AGEMA_reg_buffer_5316 ( .C (clk), .D (new_AGEMA_signal_11167), .Q (new_AGEMA_signal_11168) ) ;
    buf_clk new_AGEMA_reg_buffer_5320 ( .C (clk), .D (new_AGEMA_signal_11171), .Q (new_AGEMA_signal_11172) ) ;
    buf_clk new_AGEMA_reg_buffer_5324 ( .C (clk), .D (new_AGEMA_signal_11175), .Q (new_AGEMA_signal_11176) ) ;
    buf_clk new_AGEMA_reg_buffer_5328 ( .C (clk), .D (new_AGEMA_signal_11179), .Q (new_AGEMA_signal_11180) ) ;
    buf_clk new_AGEMA_reg_buffer_5332 ( .C (clk), .D (new_AGEMA_signal_11183), .Q (new_AGEMA_signal_11184) ) ;
    buf_clk new_AGEMA_reg_buffer_5336 ( .C (clk), .D (new_AGEMA_signal_11187), .Q (new_AGEMA_signal_11188) ) ;
    buf_clk new_AGEMA_reg_buffer_5340 ( .C (clk), .D (new_AGEMA_signal_11191), .Q (new_AGEMA_signal_11192) ) ;
    buf_clk new_AGEMA_reg_buffer_5344 ( .C (clk), .D (new_AGEMA_signal_11195), .Q (new_AGEMA_signal_11196) ) ;
    buf_clk new_AGEMA_reg_buffer_5348 ( .C (clk), .D (new_AGEMA_signal_11199), .Q (new_AGEMA_signal_11200) ) ;
    buf_clk new_AGEMA_reg_buffer_5352 ( .C (clk), .D (new_AGEMA_signal_11203), .Q (new_AGEMA_signal_11204) ) ;
    buf_clk new_AGEMA_reg_buffer_5356 ( .C (clk), .D (new_AGEMA_signal_11207), .Q (new_AGEMA_signal_11208) ) ;
    buf_clk new_AGEMA_reg_buffer_5360 ( .C (clk), .D (new_AGEMA_signal_11211), .Q (new_AGEMA_signal_11212) ) ;
    buf_clk new_AGEMA_reg_buffer_5364 ( .C (clk), .D (new_AGEMA_signal_11215), .Q (new_AGEMA_signal_11216) ) ;
    buf_clk new_AGEMA_reg_buffer_5368 ( .C (clk), .D (new_AGEMA_signal_11219), .Q (new_AGEMA_signal_11220) ) ;
    buf_clk new_AGEMA_reg_buffer_5372 ( .C (clk), .D (new_AGEMA_signal_11223), .Q (new_AGEMA_signal_11224) ) ;
    buf_clk new_AGEMA_reg_buffer_5376 ( .C (clk), .D (new_AGEMA_signal_11227), .Q (new_AGEMA_signal_11228) ) ;
    buf_clk new_AGEMA_reg_buffer_5380 ( .C (clk), .D (new_AGEMA_signal_11231), .Q (new_AGEMA_signal_11232) ) ;
    buf_clk new_AGEMA_reg_buffer_5384 ( .C (clk), .D (new_AGEMA_signal_11235), .Q (new_AGEMA_signal_11236) ) ;
    buf_clk new_AGEMA_reg_buffer_5388 ( .C (clk), .D (new_AGEMA_signal_11239), .Q (new_AGEMA_signal_11240) ) ;
    buf_clk new_AGEMA_reg_buffer_5392 ( .C (clk), .D (new_AGEMA_signal_11243), .Q (new_AGEMA_signal_11244) ) ;
    buf_clk new_AGEMA_reg_buffer_5396 ( .C (clk), .D (new_AGEMA_signal_11247), .Q (new_AGEMA_signal_11248) ) ;
    buf_clk new_AGEMA_reg_buffer_5400 ( .C (clk), .D (new_AGEMA_signal_11251), .Q (new_AGEMA_signal_11252) ) ;
    buf_clk new_AGEMA_reg_buffer_5404 ( .C (clk), .D (new_AGEMA_signal_11255), .Q (new_AGEMA_signal_11256) ) ;
    buf_clk new_AGEMA_reg_buffer_5408 ( .C (clk), .D (new_AGEMA_signal_11259), .Q (new_AGEMA_signal_11260) ) ;
    buf_clk new_AGEMA_reg_buffer_5412 ( .C (clk), .D (new_AGEMA_signal_11263), .Q (new_AGEMA_signal_11264) ) ;
    buf_clk new_AGEMA_reg_buffer_5416 ( .C (clk), .D (new_AGEMA_signal_11267), .Q (new_AGEMA_signal_11268) ) ;
    buf_clk new_AGEMA_reg_buffer_5420 ( .C (clk), .D (new_AGEMA_signal_11271), .Q (new_AGEMA_signal_11272) ) ;
    buf_clk new_AGEMA_reg_buffer_5424 ( .C (clk), .D (new_AGEMA_signal_11275), .Q (new_AGEMA_signal_11276) ) ;
    buf_clk new_AGEMA_reg_buffer_5428 ( .C (clk), .D (new_AGEMA_signal_11279), .Q (new_AGEMA_signal_11280) ) ;
    buf_clk new_AGEMA_reg_buffer_5432 ( .C (clk), .D (new_AGEMA_signal_11283), .Q (new_AGEMA_signal_11284) ) ;
    buf_clk new_AGEMA_reg_buffer_5436 ( .C (clk), .D (new_AGEMA_signal_11287), .Q (new_AGEMA_signal_11288) ) ;
    buf_clk new_AGEMA_reg_buffer_5440 ( .C (clk), .D (new_AGEMA_signal_11291), .Q (new_AGEMA_signal_11292) ) ;
    buf_clk new_AGEMA_reg_buffer_5444 ( .C (clk), .D (new_AGEMA_signal_11295), .Q (new_AGEMA_signal_11296) ) ;
    buf_clk new_AGEMA_reg_buffer_5448 ( .C (clk), .D (new_AGEMA_signal_11299), .Q (new_AGEMA_signal_11300) ) ;
    buf_clk new_AGEMA_reg_buffer_5452 ( .C (clk), .D (new_AGEMA_signal_11303), .Q (new_AGEMA_signal_11304) ) ;
    buf_clk new_AGEMA_reg_buffer_5456 ( .C (clk), .D (new_AGEMA_signal_11307), .Q (new_AGEMA_signal_11308) ) ;
    buf_clk new_AGEMA_reg_buffer_5460 ( .C (clk), .D (new_AGEMA_signal_11311), .Q (new_AGEMA_signal_11312) ) ;
    buf_clk new_AGEMA_reg_buffer_5464 ( .C (clk), .D (new_AGEMA_signal_11315), .Q (new_AGEMA_signal_11316) ) ;
    buf_clk new_AGEMA_reg_buffer_5468 ( .C (clk), .D (new_AGEMA_signal_11319), .Q (new_AGEMA_signal_11320) ) ;
    buf_clk new_AGEMA_reg_buffer_5472 ( .C (clk), .D (new_AGEMA_signal_11323), .Q (new_AGEMA_signal_11324) ) ;
    buf_clk new_AGEMA_reg_buffer_5476 ( .C (clk), .D (new_AGEMA_signal_11327), .Q (new_AGEMA_signal_11328) ) ;
    buf_clk new_AGEMA_reg_buffer_5480 ( .C (clk), .D (new_AGEMA_signal_11331), .Q (new_AGEMA_signal_11332) ) ;
    buf_clk new_AGEMA_reg_buffer_5484 ( .C (clk), .D (new_AGEMA_signal_11335), .Q (new_AGEMA_signal_11336) ) ;
    buf_clk new_AGEMA_reg_buffer_5488 ( .C (clk), .D (new_AGEMA_signal_11339), .Q (new_AGEMA_signal_11340) ) ;
    buf_clk new_AGEMA_reg_buffer_5492 ( .C (clk), .D (new_AGEMA_signal_11343), .Q (new_AGEMA_signal_11344) ) ;
    buf_clk new_AGEMA_reg_buffer_5496 ( .C (clk), .D (new_AGEMA_signal_11347), .Q (new_AGEMA_signal_11348) ) ;
    buf_clk new_AGEMA_reg_buffer_5500 ( .C (clk), .D (new_AGEMA_signal_11351), .Q (new_AGEMA_signal_11352) ) ;
    buf_clk new_AGEMA_reg_buffer_5504 ( .C (clk), .D (new_AGEMA_signal_11355), .Q (new_AGEMA_signal_11356) ) ;
    buf_clk new_AGEMA_reg_buffer_5508 ( .C (clk), .D (new_AGEMA_signal_11359), .Q (new_AGEMA_signal_11360) ) ;
    buf_clk new_AGEMA_reg_buffer_5512 ( .C (clk), .D (new_AGEMA_signal_11363), .Q (new_AGEMA_signal_11364) ) ;
    buf_clk new_AGEMA_reg_buffer_5516 ( .C (clk), .D (new_AGEMA_signal_11367), .Q (new_AGEMA_signal_11368) ) ;
    buf_clk new_AGEMA_reg_buffer_5520 ( .C (clk), .D (new_AGEMA_signal_11371), .Q (new_AGEMA_signal_11372) ) ;
    buf_clk new_AGEMA_reg_buffer_5524 ( .C (clk), .D (new_AGEMA_signal_11375), .Q (new_AGEMA_signal_11376) ) ;
    buf_clk new_AGEMA_reg_buffer_5528 ( .C (clk), .D (new_AGEMA_signal_11379), .Q (new_AGEMA_signal_11380) ) ;
    buf_clk new_AGEMA_reg_buffer_5532 ( .C (clk), .D (new_AGEMA_signal_11383), .Q (new_AGEMA_signal_11384) ) ;
    buf_clk new_AGEMA_reg_buffer_5536 ( .C (clk), .D (new_AGEMA_signal_11387), .Q (new_AGEMA_signal_11388) ) ;
    buf_clk new_AGEMA_reg_buffer_5540 ( .C (clk), .D (new_AGEMA_signal_11391), .Q (new_AGEMA_signal_11392) ) ;
    buf_clk new_AGEMA_reg_buffer_5544 ( .C (clk), .D (new_AGEMA_signal_11395), .Q (new_AGEMA_signal_11396) ) ;
    buf_clk new_AGEMA_reg_buffer_5548 ( .C (clk), .D (new_AGEMA_signal_11399), .Q (new_AGEMA_signal_11400) ) ;
    buf_clk new_AGEMA_reg_buffer_5552 ( .C (clk), .D (new_AGEMA_signal_11403), .Q (new_AGEMA_signal_11404) ) ;
    buf_clk new_AGEMA_reg_buffer_5556 ( .C (clk), .D (new_AGEMA_signal_11407), .Q (new_AGEMA_signal_11408) ) ;
    buf_clk new_AGEMA_reg_buffer_5560 ( .C (clk), .D (new_AGEMA_signal_11411), .Q (new_AGEMA_signal_11412) ) ;
    buf_clk new_AGEMA_reg_buffer_5564 ( .C (clk), .D (new_AGEMA_signal_11415), .Q (new_AGEMA_signal_11416) ) ;
    buf_clk new_AGEMA_reg_buffer_5568 ( .C (clk), .D (new_AGEMA_signal_11419), .Q (new_AGEMA_signal_11420) ) ;
    buf_clk new_AGEMA_reg_buffer_5572 ( .C (clk), .D (new_AGEMA_signal_11423), .Q (new_AGEMA_signal_11424) ) ;
    buf_clk new_AGEMA_reg_buffer_5576 ( .C (clk), .D (new_AGEMA_signal_11427), .Q (new_AGEMA_signal_11428) ) ;
    buf_clk new_AGEMA_reg_buffer_5580 ( .C (clk), .D (new_AGEMA_signal_11431), .Q (new_AGEMA_signal_11432) ) ;
    buf_clk new_AGEMA_reg_buffer_5584 ( .C (clk), .D (new_AGEMA_signal_11435), .Q (new_AGEMA_signal_11436) ) ;
    buf_clk new_AGEMA_reg_buffer_5588 ( .C (clk), .D (new_AGEMA_signal_11439), .Q (new_AGEMA_signal_11440) ) ;
    buf_clk new_AGEMA_reg_buffer_5592 ( .C (clk), .D (new_AGEMA_signal_11443), .Q (new_AGEMA_signal_11444) ) ;
    buf_clk new_AGEMA_reg_buffer_5596 ( .C (clk), .D (new_AGEMA_signal_11447), .Q (new_AGEMA_signal_11448) ) ;
    buf_clk new_AGEMA_reg_buffer_5600 ( .C (clk), .D (new_AGEMA_signal_11451), .Q (new_AGEMA_signal_11452) ) ;
    buf_clk new_AGEMA_reg_buffer_5604 ( .C (clk), .D (new_AGEMA_signal_11455), .Q (new_AGEMA_signal_11456) ) ;
    buf_clk new_AGEMA_reg_buffer_5608 ( .C (clk), .D (new_AGEMA_signal_11459), .Q (new_AGEMA_signal_11460) ) ;
    buf_clk new_AGEMA_reg_buffer_5612 ( .C (clk), .D (new_AGEMA_signal_11463), .Q (new_AGEMA_signal_11464) ) ;
    buf_clk new_AGEMA_reg_buffer_5616 ( .C (clk), .D (new_AGEMA_signal_11467), .Q (new_AGEMA_signal_11468) ) ;
    buf_clk new_AGEMA_reg_buffer_5620 ( .C (clk), .D (new_AGEMA_signal_11471), .Q (new_AGEMA_signal_11472) ) ;
    buf_clk new_AGEMA_reg_buffer_5624 ( .C (clk), .D (new_AGEMA_signal_11475), .Q (new_AGEMA_signal_11476) ) ;
    buf_clk new_AGEMA_reg_buffer_5628 ( .C (clk), .D (new_AGEMA_signal_11479), .Q (new_AGEMA_signal_11480) ) ;
    buf_clk new_AGEMA_reg_buffer_5632 ( .C (clk), .D (new_AGEMA_signal_11483), .Q (new_AGEMA_signal_11484) ) ;
    buf_clk new_AGEMA_reg_buffer_5636 ( .C (clk), .D (new_AGEMA_signal_11487), .Q (new_AGEMA_signal_11488) ) ;
    buf_clk new_AGEMA_reg_buffer_5640 ( .C (clk), .D (new_AGEMA_signal_11491), .Q (new_AGEMA_signal_11492) ) ;
    buf_clk new_AGEMA_reg_buffer_5644 ( .C (clk), .D (new_AGEMA_signal_11495), .Q (new_AGEMA_signal_11496) ) ;
    buf_clk new_AGEMA_reg_buffer_5648 ( .C (clk), .D (new_AGEMA_signal_11499), .Q (new_AGEMA_signal_11500) ) ;
    buf_clk new_AGEMA_reg_buffer_5652 ( .C (clk), .D (new_AGEMA_signal_11503), .Q (new_AGEMA_signal_11504) ) ;
    buf_clk new_AGEMA_reg_buffer_5656 ( .C (clk), .D (new_AGEMA_signal_11507), .Q (new_AGEMA_signal_11508) ) ;
    buf_clk new_AGEMA_reg_buffer_5660 ( .C (clk), .D (new_AGEMA_signal_11511), .Q (new_AGEMA_signal_11512) ) ;
    buf_clk new_AGEMA_reg_buffer_5664 ( .C (clk), .D (new_AGEMA_signal_11515), .Q (new_AGEMA_signal_11516) ) ;
    buf_clk new_AGEMA_reg_buffer_5668 ( .C (clk), .D (new_AGEMA_signal_11519), .Q (new_AGEMA_signal_11520) ) ;
    buf_clk new_AGEMA_reg_buffer_5672 ( .C (clk), .D (new_AGEMA_signal_11523), .Q (new_AGEMA_signal_11524) ) ;
    buf_clk new_AGEMA_reg_buffer_5676 ( .C (clk), .D (new_AGEMA_signal_11527), .Q (new_AGEMA_signal_11528) ) ;
    buf_clk new_AGEMA_reg_buffer_5680 ( .C (clk), .D (new_AGEMA_signal_11531), .Q (new_AGEMA_signal_11532) ) ;
    buf_clk new_AGEMA_reg_buffer_5684 ( .C (clk), .D (new_AGEMA_signal_11535), .Q (new_AGEMA_signal_11536) ) ;
    buf_clk new_AGEMA_reg_buffer_5688 ( .C (clk), .D (new_AGEMA_signal_11539), .Q (new_AGEMA_signal_11540) ) ;
    buf_clk new_AGEMA_reg_buffer_5692 ( .C (clk), .D (new_AGEMA_signal_11543), .Q (new_AGEMA_signal_11544) ) ;
    buf_clk new_AGEMA_reg_buffer_5696 ( .C (clk), .D (new_AGEMA_signal_11547), .Q (new_AGEMA_signal_11548) ) ;
    buf_clk new_AGEMA_reg_buffer_5700 ( .C (clk), .D (new_AGEMA_signal_11551), .Q (new_AGEMA_signal_11552) ) ;
    buf_clk new_AGEMA_reg_buffer_5704 ( .C (clk), .D (new_AGEMA_signal_11555), .Q (new_AGEMA_signal_11556) ) ;
    buf_clk new_AGEMA_reg_buffer_5708 ( .C (clk), .D (new_AGEMA_signal_11559), .Q (new_AGEMA_signal_11560) ) ;
    buf_clk new_AGEMA_reg_buffer_5712 ( .C (clk), .D (new_AGEMA_signal_11563), .Q (new_AGEMA_signal_11564) ) ;
    buf_clk new_AGEMA_reg_buffer_5716 ( .C (clk), .D (new_AGEMA_signal_11567), .Q (new_AGEMA_signal_11568) ) ;
    buf_clk new_AGEMA_reg_buffer_5720 ( .C (clk), .D (new_AGEMA_signal_11571), .Q (new_AGEMA_signal_11572) ) ;
    buf_clk new_AGEMA_reg_buffer_5724 ( .C (clk), .D (new_AGEMA_signal_11575), .Q (new_AGEMA_signal_11576) ) ;
    buf_clk new_AGEMA_reg_buffer_5728 ( .C (clk), .D (new_AGEMA_signal_11579), .Q (new_AGEMA_signal_11580) ) ;
    buf_clk new_AGEMA_reg_buffer_5732 ( .C (clk), .D (new_AGEMA_signal_11583), .Q (new_AGEMA_signal_11584) ) ;
    buf_clk new_AGEMA_reg_buffer_5736 ( .C (clk), .D (new_AGEMA_signal_11587), .Q (new_AGEMA_signal_11588) ) ;
    buf_clk new_AGEMA_reg_buffer_5740 ( .C (clk), .D (new_AGEMA_signal_11591), .Q (new_AGEMA_signal_11592) ) ;
    buf_clk new_AGEMA_reg_buffer_5744 ( .C (clk), .D (new_AGEMA_signal_11595), .Q (new_AGEMA_signal_11596) ) ;
    buf_clk new_AGEMA_reg_buffer_7476 ( .C (clk), .D (new_AGEMA_signal_13327), .Q (new_AGEMA_signal_13328) ) ;
    buf_clk new_AGEMA_reg_buffer_7480 ( .C (clk), .D (new_AGEMA_signal_13331), .Q (new_AGEMA_signal_13332) ) ;
    buf_clk new_AGEMA_reg_buffer_7484 ( .C (clk), .D (new_AGEMA_signal_13335), .Q (new_AGEMA_signal_13336) ) ;
    buf_clk new_AGEMA_reg_buffer_7488 ( .C (clk), .D (new_AGEMA_signal_13339), .Q (new_AGEMA_signal_13340) ) ;
    buf_clk new_AGEMA_reg_buffer_7492 ( .C (clk), .D (new_AGEMA_signal_13343), .Q (new_AGEMA_signal_13344) ) ;
    buf_clk new_AGEMA_reg_buffer_7496 ( .C (clk), .D (new_AGEMA_signal_13347), .Q (new_AGEMA_signal_13348) ) ;
    buf_clk new_AGEMA_reg_buffer_7500 ( .C (clk), .D (new_AGEMA_signal_13351), .Q (new_AGEMA_signal_13352) ) ;
    buf_clk new_AGEMA_reg_buffer_7504 ( .C (clk), .D (new_AGEMA_signal_13355), .Q (new_AGEMA_signal_13356) ) ;
    buf_clk new_AGEMA_reg_buffer_7508 ( .C (clk), .D (new_AGEMA_signal_13359), .Q (new_AGEMA_signal_13360) ) ;
    buf_clk new_AGEMA_reg_buffer_7512 ( .C (clk), .D (new_AGEMA_signal_13363), .Q (new_AGEMA_signal_13364) ) ;
    buf_clk new_AGEMA_reg_buffer_7516 ( .C (clk), .D (new_AGEMA_signal_13367), .Q (new_AGEMA_signal_13368) ) ;
    buf_clk new_AGEMA_reg_buffer_7520 ( .C (clk), .D (new_AGEMA_signal_13371), .Q (new_AGEMA_signal_13372) ) ;
    buf_clk new_AGEMA_reg_buffer_7524 ( .C (clk), .D (new_AGEMA_signal_13375), .Q (new_AGEMA_signal_13376) ) ;
    buf_clk new_AGEMA_reg_buffer_7528 ( .C (clk), .D (new_AGEMA_signal_13379), .Q (new_AGEMA_signal_13380) ) ;
    buf_clk new_AGEMA_reg_buffer_7532 ( .C (clk), .D (new_AGEMA_signal_13383), .Q (new_AGEMA_signal_13384) ) ;
    buf_clk new_AGEMA_reg_buffer_7536 ( .C (clk), .D (new_AGEMA_signal_13387), .Q (new_AGEMA_signal_13388) ) ;
    buf_clk new_AGEMA_reg_buffer_7540 ( .C (clk), .D (new_AGEMA_signal_13391), .Q (new_AGEMA_signal_13392) ) ;
    buf_clk new_AGEMA_reg_buffer_7544 ( .C (clk), .D (new_AGEMA_signal_13395), .Q (new_AGEMA_signal_13396) ) ;
    buf_clk new_AGEMA_reg_buffer_7548 ( .C (clk), .D (new_AGEMA_signal_13399), .Q (new_AGEMA_signal_13400) ) ;
    buf_clk new_AGEMA_reg_buffer_7552 ( .C (clk), .D (new_AGEMA_signal_13403), .Q (new_AGEMA_signal_13404) ) ;
    buf_clk new_AGEMA_reg_buffer_7556 ( .C (clk), .D (new_AGEMA_signal_13407), .Q (new_AGEMA_signal_13408) ) ;
    buf_clk new_AGEMA_reg_buffer_7560 ( .C (clk), .D (new_AGEMA_signal_13411), .Q (new_AGEMA_signal_13412) ) ;
    buf_clk new_AGEMA_reg_buffer_7564 ( .C (clk), .D (new_AGEMA_signal_13415), .Q (new_AGEMA_signal_13416) ) ;
    buf_clk new_AGEMA_reg_buffer_7568 ( .C (clk), .D (new_AGEMA_signal_13419), .Q (new_AGEMA_signal_13420) ) ;
    buf_clk new_AGEMA_reg_buffer_7572 ( .C (clk), .D (new_AGEMA_signal_13423), .Q (new_AGEMA_signal_13424) ) ;
    buf_clk new_AGEMA_reg_buffer_7576 ( .C (clk), .D (new_AGEMA_signal_13427), .Q (new_AGEMA_signal_13428) ) ;
    buf_clk new_AGEMA_reg_buffer_7580 ( .C (clk), .D (new_AGEMA_signal_13431), .Q (new_AGEMA_signal_13432) ) ;
    buf_clk new_AGEMA_reg_buffer_7584 ( .C (clk), .D (new_AGEMA_signal_13435), .Q (new_AGEMA_signal_13436) ) ;
    buf_clk new_AGEMA_reg_buffer_7588 ( .C (clk), .D (new_AGEMA_signal_13439), .Q (new_AGEMA_signal_13440) ) ;
    buf_clk new_AGEMA_reg_buffer_7592 ( .C (clk), .D (new_AGEMA_signal_13443), .Q (new_AGEMA_signal_13444) ) ;
    buf_clk new_AGEMA_reg_buffer_7596 ( .C (clk), .D (new_AGEMA_signal_13447), .Q (new_AGEMA_signal_13448) ) ;
    buf_clk new_AGEMA_reg_buffer_7600 ( .C (clk), .D (new_AGEMA_signal_13451), .Q (new_AGEMA_signal_13452) ) ;
    buf_clk new_AGEMA_reg_buffer_7604 ( .C (clk), .D (new_AGEMA_signal_13455), .Q (new_AGEMA_signal_13456) ) ;
    buf_clk new_AGEMA_reg_buffer_7608 ( .C (clk), .D (new_AGEMA_signal_13459), .Q (new_AGEMA_signal_13460) ) ;
    buf_clk new_AGEMA_reg_buffer_7612 ( .C (clk), .D (new_AGEMA_signal_13463), .Q (new_AGEMA_signal_13464) ) ;
    buf_clk new_AGEMA_reg_buffer_7616 ( .C (clk), .D (new_AGEMA_signal_13467), .Q (new_AGEMA_signal_13468) ) ;
    buf_clk new_AGEMA_reg_buffer_7620 ( .C (clk), .D (new_AGEMA_signal_13471), .Q (new_AGEMA_signal_13472) ) ;
    buf_clk new_AGEMA_reg_buffer_7624 ( .C (clk), .D (new_AGEMA_signal_13475), .Q (new_AGEMA_signal_13476) ) ;
    buf_clk new_AGEMA_reg_buffer_7628 ( .C (clk), .D (new_AGEMA_signal_13479), .Q (new_AGEMA_signal_13480) ) ;
    buf_clk new_AGEMA_reg_buffer_7632 ( .C (clk), .D (new_AGEMA_signal_13483), .Q (new_AGEMA_signal_13484) ) ;
    buf_clk new_AGEMA_reg_buffer_7636 ( .C (clk), .D (new_AGEMA_signal_13487), .Q (new_AGEMA_signal_13488) ) ;
    buf_clk new_AGEMA_reg_buffer_7640 ( .C (clk), .D (new_AGEMA_signal_13491), .Q (new_AGEMA_signal_13492) ) ;
    buf_clk new_AGEMA_reg_buffer_7644 ( .C (clk), .D (new_AGEMA_signal_13495), .Q (new_AGEMA_signal_13496) ) ;
    buf_clk new_AGEMA_reg_buffer_7648 ( .C (clk), .D (new_AGEMA_signal_13499), .Q (new_AGEMA_signal_13500) ) ;
    buf_clk new_AGEMA_reg_buffer_7652 ( .C (clk), .D (new_AGEMA_signal_13503), .Q (new_AGEMA_signal_13504) ) ;
    buf_clk new_AGEMA_reg_buffer_7656 ( .C (clk), .D (new_AGEMA_signal_13507), .Q (new_AGEMA_signal_13508) ) ;
    buf_clk new_AGEMA_reg_buffer_7660 ( .C (clk), .D (new_AGEMA_signal_13511), .Q (new_AGEMA_signal_13512) ) ;
    buf_clk new_AGEMA_reg_buffer_7664 ( .C (clk), .D (new_AGEMA_signal_13515), .Q (new_AGEMA_signal_13516) ) ;
    buf_clk new_AGEMA_reg_buffer_7668 ( .C (clk), .D (new_AGEMA_signal_13519), .Q (new_AGEMA_signal_13520) ) ;
    buf_clk new_AGEMA_reg_buffer_7672 ( .C (clk), .D (new_AGEMA_signal_13523), .Q (new_AGEMA_signal_13524) ) ;
    buf_clk new_AGEMA_reg_buffer_7676 ( .C (clk), .D (new_AGEMA_signal_13527), .Q (new_AGEMA_signal_13528) ) ;
    buf_clk new_AGEMA_reg_buffer_7680 ( .C (clk), .D (new_AGEMA_signal_13531), .Q (new_AGEMA_signal_13532) ) ;
    buf_clk new_AGEMA_reg_buffer_7684 ( .C (clk), .D (new_AGEMA_signal_13535), .Q (new_AGEMA_signal_13536) ) ;
    buf_clk new_AGEMA_reg_buffer_7688 ( .C (clk), .D (new_AGEMA_signal_13539), .Q (new_AGEMA_signal_13540) ) ;
    buf_clk new_AGEMA_reg_buffer_7692 ( .C (clk), .D (new_AGEMA_signal_13543), .Q (new_AGEMA_signal_13544) ) ;
    buf_clk new_AGEMA_reg_buffer_7696 ( .C (clk), .D (new_AGEMA_signal_13547), .Q (new_AGEMA_signal_13548) ) ;
    buf_clk new_AGEMA_reg_buffer_7700 ( .C (clk), .D (new_AGEMA_signal_13551), .Q (new_AGEMA_signal_13552) ) ;
    buf_clk new_AGEMA_reg_buffer_7704 ( .C (clk), .D (new_AGEMA_signal_13555), .Q (new_AGEMA_signal_13556) ) ;
    buf_clk new_AGEMA_reg_buffer_7708 ( .C (clk), .D (new_AGEMA_signal_13559), .Q (new_AGEMA_signal_13560) ) ;
    buf_clk new_AGEMA_reg_buffer_7712 ( .C (clk), .D (new_AGEMA_signal_13563), .Q (new_AGEMA_signal_13564) ) ;
    buf_clk new_AGEMA_reg_buffer_7716 ( .C (clk), .D (new_AGEMA_signal_13567), .Q (new_AGEMA_signal_13568) ) ;
    buf_clk new_AGEMA_reg_buffer_7720 ( .C (clk), .D (new_AGEMA_signal_13571), .Q (new_AGEMA_signal_13572) ) ;
    buf_clk new_AGEMA_reg_buffer_7724 ( .C (clk), .D (new_AGEMA_signal_13575), .Q (new_AGEMA_signal_13576) ) ;
    buf_clk new_AGEMA_reg_buffer_7728 ( .C (clk), .D (new_AGEMA_signal_13579), .Q (new_AGEMA_signal_13580) ) ;
    buf_clk new_AGEMA_reg_buffer_7732 ( .C (clk), .D (new_AGEMA_signal_13583), .Q (new_AGEMA_signal_13584) ) ;
    buf_clk new_AGEMA_reg_buffer_7736 ( .C (clk), .D (new_AGEMA_signal_13587), .Q (new_AGEMA_signal_13588) ) ;
    buf_clk new_AGEMA_reg_buffer_7740 ( .C (clk), .D (new_AGEMA_signal_13591), .Q (new_AGEMA_signal_13592) ) ;
    buf_clk new_AGEMA_reg_buffer_7744 ( .C (clk), .D (new_AGEMA_signal_13595), .Q (new_AGEMA_signal_13596) ) ;
    buf_clk new_AGEMA_reg_buffer_7748 ( .C (clk), .D (new_AGEMA_signal_13599), .Q (new_AGEMA_signal_13600) ) ;
    buf_clk new_AGEMA_reg_buffer_7752 ( .C (clk), .D (new_AGEMA_signal_13603), .Q (new_AGEMA_signal_13604) ) ;
    buf_clk new_AGEMA_reg_buffer_7756 ( .C (clk), .D (new_AGEMA_signal_13607), .Q (new_AGEMA_signal_13608) ) ;
    buf_clk new_AGEMA_reg_buffer_7760 ( .C (clk), .D (new_AGEMA_signal_13611), .Q (new_AGEMA_signal_13612) ) ;
    buf_clk new_AGEMA_reg_buffer_7764 ( .C (clk), .D (new_AGEMA_signal_13615), .Q (new_AGEMA_signal_13616) ) ;
    buf_clk new_AGEMA_reg_buffer_7768 ( .C (clk), .D (new_AGEMA_signal_13619), .Q (new_AGEMA_signal_13620) ) ;
    buf_clk new_AGEMA_reg_buffer_7772 ( .C (clk), .D (new_AGEMA_signal_13623), .Q (new_AGEMA_signal_13624) ) ;
    buf_clk new_AGEMA_reg_buffer_7776 ( .C (clk), .D (new_AGEMA_signal_13627), .Q (new_AGEMA_signal_13628) ) ;
    buf_clk new_AGEMA_reg_buffer_7780 ( .C (clk), .D (new_AGEMA_signal_13631), .Q (new_AGEMA_signal_13632) ) ;
    buf_clk new_AGEMA_reg_buffer_7784 ( .C (clk), .D (new_AGEMA_signal_13635), .Q (new_AGEMA_signal_13636) ) ;
    buf_clk new_AGEMA_reg_buffer_7788 ( .C (clk), .D (new_AGEMA_signal_13639), .Q (new_AGEMA_signal_13640) ) ;
    buf_clk new_AGEMA_reg_buffer_7792 ( .C (clk), .D (new_AGEMA_signal_13643), .Q (new_AGEMA_signal_13644) ) ;
    buf_clk new_AGEMA_reg_buffer_7796 ( .C (clk), .D (new_AGEMA_signal_13647), .Q (new_AGEMA_signal_13648) ) ;
    buf_clk new_AGEMA_reg_buffer_7800 ( .C (clk), .D (new_AGEMA_signal_13651), .Q (new_AGEMA_signal_13652) ) ;
    buf_clk new_AGEMA_reg_buffer_7804 ( .C (clk), .D (new_AGEMA_signal_13655), .Q (new_AGEMA_signal_13656) ) ;
    buf_clk new_AGEMA_reg_buffer_7808 ( .C (clk), .D (new_AGEMA_signal_13659), .Q (new_AGEMA_signal_13660) ) ;
    buf_clk new_AGEMA_reg_buffer_7812 ( .C (clk), .D (new_AGEMA_signal_13663), .Q (new_AGEMA_signal_13664) ) ;
    buf_clk new_AGEMA_reg_buffer_7816 ( .C (clk), .D (new_AGEMA_signal_13667), .Q (new_AGEMA_signal_13668) ) ;
    buf_clk new_AGEMA_reg_buffer_7820 ( .C (clk), .D (new_AGEMA_signal_13671), .Q (new_AGEMA_signal_13672) ) ;
    buf_clk new_AGEMA_reg_buffer_7824 ( .C (clk), .D (new_AGEMA_signal_13675), .Q (new_AGEMA_signal_13676) ) ;
    buf_clk new_AGEMA_reg_buffer_7828 ( .C (clk), .D (new_AGEMA_signal_13679), .Q (new_AGEMA_signal_13680) ) ;
    buf_clk new_AGEMA_reg_buffer_7832 ( .C (clk), .D (new_AGEMA_signal_13683), .Q (new_AGEMA_signal_13684) ) ;
    buf_clk new_AGEMA_reg_buffer_7836 ( .C (clk), .D (new_AGEMA_signal_13687), .Q (new_AGEMA_signal_13688) ) ;
    buf_clk new_AGEMA_reg_buffer_7840 ( .C (clk), .D (new_AGEMA_signal_13691), .Q (new_AGEMA_signal_13692) ) ;
    buf_clk new_AGEMA_reg_buffer_7844 ( .C (clk), .D (new_AGEMA_signal_13695), .Q (new_AGEMA_signal_13696) ) ;
    buf_clk new_AGEMA_reg_buffer_7848 ( .C (clk), .D (new_AGEMA_signal_13699), .Q (new_AGEMA_signal_13700) ) ;
    buf_clk new_AGEMA_reg_buffer_7852 ( .C (clk), .D (new_AGEMA_signal_13703), .Q (new_AGEMA_signal_13704) ) ;
    buf_clk new_AGEMA_reg_buffer_7856 ( .C (clk), .D (new_AGEMA_signal_13707), .Q (new_AGEMA_signal_13708) ) ;
    buf_clk new_AGEMA_reg_buffer_7860 ( .C (clk), .D (new_AGEMA_signal_13711), .Q (new_AGEMA_signal_13712) ) ;
    buf_clk new_AGEMA_reg_buffer_7864 ( .C (clk), .D (new_AGEMA_signal_13715), .Q (new_AGEMA_signal_13716) ) ;
    buf_clk new_AGEMA_reg_buffer_7868 ( .C (clk), .D (new_AGEMA_signal_13719), .Q (new_AGEMA_signal_13720) ) ;
    buf_clk new_AGEMA_reg_buffer_7872 ( .C (clk), .D (new_AGEMA_signal_13723), .Q (new_AGEMA_signal_13724) ) ;
    buf_clk new_AGEMA_reg_buffer_7876 ( .C (clk), .D (new_AGEMA_signal_13727), .Q (new_AGEMA_signal_13728) ) ;
    buf_clk new_AGEMA_reg_buffer_7880 ( .C (clk), .D (new_AGEMA_signal_13731), .Q (new_AGEMA_signal_13732) ) ;
    buf_clk new_AGEMA_reg_buffer_7884 ( .C (clk), .D (new_AGEMA_signal_13735), .Q (new_AGEMA_signal_13736) ) ;
    buf_clk new_AGEMA_reg_buffer_7888 ( .C (clk), .D (new_AGEMA_signal_13739), .Q (new_AGEMA_signal_13740) ) ;
    buf_clk new_AGEMA_reg_buffer_7892 ( .C (clk), .D (new_AGEMA_signal_13743), .Q (new_AGEMA_signal_13744) ) ;
    buf_clk new_AGEMA_reg_buffer_7896 ( .C (clk), .D (new_AGEMA_signal_13747), .Q (new_AGEMA_signal_13748) ) ;
    buf_clk new_AGEMA_reg_buffer_7900 ( .C (clk), .D (new_AGEMA_signal_13751), .Q (new_AGEMA_signal_13752) ) ;
    buf_clk new_AGEMA_reg_buffer_7904 ( .C (clk), .D (new_AGEMA_signal_13755), .Q (new_AGEMA_signal_13756) ) ;
    buf_clk new_AGEMA_reg_buffer_7908 ( .C (clk), .D (new_AGEMA_signal_13759), .Q (new_AGEMA_signal_13760) ) ;
    buf_clk new_AGEMA_reg_buffer_7912 ( .C (clk), .D (new_AGEMA_signal_13763), .Q (new_AGEMA_signal_13764) ) ;
    buf_clk new_AGEMA_reg_buffer_7916 ( .C (clk), .D (new_AGEMA_signal_13767), .Q (new_AGEMA_signal_13768) ) ;
    buf_clk new_AGEMA_reg_buffer_7920 ( .C (clk), .D (new_AGEMA_signal_13771), .Q (new_AGEMA_signal_13772) ) ;
    buf_clk new_AGEMA_reg_buffer_7924 ( .C (clk), .D (new_AGEMA_signal_13775), .Q (new_AGEMA_signal_13776) ) ;
    buf_clk new_AGEMA_reg_buffer_7928 ( .C (clk), .D (new_AGEMA_signal_13779), .Q (new_AGEMA_signal_13780) ) ;
    buf_clk new_AGEMA_reg_buffer_7932 ( .C (clk), .D (new_AGEMA_signal_13783), .Q (new_AGEMA_signal_13784) ) ;
    buf_clk new_AGEMA_reg_buffer_7936 ( .C (clk), .D (new_AGEMA_signal_13787), .Q (new_AGEMA_signal_13788) ) ;
    buf_clk new_AGEMA_reg_buffer_7940 ( .C (clk), .D (new_AGEMA_signal_13791), .Q (new_AGEMA_signal_13792) ) ;
    buf_clk new_AGEMA_reg_buffer_7944 ( .C (clk), .D (new_AGEMA_signal_13795), .Q (new_AGEMA_signal_13796) ) ;
    buf_clk new_AGEMA_reg_buffer_7948 ( .C (clk), .D (new_AGEMA_signal_13799), .Q (new_AGEMA_signal_13800) ) ;
    buf_clk new_AGEMA_reg_buffer_7952 ( .C (clk), .D (new_AGEMA_signal_13803), .Q (new_AGEMA_signal_13804) ) ;
    buf_clk new_AGEMA_reg_buffer_7956 ( .C (clk), .D (new_AGEMA_signal_13807), .Q (new_AGEMA_signal_13808) ) ;
    buf_clk new_AGEMA_reg_buffer_7960 ( .C (clk), .D (new_AGEMA_signal_13811), .Q (new_AGEMA_signal_13812) ) ;
    buf_clk new_AGEMA_reg_buffer_7964 ( .C (clk), .D (new_AGEMA_signal_13815), .Q (new_AGEMA_signal_13816) ) ;
    buf_clk new_AGEMA_reg_buffer_7968 ( .C (clk), .D (new_AGEMA_signal_13819), .Q (new_AGEMA_signal_13820) ) ;
    buf_clk new_AGEMA_reg_buffer_7972 ( .C (clk), .D (new_AGEMA_signal_13823), .Q (new_AGEMA_signal_13824) ) ;
    buf_clk new_AGEMA_reg_buffer_7976 ( .C (clk), .D (new_AGEMA_signal_13827), .Q (new_AGEMA_signal_13828) ) ;
    buf_clk new_AGEMA_reg_buffer_7980 ( .C (clk), .D (new_AGEMA_signal_13831), .Q (new_AGEMA_signal_13832) ) ;
    buf_clk new_AGEMA_reg_buffer_7984 ( .C (clk), .D (new_AGEMA_signal_13835), .Q (new_AGEMA_signal_13836) ) ;
    buf_clk new_AGEMA_reg_buffer_7988 ( .C (clk), .D (new_AGEMA_signal_13839), .Q (new_AGEMA_signal_13840) ) ;
    buf_clk new_AGEMA_reg_buffer_7992 ( .C (clk), .D (new_AGEMA_signal_13843), .Q (new_AGEMA_signal_13844) ) ;
    buf_clk new_AGEMA_reg_buffer_7996 ( .C (clk), .D (new_AGEMA_signal_13847), .Q (new_AGEMA_signal_13848) ) ;
    buf_clk new_AGEMA_reg_buffer_8000 ( .C (clk), .D (new_AGEMA_signal_13851), .Q (new_AGEMA_signal_13852) ) ;
    buf_clk new_AGEMA_reg_buffer_8004 ( .C (clk), .D (new_AGEMA_signal_13855), .Q (new_AGEMA_signal_13856) ) ;
    buf_clk new_AGEMA_reg_buffer_8008 ( .C (clk), .D (new_AGEMA_signal_13859), .Q (new_AGEMA_signal_13860) ) ;
    buf_clk new_AGEMA_reg_buffer_8012 ( .C (clk), .D (new_AGEMA_signal_13863), .Q (new_AGEMA_signal_13864) ) ;
    buf_clk new_AGEMA_reg_buffer_8016 ( .C (clk), .D (new_AGEMA_signal_13867), .Q (new_AGEMA_signal_13868) ) ;
    buf_clk new_AGEMA_reg_buffer_8020 ( .C (clk), .D (new_AGEMA_signal_13871), .Q (new_AGEMA_signal_13872) ) ;
    buf_clk new_AGEMA_reg_buffer_8024 ( .C (clk), .D (new_AGEMA_signal_13875), .Q (new_AGEMA_signal_13876) ) ;
    buf_clk new_AGEMA_reg_buffer_8028 ( .C (clk), .D (new_AGEMA_signal_13879), .Q (new_AGEMA_signal_13880) ) ;
    buf_clk new_AGEMA_reg_buffer_8032 ( .C (clk), .D (new_AGEMA_signal_13883), .Q (new_AGEMA_signal_13884) ) ;
    buf_clk new_AGEMA_reg_buffer_8036 ( .C (clk), .D (new_AGEMA_signal_13887), .Q (new_AGEMA_signal_13888) ) ;
    buf_clk new_AGEMA_reg_buffer_8040 ( .C (clk), .D (new_AGEMA_signal_13891), .Q (new_AGEMA_signal_13892) ) ;
    buf_clk new_AGEMA_reg_buffer_8044 ( .C (clk), .D (new_AGEMA_signal_13895), .Q (new_AGEMA_signal_13896) ) ;
    buf_clk new_AGEMA_reg_buffer_8048 ( .C (clk), .D (new_AGEMA_signal_13899), .Q (new_AGEMA_signal_13900) ) ;
    buf_clk new_AGEMA_reg_buffer_8052 ( .C (clk), .D (new_AGEMA_signal_13903), .Q (new_AGEMA_signal_13904) ) ;
    buf_clk new_AGEMA_reg_buffer_8056 ( .C (clk), .D (new_AGEMA_signal_13907), .Q (new_AGEMA_signal_13908) ) ;
    buf_clk new_AGEMA_reg_buffer_8060 ( .C (clk), .D (new_AGEMA_signal_13911), .Q (new_AGEMA_signal_13912) ) ;
    buf_clk new_AGEMA_reg_buffer_8064 ( .C (clk), .D (new_AGEMA_signal_13915), .Q (new_AGEMA_signal_13916) ) ;
    buf_clk new_AGEMA_reg_buffer_8068 ( .C (clk), .D (new_AGEMA_signal_13919), .Q (new_AGEMA_signal_13920) ) ;
    buf_clk new_AGEMA_reg_buffer_8072 ( .C (clk), .D (new_AGEMA_signal_13923), .Q (new_AGEMA_signal_13924) ) ;
    buf_clk new_AGEMA_reg_buffer_8076 ( .C (clk), .D (new_AGEMA_signal_13927), .Q (new_AGEMA_signal_13928) ) ;
    buf_clk new_AGEMA_reg_buffer_8080 ( .C (clk), .D (new_AGEMA_signal_13931), .Q (new_AGEMA_signal_13932) ) ;
    buf_clk new_AGEMA_reg_buffer_8084 ( .C (clk), .D (new_AGEMA_signal_13935), .Q (new_AGEMA_signal_13936) ) ;
    buf_clk new_AGEMA_reg_buffer_8088 ( .C (clk), .D (new_AGEMA_signal_13939), .Q (new_AGEMA_signal_13940) ) ;
    buf_clk new_AGEMA_reg_buffer_8092 ( .C (clk), .D (new_AGEMA_signal_13943), .Q (new_AGEMA_signal_13944) ) ;
    buf_clk new_AGEMA_reg_buffer_8096 ( .C (clk), .D (new_AGEMA_signal_13947), .Q (new_AGEMA_signal_13948) ) ;
    buf_clk new_AGEMA_reg_buffer_8100 ( .C (clk), .D (new_AGEMA_signal_13951), .Q (new_AGEMA_signal_13952) ) ;
    buf_clk new_AGEMA_reg_buffer_8104 ( .C (clk), .D (new_AGEMA_signal_13955), .Q (new_AGEMA_signal_13956) ) ;
    buf_clk new_AGEMA_reg_buffer_8108 ( .C (clk), .D (new_AGEMA_signal_13959), .Q (new_AGEMA_signal_13960) ) ;
    buf_clk new_AGEMA_reg_buffer_8112 ( .C (clk), .D (new_AGEMA_signal_13963), .Q (new_AGEMA_signal_13964) ) ;
    buf_clk new_AGEMA_reg_buffer_8116 ( .C (clk), .D (new_AGEMA_signal_13967), .Q (new_AGEMA_signal_13968) ) ;
    buf_clk new_AGEMA_reg_buffer_8120 ( .C (clk), .D (new_AGEMA_signal_13971), .Q (new_AGEMA_signal_13972) ) ;
    buf_clk new_AGEMA_reg_buffer_8124 ( .C (clk), .D (new_AGEMA_signal_13975), .Q (new_AGEMA_signal_13976) ) ;
    buf_clk new_AGEMA_reg_buffer_8128 ( .C (clk), .D (new_AGEMA_signal_13979), .Q (new_AGEMA_signal_13980) ) ;
    buf_clk new_AGEMA_reg_buffer_8132 ( .C (clk), .D (new_AGEMA_signal_13983), .Q (new_AGEMA_signal_13984) ) ;
    buf_clk new_AGEMA_reg_buffer_8136 ( .C (clk), .D (new_AGEMA_signal_13987), .Q (new_AGEMA_signal_13988) ) ;
    buf_clk new_AGEMA_reg_buffer_8140 ( .C (clk), .D (new_AGEMA_signal_13991), .Q (new_AGEMA_signal_13992) ) ;
    buf_clk new_AGEMA_reg_buffer_8144 ( .C (clk), .D (new_AGEMA_signal_13995), .Q (new_AGEMA_signal_13996) ) ;
    buf_clk new_AGEMA_reg_buffer_8148 ( .C (clk), .D (new_AGEMA_signal_13999), .Q (new_AGEMA_signal_14000) ) ;
    buf_clk new_AGEMA_reg_buffer_8152 ( .C (clk), .D (new_AGEMA_signal_14003), .Q (new_AGEMA_signal_14004) ) ;
    buf_clk new_AGEMA_reg_buffer_8156 ( .C (clk), .D (new_AGEMA_signal_14007), .Q (new_AGEMA_signal_14008) ) ;
    buf_clk new_AGEMA_reg_buffer_8160 ( .C (clk), .D (new_AGEMA_signal_14011), .Q (new_AGEMA_signal_14012) ) ;
    buf_clk new_AGEMA_reg_buffer_8164 ( .C (clk), .D (new_AGEMA_signal_14015), .Q (new_AGEMA_signal_14016) ) ;
    buf_clk new_AGEMA_reg_buffer_8168 ( .C (clk), .D (new_AGEMA_signal_14019), .Q (new_AGEMA_signal_14020) ) ;
    buf_clk new_AGEMA_reg_buffer_8172 ( .C (clk), .D (new_AGEMA_signal_14023), .Q (new_AGEMA_signal_14024) ) ;
    buf_clk new_AGEMA_reg_buffer_8176 ( .C (clk), .D (new_AGEMA_signal_14027), .Q (new_AGEMA_signal_14028) ) ;
    buf_clk new_AGEMA_reg_buffer_8180 ( .C (clk), .D (new_AGEMA_signal_14031), .Q (new_AGEMA_signal_14032) ) ;
    buf_clk new_AGEMA_reg_buffer_8184 ( .C (clk), .D (new_AGEMA_signal_14035), .Q (new_AGEMA_signal_14036) ) ;
    buf_clk new_AGEMA_reg_buffer_8188 ( .C (clk), .D (new_AGEMA_signal_14039), .Q (new_AGEMA_signal_14040) ) ;
    buf_clk new_AGEMA_reg_buffer_8192 ( .C (clk), .D (new_AGEMA_signal_14043), .Q (new_AGEMA_signal_14044) ) ;
    buf_clk new_AGEMA_reg_buffer_8196 ( .C (clk), .D (new_AGEMA_signal_14047), .Q (new_AGEMA_signal_14048) ) ;
    buf_clk new_AGEMA_reg_buffer_8200 ( .C (clk), .D (new_AGEMA_signal_14051), .Q (new_AGEMA_signal_14052) ) ;
    buf_clk new_AGEMA_reg_buffer_8204 ( .C (clk), .D (new_AGEMA_signal_14055), .Q (new_AGEMA_signal_14056) ) ;
    buf_clk new_AGEMA_reg_buffer_8208 ( .C (clk), .D (new_AGEMA_signal_14059), .Q (new_AGEMA_signal_14060) ) ;
    buf_clk new_AGEMA_reg_buffer_8212 ( .C (clk), .D (new_AGEMA_signal_14063), .Q (new_AGEMA_signal_14064) ) ;
    buf_clk new_AGEMA_reg_buffer_8216 ( .C (clk), .D (new_AGEMA_signal_14067), .Q (new_AGEMA_signal_14068) ) ;
    buf_clk new_AGEMA_reg_buffer_8220 ( .C (clk), .D (new_AGEMA_signal_14071), .Q (new_AGEMA_signal_14072) ) ;
    buf_clk new_AGEMA_reg_buffer_8224 ( .C (clk), .D (new_AGEMA_signal_14075), .Q (new_AGEMA_signal_14076) ) ;
    buf_clk new_AGEMA_reg_buffer_8228 ( .C (clk), .D (new_AGEMA_signal_14079), .Q (new_AGEMA_signal_14080) ) ;
    buf_clk new_AGEMA_reg_buffer_8232 ( .C (clk), .D (new_AGEMA_signal_14083), .Q (new_AGEMA_signal_14084) ) ;
    buf_clk new_AGEMA_reg_buffer_8236 ( .C (clk), .D (new_AGEMA_signal_14087), .Q (new_AGEMA_signal_14088) ) ;
    buf_clk new_AGEMA_reg_buffer_8240 ( .C (clk), .D (new_AGEMA_signal_14091), .Q (new_AGEMA_signal_14092) ) ;
    buf_clk new_AGEMA_reg_buffer_8244 ( .C (clk), .D (new_AGEMA_signal_14095), .Q (new_AGEMA_signal_14096) ) ;
    buf_clk new_AGEMA_reg_buffer_8248 ( .C (clk), .D (new_AGEMA_signal_14099), .Q (new_AGEMA_signal_14100) ) ;
    buf_clk new_AGEMA_reg_buffer_8252 ( .C (clk), .D (new_AGEMA_signal_14103), .Q (new_AGEMA_signal_14104) ) ;
    buf_clk new_AGEMA_reg_buffer_8256 ( .C (clk), .D (new_AGEMA_signal_14107), .Q (new_AGEMA_signal_14108) ) ;
    buf_clk new_AGEMA_reg_buffer_8260 ( .C (clk), .D (new_AGEMA_signal_14111), .Q (new_AGEMA_signal_14112) ) ;
    buf_clk new_AGEMA_reg_buffer_8264 ( .C (clk), .D (new_AGEMA_signal_14115), .Q (new_AGEMA_signal_14116) ) ;
    buf_clk new_AGEMA_reg_buffer_8268 ( .C (clk), .D (new_AGEMA_signal_14119), .Q (new_AGEMA_signal_14120) ) ;
    buf_clk new_AGEMA_reg_buffer_8272 ( .C (clk), .D (new_AGEMA_signal_14123), .Q (new_AGEMA_signal_14124) ) ;
    buf_clk new_AGEMA_reg_buffer_8276 ( .C (clk), .D (new_AGEMA_signal_14127), .Q (new_AGEMA_signal_14128) ) ;
    buf_clk new_AGEMA_reg_buffer_8280 ( .C (clk), .D (new_AGEMA_signal_14131), .Q (new_AGEMA_signal_14132) ) ;
    buf_clk new_AGEMA_reg_buffer_8284 ( .C (clk), .D (new_AGEMA_signal_14135), .Q (new_AGEMA_signal_14136) ) ;
    buf_clk new_AGEMA_reg_buffer_8288 ( .C (clk), .D (new_AGEMA_signal_14139), .Q (new_AGEMA_signal_14140) ) ;
    buf_clk new_AGEMA_reg_buffer_8292 ( .C (clk), .D (new_AGEMA_signal_14143), .Q (new_AGEMA_signal_14144) ) ;
    buf_clk new_AGEMA_reg_buffer_8296 ( .C (clk), .D (new_AGEMA_signal_14147), .Q (new_AGEMA_signal_14148) ) ;
    buf_clk new_AGEMA_reg_buffer_8300 ( .C (clk), .D (new_AGEMA_signal_14151), .Q (new_AGEMA_signal_14152) ) ;
    buf_clk new_AGEMA_reg_buffer_8304 ( .C (clk), .D (new_AGEMA_signal_14155), .Q (new_AGEMA_signal_14156) ) ;
    buf_clk new_AGEMA_reg_buffer_8308 ( .C (clk), .D (new_AGEMA_signal_14159), .Q (new_AGEMA_signal_14160) ) ;
    buf_clk new_AGEMA_reg_buffer_8312 ( .C (clk), .D (new_AGEMA_signal_14163), .Q (new_AGEMA_signal_14164) ) ;
    buf_clk new_AGEMA_reg_buffer_8316 ( .C (clk), .D (new_AGEMA_signal_14167), .Q (new_AGEMA_signal_14168) ) ;
    buf_clk new_AGEMA_reg_buffer_8320 ( .C (clk), .D (new_AGEMA_signal_14171), .Q (new_AGEMA_signal_14172) ) ;
    buf_clk new_AGEMA_reg_buffer_8324 ( .C (clk), .D (new_AGEMA_signal_14175), .Q (new_AGEMA_signal_14176) ) ;
    buf_clk new_AGEMA_reg_buffer_8328 ( .C (clk), .D (new_AGEMA_signal_14179), .Q (new_AGEMA_signal_14180) ) ;
    buf_clk new_AGEMA_reg_buffer_8332 ( .C (clk), .D (new_AGEMA_signal_14183), .Q (new_AGEMA_signal_14184) ) ;
    buf_clk new_AGEMA_reg_buffer_8336 ( .C (clk), .D (new_AGEMA_signal_14187), .Q (new_AGEMA_signal_14188) ) ;
    buf_clk new_AGEMA_reg_buffer_8340 ( .C (clk), .D (new_AGEMA_signal_14191), .Q (new_AGEMA_signal_14192) ) ;
    buf_clk new_AGEMA_reg_buffer_8344 ( .C (clk), .D (new_AGEMA_signal_14195), .Q (new_AGEMA_signal_14196) ) ;
    buf_clk new_AGEMA_reg_buffer_8348 ( .C (clk), .D (new_AGEMA_signal_14199), .Q (new_AGEMA_signal_14200) ) ;
    buf_clk new_AGEMA_reg_buffer_8352 ( .C (clk), .D (new_AGEMA_signal_14203), .Q (new_AGEMA_signal_14204) ) ;
    buf_clk new_AGEMA_reg_buffer_8356 ( .C (clk), .D (new_AGEMA_signal_14207), .Q (new_AGEMA_signal_14208) ) ;
    buf_clk new_AGEMA_reg_buffer_8360 ( .C (clk), .D (new_AGEMA_signal_14211), .Q (new_AGEMA_signal_14212) ) ;
    buf_clk new_AGEMA_reg_buffer_8364 ( .C (clk), .D (new_AGEMA_signal_14215), .Q (new_AGEMA_signal_14216) ) ;
    buf_clk new_AGEMA_reg_buffer_8368 ( .C (clk), .D (new_AGEMA_signal_14219), .Q (new_AGEMA_signal_14220) ) ;
    buf_clk new_AGEMA_reg_buffer_8372 ( .C (clk), .D (new_AGEMA_signal_14223), .Q (new_AGEMA_signal_14224) ) ;
    buf_clk new_AGEMA_reg_buffer_8376 ( .C (clk), .D (new_AGEMA_signal_14227), .Q (new_AGEMA_signal_14228) ) ;
    buf_clk new_AGEMA_reg_buffer_8380 ( .C (clk), .D (new_AGEMA_signal_14231), .Q (new_AGEMA_signal_14232) ) ;
    buf_clk new_AGEMA_reg_buffer_8384 ( .C (clk), .D (new_AGEMA_signal_14235), .Q (new_AGEMA_signal_14236) ) ;
    buf_clk new_AGEMA_reg_buffer_8388 ( .C (clk), .D (new_AGEMA_signal_14239), .Q (new_AGEMA_signal_14240) ) ;
    buf_clk new_AGEMA_reg_buffer_8392 ( .C (clk), .D (new_AGEMA_signal_14243), .Q (new_AGEMA_signal_14244) ) ;
    buf_clk new_AGEMA_reg_buffer_8396 ( .C (clk), .D (new_AGEMA_signal_14247), .Q (new_AGEMA_signal_14248) ) ;
    buf_clk new_AGEMA_reg_buffer_8400 ( .C (clk), .D (new_AGEMA_signal_14251), .Q (new_AGEMA_signal_14252) ) ;
    buf_clk new_AGEMA_reg_buffer_8404 ( .C (clk), .D (new_AGEMA_signal_14255), .Q (new_AGEMA_signal_14256) ) ;
    buf_clk new_AGEMA_reg_buffer_8408 ( .C (clk), .D (new_AGEMA_signal_14259), .Q (new_AGEMA_signal_14260) ) ;
    buf_clk new_AGEMA_reg_buffer_8412 ( .C (clk), .D (new_AGEMA_signal_14263), .Q (new_AGEMA_signal_14264) ) ;
    buf_clk new_AGEMA_reg_buffer_8416 ( .C (clk), .D (new_AGEMA_signal_14267), .Q (new_AGEMA_signal_14268) ) ;
    buf_clk new_AGEMA_reg_buffer_8420 ( .C (clk), .D (new_AGEMA_signal_14271), .Q (new_AGEMA_signal_14272) ) ;
    buf_clk new_AGEMA_reg_buffer_8424 ( .C (clk), .D (new_AGEMA_signal_14275), .Q (new_AGEMA_signal_14276) ) ;
    buf_clk new_AGEMA_reg_buffer_8428 ( .C (clk), .D (new_AGEMA_signal_14279), .Q (new_AGEMA_signal_14280) ) ;
    buf_clk new_AGEMA_reg_buffer_8432 ( .C (clk), .D (new_AGEMA_signal_14283), .Q (new_AGEMA_signal_14284) ) ;
    buf_clk new_AGEMA_reg_buffer_8436 ( .C (clk), .D (new_AGEMA_signal_14287), .Q (new_AGEMA_signal_14288) ) ;
    buf_clk new_AGEMA_reg_buffer_8440 ( .C (clk), .D (new_AGEMA_signal_14291), .Q (new_AGEMA_signal_14292) ) ;
    buf_clk new_AGEMA_reg_buffer_8444 ( .C (clk), .D (new_AGEMA_signal_14295), .Q (new_AGEMA_signal_14296) ) ;
    buf_clk new_AGEMA_reg_buffer_8448 ( .C (clk), .D (new_AGEMA_signal_14299), .Q (new_AGEMA_signal_14300) ) ;
    buf_clk new_AGEMA_reg_buffer_8452 ( .C (clk), .D (new_AGEMA_signal_14303), .Q (new_AGEMA_signal_14304) ) ;
    buf_clk new_AGEMA_reg_buffer_8456 ( .C (clk), .D (new_AGEMA_signal_14307), .Q (new_AGEMA_signal_14308) ) ;
    buf_clk new_AGEMA_reg_buffer_8460 ( .C (clk), .D (new_AGEMA_signal_14311), .Q (new_AGEMA_signal_14312) ) ;
    buf_clk new_AGEMA_reg_buffer_8464 ( .C (clk), .D (new_AGEMA_signal_14315), .Q (new_AGEMA_signal_14316) ) ;
    buf_clk new_AGEMA_reg_buffer_8468 ( .C (clk), .D (new_AGEMA_signal_14319), .Q (new_AGEMA_signal_14320) ) ;
    buf_clk new_AGEMA_reg_buffer_8472 ( .C (clk), .D (new_AGEMA_signal_14323), .Q (new_AGEMA_signal_14324) ) ;
    buf_clk new_AGEMA_reg_buffer_8476 ( .C (clk), .D (new_AGEMA_signal_14327), .Q (new_AGEMA_signal_14328) ) ;
    buf_clk new_AGEMA_reg_buffer_8480 ( .C (clk), .D (new_AGEMA_signal_14331), .Q (new_AGEMA_signal_14332) ) ;
    buf_clk new_AGEMA_reg_buffer_8484 ( .C (clk), .D (new_AGEMA_signal_14335), .Q (new_AGEMA_signal_14336) ) ;
    buf_clk new_AGEMA_reg_buffer_8488 ( .C (clk), .D (new_AGEMA_signal_14339), .Q (new_AGEMA_signal_14340) ) ;
    buf_clk new_AGEMA_reg_buffer_8492 ( .C (clk), .D (new_AGEMA_signal_14343), .Q (new_AGEMA_signal_14344) ) ;
    buf_clk new_AGEMA_reg_buffer_8496 ( .C (clk), .D (new_AGEMA_signal_14347), .Q (new_AGEMA_signal_14348) ) ;
    buf_clk new_AGEMA_reg_buffer_8500 ( .C (clk), .D (new_AGEMA_signal_14351), .Q (new_AGEMA_signal_14352) ) ;
    buf_clk new_AGEMA_reg_buffer_8504 ( .C (clk), .D (new_AGEMA_signal_14355), .Q (new_AGEMA_signal_14356) ) ;
    buf_clk new_AGEMA_reg_buffer_8508 ( .C (clk), .D (new_AGEMA_signal_14359), .Q (new_AGEMA_signal_14360) ) ;
    buf_clk new_AGEMA_reg_buffer_8512 ( .C (clk), .D (new_AGEMA_signal_14363), .Q (new_AGEMA_signal_14364) ) ;
    buf_clk new_AGEMA_reg_buffer_8516 ( .C (clk), .D (new_AGEMA_signal_14367), .Q (new_AGEMA_signal_14368) ) ;
    buf_clk new_AGEMA_reg_buffer_8520 ( .C (clk), .D (new_AGEMA_signal_14371), .Q (new_AGEMA_signal_14372) ) ;
    buf_clk new_AGEMA_reg_buffer_8524 ( .C (clk), .D (new_AGEMA_signal_14375), .Q (new_AGEMA_signal_14376) ) ;
    buf_clk new_AGEMA_reg_buffer_8528 ( .C (clk), .D (new_AGEMA_signal_14379), .Q (new_AGEMA_signal_14380) ) ;
    buf_clk new_AGEMA_reg_buffer_8532 ( .C (clk), .D (new_AGEMA_signal_14383), .Q (new_AGEMA_signal_14384) ) ;
    buf_clk new_AGEMA_reg_buffer_8536 ( .C (clk), .D (new_AGEMA_signal_14387), .Q (new_AGEMA_signal_14388) ) ;
    buf_clk new_AGEMA_reg_buffer_8540 ( .C (clk), .D (new_AGEMA_signal_14391), .Q (new_AGEMA_signal_14392) ) ;
    buf_clk new_AGEMA_reg_buffer_8544 ( .C (clk), .D (new_AGEMA_signal_14395), .Q (new_AGEMA_signal_14396) ) ;
    buf_clk new_AGEMA_reg_buffer_8548 ( .C (clk), .D (new_AGEMA_signal_14399), .Q (new_AGEMA_signal_14400) ) ;
    buf_clk new_AGEMA_reg_buffer_8552 ( .C (clk), .D (new_AGEMA_signal_14403), .Q (new_AGEMA_signal_14404) ) ;
    buf_clk new_AGEMA_reg_buffer_8556 ( .C (clk), .D (new_AGEMA_signal_14407), .Q (new_AGEMA_signal_14408) ) ;
    buf_clk new_AGEMA_reg_buffer_8560 ( .C (clk), .D (new_AGEMA_signal_14411), .Q (new_AGEMA_signal_14412) ) ;
    buf_clk new_AGEMA_reg_buffer_8564 ( .C (clk), .D (new_AGEMA_signal_14415), .Q (new_AGEMA_signal_14416) ) ;
    buf_clk new_AGEMA_reg_buffer_8568 ( .C (clk), .D (new_AGEMA_signal_14419), .Q (new_AGEMA_signal_14420) ) ;
    buf_clk new_AGEMA_reg_buffer_8572 ( .C (clk), .D (new_AGEMA_signal_14423), .Q (new_AGEMA_signal_14424) ) ;
    buf_clk new_AGEMA_reg_buffer_8576 ( .C (clk), .D (new_AGEMA_signal_14427), .Q (new_AGEMA_signal_14428) ) ;
    buf_clk new_AGEMA_reg_buffer_8580 ( .C (clk), .D (new_AGEMA_signal_14431), .Q (new_AGEMA_signal_14432) ) ;
    buf_clk new_AGEMA_reg_buffer_8584 ( .C (clk), .D (new_AGEMA_signal_14435), .Q (new_AGEMA_signal_14436) ) ;
    buf_clk new_AGEMA_reg_buffer_8588 ( .C (clk), .D (new_AGEMA_signal_14439), .Q (new_AGEMA_signal_14440) ) ;
    buf_clk new_AGEMA_reg_buffer_8592 ( .C (clk), .D (new_AGEMA_signal_14443), .Q (new_AGEMA_signal_14444) ) ;
    buf_clk new_AGEMA_reg_buffer_8596 ( .C (clk), .D (new_AGEMA_signal_14447), .Q (new_AGEMA_signal_14448) ) ;
    buf_clk new_AGEMA_reg_buffer_8600 ( .C (clk), .D (new_AGEMA_signal_14451), .Q (new_AGEMA_signal_14452) ) ;
    buf_clk new_AGEMA_reg_buffer_8604 ( .C (clk), .D (new_AGEMA_signal_14455), .Q (new_AGEMA_signal_14456) ) ;
    buf_clk new_AGEMA_reg_buffer_8608 ( .C (clk), .D (new_AGEMA_signal_14459), .Q (new_AGEMA_signal_14460) ) ;
    buf_clk new_AGEMA_reg_buffer_8612 ( .C (clk), .D (new_AGEMA_signal_14463), .Q (new_AGEMA_signal_14464) ) ;
    buf_clk new_AGEMA_reg_buffer_8616 ( .C (clk), .D (new_AGEMA_signal_14467), .Q (new_AGEMA_signal_14468) ) ;
    buf_clk new_AGEMA_reg_buffer_8620 ( .C (clk), .D (new_AGEMA_signal_14471), .Q (new_AGEMA_signal_14472) ) ;
    buf_clk new_AGEMA_reg_buffer_8624 ( .C (clk), .D (new_AGEMA_signal_14475), .Q (new_AGEMA_signal_14476) ) ;
    buf_clk new_AGEMA_reg_buffer_8628 ( .C (clk), .D (new_AGEMA_signal_14479), .Q (new_AGEMA_signal_14480) ) ;
    buf_clk new_AGEMA_reg_buffer_8632 ( .C (clk), .D (new_AGEMA_signal_14483), .Q (new_AGEMA_signal_14484) ) ;
    buf_clk new_AGEMA_reg_buffer_8636 ( .C (clk), .D (new_AGEMA_signal_14487), .Q (new_AGEMA_signal_14488) ) ;
    buf_clk new_AGEMA_reg_buffer_8640 ( .C (clk), .D (new_AGEMA_signal_14491), .Q (new_AGEMA_signal_14492) ) ;
    buf_clk new_AGEMA_reg_buffer_8644 ( .C (clk), .D (new_AGEMA_signal_14495), .Q (new_AGEMA_signal_14496) ) ;
    buf_clk new_AGEMA_reg_buffer_8648 ( .C (clk), .D (new_AGEMA_signal_14499), .Q (new_AGEMA_signal_14500) ) ;
    buf_clk new_AGEMA_reg_buffer_8652 ( .C (clk), .D (new_AGEMA_signal_14503), .Q (new_AGEMA_signal_14504) ) ;
    buf_clk new_AGEMA_reg_buffer_8656 ( .C (clk), .D (new_AGEMA_signal_14507), .Q (new_AGEMA_signal_14508) ) ;
    buf_clk new_AGEMA_reg_buffer_8660 ( .C (clk), .D (new_AGEMA_signal_14511), .Q (new_AGEMA_signal_14512) ) ;
    buf_clk new_AGEMA_reg_buffer_8664 ( .C (clk), .D (new_AGEMA_signal_14515), .Q (new_AGEMA_signal_14516) ) ;
    buf_clk new_AGEMA_reg_buffer_8668 ( .C (clk), .D (new_AGEMA_signal_14519), .Q (new_AGEMA_signal_14520) ) ;
    buf_clk new_AGEMA_reg_buffer_8672 ( .C (clk), .D (new_AGEMA_signal_14523), .Q (new_AGEMA_signal_14524) ) ;
    buf_clk new_AGEMA_reg_buffer_8676 ( .C (clk), .D (new_AGEMA_signal_14527), .Q (new_AGEMA_signal_14528) ) ;
    buf_clk new_AGEMA_reg_buffer_8680 ( .C (clk), .D (new_AGEMA_signal_14531), .Q (new_AGEMA_signal_14532) ) ;
    buf_clk new_AGEMA_reg_buffer_8684 ( .C (clk), .D (new_AGEMA_signal_14535), .Q (new_AGEMA_signal_14536) ) ;
    buf_clk new_AGEMA_reg_buffer_8688 ( .C (clk), .D (new_AGEMA_signal_14539), .Q (new_AGEMA_signal_14540) ) ;
    buf_clk new_AGEMA_reg_buffer_8692 ( .C (clk), .D (new_AGEMA_signal_14543), .Q (new_AGEMA_signal_14544) ) ;
    buf_clk new_AGEMA_reg_buffer_8696 ( .C (clk), .D (new_AGEMA_signal_14547), .Q (new_AGEMA_signal_14548) ) ;
    buf_clk new_AGEMA_reg_buffer_8700 ( .C (clk), .D (new_AGEMA_signal_14551), .Q (new_AGEMA_signal_14552) ) ;
    buf_clk new_AGEMA_reg_buffer_8704 ( .C (clk), .D (new_AGEMA_signal_14555), .Q (new_AGEMA_signal_14556) ) ;
    buf_clk new_AGEMA_reg_buffer_8708 ( .C (clk), .D (new_AGEMA_signal_14559), .Q (new_AGEMA_signal_14560) ) ;
    buf_clk new_AGEMA_reg_buffer_8712 ( .C (clk), .D (new_AGEMA_signal_14563), .Q (new_AGEMA_signal_14564) ) ;
    buf_clk new_AGEMA_reg_buffer_8716 ( .C (clk), .D (new_AGEMA_signal_14567), .Q (new_AGEMA_signal_14568) ) ;
    buf_clk new_AGEMA_reg_buffer_8720 ( .C (clk), .D (new_AGEMA_signal_14571), .Q (new_AGEMA_signal_14572) ) ;
    buf_clk new_AGEMA_reg_buffer_8724 ( .C (clk), .D (new_AGEMA_signal_14575), .Q (new_AGEMA_signal_14576) ) ;
    buf_clk new_AGEMA_reg_buffer_8728 ( .C (clk), .D (new_AGEMA_signal_14579), .Q (new_AGEMA_signal_14580) ) ;
    buf_clk new_AGEMA_reg_buffer_8732 ( .C (clk), .D (new_AGEMA_signal_14583), .Q (new_AGEMA_signal_14584) ) ;
    buf_clk new_AGEMA_reg_buffer_8736 ( .C (clk), .D (new_AGEMA_signal_14587), .Q (new_AGEMA_signal_14588) ) ;
    buf_clk new_AGEMA_reg_buffer_8740 ( .C (clk), .D (new_AGEMA_signal_14591), .Q (new_AGEMA_signal_14592) ) ;
    buf_clk new_AGEMA_reg_buffer_8744 ( .C (clk), .D (new_AGEMA_signal_14595), .Q (new_AGEMA_signal_14596) ) ;
    buf_clk new_AGEMA_reg_buffer_8748 ( .C (clk), .D (new_AGEMA_signal_14599), .Q (new_AGEMA_signal_14600) ) ;
    buf_clk new_AGEMA_reg_buffer_8752 ( .C (clk), .D (new_AGEMA_signal_14603), .Q (new_AGEMA_signal_14604) ) ;
    buf_clk new_AGEMA_reg_buffer_8756 ( .C (clk), .D (new_AGEMA_signal_14607), .Q (new_AGEMA_signal_14608) ) ;
    buf_clk new_AGEMA_reg_buffer_8760 ( .C (clk), .D (new_AGEMA_signal_14611), .Q (new_AGEMA_signal_14612) ) ;
    buf_clk new_AGEMA_reg_buffer_8764 ( .C (clk), .D (new_AGEMA_signal_14615), .Q (new_AGEMA_signal_14616) ) ;
    buf_clk new_AGEMA_reg_buffer_8768 ( .C (clk), .D (new_AGEMA_signal_14619), .Q (new_AGEMA_signal_14620) ) ;
    buf_clk new_AGEMA_reg_buffer_8772 ( .C (clk), .D (new_AGEMA_signal_14623), .Q (new_AGEMA_signal_14624) ) ;
    buf_clk new_AGEMA_reg_buffer_8776 ( .C (clk), .D (new_AGEMA_signal_14627), .Q (new_AGEMA_signal_14628) ) ;
    buf_clk new_AGEMA_reg_buffer_8780 ( .C (clk), .D (new_AGEMA_signal_14631), .Q (new_AGEMA_signal_14632) ) ;
    buf_clk new_AGEMA_reg_buffer_8784 ( .C (clk), .D (new_AGEMA_signal_14635), .Q (new_AGEMA_signal_14636) ) ;
    buf_clk new_AGEMA_reg_buffer_8788 ( .C (clk), .D (new_AGEMA_signal_14639), .Q (new_AGEMA_signal_14640) ) ;
    buf_clk new_AGEMA_reg_buffer_8792 ( .C (clk), .D (new_AGEMA_signal_14643), .Q (new_AGEMA_signal_14644) ) ;
    buf_clk new_AGEMA_reg_buffer_8796 ( .C (clk), .D (new_AGEMA_signal_14647), .Q (new_AGEMA_signal_14648) ) ;
    buf_clk new_AGEMA_reg_buffer_8800 ( .C (clk), .D (new_AGEMA_signal_14651), .Q (new_AGEMA_signal_14652) ) ;
    buf_clk new_AGEMA_reg_buffer_8804 ( .C (clk), .D (new_AGEMA_signal_14655), .Q (new_AGEMA_signal_14656) ) ;
    buf_clk new_AGEMA_reg_buffer_8808 ( .C (clk), .D (new_AGEMA_signal_14659), .Q (new_AGEMA_signal_14660) ) ;
    buf_clk new_AGEMA_reg_buffer_8812 ( .C (clk), .D (new_AGEMA_signal_14663), .Q (new_AGEMA_signal_14664) ) ;
    buf_clk new_AGEMA_reg_buffer_8816 ( .C (clk), .D (new_AGEMA_signal_14667), .Q (new_AGEMA_signal_14668) ) ;
    buf_clk new_AGEMA_reg_buffer_8820 ( .C (clk), .D (new_AGEMA_signal_14671), .Q (new_AGEMA_signal_14672) ) ;
    buf_clk new_AGEMA_reg_buffer_8824 ( .C (clk), .D (new_AGEMA_signal_14675), .Q (new_AGEMA_signal_14676) ) ;
    buf_clk new_AGEMA_reg_buffer_8828 ( .C (clk), .D (new_AGEMA_signal_14679), .Q (new_AGEMA_signal_14680) ) ;
    buf_clk new_AGEMA_reg_buffer_8832 ( .C (clk), .D (new_AGEMA_signal_14683), .Q (new_AGEMA_signal_14684) ) ;
    buf_clk new_AGEMA_reg_buffer_8836 ( .C (clk), .D (new_AGEMA_signal_14687), .Q (new_AGEMA_signal_14688) ) ;
    buf_clk new_AGEMA_reg_buffer_8840 ( .C (clk), .D (new_AGEMA_signal_14691), .Q (new_AGEMA_signal_14692) ) ;
    buf_clk new_AGEMA_reg_buffer_8844 ( .C (clk), .D (new_AGEMA_signal_14695), .Q (new_AGEMA_signal_14696) ) ;
    buf_clk new_AGEMA_reg_buffer_8848 ( .C (clk), .D (new_AGEMA_signal_14699), .Q (new_AGEMA_signal_14700) ) ;
    buf_clk new_AGEMA_reg_buffer_8852 ( .C (clk), .D (new_AGEMA_signal_14703), .Q (new_AGEMA_signal_14704) ) ;
    buf_clk new_AGEMA_reg_buffer_8856 ( .C (clk), .D (new_AGEMA_signal_14707), .Q (new_AGEMA_signal_14708) ) ;
    buf_clk new_AGEMA_reg_buffer_8860 ( .C (clk), .D (new_AGEMA_signal_14711), .Q (new_AGEMA_signal_14712) ) ;
    buf_clk new_AGEMA_reg_buffer_8864 ( .C (clk), .D (new_AGEMA_signal_14715), .Q (new_AGEMA_signal_14716) ) ;
    buf_clk new_AGEMA_reg_buffer_8868 ( .C (clk), .D (new_AGEMA_signal_14719), .Q (new_AGEMA_signal_14720) ) ;
    buf_clk new_AGEMA_reg_buffer_8872 ( .C (clk), .D (new_AGEMA_signal_14723), .Q (new_AGEMA_signal_14724) ) ;
    buf_clk new_AGEMA_reg_buffer_8876 ( .C (clk), .D (new_AGEMA_signal_14727), .Q (new_AGEMA_signal_14728) ) ;
    buf_clk new_AGEMA_reg_buffer_8880 ( .C (clk), .D (new_AGEMA_signal_14731), .Q (new_AGEMA_signal_14732) ) ;
    buf_clk new_AGEMA_reg_buffer_8884 ( .C (clk), .D (new_AGEMA_signal_14735), .Q (new_AGEMA_signal_14736) ) ;
    buf_clk new_AGEMA_reg_buffer_8888 ( .C (clk), .D (new_AGEMA_signal_14739), .Q (new_AGEMA_signal_14740) ) ;
    buf_clk new_AGEMA_reg_buffer_8892 ( .C (clk), .D (new_AGEMA_signal_14743), .Q (new_AGEMA_signal_14744) ) ;
    buf_clk new_AGEMA_reg_buffer_8896 ( .C (clk), .D (new_AGEMA_signal_14747), .Q (new_AGEMA_signal_14748) ) ;
    buf_clk new_AGEMA_reg_buffer_8900 ( .C (clk), .D (new_AGEMA_signal_14751), .Q (new_AGEMA_signal_14752) ) ;
    buf_clk new_AGEMA_reg_buffer_8904 ( .C (clk), .D (new_AGEMA_signal_14755), .Q (new_AGEMA_signal_14756) ) ;
    buf_clk new_AGEMA_reg_buffer_8908 ( .C (clk), .D (new_AGEMA_signal_14759), .Q (new_AGEMA_signal_14760) ) ;
    buf_clk new_AGEMA_reg_buffer_8912 ( .C (clk), .D (new_AGEMA_signal_14763), .Q (new_AGEMA_signal_14764) ) ;
    buf_clk new_AGEMA_reg_buffer_8916 ( .C (clk), .D (new_AGEMA_signal_14767), .Q (new_AGEMA_signal_14768) ) ;
    buf_clk new_AGEMA_reg_buffer_8920 ( .C (clk), .D (new_AGEMA_signal_14771), .Q (new_AGEMA_signal_14772) ) ;
    buf_clk new_AGEMA_reg_buffer_8924 ( .C (clk), .D (new_AGEMA_signal_14775), .Q (new_AGEMA_signal_14776) ) ;
    buf_clk new_AGEMA_reg_buffer_8928 ( .C (clk), .D (new_AGEMA_signal_14779), .Q (new_AGEMA_signal_14780) ) ;
    buf_clk new_AGEMA_reg_buffer_8932 ( .C (clk), .D (new_AGEMA_signal_14783), .Q (new_AGEMA_signal_14784) ) ;
    buf_clk new_AGEMA_reg_buffer_8936 ( .C (clk), .D (new_AGEMA_signal_14787), .Q (new_AGEMA_signal_14788) ) ;
    buf_clk new_AGEMA_reg_buffer_8940 ( .C (clk), .D (new_AGEMA_signal_14791), .Q (new_AGEMA_signal_14792) ) ;
    buf_clk new_AGEMA_reg_buffer_8944 ( .C (clk), .D (new_AGEMA_signal_14795), .Q (new_AGEMA_signal_14796) ) ;
    buf_clk new_AGEMA_reg_buffer_8948 ( .C (clk), .D (new_AGEMA_signal_14799), .Q (new_AGEMA_signal_14800) ) ;
    buf_clk new_AGEMA_reg_buffer_8952 ( .C (clk), .D (new_AGEMA_signal_14803), .Q (new_AGEMA_signal_14804) ) ;
    buf_clk new_AGEMA_reg_buffer_8956 ( .C (clk), .D (new_AGEMA_signal_14807), .Q (new_AGEMA_signal_14808) ) ;
    buf_clk new_AGEMA_reg_buffer_8960 ( .C (clk), .D (new_AGEMA_signal_14811), .Q (new_AGEMA_signal_14812) ) ;
    buf_clk new_AGEMA_reg_buffer_8964 ( .C (clk), .D (new_AGEMA_signal_14815), .Q (new_AGEMA_signal_14816) ) ;
    buf_clk new_AGEMA_reg_buffer_8968 ( .C (clk), .D (new_AGEMA_signal_14819), .Q (new_AGEMA_signal_14820) ) ;
    buf_clk new_AGEMA_reg_buffer_8972 ( .C (clk), .D (new_AGEMA_signal_14823), .Q (new_AGEMA_signal_14824) ) ;
    buf_clk new_AGEMA_reg_buffer_8976 ( .C (clk), .D (new_AGEMA_signal_14827), .Q (new_AGEMA_signal_14828) ) ;
    buf_clk new_AGEMA_reg_buffer_8980 ( .C (clk), .D (new_AGEMA_signal_14831), .Q (new_AGEMA_signal_14832) ) ;
    buf_clk new_AGEMA_reg_buffer_8984 ( .C (clk), .D (new_AGEMA_signal_14835), .Q (new_AGEMA_signal_14836) ) ;
    buf_clk new_AGEMA_reg_buffer_8988 ( .C (clk), .D (new_AGEMA_signal_14839), .Q (new_AGEMA_signal_14840) ) ;
    buf_clk new_AGEMA_reg_buffer_8992 ( .C (clk), .D (new_AGEMA_signal_14843), .Q (new_AGEMA_signal_14844) ) ;
    buf_clk new_AGEMA_reg_buffer_8996 ( .C (clk), .D (new_AGEMA_signal_14847), .Q (new_AGEMA_signal_14848) ) ;
    buf_clk new_AGEMA_reg_buffer_9000 ( .C (clk), .D (new_AGEMA_signal_14851), .Q (new_AGEMA_signal_14852) ) ;
    buf_clk new_AGEMA_reg_buffer_9004 ( .C (clk), .D (new_AGEMA_signal_14855), .Q (new_AGEMA_signal_14856) ) ;
    buf_clk new_AGEMA_reg_buffer_9008 ( .C (clk), .D (new_AGEMA_signal_14859), .Q (new_AGEMA_signal_14860) ) ;
    buf_clk new_AGEMA_reg_buffer_9012 ( .C (clk), .D (new_AGEMA_signal_14863), .Q (new_AGEMA_signal_14864) ) ;
    buf_clk new_AGEMA_reg_buffer_9016 ( .C (clk), .D (new_AGEMA_signal_14867), .Q (new_AGEMA_signal_14868) ) ;
    buf_clk new_AGEMA_reg_buffer_9020 ( .C (clk), .D (new_AGEMA_signal_14871), .Q (new_AGEMA_signal_14872) ) ;
    buf_clk new_AGEMA_reg_buffer_9024 ( .C (clk), .D (new_AGEMA_signal_14875), .Q (new_AGEMA_signal_14876) ) ;
    buf_clk new_AGEMA_reg_buffer_9028 ( .C (clk), .D (new_AGEMA_signal_14879), .Q (new_AGEMA_signal_14880) ) ;
    buf_clk new_AGEMA_reg_buffer_9032 ( .C (clk), .D (new_AGEMA_signal_14883), .Q (new_AGEMA_signal_14884) ) ;
    buf_clk new_AGEMA_reg_buffer_9036 ( .C (clk), .D (new_AGEMA_signal_14887), .Q (new_AGEMA_signal_14888) ) ;
    buf_clk new_AGEMA_reg_buffer_9040 ( .C (clk), .D (new_AGEMA_signal_14891), .Q (new_AGEMA_signal_14892) ) ;
    buf_clk new_AGEMA_reg_buffer_9044 ( .C (clk), .D (new_AGEMA_signal_14895), .Q (new_AGEMA_signal_14896) ) ;
    buf_clk new_AGEMA_reg_buffer_9048 ( .C (clk), .D (new_AGEMA_signal_14899), .Q (new_AGEMA_signal_14900) ) ;
    buf_clk new_AGEMA_reg_buffer_9052 ( .C (clk), .D (new_AGEMA_signal_14903), .Q (new_AGEMA_signal_14904) ) ;
    buf_clk new_AGEMA_reg_buffer_9056 ( .C (clk), .D (new_AGEMA_signal_14907), .Q (new_AGEMA_signal_14908) ) ;
    buf_clk new_AGEMA_reg_buffer_9060 ( .C (clk), .D (new_AGEMA_signal_14911), .Q (new_AGEMA_signal_14912) ) ;
    buf_clk new_AGEMA_reg_buffer_9064 ( .C (clk), .D (new_AGEMA_signal_14915), .Q (new_AGEMA_signal_14916) ) ;
    buf_clk new_AGEMA_reg_buffer_9068 ( .C (clk), .D (new_AGEMA_signal_14919), .Q (new_AGEMA_signal_14920) ) ;
    buf_clk new_AGEMA_reg_buffer_9072 ( .C (clk), .D (new_AGEMA_signal_14923), .Q (new_AGEMA_signal_14924) ) ;
    buf_clk new_AGEMA_reg_buffer_9076 ( .C (clk), .D (new_AGEMA_signal_14927), .Q (new_AGEMA_signal_14928) ) ;
    buf_clk new_AGEMA_reg_buffer_9080 ( .C (clk), .D (new_AGEMA_signal_14931), .Q (new_AGEMA_signal_14932) ) ;
    buf_clk new_AGEMA_reg_buffer_9084 ( .C (clk), .D (new_AGEMA_signal_14935), .Q (new_AGEMA_signal_14936) ) ;
    buf_clk new_AGEMA_reg_buffer_9088 ( .C (clk), .D (new_AGEMA_signal_14939), .Q (new_AGEMA_signal_14940) ) ;
    buf_clk new_AGEMA_reg_buffer_9092 ( .C (clk), .D (new_AGEMA_signal_14943), .Q (new_AGEMA_signal_14944) ) ;
    buf_clk new_AGEMA_reg_buffer_9096 ( .C (clk), .D (new_AGEMA_signal_14947), .Q (new_AGEMA_signal_14948) ) ;
    buf_clk new_AGEMA_reg_buffer_9100 ( .C (clk), .D (new_AGEMA_signal_14951), .Q (new_AGEMA_signal_14952) ) ;
    buf_clk new_AGEMA_reg_buffer_9104 ( .C (clk), .D (new_AGEMA_signal_14955), .Q (new_AGEMA_signal_14956) ) ;
    buf_clk new_AGEMA_reg_buffer_9108 ( .C (clk), .D (new_AGEMA_signal_14959), .Q (new_AGEMA_signal_14960) ) ;
    buf_clk new_AGEMA_reg_buffer_9112 ( .C (clk), .D (new_AGEMA_signal_14963), .Q (new_AGEMA_signal_14964) ) ;
    buf_clk new_AGEMA_reg_buffer_9116 ( .C (clk), .D (new_AGEMA_signal_14967), .Q (new_AGEMA_signal_14968) ) ;
    buf_clk new_AGEMA_reg_buffer_9120 ( .C (clk), .D (new_AGEMA_signal_14971), .Q (new_AGEMA_signal_14972) ) ;
    buf_clk new_AGEMA_reg_buffer_9124 ( .C (clk), .D (new_AGEMA_signal_14975), .Q (new_AGEMA_signal_14976) ) ;
    buf_clk new_AGEMA_reg_buffer_9128 ( .C (clk), .D (new_AGEMA_signal_14979), .Q (new_AGEMA_signal_14980) ) ;
    buf_clk new_AGEMA_reg_buffer_9132 ( .C (clk), .D (new_AGEMA_signal_14983), .Q (new_AGEMA_signal_14984) ) ;
    buf_clk new_AGEMA_reg_buffer_9136 ( .C (clk), .D (new_AGEMA_signal_14987), .Q (new_AGEMA_signal_14988) ) ;
    buf_clk new_AGEMA_reg_buffer_9140 ( .C (clk), .D (new_AGEMA_signal_14991), .Q (new_AGEMA_signal_14992) ) ;
    buf_clk new_AGEMA_reg_buffer_9144 ( .C (clk), .D (new_AGEMA_signal_14995), .Q (new_AGEMA_signal_14996) ) ;
    buf_clk new_AGEMA_reg_buffer_9148 ( .C (clk), .D (new_AGEMA_signal_14999), .Q (new_AGEMA_signal_15000) ) ;
    buf_clk new_AGEMA_reg_buffer_9152 ( .C (clk), .D (new_AGEMA_signal_15003), .Q (new_AGEMA_signal_15004) ) ;
    buf_clk new_AGEMA_reg_buffer_9156 ( .C (clk), .D (new_AGEMA_signal_15007), .Q (new_AGEMA_signal_15008) ) ;
    buf_clk new_AGEMA_reg_buffer_9160 ( .C (clk), .D (new_AGEMA_signal_15011), .Q (new_AGEMA_signal_15012) ) ;
    buf_clk new_AGEMA_reg_buffer_9164 ( .C (clk), .D (new_AGEMA_signal_15015), .Q (new_AGEMA_signal_15016) ) ;
    buf_clk new_AGEMA_reg_buffer_9168 ( .C (clk), .D (new_AGEMA_signal_15019), .Q (new_AGEMA_signal_15020) ) ;
    buf_clk new_AGEMA_reg_buffer_9172 ( .C (clk), .D (new_AGEMA_signal_15023), .Q (new_AGEMA_signal_15024) ) ;
    buf_clk new_AGEMA_reg_buffer_9176 ( .C (clk), .D (new_AGEMA_signal_15027), .Q (new_AGEMA_signal_15028) ) ;
    buf_clk new_AGEMA_reg_buffer_9180 ( .C (clk), .D (new_AGEMA_signal_15031), .Q (new_AGEMA_signal_15032) ) ;
    buf_clk new_AGEMA_reg_buffer_9184 ( .C (clk), .D (new_AGEMA_signal_15035), .Q (new_AGEMA_signal_15036) ) ;
    buf_clk new_AGEMA_reg_buffer_9188 ( .C (clk), .D (new_AGEMA_signal_15039), .Q (new_AGEMA_signal_15040) ) ;
    buf_clk new_AGEMA_reg_buffer_9192 ( .C (clk), .D (new_AGEMA_signal_15043), .Q (new_AGEMA_signal_15044) ) ;
    buf_clk new_AGEMA_reg_buffer_9196 ( .C (clk), .D (new_AGEMA_signal_15047), .Q (new_AGEMA_signal_15048) ) ;
    buf_clk new_AGEMA_reg_buffer_9200 ( .C (clk), .D (new_AGEMA_signal_15051), .Q (new_AGEMA_signal_15052) ) ;
    buf_clk new_AGEMA_reg_buffer_9204 ( .C (clk), .D (new_AGEMA_signal_15055), .Q (new_AGEMA_signal_15056) ) ;
    buf_clk new_AGEMA_reg_buffer_9208 ( .C (clk), .D (new_AGEMA_signal_15059), .Q (new_AGEMA_signal_15060) ) ;
    buf_clk new_AGEMA_reg_buffer_9212 ( .C (clk), .D (new_AGEMA_signal_15063), .Q (new_AGEMA_signal_15064) ) ;
    buf_clk new_AGEMA_reg_buffer_9216 ( .C (clk), .D (new_AGEMA_signal_15067), .Q (new_AGEMA_signal_15068) ) ;
    buf_clk new_AGEMA_reg_buffer_9220 ( .C (clk), .D (new_AGEMA_signal_15071), .Q (new_AGEMA_signal_15072) ) ;
    buf_clk new_AGEMA_reg_buffer_9224 ( .C (clk), .D (new_AGEMA_signal_15075), .Q (new_AGEMA_signal_15076) ) ;
    buf_clk new_AGEMA_reg_buffer_9228 ( .C (clk), .D (new_AGEMA_signal_15079), .Q (new_AGEMA_signal_15080) ) ;
    buf_clk new_AGEMA_reg_buffer_9232 ( .C (clk), .D (new_AGEMA_signal_15083), .Q (new_AGEMA_signal_15084) ) ;
    buf_clk new_AGEMA_reg_buffer_9236 ( .C (clk), .D (new_AGEMA_signal_15087), .Q (new_AGEMA_signal_15088) ) ;
    buf_clk new_AGEMA_reg_buffer_9240 ( .C (clk), .D (new_AGEMA_signal_15091), .Q (new_AGEMA_signal_15092) ) ;
    buf_clk new_AGEMA_reg_buffer_9244 ( .C (clk), .D (new_AGEMA_signal_15095), .Q (new_AGEMA_signal_15096) ) ;
    buf_clk new_AGEMA_reg_buffer_9248 ( .C (clk), .D (new_AGEMA_signal_15099), .Q (new_AGEMA_signal_15100) ) ;
    buf_clk new_AGEMA_reg_buffer_9252 ( .C (clk), .D (new_AGEMA_signal_15103), .Q (new_AGEMA_signal_15104) ) ;
    buf_clk new_AGEMA_reg_buffer_9256 ( .C (clk), .D (new_AGEMA_signal_15107), .Q (new_AGEMA_signal_15108) ) ;
    buf_clk new_AGEMA_reg_buffer_9260 ( .C (clk), .D (new_AGEMA_signal_15111), .Q (new_AGEMA_signal_15112) ) ;
    buf_clk new_AGEMA_reg_buffer_9264 ( .C (clk), .D (new_AGEMA_signal_15115), .Q (new_AGEMA_signal_15116) ) ;
    buf_clk new_AGEMA_reg_buffer_9268 ( .C (clk), .D (new_AGEMA_signal_15119), .Q (new_AGEMA_signal_15120) ) ;
    buf_clk new_AGEMA_reg_buffer_9272 ( .C (clk), .D (new_AGEMA_signal_15123), .Q (new_AGEMA_signal_15124) ) ;
    buf_clk new_AGEMA_reg_buffer_9276 ( .C (clk), .D (new_AGEMA_signal_15127), .Q (new_AGEMA_signal_15128) ) ;
    buf_clk new_AGEMA_reg_buffer_9280 ( .C (clk), .D (new_AGEMA_signal_15131), .Q (new_AGEMA_signal_15132) ) ;
    buf_clk new_AGEMA_reg_buffer_9284 ( .C (clk), .D (new_AGEMA_signal_15135), .Q (new_AGEMA_signal_15136) ) ;
    buf_clk new_AGEMA_reg_buffer_9288 ( .C (clk), .D (new_AGEMA_signal_15139), .Q (new_AGEMA_signal_15140) ) ;
    buf_clk new_AGEMA_reg_buffer_9292 ( .C (clk), .D (new_AGEMA_signal_15143), .Q (new_AGEMA_signal_15144) ) ;
    buf_clk new_AGEMA_reg_buffer_9296 ( .C (clk), .D (new_AGEMA_signal_15147), .Q (new_AGEMA_signal_15148) ) ;
    buf_clk new_AGEMA_reg_buffer_9300 ( .C (clk), .D (new_AGEMA_signal_15151), .Q (new_AGEMA_signal_15152) ) ;
    buf_clk new_AGEMA_reg_buffer_9304 ( .C (clk), .D (new_AGEMA_signal_15155), .Q (new_AGEMA_signal_15156) ) ;
    buf_clk new_AGEMA_reg_buffer_9308 ( .C (clk), .D (new_AGEMA_signal_15159), .Q (new_AGEMA_signal_15160) ) ;
    buf_clk new_AGEMA_reg_buffer_9312 ( .C (clk), .D (new_AGEMA_signal_15163), .Q (new_AGEMA_signal_15164) ) ;
    buf_clk new_AGEMA_reg_buffer_9316 ( .C (clk), .D (new_AGEMA_signal_15167), .Q (new_AGEMA_signal_15168) ) ;
    buf_clk new_AGEMA_reg_buffer_9320 ( .C (clk), .D (new_AGEMA_signal_15171), .Q (new_AGEMA_signal_15172) ) ;
    buf_clk new_AGEMA_reg_buffer_9324 ( .C (clk), .D (new_AGEMA_signal_15175), .Q (new_AGEMA_signal_15176) ) ;
    buf_clk new_AGEMA_reg_buffer_9328 ( .C (clk), .D (new_AGEMA_signal_15179), .Q (new_AGEMA_signal_15180) ) ;
    buf_clk new_AGEMA_reg_buffer_9332 ( .C (clk), .D (new_AGEMA_signal_15183), .Q (new_AGEMA_signal_15184) ) ;
    buf_clk new_AGEMA_reg_buffer_9336 ( .C (clk), .D (new_AGEMA_signal_15187), .Q (new_AGEMA_signal_15188) ) ;
    buf_clk new_AGEMA_reg_buffer_9340 ( .C (clk), .D (new_AGEMA_signal_15191), .Q (new_AGEMA_signal_15192) ) ;
    buf_clk new_AGEMA_reg_buffer_9344 ( .C (clk), .D (new_AGEMA_signal_15195), .Q (new_AGEMA_signal_15196) ) ;
    buf_clk new_AGEMA_reg_buffer_9348 ( .C (clk), .D (new_AGEMA_signal_15199), .Q (new_AGEMA_signal_15200) ) ;
    buf_clk new_AGEMA_reg_buffer_9352 ( .C (clk), .D (new_AGEMA_signal_15203), .Q (new_AGEMA_signal_15204) ) ;
    buf_clk new_AGEMA_reg_buffer_9356 ( .C (clk), .D (new_AGEMA_signal_15207), .Q (new_AGEMA_signal_15208) ) ;
    buf_clk new_AGEMA_reg_buffer_9360 ( .C (clk), .D (new_AGEMA_signal_15211), .Q (new_AGEMA_signal_15212) ) ;
    buf_clk new_AGEMA_reg_buffer_9364 ( .C (clk), .D (new_AGEMA_signal_15215), .Q (new_AGEMA_signal_15216) ) ;
    buf_clk new_AGEMA_reg_buffer_9368 ( .C (clk), .D (new_AGEMA_signal_15219), .Q (new_AGEMA_signal_15220) ) ;
    buf_clk new_AGEMA_reg_buffer_9372 ( .C (clk), .D (new_AGEMA_signal_15223), .Q (new_AGEMA_signal_15224) ) ;
    buf_clk new_AGEMA_reg_buffer_9376 ( .C (clk), .D (new_AGEMA_signal_15227), .Q (new_AGEMA_signal_15228) ) ;
    buf_clk new_AGEMA_reg_buffer_9380 ( .C (clk), .D (new_AGEMA_signal_15231), .Q (new_AGEMA_signal_15232) ) ;
    buf_clk new_AGEMA_reg_buffer_9384 ( .C (clk), .D (new_AGEMA_signal_15235), .Q (new_AGEMA_signal_15236) ) ;
    buf_clk new_AGEMA_reg_buffer_9388 ( .C (clk), .D (new_AGEMA_signal_15239), .Q (new_AGEMA_signal_15240) ) ;
    buf_clk new_AGEMA_reg_buffer_9392 ( .C (clk), .D (new_AGEMA_signal_15243), .Q (new_AGEMA_signal_15244) ) ;
    buf_clk new_AGEMA_reg_buffer_9396 ( .C (clk), .D (new_AGEMA_signal_15247), .Q (new_AGEMA_signal_15248) ) ;
    buf_clk new_AGEMA_reg_buffer_9400 ( .C (clk), .D (new_AGEMA_signal_15251), .Q (new_AGEMA_signal_15252) ) ;
    buf_clk new_AGEMA_reg_buffer_9404 ( .C (clk), .D (new_AGEMA_signal_15255), .Q (new_AGEMA_signal_15256) ) ;
    buf_clk new_AGEMA_reg_buffer_9408 ( .C (clk), .D (new_AGEMA_signal_15259), .Q (new_AGEMA_signal_15260) ) ;
    buf_clk new_AGEMA_reg_buffer_9412 ( .C (clk), .D (new_AGEMA_signal_15263), .Q (new_AGEMA_signal_15264) ) ;
    buf_clk new_AGEMA_reg_buffer_9416 ( .C (clk), .D (new_AGEMA_signal_15267), .Q (new_AGEMA_signal_15268) ) ;
    buf_clk new_AGEMA_reg_buffer_9420 ( .C (clk), .D (new_AGEMA_signal_15271), .Q (new_AGEMA_signal_15272) ) ;
    buf_clk new_AGEMA_reg_buffer_9424 ( .C (clk), .D (new_AGEMA_signal_15275), .Q (new_AGEMA_signal_15276) ) ;
    buf_clk new_AGEMA_reg_buffer_9428 ( .C (clk), .D (new_AGEMA_signal_15279), .Q (new_AGEMA_signal_15280) ) ;
    buf_clk new_AGEMA_reg_buffer_9432 ( .C (clk), .D (new_AGEMA_signal_15283), .Q (new_AGEMA_signal_15284) ) ;
    buf_clk new_AGEMA_reg_buffer_9436 ( .C (clk), .D (new_AGEMA_signal_15287), .Q (new_AGEMA_signal_15288) ) ;
    buf_clk new_AGEMA_reg_buffer_9440 ( .C (clk), .D (new_AGEMA_signal_15291), .Q (new_AGEMA_signal_15292) ) ;
    buf_clk new_AGEMA_reg_buffer_9444 ( .C (clk), .D (new_AGEMA_signal_15295), .Q (new_AGEMA_signal_15296) ) ;
    buf_clk new_AGEMA_reg_buffer_9448 ( .C (clk), .D (new_AGEMA_signal_15299), .Q (new_AGEMA_signal_15300) ) ;
    buf_clk new_AGEMA_reg_buffer_9452 ( .C (clk), .D (new_AGEMA_signal_15303), .Q (new_AGEMA_signal_15304) ) ;
    buf_clk new_AGEMA_reg_buffer_9456 ( .C (clk), .D (new_AGEMA_signal_15307), .Q (new_AGEMA_signal_15308) ) ;
    buf_clk new_AGEMA_reg_buffer_9460 ( .C (clk), .D (new_AGEMA_signal_15311), .Q (new_AGEMA_signal_15312) ) ;
    buf_clk new_AGEMA_reg_buffer_9464 ( .C (clk), .D (new_AGEMA_signal_15315), .Q (new_AGEMA_signal_15316) ) ;
    buf_clk new_AGEMA_reg_buffer_9468 ( .C (clk), .D (new_AGEMA_signal_15319), .Q (new_AGEMA_signal_15320) ) ;
    buf_clk new_AGEMA_reg_buffer_9472 ( .C (clk), .D (new_AGEMA_signal_15323), .Q (new_AGEMA_signal_15324) ) ;
    buf_clk new_AGEMA_reg_buffer_9476 ( .C (clk), .D (new_AGEMA_signal_15327), .Q (new_AGEMA_signal_15328) ) ;
    buf_clk new_AGEMA_reg_buffer_9480 ( .C (clk), .D (new_AGEMA_signal_15331), .Q (new_AGEMA_signal_15332) ) ;
    buf_clk new_AGEMA_reg_buffer_9484 ( .C (clk), .D (new_AGEMA_signal_15335), .Q (new_AGEMA_signal_15336) ) ;
    buf_clk new_AGEMA_reg_buffer_9488 ( .C (clk), .D (new_AGEMA_signal_15339), .Q (new_AGEMA_signal_15340) ) ;
    buf_clk new_AGEMA_reg_buffer_9492 ( .C (clk), .D (new_AGEMA_signal_15343), .Q (new_AGEMA_signal_15344) ) ;
    buf_clk new_AGEMA_reg_buffer_9496 ( .C (clk), .D (new_AGEMA_signal_15347), .Q (new_AGEMA_signal_15348) ) ;
    buf_clk new_AGEMA_reg_buffer_9500 ( .C (clk), .D (new_AGEMA_signal_15351), .Q (new_AGEMA_signal_15352) ) ;
    buf_clk new_AGEMA_reg_buffer_9504 ( .C (clk), .D (new_AGEMA_signal_15355), .Q (new_AGEMA_signal_15356) ) ;
    buf_clk new_AGEMA_reg_buffer_9508 ( .C (clk), .D (new_AGEMA_signal_15359), .Q (new_AGEMA_signal_15360) ) ;
    buf_clk new_AGEMA_reg_buffer_9512 ( .C (clk), .D (new_AGEMA_signal_15363), .Q (new_AGEMA_signal_15364) ) ;
    buf_clk new_AGEMA_reg_buffer_9516 ( .C (clk), .D (new_AGEMA_signal_15367), .Q (new_AGEMA_signal_15368) ) ;
    buf_clk new_AGEMA_reg_buffer_9520 ( .C (clk), .D (new_AGEMA_signal_15371), .Q (new_AGEMA_signal_15372) ) ;
    buf_clk new_AGEMA_reg_buffer_9524 ( .C (clk), .D (new_AGEMA_signal_15375), .Q (new_AGEMA_signal_15376) ) ;
    buf_clk new_AGEMA_reg_buffer_9528 ( .C (clk), .D (new_AGEMA_signal_15379), .Q (new_AGEMA_signal_15380) ) ;
    buf_clk new_AGEMA_reg_buffer_9532 ( .C (clk), .D (new_AGEMA_signal_15383), .Q (new_AGEMA_signal_15384) ) ;
    buf_clk new_AGEMA_reg_buffer_9536 ( .C (clk), .D (new_AGEMA_signal_15387), .Q (new_AGEMA_signal_15388) ) ;
    buf_clk new_AGEMA_reg_buffer_9540 ( .C (clk), .D (new_AGEMA_signal_15391), .Q (new_AGEMA_signal_15392) ) ;
    buf_clk new_AGEMA_reg_buffer_9544 ( .C (clk), .D (new_AGEMA_signal_15395), .Q (new_AGEMA_signal_15396) ) ;
    buf_clk new_AGEMA_reg_buffer_9548 ( .C (clk), .D (new_AGEMA_signal_15399), .Q (new_AGEMA_signal_15400) ) ;
    buf_clk new_AGEMA_reg_buffer_9552 ( .C (clk), .D (new_AGEMA_signal_15403), .Q (new_AGEMA_signal_15404) ) ;
    buf_clk new_AGEMA_reg_buffer_9964 ( .C (clk), .D (new_AGEMA_signal_15815), .Q (new_AGEMA_signal_15816) ) ;
    buf_clk new_AGEMA_reg_buffer_9968 ( .C (clk), .D (new_AGEMA_signal_15819), .Q (new_AGEMA_signal_15820) ) ;
    buf_clk new_AGEMA_reg_buffer_9972 ( .C (clk), .D (new_AGEMA_signal_15823), .Q (new_AGEMA_signal_15824) ) ;
    buf_clk new_AGEMA_reg_buffer_9976 ( .C (clk), .D (new_AGEMA_signal_15827), .Q (new_AGEMA_signal_15828) ) ;

    /* register cells */
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_0_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8432, RoundReg_Inst_ff_SDE_0_next_state}), .Q ({new_AGEMA_signal_4549, RoundInput[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_1_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8606, RoundReg_Inst_ff_SDE_1_next_state}), .Q ({new_AGEMA_signal_4666, RoundInput[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_2_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8434, RoundReg_Inst_ff_SDE_2_next_state}), .Q ({new_AGEMA_signal_4699, RoundInput[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_3_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8608, RoundReg_Inst_ff_SDE_3_next_state}), .Q ({new_AGEMA_signal_4732, RoundInput[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_4_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8610, RoundReg_Inst_ff_SDE_4_next_state}), .Q ({new_AGEMA_signal_4765, RoundInput[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_5_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8436, RoundReg_Inst_ff_SDE_5_next_state}), .Q ({new_AGEMA_signal_4798, RoundInput[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_6_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8438, RoundReg_Inst_ff_SDE_6_next_state}), .Q ({new_AGEMA_signal_4831, RoundInput[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_7_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8440, RoundReg_Inst_ff_SDE_7_next_state}), .Q ({new_AGEMA_signal_4864, RoundInput[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_8_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8442, RoundReg_Inst_ff_SDE_8_next_state}), .Q ({new_AGEMA_signal_4897, RoundInput[8]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_9_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8612, RoundReg_Inst_ff_SDE_9_next_state}), .Q ({new_AGEMA_signal_4930, RoundInput[9]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_10_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8444, RoundReg_Inst_ff_SDE_10_next_state}), .Q ({new_AGEMA_signal_4582, RoundInput[10]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_11_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8614, RoundReg_Inst_ff_SDE_11_next_state}), .Q ({new_AGEMA_signal_4615, RoundInput[11]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_12_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8616, RoundReg_Inst_ff_SDE_12_next_state}), .Q ({new_AGEMA_signal_4642, RoundInput[12]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_13_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8446, RoundReg_Inst_ff_SDE_13_next_state}), .Q ({new_AGEMA_signal_4645, RoundInput[13]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_14_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8448, RoundReg_Inst_ff_SDE_14_next_state}), .Q ({new_AGEMA_signal_4648, RoundInput[14]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_15_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8450, RoundReg_Inst_ff_SDE_15_next_state}), .Q ({new_AGEMA_signal_4651, RoundInput[15]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_16_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8452, RoundReg_Inst_ff_SDE_16_next_state}), .Q ({new_AGEMA_signal_4654, RoundInput[16]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_17_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8618, RoundReg_Inst_ff_SDE_17_next_state}), .Q ({new_AGEMA_signal_4657, RoundInput[17]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_18_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8454, RoundReg_Inst_ff_SDE_18_next_state}), .Q ({new_AGEMA_signal_4660, RoundInput[18]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_19_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8620, RoundReg_Inst_ff_SDE_19_next_state}), .Q ({new_AGEMA_signal_4663, RoundInput[19]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_20_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8622, RoundReg_Inst_ff_SDE_20_next_state}), .Q ({new_AGEMA_signal_4669, RoundInput[20]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_21_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8456, RoundReg_Inst_ff_SDE_21_next_state}), .Q ({new_AGEMA_signal_4672, RoundInput[21]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_22_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8458, RoundReg_Inst_ff_SDE_22_next_state}), .Q ({new_AGEMA_signal_4675, RoundInput[22]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_23_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8460, RoundReg_Inst_ff_SDE_23_next_state}), .Q ({new_AGEMA_signal_4678, RoundInput[23]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_24_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8462, RoundReg_Inst_ff_SDE_24_next_state}), .Q ({new_AGEMA_signal_4681, RoundInput[24]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_25_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8624, RoundReg_Inst_ff_SDE_25_next_state}), .Q ({new_AGEMA_signal_4684, RoundInput[25]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_26_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8464, RoundReg_Inst_ff_SDE_26_next_state}), .Q ({new_AGEMA_signal_4687, RoundInput[26]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_27_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8626, RoundReg_Inst_ff_SDE_27_next_state}), .Q ({new_AGEMA_signal_4690, RoundInput[27]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_28_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8628, RoundReg_Inst_ff_SDE_28_next_state}), .Q ({new_AGEMA_signal_4693, RoundInput[28]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_29_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8466, RoundReg_Inst_ff_SDE_29_next_state}), .Q ({new_AGEMA_signal_4696, RoundInput[29]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_30_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8468, RoundReg_Inst_ff_SDE_30_next_state}), .Q ({new_AGEMA_signal_4702, RoundInput[30]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_31_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8470, RoundReg_Inst_ff_SDE_31_next_state}), .Q ({new_AGEMA_signal_4705, RoundInput[31]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_32_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8472, RoundReg_Inst_ff_SDE_32_next_state}), .Q ({new_AGEMA_signal_4708, RoundInput[32]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_33_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8630, RoundReg_Inst_ff_SDE_33_next_state}), .Q ({new_AGEMA_signal_4711, RoundInput[33]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_34_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8474, RoundReg_Inst_ff_SDE_34_next_state}), .Q ({new_AGEMA_signal_4714, RoundInput[34]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_35_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8632, RoundReg_Inst_ff_SDE_35_next_state}), .Q ({new_AGEMA_signal_4717, RoundInput[35]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_36_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8634, RoundReg_Inst_ff_SDE_36_next_state}), .Q ({new_AGEMA_signal_4720, RoundInput[36]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_37_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8476, RoundReg_Inst_ff_SDE_37_next_state}), .Q ({new_AGEMA_signal_4723, RoundInput[37]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_38_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8478, RoundReg_Inst_ff_SDE_38_next_state}), .Q ({new_AGEMA_signal_4726, RoundInput[38]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_39_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8480, RoundReg_Inst_ff_SDE_39_next_state}), .Q ({new_AGEMA_signal_4729, RoundInput[39]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_40_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8482, RoundReg_Inst_ff_SDE_40_next_state}), .Q ({new_AGEMA_signal_4735, RoundInput[40]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_41_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8636, RoundReg_Inst_ff_SDE_41_next_state}), .Q ({new_AGEMA_signal_4738, RoundInput[41]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_42_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8484, RoundReg_Inst_ff_SDE_42_next_state}), .Q ({new_AGEMA_signal_4741, RoundInput[42]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_43_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8638, RoundReg_Inst_ff_SDE_43_next_state}), .Q ({new_AGEMA_signal_4744, RoundInput[43]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_44_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8640, RoundReg_Inst_ff_SDE_44_next_state}), .Q ({new_AGEMA_signal_4747, RoundInput[44]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_45_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8486, RoundReg_Inst_ff_SDE_45_next_state}), .Q ({new_AGEMA_signal_4750, RoundInput[45]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_46_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8488, RoundReg_Inst_ff_SDE_46_next_state}), .Q ({new_AGEMA_signal_4753, RoundInput[46]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_47_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8490, RoundReg_Inst_ff_SDE_47_next_state}), .Q ({new_AGEMA_signal_4756, RoundInput[47]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_48_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8492, RoundReg_Inst_ff_SDE_48_next_state}), .Q ({new_AGEMA_signal_4759, RoundInput[48]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_49_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8642, RoundReg_Inst_ff_SDE_49_next_state}), .Q ({new_AGEMA_signal_4762, RoundInput[49]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_50_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8494, RoundReg_Inst_ff_SDE_50_next_state}), .Q ({new_AGEMA_signal_4768, RoundInput[50]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_51_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8644, RoundReg_Inst_ff_SDE_51_next_state}), .Q ({new_AGEMA_signal_4771, RoundInput[51]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_52_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8646, RoundReg_Inst_ff_SDE_52_next_state}), .Q ({new_AGEMA_signal_4774, RoundInput[52]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_53_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8496, RoundReg_Inst_ff_SDE_53_next_state}), .Q ({new_AGEMA_signal_4777, RoundInput[53]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_54_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8498, RoundReg_Inst_ff_SDE_54_next_state}), .Q ({new_AGEMA_signal_4780, RoundInput[54]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_55_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8500, RoundReg_Inst_ff_SDE_55_next_state}), .Q ({new_AGEMA_signal_4783, RoundInput[55]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_56_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8502, RoundReg_Inst_ff_SDE_56_next_state}), .Q ({new_AGEMA_signal_4786, RoundInput[56]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_57_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8648, RoundReg_Inst_ff_SDE_57_next_state}), .Q ({new_AGEMA_signal_4789, RoundInput[57]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_58_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8504, RoundReg_Inst_ff_SDE_58_next_state}), .Q ({new_AGEMA_signal_4792, RoundInput[58]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_59_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8650, RoundReg_Inst_ff_SDE_59_next_state}), .Q ({new_AGEMA_signal_4795, RoundInput[59]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_60_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8652, RoundReg_Inst_ff_SDE_60_next_state}), .Q ({new_AGEMA_signal_4801, RoundInput[60]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_61_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8506, RoundReg_Inst_ff_SDE_61_next_state}), .Q ({new_AGEMA_signal_4804, RoundInput[61]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_62_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8508, RoundReg_Inst_ff_SDE_62_next_state}), .Q ({new_AGEMA_signal_4807, RoundInput[62]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_63_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8510, RoundReg_Inst_ff_SDE_63_next_state}), .Q ({new_AGEMA_signal_4810, RoundInput[63]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_64_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8512, RoundReg_Inst_ff_SDE_64_next_state}), .Q ({new_AGEMA_signal_4813, RoundInput[64]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_65_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8654, RoundReg_Inst_ff_SDE_65_next_state}), .Q ({new_AGEMA_signal_4816, RoundInput[65]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_66_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8514, RoundReg_Inst_ff_SDE_66_next_state}), .Q ({new_AGEMA_signal_4819, RoundInput[66]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_67_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8656, RoundReg_Inst_ff_SDE_67_next_state}), .Q ({new_AGEMA_signal_4822, RoundInput[67]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_68_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8658, RoundReg_Inst_ff_SDE_68_next_state}), .Q ({new_AGEMA_signal_4825, RoundInput[68]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_69_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8516, RoundReg_Inst_ff_SDE_69_next_state}), .Q ({new_AGEMA_signal_4828, RoundInput[69]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_70_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8518, RoundReg_Inst_ff_SDE_70_next_state}), .Q ({new_AGEMA_signal_4834, RoundInput[70]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_71_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8520, RoundReg_Inst_ff_SDE_71_next_state}), .Q ({new_AGEMA_signal_4837, RoundInput[71]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_72_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8522, RoundReg_Inst_ff_SDE_72_next_state}), .Q ({new_AGEMA_signal_4840, RoundInput[72]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_73_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8660, RoundReg_Inst_ff_SDE_73_next_state}), .Q ({new_AGEMA_signal_4843, RoundInput[73]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_74_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8524, RoundReg_Inst_ff_SDE_74_next_state}), .Q ({new_AGEMA_signal_4846, RoundInput[74]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_75_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8662, RoundReg_Inst_ff_SDE_75_next_state}), .Q ({new_AGEMA_signal_4849, RoundInput[75]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_76_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8664, RoundReg_Inst_ff_SDE_76_next_state}), .Q ({new_AGEMA_signal_4852, RoundInput[76]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_77_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8526, RoundReg_Inst_ff_SDE_77_next_state}), .Q ({new_AGEMA_signal_4855, RoundInput[77]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_78_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8528, RoundReg_Inst_ff_SDE_78_next_state}), .Q ({new_AGEMA_signal_4858, RoundInput[78]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_79_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8530, RoundReg_Inst_ff_SDE_79_next_state}), .Q ({new_AGEMA_signal_4861, RoundInput[79]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_80_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8532, RoundReg_Inst_ff_SDE_80_next_state}), .Q ({new_AGEMA_signal_4867, RoundInput[80]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_81_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8666, RoundReg_Inst_ff_SDE_81_next_state}), .Q ({new_AGEMA_signal_4870, RoundInput[81]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_82_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8534, RoundReg_Inst_ff_SDE_82_next_state}), .Q ({new_AGEMA_signal_4873, RoundInput[82]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_83_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8668, RoundReg_Inst_ff_SDE_83_next_state}), .Q ({new_AGEMA_signal_4876, RoundInput[83]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_84_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8670, RoundReg_Inst_ff_SDE_84_next_state}), .Q ({new_AGEMA_signal_4879, RoundInput[84]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_85_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8536, RoundReg_Inst_ff_SDE_85_next_state}), .Q ({new_AGEMA_signal_4882, RoundInput[85]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_86_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8538, RoundReg_Inst_ff_SDE_86_next_state}), .Q ({new_AGEMA_signal_4885, RoundInput[86]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_87_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8540, RoundReg_Inst_ff_SDE_87_next_state}), .Q ({new_AGEMA_signal_4888, RoundInput[87]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_88_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8542, RoundReg_Inst_ff_SDE_88_next_state}), .Q ({new_AGEMA_signal_4891, RoundInput[88]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_89_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8672, RoundReg_Inst_ff_SDE_89_next_state}), .Q ({new_AGEMA_signal_4894, RoundInput[89]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_90_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8544, RoundReg_Inst_ff_SDE_90_next_state}), .Q ({new_AGEMA_signal_4900, RoundInput[90]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_91_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8674, RoundReg_Inst_ff_SDE_91_next_state}), .Q ({new_AGEMA_signal_4903, RoundInput[91]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_92_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8676, RoundReg_Inst_ff_SDE_92_next_state}), .Q ({new_AGEMA_signal_4906, RoundInput[92]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_93_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8546, RoundReg_Inst_ff_SDE_93_next_state}), .Q ({new_AGEMA_signal_4909, RoundInput[93]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_94_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8548, RoundReg_Inst_ff_SDE_94_next_state}), .Q ({new_AGEMA_signal_4912, RoundInput[94]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_95_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8550, RoundReg_Inst_ff_SDE_95_next_state}), .Q ({new_AGEMA_signal_4915, RoundInput[95]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_96_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8552, RoundReg_Inst_ff_SDE_96_next_state}), .Q ({new_AGEMA_signal_4918, RoundInput[96]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_97_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8678, RoundReg_Inst_ff_SDE_97_next_state}), .Q ({new_AGEMA_signal_4921, RoundInput[97]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_98_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8554, RoundReg_Inst_ff_SDE_98_next_state}), .Q ({new_AGEMA_signal_4924, RoundInput[98]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_99_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8680, RoundReg_Inst_ff_SDE_99_next_state}), .Q ({new_AGEMA_signal_4927, RoundInput[99]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_100_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8682, RoundReg_Inst_ff_SDE_100_next_state}), .Q ({new_AGEMA_signal_4552, RoundInput[100]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_101_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8556, RoundReg_Inst_ff_SDE_101_next_state}), .Q ({new_AGEMA_signal_4555, RoundInput[101]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_102_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8558, RoundReg_Inst_ff_SDE_102_next_state}), .Q ({new_AGEMA_signal_4558, RoundInput[102]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_103_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8560, RoundReg_Inst_ff_SDE_103_next_state}), .Q ({new_AGEMA_signal_4561, RoundInput[103]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_104_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8562, RoundReg_Inst_ff_SDE_104_next_state}), .Q ({new_AGEMA_signal_4564, RoundInput[104]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_105_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8684, RoundReg_Inst_ff_SDE_105_next_state}), .Q ({new_AGEMA_signal_4567, RoundInput[105]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_106_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8564, RoundReg_Inst_ff_SDE_106_next_state}), .Q ({new_AGEMA_signal_4570, RoundInput[106]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_107_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8686, RoundReg_Inst_ff_SDE_107_next_state}), .Q ({new_AGEMA_signal_4573, RoundInput[107]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_108_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8688, RoundReg_Inst_ff_SDE_108_next_state}), .Q ({new_AGEMA_signal_4576, RoundInput[108]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_109_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8566, RoundReg_Inst_ff_SDE_109_next_state}), .Q ({new_AGEMA_signal_4579, RoundInput[109]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_110_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8568, RoundReg_Inst_ff_SDE_110_next_state}), .Q ({new_AGEMA_signal_4585, RoundInput[110]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_111_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8570, RoundReg_Inst_ff_SDE_111_next_state}), .Q ({new_AGEMA_signal_4588, RoundInput[111]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_112_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8572, RoundReg_Inst_ff_SDE_112_next_state}), .Q ({new_AGEMA_signal_4591, RoundInput[112]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_113_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8690, RoundReg_Inst_ff_SDE_113_next_state}), .Q ({new_AGEMA_signal_4594, RoundInput[113]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_114_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8574, RoundReg_Inst_ff_SDE_114_next_state}), .Q ({new_AGEMA_signal_4597, RoundInput[114]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_115_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8692, RoundReg_Inst_ff_SDE_115_next_state}), .Q ({new_AGEMA_signal_4600, RoundInput[115]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_116_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8694, RoundReg_Inst_ff_SDE_116_next_state}), .Q ({new_AGEMA_signal_4603, RoundInput[116]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_117_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8576, RoundReg_Inst_ff_SDE_117_next_state}), .Q ({new_AGEMA_signal_4606, RoundInput[117]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_118_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8578, RoundReg_Inst_ff_SDE_118_next_state}), .Q ({new_AGEMA_signal_4609, RoundInput[118]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_119_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8580, RoundReg_Inst_ff_SDE_119_next_state}), .Q ({new_AGEMA_signal_4612, RoundInput[119]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_120_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8582, RoundReg_Inst_ff_SDE_120_next_state}), .Q ({new_AGEMA_signal_4618, RoundInput[120]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_121_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8696, RoundReg_Inst_ff_SDE_121_next_state}), .Q ({new_AGEMA_signal_4621, RoundInput[121]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_122_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8584, RoundReg_Inst_ff_SDE_122_next_state}), .Q ({new_AGEMA_signal_4624, RoundInput[122]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_123_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8698, RoundReg_Inst_ff_SDE_123_next_state}), .Q ({new_AGEMA_signal_4627, RoundInput[123]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_124_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8700, RoundReg_Inst_ff_SDE_124_next_state}), .Q ({new_AGEMA_signal_4630, RoundInput[124]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_125_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8586, RoundReg_Inst_ff_SDE_125_next_state}), .Q ({new_AGEMA_signal_4633, RoundInput[125]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_126_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8588, RoundReg_Inst_ff_SDE_126_next_state}), .Q ({new_AGEMA_signal_4636, RoundInput[126]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_127_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8590, RoundReg_Inst_ff_SDE_127_next_state}), .Q ({new_AGEMA_signal_4639, RoundInput[127]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_0_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8098, KeyReg_Inst_ff_SDE_0_next_state}), .Q ({new_AGEMA_signal_4550, RoundKey[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_1_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8319, KeyReg_Inst_ff_SDE_1_next_state}), .Q ({new_AGEMA_signal_4667, RoundKey[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_2_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8321, KeyReg_Inst_ff_SDE_2_next_state}), .Q ({new_AGEMA_signal_4700, RoundKey[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_3_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8323, KeyReg_Inst_ff_SDE_3_next_state}), .Q ({new_AGEMA_signal_4733, RoundKey[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_4_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8325, KeyReg_Inst_ff_SDE_4_next_state}), .Q ({new_AGEMA_signal_4766, RoundKey[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_5_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8327, KeyReg_Inst_ff_SDE_5_next_state}), .Q ({new_AGEMA_signal_4799, RoundKey[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_6_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8329, KeyReg_Inst_ff_SDE_6_next_state}), .Q ({new_AGEMA_signal_4832, RoundKey[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_7_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8331, KeyReg_Inst_ff_SDE_7_next_state}), .Q ({new_AGEMA_signal_4865, RoundKey[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_8_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8100, KeyReg_Inst_ff_SDE_8_next_state}), .Q ({new_AGEMA_signal_4898, RoundKey[8]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_9_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8333, KeyReg_Inst_ff_SDE_9_next_state}), .Q ({new_AGEMA_signal_4931, RoundKey[9]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_10_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8335, KeyReg_Inst_ff_SDE_10_next_state}), .Q ({new_AGEMA_signal_4583, RoundKey[10]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_11_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8337, KeyReg_Inst_ff_SDE_11_next_state}), .Q ({new_AGEMA_signal_4616, RoundKey[11]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_12_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8339, KeyReg_Inst_ff_SDE_12_next_state}), .Q ({new_AGEMA_signal_4643, RoundKey[12]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_13_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8341, KeyReg_Inst_ff_SDE_13_next_state}), .Q ({new_AGEMA_signal_4646, RoundKey[13]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_14_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8343, KeyReg_Inst_ff_SDE_14_next_state}), .Q ({new_AGEMA_signal_4649, RoundKey[14]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_15_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8345, KeyReg_Inst_ff_SDE_15_next_state}), .Q ({new_AGEMA_signal_4652, RoundKey[15]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_16_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8102, KeyReg_Inst_ff_SDE_16_next_state}), .Q ({new_AGEMA_signal_4655, RoundKey[16]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_17_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8347, KeyReg_Inst_ff_SDE_17_next_state}), .Q ({new_AGEMA_signal_4658, RoundKey[17]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_18_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8349, KeyReg_Inst_ff_SDE_18_next_state}), .Q ({new_AGEMA_signal_4661, RoundKey[18]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_19_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8351, KeyReg_Inst_ff_SDE_19_next_state}), .Q ({new_AGEMA_signal_4664, RoundKey[19]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_20_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8353, KeyReg_Inst_ff_SDE_20_next_state}), .Q ({new_AGEMA_signal_4670, RoundKey[20]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_21_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8355, KeyReg_Inst_ff_SDE_21_next_state}), .Q ({new_AGEMA_signal_4673, RoundKey[21]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_22_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8357, KeyReg_Inst_ff_SDE_22_next_state}), .Q ({new_AGEMA_signal_4676, RoundKey[22]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_23_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8359, KeyReg_Inst_ff_SDE_23_next_state}), .Q ({new_AGEMA_signal_4679, RoundKey[23]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_24_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8361, KeyReg_Inst_ff_SDE_24_next_state}), .Q ({new_AGEMA_signal_4682, RoundKey[24]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_25_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8592, KeyReg_Inst_ff_SDE_25_next_state}), .Q ({new_AGEMA_signal_4685, RoundKey[25]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_26_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8594, KeyReg_Inst_ff_SDE_26_next_state}), .Q ({new_AGEMA_signal_4688, RoundKey[26]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_27_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8596, KeyReg_Inst_ff_SDE_27_next_state}), .Q ({new_AGEMA_signal_4691, RoundKey[27]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_28_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8598, KeyReg_Inst_ff_SDE_28_next_state}), .Q ({new_AGEMA_signal_4694, RoundKey[28]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_29_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8600, KeyReg_Inst_ff_SDE_29_next_state}), .Q ({new_AGEMA_signal_4697, RoundKey[29]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_30_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8602, KeyReg_Inst_ff_SDE_30_next_state}), .Q ({new_AGEMA_signal_4703, RoundKey[30]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_31_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8604, KeyReg_Inst_ff_SDE_31_next_state}), .Q ({new_AGEMA_signal_4706, RoundKey[31]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_32_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7874, KeyReg_Inst_ff_SDE_32_next_state}), .Q ({new_AGEMA_signal_4709, RoundKey[32]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_33_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8104, KeyReg_Inst_ff_SDE_33_next_state}), .Q ({new_AGEMA_signal_4712, RoundKey[33]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_34_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8106, KeyReg_Inst_ff_SDE_34_next_state}), .Q ({new_AGEMA_signal_4715, RoundKey[34]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_35_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8108, KeyReg_Inst_ff_SDE_35_next_state}), .Q ({new_AGEMA_signal_4718, RoundKey[35]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_36_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8110, KeyReg_Inst_ff_SDE_36_next_state}), .Q ({new_AGEMA_signal_4721, RoundKey[36]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_37_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8112, KeyReg_Inst_ff_SDE_37_next_state}), .Q ({new_AGEMA_signal_4724, RoundKey[37]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_38_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8114, KeyReg_Inst_ff_SDE_38_next_state}), .Q ({new_AGEMA_signal_4727, RoundKey[38]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_39_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8116, KeyReg_Inst_ff_SDE_39_next_state}), .Q ({new_AGEMA_signal_4730, RoundKey[39]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_40_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7876, KeyReg_Inst_ff_SDE_40_next_state}), .Q ({new_AGEMA_signal_4736, RoundKey[40]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_41_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8118, KeyReg_Inst_ff_SDE_41_next_state}), .Q ({new_AGEMA_signal_4739, RoundKey[41]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_42_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8120, KeyReg_Inst_ff_SDE_42_next_state}), .Q ({new_AGEMA_signal_4742, RoundKey[42]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_43_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8122, KeyReg_Inst_ff_SDE_43_next_state}), .Q ({new_AGEMA_signal_4745, RoundKey[43]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_44_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8124, KeyReg_Inst_ff_SDE_44_next_state}), .Q ({new_AGEMA_signal_4748, RoundKey[44]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_45_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8126, KeyReg_Inst_ff_SDE_45_next_state}), .Q ({new_AGEMA_signal_4751, RoundKey[45]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_46_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8128, KeyReg_Inst_ff_SDE_46_next_state}), .Q ({new_AGEMA_signal_4754, RoundKey[46]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_47_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8130, KeyReg_Inst_ff_SDE_47_next_state}), .Q ({new_AGEMA_signal_4757, RoundKey[47]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_48_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7878, KeyReg_Inst_ff_SDE_48_next_state}), .Q ({new_AGEMA_signal_4760, RoundKey[48]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_49_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8132, KeyReg_Inst_ff_SDE_49_next_state}), .Q ({new_AGEMA_signal_4763, RoundKey[49]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_50_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8134, KeyReg_Inst_ff_SDE_50_next_state}), .Q ({new_AGEMA_signal_4769, RoundKey[50]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_51_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8136, KeyReg_Inst_ff_SDE_51_next_state}), .Q ({new_AGEMA_signal_4772, RoundKey[51]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_52_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8138, KeyReg_Inst_ff_SDE_52_next_state}), .Q ({new_AGEMA_signal_4775, RoundKey[52]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_53_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8140, KeyReg_Inst_ff_SDE_53_next_state}), .Q ({new_AGEMA_signal_4778, RoundKey[53]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_54_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8142, KeyReg_Inst_ff_SDE_54_next_state}), .Q ({new_AGEMA_signal_4781, RoundKey[54]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_55_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8144, KeyReg_Inst_ff_SDE_55_next_state}), .Q ({new_AGEMA_signal_4784, RoundKey[55]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_56_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8146, KeyReg_Inst_ff_SDE_56_next_state}), .Q ({new_AGEMA_signal_4787, RoundKey[56]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_57_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8363, KeyReg_Inst_ff_SDE_57_next_state}), .Q ({new_AGEMA_signal_4790, RoundKey[57]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_58_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8365, KeyReg_Inst_ff_SDE_58_next_state}), .Q ({new_AGEMA_signal_4793, RoundKey[58]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_59_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8367, KeyReg_Inst_ff_SDE_59_next_state}), .Q ({new_AGEMA_signal_4796, RoundKey[59]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_60_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8369, KeyReg_Inst_ff_SDE_60_next_state}), .Q ({new_AGEMA_signal_4802, RoundKey[60]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_61_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8371, KeyReg_Inst_ff_SDE_61_next_state}), .Q ({new_AGEMA_signal_4805, RoundKey[61]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_62_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8373, KeyReg_Inst_ff_SDE_62_next_state}), .Q ({new_AGEMA_signal_4808, RoundKey[62]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_63_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8375, KeyReg_Inst_ff_SDE_63_next_state}), .Q ({new_AGEMA_signal_4811, RoundKey[63]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_64_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7664, KeyReg_Inst_ff_SDE_64_next_state}), .Q ({new_AGEMA_signal_4814, RoundKey[64]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_65_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7880, KeyReg_Inst_ff_SDE_65_next_state}), .Q ({new_AGEMA_signal_4817, RoundKey[65]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_66_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7882, KeyReg_Inst_ff_SDE_66_next_state}), .Q ({new_AGEMA_signal_4820, RoundKey[66]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_67_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7884, KeyReg_Inst_ff_SDE_67_next_state}), .Q ({new_AGEMA_signal_4823, RoundKey[67]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_68_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7886, KeyReg_Inst_ff_SDE_68_next_state}), .Q ({new_AGEMA_signal_4826, RoundKey[68]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_69_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7888, KeyReg_Inst_ff_SDE_69_next_state}), .Q ({new_AGEMA_signal_4829, RoundKey[69]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_70_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7890, KeyReg_Inst_ff_SDE_70_next_state}), .Q ({new_AGEMA_signal_4835, RoundKey[70]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_71_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7892, KeyReg_Inst_ff_SDE_71_next_state}), .Q ({new_AGEMA_signal_4838, RoundKey[71]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_72_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7666, KeyReg_Inst_ff_SDE_72_next_state}), .Q ({new_AGEMA_signal_4841, RoundKey[72]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_73_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7894, KeyReg_Inst_ff_SDE_73_next_state}), .Q ({new_AGEMA_signal_4844, RoundKey[73]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_74_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7896, KeyReg_Inst_ff_SDE_74_next_state}), .Q ({new_AGEMA_signal_4847, RoundKey[74]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_75_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7898, KeyReg_Inst_ff_SDE_75_next_state}), .Q ({new_AGEMA_signal_4850, RoundKey[75]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_76_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7900, KeyReg_Inst_ff_SDE_76_next_state}), .Q ({new_AGEMA_signal_4853, RoundKey[76]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_77_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7902, KeyReg_Inst_ff_SDE_77_next_state}), .Q ({new_AGEMA_signal_4856, RoundKey[77]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_78_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7904, KeyReg_Inst_ff_SDE_78_next_state}), .Q ({new_AGEMA_signal_4859, RoundKey[78]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_79_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7906, KeyReg_Inst_ff_SDE_79_next_state}), .Q ({new_AGEMA_signal_4862, RoundKey[79]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_80_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7668, KeyReg_Inst_ff_SDE_80_next_state}), .Q ({new_AGEMA_signal_4868, RoundKey[80]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_81_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7908, KeyReg_Inst_ff_SDE_81_next_state}), .Q ({new_AGEMA_signal_4871, RoundKey[81]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_82_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7910, KeyReg_Inst_ff_SDE_82_next_state}), .Q ({new_AGEMA_signal_4874, RoundKey[82]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_83_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7912, KeyReg_Inst_ff_SDE_83_next_state}), .Q ({new_AGEMA_signal_4877, RoundKey[83]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_84_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7914, KeyReg_Inst_ff_SDE_84_next_state}), .Q ({new_AGEMA_signal_4880, RoundKey[84]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_85_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7916, KeyReg_Inst_ff_SDE_85_next_state}), .Q ({new_AGEMA_signal_4883, RoundKey[85]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_86_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7918, KeyReg_Inst_ff_SDE_86_next_state}), .Q ({new_AGEMA_signal_4886, RoundKey[86]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_87_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7920, KeyReg_Inst_ff_SDE_87_next_state}), .Q ({new_AGEMA_signal_4889, RoundKey[87]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_88_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7922, KeyReg_Inst_ff_SDE_88_next_state}), .Q ({new_AGEMA_signal_4892, RoundKey[88]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_89_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8148, KeyReg_Inst_ff_SDE_89_next_state}), .Q ({new_AGEMA_signal_4895, RoundKey[89]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_90_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8150, KeyReg_Inst_ff_SDE_90_next_state}), .Q ({new_AGEMA_signal_4901, RoundKey[90]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_91_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8152, KeyReg_Inst_ff_SDE_91_next_state}), .Q ({new_AGEMA_signal_4904, RoundKey[91]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_92_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8154, KeyReg_Inst_ff_SDE_92_next_state}), .Q ({new_AGEMA_signal_4907, RoundKey[92]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_93_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8156, KeyReg_Inst_ff_SDE_93_next_state}), .Q ({new_AGEMA_signal_4910, RoundKey[93]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_94_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8158, KeyReg_Inst_ff_SDE_94_next_state}), .Q ({new_AGEMA_signal_4913, RoundKey[94]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_95_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8160, KeyReg_Inst_ff_SDE_95_next_state}), .Q ({new_AGEMA_signal_4916, RoundKey[95]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_96_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7498, KeyReg_Inst_ff_SDE_96_next_state}), .Q ({new_AGEMA_signal_4919, RoundKey[96]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_97_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7670, KeyReg_Inst_ff_SDE_97_next_state}), .Q ({new_AGEMA_signal_4922, RoundKey[97]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_98_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7672, KeyReg_Inst_ff_SDE_98_next_state}), .Q ({new_AGEMA_signal_4925, RoundKey[98]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_99_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7674, KeyReg_Inst_ff_SDE_99_next_state}), .Q ({new_AGEMA_signal_4928, RoundKey[99]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_100_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7676, KeyReg_Inst_ff_SDE_100_next_state}), .Q ({new_AGEMA_signal_4553, RoundKey[100]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_101_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7678, KeyReg_Inst_ff_SDE_101_next_state}), .Q ({new_AGEMA_signal_4556, RoundKey[101]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_102_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7680, KeyReg_Inst_ff_SDE_102_next_state}), .Q ({new_AGEMA_signal_4559, RoundKey[102]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_103_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7682, KeyReg_Inst_ff_SDE_103_next_state}), .Q ({new_AGEMA_signal_4562, RoundKey[103]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_104_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7500, KeyReg_Inst_ff_SDE_104_next_state}), .Q ({new_AGEMA_signal_4565, RoundKey[104]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_105_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7684, KeyReg_Inst_ff_SDE_105_next_state}), .Q ({new_AGEMA_signal_4568, RoundKey[105]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_106_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7686, KeyReg_Inst_ff_SDE_106_next_state}), .Q ({new_AGEMA_signal_4571, RoundKey[106]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_107_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7688, KeyReg_Inst_ff_SDE_107_next_state}), .Q ({new_AGEMA_signal_4574, RoundKey[107]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_108_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7690, KeyReg_Inst_ff_SDE_108_next_state}), .Q ({new_AGEMA_signal_4577, RoundKey[108]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_109_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7692, KeyReg_Inst_ff_SDE_109_next_state}), .Q ({new_AGEMA_signal_4580, RoundKey[109]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_110_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7694, KeyReg_Inst_ff_SDE_110_next_state}), .Q ({new_AGEMA_signal_4586, RoundKey[110]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_111_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7696, KeyReg_Inst_ff_SDE_111_next_state}), .Q ({new_AGEMA_signal_4589, RoundKey[111]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_112_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7502, KeyReg_Inst_ff_SDE_112_next_state}), .Q ({new_AGEMA_signal_4592, RoundKey[112]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_113_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7698, KeyReg_Inst_ff_SDE_113_next_state}), .Q ({new_AGEMA_signal_4595, RoundKey[113]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_114_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7700, KeyReg_Inst_ff_SDE_114_next_state}), .Q ({new_AGEMA_signal_4598, RoundKey[114]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_115_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7702, KeyReg_Inst_ff_SDE_115_next_state}), .Q ({new_AGEMA_signal_4601, RoundKey[115]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_116_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7704, KeyReg_Inst_ff_SDE_116_next_state}), .Q ({new_AGEMA_signal_4604, RoundKey[116]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_117_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7706, KeyReg_Inst_ff_SDE_117_next_state}), .Q ({new_AGEMA_signal_4607, RoundKey[117]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_118_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7708, KeyReg_Inst_ff_SDE_118_next_state}), .Q ({new_AGEMA_signal_4610, RoundKey[118]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_119_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7710, KeyReg_Inst_ff_SDE_119_next_state}), .Q ({new_AGEMA_signal_4613, RoundKey[119]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_120_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7712, KeyReg_Inst_ff_SDE_120_next_state}), .Q ({new_AGEMA_signal_4619, RoundKey[120]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_121_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7924, KeyReg_Inst_ff_SDE_121_next_state}), .Q ({new_AGEMA_signal_4622, RoundKey[121]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_122_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7926, KeyReg_Inst_ff_SDE_122_next_state}), .Q ({new_AGEMA_signal_4625, RoundKey[122]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_123_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7928, KeyReg_Inst_ff_SDE_123_next_state}), .Q ({new_AGEMA_signal_4628, RoundKey[123]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_124_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7930, KeyReg_Inst_ff_SDE_124_next_state}), .Q ({new_AGEMA_signal_4631, RoundKey[124]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_125_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7932, KeyReg_Inst_ff_SDE_125_next_state}), .Q ({new_AGEMA_signal_4634, RoundKey[125]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_126_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7934, KeyReg_Inst_ff_SDE_126_next_state}), .Q ({new_AGEMA_signal_4637, RoundKey[126]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_127_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_7936, KeyReg_Inst_ff_SDE_127_next_state}), .Q ({new_AGEMA_signal_4640, RoundKey[127]}) ) ;
    DFF_X1 RoundCounterIns_count_reg_0__FF_FF ( .CK (clk), .D (new_AGEMA_signal_15816), .Q (RoundCounter[0]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_1__FF_FF ( .CK (clk), .D (new_AGEMA_signal_15820), .Q (RoundCounter[1]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_2__FF_FF ( .CK (clk), .D (new_AGEMA_signal_15824), .Q (RoundCounter[2]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_3__FF_FF ( .CK (clk), .D (new_AGEMA_signal_15828), .Q (RoundCounter[3]), .QN () ) ;
endmodule
