module sbox (SI, clk, SO);
   
   /* Inputs */
   input      [7:0] SI;
   input      clk;
   
   /* Outputs */
   output reg [7:0] SO;   
   
   /* Always blocks */
   always @(posedge clk)
   begin
      case(SI)
	8'h00 :  SO = 8'h63;
	8'h01 :  SO = 8'h7C;
	8'h02 :  SO = 8'h77;
	8'h03 :  SO = 8'h7B;
	8'h04 :  SO = 8'hF2;
	8'h05 :  SO = 8'h6B;
	8'h06 :  SO = 8'h6F;
	8'h07 :  SO = 8'hC5;
	8'h08 :  SO = 8'h30;
	8'h09 :  SO = 8'h01;
	8'h0A :  SO = 8'h67;
	8'h0B :  SO = 8'h2B;
	8'h0C :  SO = 8'hFE;
	8'h0D :  SO = 8'hD7;
	8'h0E :  SO = 8'hAB;
	8'h0F :  SO = 8'h76;
	8'h10 :  SO = 8'hCA;
	8'h11 :  SO = 8'h82;
	8'h12 :  SO = 8'hC9;
	8'h13 :  SO = 8'h7D;
	8'h14 :  SO = 8'hFA;
	8'h15 :  SO = 8'h59;
	8'h16 :  SO = 8'h47;
	8'h17 :  SO = 8'hF0;
	8'h18 :  SO = 8'hAD;
	8'h19 :  SO = 8'hD4;
	8'h1A :  SO = 8'hA2;
	8'h1B :  SO = 8'hAF;
	8'h1C :  SO = 8'h9C;
	8'h1D :  SO = 8'hA4;
	8'h1E :  SO = 8'h72;
	8'h1F :  SO = 8'hC0;
	8'h20 :  SO = 8'hB7;
	8'h21 :  SO = 8'hFD;
	8'h22 :  SO = 8'h93;
	8'h23 :  SO = 8'h26;
	8'h24 :  SO = 8'h36;
	8'h25 :  SO = 8'h3F;
	8'h26 :  SO = 8'hF7;
	8'h27 :  SO = 8'hCC;
	8'h28 :  SO = 8'h34;
	8'h29 :  SO = 8'hA5;
	8'h2A :  SO = 8'hE5;
	8'h2B :  SO = 8'hF1;
	8'h2C :  SO = 8'h71;
	8'h2D :  SO = 8'hD8;
	8'h2E :  SO = 8'h31;
	8'h2F :  SO = 8'h15;
	8'h30 :  SO = 8'h04;
	8'h31 :  SO = 8'hC7;
	8'h32 :  SO = 8'h23;
	8'h33 :  SO = 8'hC3;
	8'h34 :  SO = 8'h18;
	8'h35 :  SO = 8'h96;
	8'h36 :  SO = 8'h05;
	8'h37 :  SO = 8'h9A;
	8'h38 :  SO = 8'h07;
	8'h39 :  SO = 8'h12;
	8'h3A :  SO = 8'h80;
	8'h3B :  SO = 8'hE2;
	8'h3C :  SO = 8'hEB;
	8'h3D :  SO = 8'h27;
	8'h3E :  SO = 8'hB2;
	8'h3F :  SO = 8'h75;
	8'h40 :  SO = 8'h09;
	8'h41 :  SO = 8'h83;
	8'h42 :  SO = 8'h2C;
	8'h43 :  SO = 8'h1A;
	8'h44 :  SO = 8'h1B;
	8'h45 :  SO = 8'h6E;
	8'h46 :  SO = 8'h5A;
	8'h47 :  SO = 8'hA0;
	8'h48 :  SO = 8'h52;
	8'h49 :  SO = 8'h3B;
	8'h4A :  SO = 8'hD6;
	8'h4B :  SO = 8'hB3;
	8'h4C :  SO = 8'h29;
	8'h4D :  SO = 8'hE3;
	8'h4E :  SO = 8'h2F;
	8'h4F :  SO = 8'h84;
	8'h50 :  SO = 8'h53;
	8'h51 :  SO = 8'hD1;
	8'h52 :  SO = 8'h00;
	8'h53 :  SO = 8'hED;
	8'h54 :  SO = 8'h20;
	8'h55 :  SO = 8'hFC;
	8'h56 :  SO = 8'hB1;
	8'h57 :  SO = 8'h5B;
	8'h58 :  SO = 8'h6A;
	8'h59 :  SO = 8'hCB;
	8'h5A :  SO = 8'hBE;
	8'h5B :  SO = 8'h39;
	8'h5C :  SO = 8'h4A;
	8'h5D :  SO = 8'h4C;
	8'h5E :  SO = 8'h58;
	8'h5F :  SO = 8'hCF;
	8'h60 :  SO = 8'hD0;
	8'h61 :  SO = 8'hEF;
	8'h62 :  SO = 8'hAA;
	8'h63 :  SO = 8'hFB;
	8'h64 :  SO = 8'h43;
	8'h65 :  SO = 8'h4D;
	8'h66 :  SO = 8'h33;
	8'h67 :  SO = 8'h85;
	8'h68 :  SO = 8'h45;
	8'h69 :  SO = 8'hF9;
	8'h6A :  SO = 8'h02;
	8'h6B :  SO = 8'h7F;
	8'h6C :  SO = 8'h50;
	8'h6D :  SO = 8'h3C;
	8'h6E :  SO = 8'h9F;
	8'h6F :  SO = 8'hA8;
	8'h70 :  SO = 8'h51;
	8'h71 :  SO = 8'hA3;
	8'h72 :  SO = 8'h40;
	8'h73 :  SO = 8'h8F;
	8'h74 :  SO = 8'h92;
	8'h75 :  SO = 8'h9D;
	8'h76 :  SO = 8'h38;
	8'h77 :  SO = 8'hF5;
	8'h78 :  SO = 8'hBC;
	8'h79 :  SO = 8'hB6;
	8'h7A :  SO = 8'hDA;
	8'h7B :  SO = 8'h21;
	8'h7C :  SO = 8'h10;
	8'h7D :  SO = 8'hFF;
	8'h7E :  SO = 8'hF3;
	8'h7F :  SO = 8'hD2;
	8'h80 :  SO = 8'hCD;
	8'h81 :  SO = 8'h0C;
	8'h82 :  SO = 8'h13;
	8'h83 :  SO = 8'hEC;
	8'h84 :  SO = 8'h5F;
	8'h85 :  SO = 8'h97;
	8'h86 :  SO = 8'h44;
	8'h87 :  SO = 8'h17;
	8'h88 :  SO = 8'hC4;
	8'h89 :  SO = 8'hA7;
	8'h8A :  SO = 8'h7E;
	8'h8B :  SO = 8'h3D;
	8'h8C :  SO = 8'h64;
	8'h8D :  SO = 8'h5D;
	8'h8E :  SO = 8'h19;
	8'h8F :  SO = 8'h73;
	8'h90 :  SO = 8'h60;
	8'h91 :  SO = 8'h81;
	8'h92 :  SO = 8'h4F;
	8'h93 :  SO = 8'hDC;
	8'h94 :  SO = 8'h22;
	8'h95 :  SO = 8'h2A;
	8'h96 :  SO = 8'h90;
	8'h97 :  SO = 8'h88;
	8'h98 :  SO = 8'h46;
	8'h99 :  SO = 8'hEE;
	8'h9A :  SO = 8'hB8;
	8'h9B :  SO = 8'h14;
	8'h9C :  SO = 8'hDE;
	8'h9D :  SO = 8'h5E;
	8'h9E :  SO = 8'h0B;
	8'h9F :  SO = 8'hDB;
	8'hA0 :  SO = 8'hE0;
	8'hA1 :  SO = 8'h32;
	8'hA2 :  SO = 8'h3A;
	8'hA3 :  SO = 8'h0A;
	8'hA4 :  SO = 8'h49;
	8'hA5 :  SO = 8'h06;
	8'hA6 :  SO = 8'h24;
	8'hA7 :  SO = 8'h5C;
	8'hA8 :  SO = 8'hC2;
	8'hA9 :  SO = 8'hD3;
	8'hAA :  SO = 8'hAC;
	8'hAB :  SO = 8'h62;
	8'hAC :  SO = 8'h91;
	8'hAD :  SO = 8'h95;
	8'hAE :  SO = 8'hE4;
	8'hAF :  SO = 8'h79;
	8'hB0 :  SO = 8'hE7;
	8'hB1 :  SO = 8'hC8;
	8'hB2 :  SO = 8'h37;
	8'hB3 :  SO = 8'h6D;
	8'hB4 :  SO = 8'h8D;
	8'hB5 :  SO = 8'hD5;
	8'hB6 :  SO = 8'h4E;
	8'hB7 :  SO = 8'hA9;
	8'hB8 :  SO = 8'h6C;
	8'hB9 :  SO = 8'h56;
	8'hBA :  SO = 8'hF4;
	8'hBB :  SO = 8'hEA;
	8'hBC :  SO = 8'h65;
	8'hBD :  SO = 8'h7A;
	8'hBE :  SO = 8'hAE;
	8'hBF :  SO = 8'h08;
	8'hC0 :  SO = 8'hBA;
	8'hC1 :  SO = 8'h78;
	8'hC2 :  SO = 8'h25;
	8'hC3 :  SO = 8'h2E;
	8'hC4 :  SO = 8'h1C;
	8'hC5 :  SO = 8'hA6;
	8'hC6 :  SO = 8'hB4;
	8'hC7 :  SO = 8'hC6;
	8'hC8 :  SO = 8'hE8;
	8'hC9 :  SO = 8'hDD;
	8'hCA :  SO = 8'h74;
	8'hCB :  SO = 8'h1F;
	8'hCC :  SO = 8'h4B;
	8'hCD :  SO = 8'hBD;
	8'hCE :  SO = 8'h8B;
	8'hCF :  SO = 8'h8A;
	8'hD0 :  SO = 8'h70;
	8'hD1 :  SO = 8'h3E;
	8'hD2 :  SO = 8'hB5;
	8'hD3 :  SO = 8'h66;
	8'hD4 :  SO = 8'h48;
	8'hD5 :  SO = 8'h03;
	8'hD6 :  SO = 8'hF6;
	8'hD7 :  SO = 8'h0E;
	8'hD8 :  SO = 8'h61;
	8'hD9 :  SO = 8'h35;
	8'hDA :  SO = 8'h57;
	8'hDB :  SO = 8'hB9;
	8'hDC :  SO = 8'h86;
	8'hDD :  SO = 8'hC1;
	8'hDE :  SO = 8'h1D;
	8'hDF :  SO = 8'h9E;
	8'hE0 :  SO = 8'hE1;
	8'hE1 :  SO = 8'hF8;
	8'hE2 :  SO = 8'h98;
	8'hE3 :  SO = 8'h11;
	8'hE4 :  SO = 8'h69;
	8'hE5 :  SO = 8'hD9;
	8'hE6 :  SO = 8'h8E;
	8'hE7 :  SO = 8'h94;
	8'hE8 :  SO = 8'h9B;
	8'hE9 :  SO = 8'h1E;
	8'hEA :  SO = 8'h87;
	8'hEB :  SO = 8'hE9;
	8'hEC :  SO = 8'hCE;
	8'hED :  SO = 8'h55;
	8'hEE :  SO = 8'h28;
	8'hEF :  SO = 8'hDF;
	8'hF0 :  SO = 8'h8C;
	8'hF1 :  SO = 8'hA1;
	8'hF2 :  SO = 8'h89;
	8'hF3 :  SO = 8'h0D;
	8'hF4 :  SO = 8'hBF;
	8'hF5 :  SO = 8'hE6;
	8'hF6 :  SO = 8'h42;
	8'hF7 :  SO = 8'h68;
	8'hF8 :  SO = 8'h41;
	8'hF9 :  SO = 8'h99;
	8'hFA :  SO = 8'h2D;
	8'hFB :  SO = 8'h0F;
	8'hFC :  SO = 8'hB0;
	8'hFD :  SO = 8'h54;
	8'hFE :  SO = 8'hBB;
	8'hFF :  SO = 8'h16;
      endcase
   end

endmodule


			
