/* modified netlist. Source: module CRAFT in file /mnt/c/Users/Amir/Desktop/Papers_in_progress/AGEMA/Designs/CRAFT_round-based/AGEMA/CRAFT.v */
/* clock gating is added to the circuit, the latency increased 8 time(s)  */

module CRAFT_HPC2_AIG_ClockGating_d1 (plaintext_s0, key_s0, clk, rst, key_s1, plaintext_s1, Fresh, ciphertext_s0, done, ciphertext_s1, Synch);
    input [63:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input rst ;
    input [127:0] key_s1 ;
    input [63:0] plaintext_s1 ;
    input [255:0] Fresh ;
    output [63:0] ciphertext_s0 ;
    output done ;
    output [63:0] ciphertext_s1 ;
    output Synch ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_285 ;
    wire signal_286 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_295 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_352 ;
    wire signal_353 ;
    wire signal_354 ;
    wire signal_355 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_359 ;
    wire signal_360 ;
    wire signal_361 ;
    wire signal_362 ;
    wire signal_363 ;
    wire signal_364 ;
    wire signal_365 ;
    wire signal_366 ;
    wire signal_367 ;
    wire signal_368 ;
    wire signal_369 ;
    wire signal_370 ;
    wire signal_371 ;
    wire signal_372 ;
    wire signal_373 ;
    wire signal_374 ;
    wire signal_375 ;
    wire signal_376 ;
    wire signal_377 ;
    wire signal_378 ;
    wire signal_379 ;
    wire signal_380 ;
    wire signal_381 ;
    wire signal_382 ;
    wire signal_383 ;
    wire signal_384 ;
    wire signal_385 ;
    wire signal_386 ;
    wire signal_387 ;
    wire signal_692 ;
    wire signal_693 ;
    wire signal_694 ;
    wire signal_702 ;
    wire signal_703 ;
    wire signal_704 ;
    wire signal_705 ;
    wire signal_706 ;
    wire signal_707 ;
    wire signal_711 ;
    wire signal_712 ;
    wire signal_713 ;
    wire signal_714 ;
    wire signal_715 ;
    wire signal_716 ;
    wire signal_717 ;
    wire signal_718 ;
    wire signal_719 ;
    wire signal_720 ;
    wire signal_721 ;
    wire signal_722 ;
    wire signal_723 ;
    wire signal_724 ;
    wire signal_725 ;
    wire signal_726 ;
    wire signal_727 ;
    wire signal_728 ;
    wire signal_729 ;
    wire signal_730 ;
    wire signal_731 ;
    wire signal_732 ;
    wire signal_733 ;
    wire signal_734 ;
    wire signal_735 ;
    wire signal_736 ;
    wire signal_737 ;
    wire signal_738 ;
    wire signal_739 ;
    wire signal_740 ;
    wire signal_741 ;
    wire signal_742 ;
    wire signal_743 ;
    wire signal_744 ;
    wire signal_745 ;
    wire signal_746 ;
    wire signal_747 ;
    wire signal_748 ;
    wire signal_749 ;
    wire signal_750 ;
    wire signal_751 ;
    wire signal_752 ;
    wire signal_753 ;
    wire signal_754 ;
    wire signal_755 ;
    wire signal_756 ;
    wire signal_757 ;
    wire signal_758 ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_768 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_771 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_774 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_777 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_780 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_783 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_786 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_789 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_792 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_809 ;
    wire signal_810 ;
    wire signal_811 ;
    wire signal_812 ;
    wire signal_813 ;
    wire signal_814 ;
    wire signal_815 ;
    wire signal_816 ;
    wire signal_817 ;
    wire signal_818 ;
    wire signal_819 ;
    wire signal_820 ;
    wire signal_821 ;
    wire signal_822 ;
    wire signal_823 ;
    wire signal_824 ;
    wire signal_825 ;
    wire signal_826 ;
    wire signal_827 ;
    wire signal_828 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_831 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_834 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_837 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_840 ;
    wire signal_841 ;
    wire signal_842 ;
    wire signal_843 ;
    wire signal_844 ;
    wire signal_845 ;
    wire signal_846 ;
    wire signal_847 ;
    wire signal_848 ;
    wire signal_849 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_852 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_855 ;
    wire signal_856 ;
    wire signal_857 ;
    wire signal_858 ;
    wire signal_859 ;
    wire signal_860 ;
    wire signal_861 ;
    wire signal_862 ;
    wire signal_863 ;
    wire signal_864 ;
    wire signal_865 ;
    wire signal_866 ;
    wire signal_867 ;
    wire signal_868 ;
    wire signal_869 ;
    wire signal_870 ;
    wire signal_871 ;
    wire signal_872 ;
    wire signal_873 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_879 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_885 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_888 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_891 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_894 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_897 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_900 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_903 ;
    wire signal_904 ;
    wire signal_905 ;
    wire signal_906 ;
    wire signal_907 ;
    wire signal_908 ;
    wire signal_909 ;
    wire signal_910 ;
    wire signal_911 ;
    wire signal_912 ;
    wire signal_913 ;
    wire signal_914 ;
    wire signal_915 ;
    wire signal_916 ;
    wire signal_917 ;
    wire signal_918 ;
    wire signal_919 ;
    wire signal_920 ;
    wire signal_921 ;
    wire signal_922 ;
    wire signal_923 ;
    wire signal_924 ;
    wire signal_925 ;
    wire signal_926 ;
    wire signal_927 ;
    wire signal_928 ;
    wire signal_929 ;
    wire signal_930 ;
    wire signal_931 ;
    wire signal_932 ;
    wire signal_933 ;
    wire signal_934 ;
    wire signal_935 ;
    wire signal_936 ;
    wire signal_937 ;
    wire signal_938 ;
    wire signal_939 ;
    wire signal_940 ;
    wire signal_941 ;
    wire signal_942 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1020 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1023 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1276 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1279 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1282 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1285 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1288 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1294 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1297 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1300 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1303 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1309 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1494 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1499 ;
    wire signal_1500 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1503 ;
    wire signal_1504 ;
    wire signal_1505 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1509 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1512 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1516 ;
    wire signal_1518 ;
    wire signal_1520 ;
    wire signal_1522 ;
    wire signal_1524 ;
    wire signal_1526 ;
    wire signal_1528 ;
    wire signal_1530 ;
    wire signal_1532 ;
    wire signal_1534 ;
    wire signal_1536 ;
    wire signal_1538 ;
    wire signal_1540 ;
    wire signal_1542 ;
    wire signal_1544 ;
    wire signal_1546 ;
    wire signal_1548 ;
    wire signal_1550 ;
    wire signal_1552 ;
    wire signal_1554 ;
    wire signal_1556 ;
    wire signal_1558 ;
    wire signal_1560 ;
    wire signal_1562 ;
    wire signal_1564 ;
    wire signal_1566 ;
    wire signal_1568 ;
    wire signal_1570 ;
    wire signal_1572 ;
    wire signal_1574 ;
    wire signal_1576 ;
    wire signal_1578 ;
    wire signal_1580 ;
    wire signal_1582 ;
    wire signal_1584 ;
    wire signal_1586 ;
    wire signal_1588 ;
    wire signal_1590 ;
    wire signal_1592 ;
    wire signal_1594 ;
    wire signal_1596 ;
    wire signal_1598 ;
    wire signal_1600 ;
    wire signal_1602 ;
    wire signal_1604 ;
    wire signal_1606 ;
    wire signal_1608 ;
    wire signal_1610 ;
    wire signal_1612 ;
    wire signal_1614 ;
    wire signal_1616 ;
    wire signal_1618 ;
    wire signal_1620 ;
    wire signal_1622 ;
    wire signal_1624 ;
    wire signal_1626 ;
    wire signal_1628 ;
    wire signal_1630 ;
    wire signal_1632 ;
    wire signal_1634 ;
    wire signal_1636 ;
    wire signal_1638 ;
    wire signal_1640 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1657 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1660 ;
    wire signal_1661 ;
    wire signal_1662 ;
    wire signal_1663 ;
    wire signal_1664 ;
    wire signal_1665 ;
    wire signal_1666 ;
    wire signal_1667 ;
    wire signal_1668 ;
    wire signal_1669 ;
    wire signal_1670 ;
    wire signal_1671 ;
    wire signal_1672 ;
    wire signal_1673 ;
    wire signal_1674 ;
    wire signal_1677 ;
    wire signal_1680 ;
    wire signal_1683 ;
    wire signal_1686 ;
    wire signal_1689 ;
    wire signal_1692 ;
    wire signal_1695 ;
    wire signal_1698 ;
    wire signal_1701 ;
    wire signal_1704 ;
    wire signal_1707 ;
    wire signal_1710 ;
    wire signal_1713 ;
    wire signal_1716 ;
    wire signal_1719 ;
    wire signal_1722 ;
    wire signal_1723 ;
    wire signal_1724 ;
    wire signal_1725 ;
    wire signal_1726 ;
    wire signal_1727 ;
    wire signal_1728 ;
    wire signal_1729 ;
    wire signal_1730 ;
    wire signal_1731 ;
    wire signal_1732 ;
    wire signal_1733 ;
    wire signal_1734 ;
    wire signal_1735 ;
    wire signal_1736 ;
    wire signal_1737 ;
    wire signal_1738 ;
    wire signal_1739 ;
    wire signal_1740 ;
    wire signal_1741 ;
    wire signal_1742 ;
    wire signal_1743 ;
    wire signal_1744 ;
    wire signal_1745 ;
    wire signal_1746 ;
    wire signal_1747 ;
    wire signal_1748 ;
    wire signal_1749 ;
    wire signal_1750 ;
    wire signal_1751 ;
    wire signal_1752 ;
    wire signal_1753 ;
    wire signal_1754 ;
    wire signal_1755 ;
    wire signal_1756 ;
    wire signal_1757 ;
    wire signal_1758 ;
    wire signal_1759 ;
    wire signal_1760 ;
    wire signal_1761 ;
    wire signal_1762 ;
    wire signal_1763 ;
    wire signal_1764 ;
    wire signal_1765 ;
    wire signal_1766 ;
    wire signal_1767 ;
    wire signal_1768 ;
    wire signal_1769 ;
    wire signal_1770 ;
    wire signal_1771 ;
    wire signal_1772 ;
    wire signal_1773 ;
    wire signal_1774 ;
    wire signal_1775 ;
    wire signal_1776 ;
    wire signal_1777 ;
    wire signal_1778 ;
    wire signal_1779 ;
    wire signal_1780 ;
    wire signal_1781 ;
    wire signal_1782 ;
    wire signal_1783 ;
    wire signal_1784 ;
    wire signal_1785 ;
    wire signal_1786 ;
    wire signal_1787 ;
    wire signal_1788 ;
    wire signal_1789 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1792 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1795 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1813 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1844 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1854 ;
    wire signal_1855 ;
    wire signal_1856 ;
    wire signal_1857 ;
    wire signal_1858 ;
    wire signal_1859 ;
    wire signal_1860 ;
    wire signal_1861 ;
    wire signal_1862 ;
    wire signal_1863 ;
    wire signal_1864 ;
    wire signal_1865 ;
    wire signal_1866 ;
    wire signal_1867 ;
    wire signal_1868 ;
    wire signal_1869 ;
    wire signal_1870 ;
    wire signal_1871 ;
    wire signal_1872 ;
    wire signal_1873 ;
    wire signal_1874 ;
    wire signal_1875 ;
    wire signal_1876 ;
    wire signal_1877 ;
    wire signal_1878 ;
    wire signal_1879 ;
    wire signal_1880 ;
    wire signal_1881 ;
    wire signal_1882 ;
    wire signal_1883 ;
    wire signal_1884 ;
    wire signal_1885 ;
    wire signal_1886 ;
    wire signal_1887 ;
    wire signal_1888 ;
    wire signal_1889 ;
    wire signal_1890 ;
    wire signal_1891 ;
    wire signal_1892 ;
    wire signal_1893 ;
    wire signal_1894 ;
    wire signal_1895 ;
    wire signal_1896 ;
    wire signal_1897 ;
    wire signal_1898 ;
    wire signal_1899 ;
    wire signal_1900 ;
    wire signal_1901 ;
    wire signal_1902 ;
    wire signal_1903 ;
    wire signal_1904 ;
    wire signal_1905 ;
    wire signal_1906 ;
    wire signal_1907 ;
    wire signal_1908 ;
    wire signal_1909 ;
    wire signal_1910 ;
    wire signal_1911 ;
    wire signal_1912 ;
    wire signal_1913 ;
    wire signal_1914 ;
    wire signal_1917 ;
    wire signal_1920 ;
    wire signal_1923 ;
    wire signal_1926 ;
    wire signal_1929 ;
    wire signal_1932 ;
    wire signal_1935 ;
    wire signal_1938 ;
    wire signal_1941 ;
    wire signal_1944 ;
    wire signal_1947 ;
    wire signal_1950 ;
    wire signal_1953 ;
    wire signal_1956 ;
    wire signal_1959 ;
    wire signal_1962 ;
    wire signal_1965 ;
    wire signal_1968 ;
    wire signal_1971 ;
    wire signal_1974 ;
    wire signal_1977 ;
    wire signal_1980 ;
    wire signal_1983 ;
    wire signal_1986 ;
    wire signal_1989 ;
    wire signal_1992 ;
    wire signal_1995 ;
    wire signal_1998 ;
    wire signal_2001 ;
    wire signal_2004 ;
    wire signal_2007 ;
    wire signal_2010 ;
    wire signal_2013 ;
    wire signal_2016 ;
    wire signal_2019 ;
    wire signal_2022 ;
    wire signal_2025 ;
    wire signal_2028 ;
    wire signal_2031 ;
    wire signal_2034 ;
    wire signal_2037 ;
    wire signal_2040 ;
    wire signal_2043 ;
    wire signal_2046 ;
    wire signal_2049 ;
    wire signal_2052 ;
    wire signal_2055 ;
    wire signal_2058 ;
    wire signal_2059 ;
    wire signal_2060 ;
    wire signal_2061 ;
    wire signal_2062 ;
    wire signal_2063 ;
    wire signal_2064 ;
    wire signal_2065 ;
    wire signal_2066 ;
    wire signal_2067 ;
    wire signal_2068 ;
    wire signal_2069 ;
    wire signal_2070 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2079 ;
    wire signal_2080 ;
    wire signal_2081 ;
    wire signal_2082 ;
    wire signal_2083 ;
    wire signal_2084 ;
    wire signal_2085 ;
    wire signal_2086 ;
    wire signal_2087 ;
    wire signal_2088 ;
    wire signal_2089 ;
    wire signal_2090 ;
    wire signal_2091 ;
    wire signal_2092 ;
    wire signal_2093 ;
    wire signal_2094 ;
    wire signal_2095 ;
    wire signal_2096 ;
    wire signal_2097 ;
    wire signal_2098 ;
    wire signal_2099 ;
    wire signal_2100 ;
    wire signal_2101 ;
    wire signal_2102 ;
    wire signal_2103 ;
    wire signal_2104 ;
    wire signal_2105 ;
    wire signal_2106 ;
    wire signal_2107 ;
    wire signal_2108 ;
    wire signal_2109 ;
    wire signal_2110 ;
    wire signal_2111 ;
    wire signal_2112 ;
    wire signal_2113 ;
    wire signal_2114 ;
    wire signal_2115 ;
    wire signal_2116 ;
    wire signal_2117 ;
    wire signal_2118 ;
    wire signal_2119 ;
    wire signal_2120 ;
    wire signal_2121 ;
    wire signal_2122 ;
    wire signal_2123 ;
    wire signal_2124 ;
    wire signal_2125 ;
    wire signal_2126 ;
    wire signal_2127 ;
    wire signal_2128 ;
    wire signal_2129 ;
    wire signal_2130 ;
    wire signal_2131 ;
    wire signal_2132 ;
    wire signal_2133 ;
    wire signal_2134 ;
    wire signal_2135 ;
    wire signal_2136 ;
    wire signal_2137 ;
    wire signal_2138 ;
    wire signal_2139 ;
    wire signal_2140 ;
    wire signal_2141 ;
    wire signal_2142 ;
    wire signal_2143 ;
    wire signal_2144 ;
    wire signal_2145 ;
    wire signal_2146 ;
    wire signal_2147 ;
    wire signal_2148 ;
    wire signal_2149 ;
    wire signal_2150 ;
    wire signal_2151 ;
    wire signal_2152 ;
    wire signal_2153 ;
    wire signal_2154 ;
    wire signal_2155 ;
    wire signal_2156 ;
    wire signal_2157 ;
    wire signal_2158 ;
    wire signal_2159 ;
    wire signal_2160 ;
    wire signal_2161 ;
    wire signal_2162 ;
    wire signal_2163 ;
    wire signal_2164 ;
    wire signal_2165 ;
    wire signal_2166 ;
    wire signal_2167 ;
    wire signal_2168 ;
    wire signal_2169 ;
    wire signal_2170 ;
    wire signal_2171 ;
    wire signal_2172 ;
    wire signal_2173 ;
    wire signal_2174 ;
    wire signal_2175 ;
    wire signal_2176 ;
    wire signal_2177 ;
    wire signal_2178 ;
    wire signal_2179 ;
    wire signal_2180 ;
    wire signal_2181 ;
    wire signal_2182 ;
    wire signal_2183 ;
    wire signal_2184 ;
    wire signal_2185 ;
    wire signal_2186 ;
    wire signal_2187 ;
    wire signal_2188 ;
    wire signal_2189 ;
    wire signal_2190 ;
    wire signal_2191 ;
    wire signal_2192 ;
    wire signal_2193 ;
    wire signal_2194 ;
    wire signal_2195 ;
    wire signal_2196 ;
    wire signal_2197 ;
    wire signal_2198 ;
    wire signal_2199 ;
    wire signal_2200 ;
    wire signal_2201 ;
    wire signal_2202 ;
    wire signal_2203 ;
    wire signal_2204 ;
    wire signal_2205 ;
    wire signal_2206 ;
    wire signal_2207 ;
    wire signal_2208 ;
    wire signal_2209 ;
    wire signal_2210 ;
    wire signal_2211 ;
    wire signal_2212 ;
    wire signal_2213 ;
    wire signal_2214 ;
    wire signal_2215 ;
    wire signal_2216 ;
    wire signal_2217 ;
    wire signal_2218 ;
    wire signal_2219 ;
    wire signal_2220 ;
    wire signal_2221 ;
    wire signal_2222 ;
    wire signal_2223 ;
    wire signal_2224 ;
    wire signal_2225 ;
    wire signal_2226 ;
    wire signal_2227 ;
    wire signal_2228 ;
    wire signal_2229 ;
    wire signal_2230 ;
    wire signal_2231 ;
    wire signal_2232 ;
    wire signal_2233 ;
    wire signal_2234 ;
    wire signal_2235 ;
    wire signal_2236 ;
    wire signal_2237 ;
    wire signal_2238 ;
    wire signal_2239 ;
    wire signal_2240 ;
    wire signal_2241 ;
    wire signal_2242 ;
    wire signal_2243 ;
    wire signal_2244 ;
    wire signal_2245 ;
    wire signal_2246 ;
    wire signal_2247 ;
    wire signal_2248 ;
    wire signal_2249 ;
    wire signal_2250 ;
    wire signal_2251 ;
    wire signal_2252 ;
    wire signal_2253 ;
    wire signal_2254 ;
    wire signal_2255 ;
    wire signal_2256 ;
    wire signal_2257 ;
    wire signal_2258 ;
    wire signal_2260 ;
    wire signal_2262 ;
    wire signal_2264 ;
    wire signal_2266 ;
    wire signal_2268 ;
    wire signal_2270 ;
    wire signal_2272 ;
    wire signal_2274 ;
    wire signal_2276 ;
    wire signal_2278 ;
    wire signal_2280 ;
    wire signal_2282 ;
    wire signal_2284 ;
    wire signal_2286 ;
    wire signal_2288 ;
    wire signal_2290 ;
    wire signal_2291 ;
    wire signal_2292 ;
    wire signal_2293 ;
    wire signal_2294 ;
    wire signal_2295 ;
    wire signal_2296 ;
    wire signal_2297 ;
    wire signal_2298 ;
    wire signal_2299 ;
    wire signal_2300 ;
    wire signal_2301 ;
    wire signal_2302 ;
    wire signal_2303 ;
    wire signal_2304 ;
    wire signal_2305 ;
    wire signal_2306 ;
    wire signal_2307 ;
    wire signal_2308 ;
    wire signal_2309 ;
    wire signal_2310 ;
    wire signal_2311 ;
    wire signal_2312 ;
    wire signal_2313 ;
    wire signal_2314 ;
    wire signal_2315 ;
    wire signal_2316 ;
    wire signal_2317 ;
    wire signal_2318 ;
    wire signal_2319 ;
    wire signal_2320 ;
    wire signal_2321 ;
    wire signal_2322 ;
    wire signal_2323 ;
    wire signal_2324 ;
    wire signal_2325 ;
    wire signal_2326 ;
    wire signal_2327 ;
    wire signal_2328 ;
    wire signal_2329 ;
    wire signal_2330 ;
    wire signal_2331 ;
    wire signal_2332 ;
    wire signal_2333 ;
    wire signal_2334 ;
    wire signal_2335 ;
    wire signal_2336 ;
    wire signal_2337 ;
    wire signal_2338 ;
    wire signal_2340 ;
    wire signal_2342 ;
    wire signal_2344 ;
    wire signal_2346 ;
    wire signal_2348 ;
    wire signal_2350 ;
    wire signal_2352 ;
    wire signal_2354 ;
    wire signal_2356 ;
    wire signal_2358 ;
    wire signal_2360 ;
    wire signal_2362 ;
    wire signal_2364 ;
    wire signal_2366 ;
    wire signal_2368 ;
    wire signal_2370 ;
    wire signal_2371 ;
    wire signal_2372 ;
    wire signal_2373 ;
    wire signal_2374 ;
    wire signal_2375 ;
    wire signal_2376 ;
    wire signal_2377 ;
    wire signal_2378 ;
    wire signal_2379 ;
    wire signal_2380 ;
    wire signal_2381 ;
    wire signal_2382 ;
    wire signal_2383 ;
    wire signal_2384 ;
    wire signal_2385 ;
    wire signal_2386 ;
    wire signal_2387 ;
    wire signal_2388 ;
    wire signal_2389 ;
    wire signal_2390 ;
    wire signal_2391 ;
    wire signal_2392 ;
    wire signal_2393 ;
    wire signal_2394 ;
    wire signal_2395 ;
    wire signal_2396 ;
    wire signal_2397 ;
    wire signal_2398 ;
    wire signal_2399 ;
    wire signal_2400 ;
    wire signal_2401 ;
    wire signal_2402 ;
    wire signal_2403 ;
    wire signal_2404 ;
    wire signal_2405 ;
    wire signal_2406 ;
    wire signal_2407 ;
    wire signal_2408 ;
    wire signal_2409 ;
    wire signal_2410 ;
    wire signal_2411 ;
    wire signal_2412 ;
    wire signal_2413 ;
    wire signal_2414 ;
    wire signal_2415 ;
    wire signal_2416 ;
    wire signal_2417 ;
    wire signal_2418 ;
    wire signal_2419 ;
    wire signal_2420 ;
    wire signal_2421 ;
    wire signal_2422 ;
    wire signal_2424 ;
    wire signal_2426 ;
    wire signal_2428 ;
    wire signal_2430 ;
    wire signal_2432 ;
    wire signal_2434 ;
    wire signal_2436 ;
    wire signal_2438 ;
    wire signal_2440 ;
    wire signal_2442 ;
    wire signal_2444 ;
    wire signal_2446 ;
    wire signal_2448 ;
    wire signal_2450 ;
    wire signal_2452 ;
    wire signal_2454 ;
    wire signal_2456 ;
    wire signal_2458 ;
    wire signal_2460 ;
    wire signal_2462 ;
    wire signal_2464 ;
    wire signal_2466 ;
    wire signal_2468 ;
    wire signal_2470 ;
    wire signal_2472 ;
    wire signal_2474 ;
    wire signal_2476 ;
    wire signal_2478 ;
    wire signal_2480 ;
    wire signal_2482 ;
    wire signal_2484 ;
    wire signal_2486 ;
    wire signal_2487 ;
    wire signal_2488 ;
    wire signal_2489 ;
    wire signal_2490 ;
    wire signal_2491 ;
    wire signal_2492 ;
    wire signal_2493 ;
    wire signal_2494 ;
    wire signal_2495 ;
    wire signal_2496 ;
    wire signal_2497 ;
    wire signal_2498 ;
    wire signal_2499 ;
    wire signal_2500 ;
    wire signal_2501 ;
    wire signal_2502 ;
    wire signal_2503 ;
    wire signal_2504 ;
    wire signal_2505 ;
    wire signal_2506 ;
    wire signal_2507 ;
    wire signal_2508 ;
    wire signal_2509 ;
    wire signal_2510 ;
    wire signal_2511 ;
    wire signal_2512 ;
    wire signal_2513 ;
    wire signal_2514 ;
    wire signal_2515 ;
    wire signal_2516 ;
    wire signal_2517 ;
    wire signal_2518 ;
    wire signal_2519 ;
    wire signal_2520 ;
    wire signal_2521 ;
    wire signal_2522 ;
    wire signal_2523 ;
    wire signal_2524 ;
    wire signal_2525 ;
    wire signal_2526 ;
    wire signal_2527 ;
    wire signal_2528 ;
    wire signal_2529 ;
    wire signal_2530 ;
    wire signal_2531 ;
    wire signal_2532 ;
    wire signal_2533 ;
    wire signal_2534 ;
    wire signal_2535 ;
    wire signal_2536 ;
    wire signal_2537 ;
    wire signal_2538 ;
    wire signal_2539 ;
    wire signal_2540 ;
    wire signal_2541 ;
    wire signal_2542 ;
    wire signal_2543 ;
    wire signal_2544 ;
    wire signal_2545 ;
    wire signal_2546 ;
    wire signal_2547 ;
    wire signal_2548 ;
    wire signal_2549 ;
    wire signal_2550 ;
    wire signal_2551 ;
    wire signal_2552 ;
    wire signal_2553 ;
    wire signal_2554 ;
    wire signal_2555 ;
    wire signal_2556 ;
    wire signal_2557 ;
    wire signal_2558 ;
    wire signal_2559 ;
    wire signal_2560 ;
    wire signal_2561 ;
    wire signal_2562 ;
    wire signal_2563 ;
    wire signal_2564 ;
    wire signal_2565 ;
    wire signal_2566 ;
    wire signal_2567 ;
    wire signal_2568 ;
    wire signal_2569 ;
    wire signal_2570 ;
    wire signal_2571 ;
    wire signal_2572 ;
    wire signal_2573 ;
    wire signal_2574 ;
    wire signal_2575 ;
    wire signal_2576 ;
    wire signal_2577 ;
    wire signal_2578 ;
    wire signal_2579 ;
    wire signal_2580 ;
    wire signal_2581 ;
    wire signal_2582 ;
    wire signal_2583 ;
    wire signal_2584 ;
    wire signal_2585 ;
    wire signal_2586 ;
    wire signal_2587 ;
    wire signal_2588 ;
    wire signal_2589 ;
    wire signal_2590 ;
    wire signal_2591 ;
    wire signal_2592 ;
    wire signal_2593 ;
    wire signal_2594 ;
    wire signal_2595 ;
    wire signal_2596 ;
    wire signal_2597 ;
    wire signal_2598 ;
    wire signal_2599 ;
    wire signal_2600 ;
    wire signal_2601 ;
    wire signal_2602 ;
    wire signal_2603 ;
    wire signal_2604 ;
    wire signal_2605 ;
    wire signal_2606 ;
    wire signal_2607 ;
    wire signal_2608 ;
    wire signal_2609 ;
    wire signal_2610 ;
    wire signal_2611 ;
    wire signal_2612 ;
    wire signal_2613 ;
    wire signal_2614 ;
    wire signal_2615 ;
    wire signal_2616 ;
    wire signal_2617 ;
    wire signal_2618 ;
    wire signal_2619 ;
    wire signal_2620 ;
    wire signal_2621 ;
    wire signal_2622 ;
    wire signal_2623 ;
    wire signal_2624 ;
    wire signal_2625 ;
    wire signal_2626 ;
    wire signal_2627 ;
    wire signal_2628 ;
    wire signal_2629 ;
    wire signal_2630 ;
    wire signal_2631 ;
    wire signal_2632 ;
    wire signal_2633 ;
    wire signal_2634 ;
    wire signal_2635 ;
    wire signal_2636 ;
    wire signal_2637 ;
    wire signal_2638 ;
    wire signal_2639 ;
    wire signal_2640 ;
    wire signal_2641 ;
    wire signal_2642 ;
    wire signal_2643 ;
    wire signal_2644 ;
    wire signal_2645 ;
    wire signal_2646 ;
    wire signal_2647 ;
    wire signal_2648 ;
    wire signal_2649 ;
    wire signal_2650 ;
    wire signal_2651 ;
    wire signal_2652 ;
    wire signal_2653 ;
    wire signal_2654 ;
    wire signal_2655 ;
    wire signal_2656 ;
    wire signal_2657 ;
    wire signal_2658 ;
    wire signal_2659 ;
    wire signal_2660 ;
    wire signal_2661 ;
    wire signal_2662 ;
    wire signal_2663 ;
    wire signal_2664 ;
    wire signal_2665 ;
    wire signal_2666 ;
    wire signal_2667 ;
    wire signal_2668 ;
    wire signal_2669 ;
    wire signal_2670 ;
    wire signal_2671 ;
    wire signal_2672 ;
    wire signal_2673 ;
    wire signal_2674 ;
    wire signal_2931 ;

    /* cells in depth 0 */
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_177 ( .a ({signal_2004, signal_894}), .b ({1'b0, signal_266}), .c ({signal_2123, signal_333}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_180 ( .a ({signal_2007, signal_893}), .b ({1'b0, signal_1014}), .c ({signal_2124, signal_335}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_183 ( .a ({signal_2010, signal_892}), .b ({1'b0, signal_1013}), .c ({signal_2125, signal_337}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_186 ( .a ({signal_2013, signal_891}), .b ({1'b0, 1'b0}), .c ({signal_2126, signal_339}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_189 ( .a ({signal_2016, signal_890}), .b ({1'b0, signal_265}), .c ({signal_2127, signal_341}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_192 ( .a ({signal_2019, signal_889}), .b ({1'b0, signal_1011}), .c ({signal_2128, signal_343}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_195 ( .a ({signal_2022, signal_888}), .b ({1'b0, signal_1010}), .c ({signal_2129, signal_345}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_198 ( .a ({signal_2025, signal_887}), .b ({1'b0, signal_1009}), .c ({signal_2130, signal_347}) ) ;
    INV_X1 cell_712 ( .A (signal_1000), .ZN (signal_692) ) ;
    INV_X1 cell_713 ( .A (signal_692), .ZN (signal_693) ) ;
    INV_X1 cell_714 ( .A (signal_692), .ZN (signal_694) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_715 ( .s (signal_1000), .b ({key_s1[64], key_s0[64]}), .a ({key_s1[0], key_s0[0]}), .c ({signal_1677, signal_934}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_716 ( .s (signal_693), .b ({key_s1[65], key_s0[65]}), .a ({key_s1[1], key_s0[1]}), .c ({signal_1917, signal_933}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_717 ( .s (signal_1000), .b ({key_s1[66], key_s0[66]}), .a ({key_s1[2], key_s0[2]}), .c ({signal_1680, signal_932}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_718 ( .s (signal_693), .b ({key_s1[67], key_s0[67]}), .a ({key_s1[3], key_s0[3]}), .c ({signal_1920, signal_931}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_719 ( .s (signal_693), .b ({key_s1[68], key_s0[68]}), .a ({key_s1[4], key_s0[4]}), .c ({signal_1923, signal_930}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_720 ( .s (signal_693), .b ({key_s1[69], key_s0[69]}), .a ({key_s1[5], key_s0[5]}), .c ({signal_1926, signal_929}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_721 ( .s (signal_693), .b ({key_s1[70], key_s0[70]}), .a ({key_s1[6], key_s0[6]}), .c ({signal_1929, signal_928}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_722 ( .s (signal_693), .b ({key_s1[71], key_s0[71]}), .a ({key_s1[7], key_s0[7]}), .c ({signal_1932, signal_927}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_723 ( .s (signal_693), .b ({key_s1[72], key_s0[72]}), .a ({key_s1[8], key_s0[8]}), .c ({signal_1935, signal_926}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_724 ( .s (signal_693), .b ({key_s1[73], key_s0[73]}), .a ({key_s1[9], key_s0[9]}), .c ({signal_1938, signal_925}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_725 ( .s (signal_693), .b ({key_s1[74], key_s0[74]}), .a ({key_s1[10], key_s0[10]}), .c ({signal_1941, signal_924}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_726 ( .s (signal_693), .b ({key_s1[75], key_s0[75]}), .a ({key_s1[11], key_s0[11]}), .c ({signal_1944, signal_923}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_727 ( .s (signal_693), .b ({key_s1[76], key_s0[76]}), .a ({key_s1[12], key_s0[12]}), .c ({signal_1947, signal_922}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_728 ( .s (signal_693), .b ({key_s1[77], key_s0[77]}), .a ({key_s1[13], key_s0[13]}), .c ({signal_1950, signal_921}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_729 ( .s (signal_693), .b ({key_s1[78], key_s0[78]}), .a ({key_s1[14], key_s0[14]}), .c ({signal_1953, signal_920}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_730 ( .s (signal_693), .b ({key_s1[79], key_s0[79]}), .a ({key_s1[15], key_s0[15]}), .c ({signal_1956, signal_919}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_731 ( .s (signal_693), .b ({key_s1[80], key_s0[80]}), .a ({key_s1[16], key_s0[16]}), .c ({signal_1959, signal_918}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_732 ( .s (signal_693), .b ({key_s1[81], key_s0[81]}), .a ({key_s1[17], key_s0[17]}), .c ({signal_1962, signal_917}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_733 ( .s (signal_693), .b ({key_s1[82], key_s0[82]}), .a ({key_s1[18], key_s0[18]}), .c ({signal_1965, signal_916}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_734 ( .s (signal_693), .b ({key_s1[83], key_s0[83]}), .a ({key_s1[19], key_s0[19]}), .c ({signal_1968, signal_915}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_735 ( .s (signal_693), .b ({key_s1[84], key_s0[84]}), .a ({key_s1[20], key_s0[20]}), .c ({signal_1971, signal_914}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_736 ( .s (signal_693), .b ({key_s1[85], key_s0[85]}), .a ({key_s1[21], key_s0[21]}), .c ({signal_1974, signal_913}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_737 ( .s (signal_1000), .b ({key_s1[86], key_s0[86]}), .a ({key_s1[22], key_s0[22]}), .c ({signal_1683, signal_912}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_738 ( .s (signal_1000), .b ({key_s1[87], key_s0[87]}), .a ({key_s1[23], key_s0[23]}), .c ({signal_1686, signal_911}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_739 ( .s (signal_1000), .b ({key_s1[88], key_s0[88]}), .a ({key_s1[24], key_s0[24]}), .c ({signal_1689, signal_910}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_740 ( .s (signal_1000), .b ({key_s1[89], key_s0[89]}), .a ({key_s1[25], key_s0[25]}), .c ({signal_1692, signal_909}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_741 ( .s (signal_1000), .b ({key_s1[90], key_s0[90]}), .a ({key_s1[26], key_s0[26]}), .c ({signal_1695, signal_908}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_742 ( .s (signal_1000), .b ({key_s1[91], key_s0[91]}), .a ({key_s1[27], key_s0[27]}), .c ({signal_1698, signal_907}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_743 ( .s (signal_694), .b ({key_s1[92], key_s0[92]}), .a ({key_s1[28], key_s0[28]}), .c ({signal_1977, signal_906}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_744 ( .s (signal_694), .b ({key_s1[93], key_s0[93]}), .a ({key_s1[29], key_s0[29]}), .c ({signal_1980, signal_905}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_745 ( .s (signal_694), .b ({key_s1[94], key_s0[94]}), .a ({key_s1[30], key_s0[30]}), .c ({signal_1983, signal_904}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_746 ( .s (signal_694), .b ({key_s1[95], key_s0[95]}), .a ({key_s1[31], key_s0[31]}), .c ({signal_1986, signal_903}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_747 ( .s (signal_694), .b ({key_s1[96], key_s0[96]}), .a ({key_s1[32], key_s0[32]}), .c ({signal_1989, signal_902}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_748 ( .s (signal_1000), .b ({key_s1[97], key_s0[97]}), .a ({key_s1[33], key_s0[33]}), .c ({signal_1701, signal_901}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_749 ( .s (signal_694), .b ({key_s1[98], key_s0[98]}), .a ({key_s1[34], key_s0[34]}), .c ({signal_1992, signal_900}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_750 ( .s (signal_694), .b ({key_s1[99], key_s0[99]}), .a ({key_s1[35], key_s0[35]}), .c ({signal_1995, signal_899}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_751 ( .s (signal_1000), .b ({key_s1[100], key_s0[100]}), .a ({key_s1[36], key_s0[36]}), .c ({signal_1704, signal_898}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_752 ( .s (signal_694), .b ({key_s1[101], key_s0[101]}), .a ({key_s1[37], key_s0[37]}), .c ({signal_1998, signal_897}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_753 ( .s (signal_694), .b ({key_s1[102], key_s0[102]}), .a ({key_s1[38], key_s0[38]}), .c ({signal_2001, signal_896}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_754 ( .s (signal_1000), .b ({key_s1[103], key_s0[103]}), .a ({key_s1[39], key_s0[39]}), .c ({signal_1707, signal_895}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_755 ( .s (signal_694), .b ({key_s1[104], key_s0[104]}), .a ({key_s1[40], key_s0[40]}), .c ({signal_2004, signal_894}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_756 ( .s (signal_694), .b ({key_s1[105], key_s0[105]}), .a ({key_s1[41], key_s0[41]}), .c ({signal_2007, signal_893}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_757 ( .s (signal_694), .b ({key_s1[106], key_s0[106]}), .a ({key_s1[42], key_s0[42]}), .c ({signal_2010, signal_892}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_758 ( .s (signal_694), .b ({key_s1[107], key_s0[107]}), .a ({key_s1[43], key_s0[43]}), .c ({signal_2013, signal_891}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_759 ( .s (signal_694), .b ({key_s1[108], key_s0[108]}), .a ({key_s1[44], key_s0[44]}), .c ({signal_2016, signal_890}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_760 ( .s (signal_694), .b ({key_s1[109], key_s0[109]}), .a ({key_s1[45], key_s0[45]}), .c ({signal_2019, signal_889}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_761 ( .s (signal_694), .b ({key_s1[110], key_s0[110]}), .a ({key_s1[46], key_s0[46]}), .c ({signal_2022, signal_888}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_762 ( .s (signal_694), .b ({key_s1[111], key_s0[111]}), .a ({key_s1[47], key_s0[47]}), .c ({signal_2025, signal_887}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_763 ( .s (signal_694), .b ({key_s1[112], key_s0[112]}), .a ({key_s1[48], key_s0[48]}), .c ({signal_2028, signal_886}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_764 ( .s (signal_694), .b ({key_s1[113], key_s0[113]}), .a ({key_s1[49], key_s0[49]}), .c ({signal_2031, signal_885}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_765 ( .s (signal_694), .b ({key_s1[114], key_s0[114]}), .a ({key_s1[50], key_s0[50]}), .c ({signal_2034, signal_884}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_766 ( .s (signal_694), .b ({key_s1[115], key_s0[115]}), .a ({key_s1[51], key_s0[51]}), .c ({signal_2037, signal_883}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_767 ( .s (signal_694), .b ({key_s1[116], key_s0[116]}), .a ({key_s1[52], key_s0[52]}), .c ({signal_2040, signal_882}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_768 ( .s (signal_1000), .b ({key_s1[117], key_s0[117]}), .a ({key_s1[53], key_s0[53]}), .c ({signal_1710, signal_881}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_769 ( .s (signal_1000), .b ({key_s1[118], key_s0[118]}), .a ({key_s1[54], key_s0[54]}), .c ({signal_1713, signal_880}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_770 ( .s (signal_694), .b ({key_s1[119], key_s0[119]}), .a ({key_s1[55], key_s0[55]}), .c ({signal_2043, signal_879}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_771 ( .s (signal_1000), .b ({key_s1[120], key_s0[120]}), .a ({key_s1[56], key_s0[56]}), .c ({signal_1716, signal_878}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_772 ( .s (signal_694), .b ({key_s1[121], key_s0[121]}), .a ({key_s1[57], key_s0[57]}), .c ({signal_2046, signal_877}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_773 ( .s (signal_694), .b ({key_s1[122], key_s0[122]}), .a ({key_s1[58], key_s0[58]}), .c ({signal_2049, signal_876}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_774 ( .s (signal_1000), .b ({key_s1[123], key_s0[123]}), .a ({key_s1[59], key_s0[59]}), .c ({signal_1719, signal_875}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_775 ( .s (signal_694), .b ({key_s1[124], key_s0[124]}), .a ({key_s1[60], key_s0[60]}), .c ({signal_2052, signal_874}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_776 ( .s (signal_694), .b ({key_s1[125], key_s0[125]}), .a ({key_s1[61], key_s0[61]}), .c ({signal_2055, signal_873}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_777 ( .s (signal_1000), .b ({key_s1[126], key_s0[126]}), .a ({key_s1[62], key_s0[62]}), .c ({signal_1722, signal_872}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_778 ( .s (signal_694), .b ({key_s1[127], key_s0[127]}), .a ({key_s1[63], key_s0[63]}), .c ({signal_2058, signal_871}) ) ;
    MUX2_X1 cell_779 ( .S (rst), .A (signal_1007), .B (1'b1), .Z (signal_266) ) ;
    MUX2_X1 cell_780 ( .S (rst), .A (signal_1006), .B (1'b0), .Z (signal_1014) ) ;
    MUX2_X1 cell_781 ( .S (rst), .A (signal_1005), .B (1'b0), .Z (signal_1013) ) ;
    MUX2_X1 cell_782 ( .S (rst), .A (signal_1004), .B (1'b1), .Z (signal_265) ) ;
    MUX2_X1 cell_783 ( .S (rst), .A (signal_1003), .B (1'b0), .Z (signal_1011) ) ;
    MUX2_X1 cell_784 ( .S (rst), .A (signal_1002), .B (1'b0), .Z (signal_1010) ) ;
    MUX2_X1 cell_785 ( .S (rst), .A (signal_1001), .B (1'b0), .Z (signal_1009) ) ;
    XOR2_X1 cell_786 ( .A (signal_265), .B (signal_1011), .Z (signal_1008) ) ;
    XOR2_X1 cell_787 ( .A (signal_1014), .B (signal_266), .Z (signal_1012) ) ;
    AND2_X1 cell_802 ( .A1 (signal_1009), .A2 (signal_702), .ZN (signal_267) ) ;
    NOR2_X1 cell_803 ( .A1 (signal_703), .A2 (signal_704), .ZN (signal_702) ) ;
    NAND2_X1 cell_804 ( .A1 (signal_705), .A2 (signal_706), .ZN (signal_704) ) ;
    NOR2_X1 cell_805 ( .A1 (signal_1011), .A2 (signal_1010), .ZN (signal_706) ) ;
    NOR2_X1 cell_806 ( .A1 (signal_1014), .A2 (signal_265), .ZN (signal_705) ) ;
    NAND2_X1 cell_807 ( .A1 (signal_266), .A2 (signal_1013), .ZN (signal_703) ) ;
    MUX2_X1 cell_808 ( .S (rst), .A (signal_1016), .B (1'b0), .Z (signal_1000) ) ;
    MUX2_X1 cell_809 ( .S (rst), .A (signal_1015), .B (1'b0), .Z (signal_999) ) ;
    XNOR2_X1 cell_810 ( .A (signal_707), .B (signal_999), .ZN (signal_1017) ) ;
    XNOR2_X1 cell_811 ( .A (signal_1000), .B (1'b0), .ZN (signal_707) ) ;
    INV_X1 cell_812 ( .A (signal_1000), .ZN (signal_1018) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_819 ( .a ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({signal_1516, signal_1019}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_820 ( .a ({ciphertext_s1[1], ciphertext_s0[1]}), .b ({signal_1518, signal_1020}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_821 ( .a ({ciphertext_s1[2], ciphertext_s0[2]}), .b ({signal_1520, signal_1021}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_822 ( .a ({ciphertext_s1[3], ciphertext_s0[3]}), .b ({signal_1522, signal_1022}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_823 ( .a ({ciphertext_s1[4], ciphertext_s0[4]}), .b ({signal_1524, signal_1023}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_824 ( .a ({ciphertext_s1[5], ciphertext_s0[5]}), .b ({signal_1526, signal_1024}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_825 ( .a ({ciphertext_s1[6], ciphertext_s0[6]}), .b ({signal_1528, signal_1025}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_826 ( .a ({ciphertext_s1[7], ciphertext_s0[7]}), .b ({signal_1530, signal_1026}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_827 ( .a ({ciphertext_s1[8], ciphertext_s0[8]}), .b ({signal_1532, signal_1027}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_828 ( .a ({ciphertext_s1[9], ciphertext_s0[9]}), .b ({signal_1534, signal_1028}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_829 ( .a ({ciphertext_s1[10], ciphertext_s0[10]}), .b ({signal_1536, signal_1029}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_830 ( .a ({ciphertext_s1[11], ciphertext_s0[11]}), .b ({signal_1538, signal_1030}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_831 ( .a ({ciphertext_s1[12], ciphertext_s0[12]}), .b ({signal_1540, signal_1031}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_832 ( .a ({ciphertext_s1[13], ciphertext_s0[13]}), .b ({signal_1542, signal_1032}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_833 ( .a ({ciphertext_s1[14], ciphertext_s0[14]}), .b ({signal_1544, signal_1033}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_834 ( .a ({ciphertext_s1[15], ciphertext_s0[15]}), .b ({signal_1546, signal_1034}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_835 ( .a ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({signal_1548, signal_1035}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_836 ( .a ({ciphertext_s1[17], ciphertext_s0[17]}), .b ({signal_1550, signal_1036}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_837 ( .a ({ciphertext_s1[18], ciphertext_s0[18]}), .b ({signal_1552, signal_1037}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_838 ( .a ({ciphertext_s1[19], ciphertext_s0[19]}), .b ({signal_1554, signal_1038}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_839 ( .a ({ciphertext_s1[20], ciphertext_s0[20]}), .b ({signal_1556, signal_1039}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_840 ( .a ({ciphertext_s1[21], ciphertext_s0[21]}), .b ({signal_1558, signal_1040}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_841 ( .a ({ciphertext_s1[22], ciphertext_s0[22]}), .b ({signal_1560, signal_1041}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_842 ( .a ({ciphertext_s1[23], ciphertext_s0[23]}), .b ({signal_1562, signal_1042}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_843 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({signal_1564, signal_1043}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_844 ( .a ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({signal_1566, signal_1044}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_845 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({signal_1568, signal_1045}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_846 ( .a ({ciphertext_s1[27], ciphertext_s0[27]}), .b ({signal_1570, signal_1046}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_847 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({signal_1572, signal_1047}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_848 ( .a ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({signal_1574, signal_1048}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_849 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({signal_1576, signal_1049}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_850 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({signal_1578, signal_1050}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_851 ( .a ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({signal_1580, signal_1051}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_852 ( .a ({ciphertext_s1[33], ciphertext_s0[33]}), .b ({signal_1582, signal_1052}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_853 ( .a ({ciphertext_s1[34], ciphertext_s0[34]}), .b ({signal_1584, signal_1053}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_854 ( .a ({ciphertext_s1[35], ciphertext_s0[35]}), .b ({signal_1586, signal_1054}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_855 ( .a ({ciphertext_s1[36], ciphertext_s0[36]}), .b ({signal_1588, signal_1055}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_856 ( .a ({ciphertext_s1[37], ciphertext_s0[37]}), .b ({signal_1590, signal_1056}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_857 ( .a ({ciphertext_s1[38], ciphertext_s0[38]}), .b ({signal_1592, signal_1057}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_858 ( .a ({ciphertext_s1[39], ciphertext_s0[39]}), .b ({signal_1594, signal_1058}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_859 ( .a ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({signal_1596, signal_1059}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_860 ( .a ({ciphertext_s1[41], ciphertext_s0[41]}), .b ({signal_1598, signal_1060}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_861 ( .a ({ciphertext_s1[42], ciphertext_s0[42]}), .b ({signal_1600, signal_1061}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_862 ( .a ({ciphertext_s1[43], ciphertext_s0[43]}), .b ({signal_1602, signal_1062}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_863 ( .a ({ciphertext_s1[44], ciphertext_s0[44]}), .b ({signal_1604, signal_1063}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_864 ( .a ({ciphertext_s1[45], ciphertext_s0[45]}), .b ({signal_1606, signal_1064}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_865 ( .a ({ciphertext_s1[46], ciphertext_s0[46]}), .b ({signal_1608, signal_1065}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_866 ( .a ({ciphertext_s1[47], ciphertext_s0[47]}), .b ({signal_1610, signal_1066}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_867 ( .a ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({signal_1612, signal_1067}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_868 ( .a ({ciphertext_s1[49], ciphertext_s0[49]}), .b ({signal_1614, signal_1068}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_869 ( .a ({ciphertext_s1[50], ciphertext_s0[50]}), .b ({signal_1616, signal_1069}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_870 ( .a ({ciphertext_s1[51], ciphertext_s0[51]}), .b ({signal_1618, signal_1070}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_871 ( .a ({ciphertext_s1[52], ciphertext_s0[52]}), .b ({signal_1620, signal_1071}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_872 ( .a ({ciphertext_s1[53], ciphertext_s0[53]}), .b ({signal_1622, signal_1072}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_873 ( .a ({ciphertext_s1[54], ciphertext_s0[54]}), .b ({signal_1624, signal_1073}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_874 ( .a ({ciphertext_s1[55], ciphertext_s0[55]}), .b ({signal_1626, signal_1074}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_875 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({signal_1628, signal_1075}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_876 ( .a ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({signal_1630, signal_1076}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_877 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({signal_1632, signal_1077}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_878 ( .a ({ciphertext_s1[59], ciphertext_s0[59]}), .b ({signal_1634, signal_1078}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_879 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({signal_1636, signal_1079}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_880 ( .a ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({signal_1638, signal_1080}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_881 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({signal_1640, signal_1081}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_882 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({signal_1642, signal_1082}) ) ;
    ClockGatingController #(9) cell_1379 ( .clk (clk), .rst (rst), .GatedClk (signal_2931), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_883 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .clk (clk), .r (Fresh[0]), .c ({signal_1643, signal_1083}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_884 ( .a ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({ciphertext_s1[51], ciphertext_s0[51]}), .clk (clk), .r (Fresh[1]), .c ({signal_1644, signal_1084}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_885 ( .a ({ciphertext_s1[52], ciphertext_s0[52]}), .b ({ciphertext_s1[55], ciphertext_s0[55]}), .clk (clk), .r (Fresh[2]), .c ({signal_1645, signal_1085}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_886 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .clk (clk), .r (Fresh[3]), .c ({signal_1646, signal_1086}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_887 ( .a ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({ciphertext_s1[35], ciphertext_s0[35]}), .clk (clk), .r (Fresh[4]), .c ({signal_1647, signal_1087}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_888 ( .a ({ciphertext_s1[44], ciphertext_s0[44]}), .b ({ciphertext_s1[47], ciphertext_s0[47]}), .clk (clk), .r (Fresh[5]), .c ({signal_1648, signal_1088}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_889 ( .a ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({ciphertext_s1[43], ciphertext_s0[43]}), .clk (clk), .r (Fresh[6]), .c ({signal_1649, signal_1089}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_890 ( .a ({ciphertext_s1[36], ciphertext_s0[36]}), .b ({ciphertext_s1[39], ciphertext_s0[39]}), .clk (clk), .r (Fresh[7]), .c ({signal_1650, signal_1090}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_891 ( .a ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({ciphertext_s1[19], ciphertext_s0[19]}), .clk (clk), .r (Fresh[8]), .c ({signal_1651, signal_1091}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_892 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .clk (clk), .r (Fresh[9]), .c ({signal_1652, signal_1092}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_893 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .clk (clk), .r (Fresh[10]), .c ({signal_1653, signal_1093}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_894 ( .a ({ciphertext_s1[20], ciphertext_s0[20]}), .b ({ciphertext_s1[23], ciphertext_s0[23]}), .clk (clk), .r (Fresh[11]), .c ({signal_1654, signal_1094}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_895 ( .a ({ciphertext_s1[4], ciphertext_s0[4]}), .b ({ciphertext_s1[7], ciphertext_s0[7]}), .clk (clk), .r (Fresh[12]), .c ({signal_1655, signal_1095}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_896 ( .a ({ciphertext_s1[8], ciphertext_s0[8]}), .b ({ciphertext_s1[11], ciphertext_s0[11]}), .clk (clk), .r (Fresh[13]), .c ({signal_1656, signal_1096}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_897 ( .a ({ciphertext_s1[12], ciphertext_s0[12]}), .b ({ciphertext_s1[15], ciphertext_s0[15]}), .clk (clk), .r (Fresh[14]), .c ({signal_1657, signal_1097}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_898 ( .a ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({ciphertext_s1[3], ciphertext_s0[3]}), .clk (clk), .r (Fresh[15]), .c ({signal_1658, signal_1098}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_899 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .clk (clk), .r (Fresh[16]), .c ({signal_1659, signal_1099}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_900 ( .a ({ciphertext_s1[50], ciphertext_s0[50]}), .b ({ciphertext_s1[51], ciphertext_s0[51]}), .clk (clk), .r (Fresh[17]), .c ({signal_1660, signal_1100}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_901 ( .a ({ciphertext_s1[54], ciphertext_s0[54]}), .b ({ciphertext_s1[55], ciphertext_s0[55]}), .clk (clk), .r (Fresh[18]), .c ({signal_1661, signal_1101}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_902 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .clk (clk), .r (Fresh[19]), .c ({signal_1662, signal_1102}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_903 ( .a ({ciphertext_s1[34], ciphertext_s0[34]}), .b ({ciphertext_s1[35], ciphertext_s0[35]}), .clk (clk), .r (Fresh[20]), .c ({signal_1663, signal_1103}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_904 ( .a ({ciphertext_s1[46], ciphertext_s0[46]}), .b ({ciphertext_s1[47], ciphertext_s0[47]}), .clk (clk), .r (Fresh[21]), .c ({signal_1664, signal_1104}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_905 ( .a ({ciphertext_s1[42], ciphertext_s0[42]}), .b ({ciphertext_s1[43], ciphertext_s0[43]}), .clk (clk), .r (Fresh[22]), .c ({signal_1665, signal_1105}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_906 ( .a ({ciphertext_s1[38], ciphertext_s0[38]}), .b ({ciphertext_s1[39], ciphertext_s0[39]}), .clk (clk), .r (Fresh[23]), .c ({signal_1666, signal_1106}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_907 ( .a ({ciphertext_s1[18], ciphertext_s0[18]}), .b ({ciphertext_s1[19], ciphertext_s0[19]}), .clk (clk), .r (Fresh[24]), .c ({signal_1667, signal_1107}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_908 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .clk (clk), .r (Fresh[25]), .c ({signal_1668, signal_1108}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_909 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .clk (clk), .r (Fresh[26]), .c ({signal_1669, signal_1109}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_910 ( .a ({ciphertext_s1[22], ciphertext_s0[22]}), .b ({ciphertext_s1[23], ciphertext_s0[23]}), .clk (clk), .r (Fresh[27]), .c ({signal_1670, signal_1110}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_911 ( .a ({ciphertext_s1[6], ciphertext_s0[6]}), .b ({ciphertext_s1[7], ciphertext_s0[7]}), .clk (clk), .r (Fresh[28]), .c ({signal_1671, signal_1111}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_912 ( .a ({ciphertext_s1[10], ciphertext_s0[10]}), .b ({ciphertext_s1[11], ciphertext_s0[11]}), .clk (clk), .r (Fresh[29]), .c ({signal_1672, signal_1112}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_913 ( .a ({ciphertext_s1[14], ciphertext_s0[14]}), .b ({ciphertext_s1[15], ciphertext_s0[15]}), .clk (clk), .r (Fresh[30]), .c ({signal_1673, signal_1113}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_914 ( .a ({ciphertext_s1[2], ciphertext_s0[2]}), .b ({ciphertext_s1[3], ciphertext_s0[3]}), .clk (clk), .r (Fresh[31]), .c ({signal_1674, signal_1114}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_915 ( .a ({signal_1643, signal_1083}), .b ({signal_1723, signal_1115}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_916 ( .a ({signal_1644, signal_1084}), .b ({signal_1724, signal_1116}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_917 ( .a ({signal_1645, signal_1085}), .b ({signal_1725, signal_1117}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_918 ( .a ({signal_1646, signal_1086}), .b ({signal_1726, signal_1118}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_919 ( .a ({signal_1647, signal_1087}), .b ({signal_1727, signal_1119}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_920 ( .a ({signal_1648, signal_1088}), .b ({signal_1728, signal_1120}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_921 ( .a ({signal_1649, signal_1089}), .b ({signal_1729, signal_1121}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_922 ( .a ({signal_1650, signal_1090}), .b ({signal_1730, signal_1122}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_923 ( .a ({signal_1651, signal_1091}), .b ({signal_1731, signal_1123}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_924 ( .a ({signal_1652, signal_1092}), .b ({signal_1732, signal_1124}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_925 ( .a ({signal_1653, signal_1093}), .b ({signal_1733, signal_1125}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_926 ( .a ({signal_1654, signal_1094}), .b ({signal_1734, signal_1126}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_927 ( .a ({signal_1655, signal_1095}), .b ({signal_1735, signal_1127}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_928 ( .a ({signal_1656, signal_1096}), .b ({signal_1736, signal_1128}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_929 ( .a ({signal_1657, signal_1097}), .b ({signal_1737, signal_1129}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_930 ( .a ({signal_1658, signal_1098}), .b ({signal_1738, signal_1130}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_931 ( .a ({signal_1659, signal_1099}), .b ({signal_1739, signal_1131}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_932 ( .a ({signal_1660, signal_1100}), .b ({signal_1740, signal_1132}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_933 ( .a ({signal_1661, signal_1101}), .b ({signal_1741, signal_1133}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_934 ( .a ({signal_1662, signal_1102}), .b ({signal_1742, signal_1134}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_935 ( .a ({signal_1663, signal_1103}), .b ({signal_1743, signal_1135}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_936 ( .a ({signal_1664, signal_1104}), .b ({signal_1744, signal_1136}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_937 ( .a ({signal_1665, signal_1105}), .b ({signal_1745, signal_1137}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_938 ( .a ({signal_1666, signal_1106}), .b ({signal_1746, signal_1138}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_939 ( .a ({signal_1667, signal_1107}), .b ({signal_1747, signal_1139}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_940 ( .a ({signal_1668, signal_1108}), .b ({signal_1748, signal_1140}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_941 ( .a ({signal_1669, signal_1109}), .b ({signal_1749, signal_1141}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_942 ( .a ({signal_1670, signal_1110}), .b ({signal_1750, signal_1142}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_943 ( .a ({signal_1671, signal_1111}), .b ({signal_1751, signal_1143}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_944 ( .a ({signal_1672, signal_1112}), .b ({signal_1752, signal_1144}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_945 ( .a ({signal_1673, signal_1113}), .b ({signal_1753, signal_1145}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_946 ( .a ({signal_1674, signal_1114}), .b ({signal_1754, signal_1146}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_947 ( .a ({signal_1640, signal_1081}), .b ({signal_1642, signal_1082}), .clk (clk), .r (Fresh[32]), .c ({signal_1755, signal_1147}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_948 ( .a ({signal_1616, signal_1069}), .b ({signal_1618, signal_1070}), .clk (clk), .r (Fresh[33]), .c ({signal_1756, signal_1148}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_949 ( .a ({signal_1624, signal_1073}), .b ({signal_1626, signal_1074}), .clk (clk), .r (Fresh[34]), .c ({signal_1757, signal_1149}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_950 ( .a ({signal_1632, signal_1077}), .b ({signal_1634, signal_1078}), .clk (clk), .r (Fresh[35]), .c ({signal_1758, signal_1150}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_951 ( .a ({signal_1584, signal_1053}), .b ({signal_1586, signal_1054}), .clk (clk), .r (Fresh[36]), .c ({signal_1759, signal_1151}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_952 ( .a ({signal_1608, signal_1065}), .b ({signal_1610, signal_1066}), .clk (clk), .r (Fresh[37]), .c ({signal_1760, signal_1152}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_953 ( .a ({signal_1600, signal_1061}), .b ({signal_1602, signal_1062}), .clk (clk), .r (Fresh[38]), .c ({signal_1761, signal_1153}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_954 ( .a ({signal_1592, signal_1057}), .b ({signal_1594, signal_1058}), .clk (clk), .r (Fresh[39]), .c ({signal_1762, signal_1154}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_955 ( .a ({signal_1552, signal_1037}), .b ({signal_1554, signal_1038}), .clk (clk), .r (Fresh[40]), .c ({signal_1763, signal_1155}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_956 ( .a ({signal_1576, signal_1049}), .b ({signal_1578, signal_1050}), .clk (clk), .r (Fresh[41]), .c ({signal_1764, signal_1156}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_957 ( .a ({signal_1568, signal_1045}), .b ({signal_1570, signal_1046}), .clk (clk), .r (Fresh[42]), .c ({signal_1765, signal_1157}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_958 ( .a ({signal_1560, signal_1041}), .b ({signal_1562, signal_1042}), .clk (clk), .r (Fresh[43]), .c ({signal_1766, signal_1158}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_959 ( .a ({signal_1528, signal_1025}), .b ({signal_1530, signal_1026}), .clk (clk), .r (Fresh[44]), .c ({signal_1767, signal_1159}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_960 ( .a ({signal_1536, signal_1029}), .b ({signal_1538, signal_1030}), .clk (clk), .r (Fresh[45]), .c ({signal_1768, signal_1160}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_961 ( .a ({signal_1544, signal_1033}), .b ({signal_1546, signal_1034}), .clk (clk), .r (Fresh[46]), .c ({signal_1769, signal_1161}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_962 ( .a ({signal_1520, signal_1021}), .b ({signal_1522, signal_1022}), .clk (clk), .r (Fresh[47]), .c ({signal_1770, signal_1162}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_963 ( .a ({signal_1636, signal_1079}), .b ({signal_1642, signal_1082}), .clk (clk), .r (Fresh[48]), .c ({signal_1771, signal_1163}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_964 ( .a ({signal_1640, signal_1081}), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .clk (clk), .r (Fresh[49]), .c ({signal_1772, signal_1164}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_965 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({signal_1642, signal_1082}), .clk (clk), .r (Fresh[50]), .c ({signal_1773, signal_1165}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_966 ( .a ({signal_1612, signal_1067}), .b ({signal_1618, signal_1070}), .clk (clk), .r (Fresh[51]), .c ({signal_1774, signal_1166}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_967 ( .a ({signal_1616, signal_1069}), .b ({ciphertext_s1[51], ciphertext_s0[51]}), .clk (clk), .r (Fresh[52]), .c ({signal_1775, signal_1167}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_968 ( .a ({ciphertext_s1[50], ciphertext_s0[50]}), .b ({signal_1618, signal_1070}), .clk (clk), .r (Fresh[53]), .c ({signal_1776, signal_1168}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_969 ( .a ({signal_1620, signal_1071}), .b ({signal_1626, signal_1074}), .clk (clk), .r (Fresh[54]), .c ({signal_1777, signal_1169}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_970 ( .a ({signal_1624, signal_1073}), .b ({ciphertext_s1[55], ciphertext_s0[55]}), .clk (clk), .r (Fresh[55]), .c ({signal_1778, signal_1170}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_971 ( .a ({ciphertext_s1[54], ciphertext_s0[54]}), .b ({signal_1626, signal_1074}), .clk (clk), .r (Fresh[56]), .c ({signal_1779, signal_1171}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_972 ( .a ({signal_1628, signal_1075}), .b ({signal_1634, signal_1078}), .clk (clk), .r (Fresh[57]), .c ({signal_1780, signal_1172}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_973 ( .a ({signal_1632, signal_1077}), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .clk (clk), .r (Fresh[58]), .c ({signal_1781, signal_1173}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_974 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({signal_1634, signal_1078}), .clk (clk), .r (Fresh[59]), .c ({signal_1782, signal_1174}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_975 ( .a ({signal_1580, signal_1051}), .b ({signal_1586, signal_1054}), .clk (clk), .r (Fresh[60]), .c ({signal_1783, signal_1175}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_976 ( .a ({signal_1584, signal_1053}), .b ({ciphertext_s1[35], ciphertext_s0[35]}), .clk (clk), .r (Fresh[61]), .c ({signal_1784, signal_1176}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_977 ( .a ({ciphertext_s1[34], ciphertext_s0[34]}), .b ({signal_1586, signal_1054}), .clk (clk), .r (Fresh[62]), .c ({signal_1785, signal_1177}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_978 ( .a ({signal_1604, signal_1063}), .b ({signal_1610, signal_1066}), .clk (clk), .r (Fresh[63]), .c ({signal_1786, signal_1178}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_979 ( .a ({signal_1608, signal_1065}), .b ({ciphertext_s1[47], ciphertext_s0[47]}), .clk (clk), .r (Fresh[64]), .c ({signal_1787, signal_1179}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_980 ( .a ({ciphertext_s1[46], ciphertext_s0[46]}), .b ({signal_1610, signal_1066}), .clk (clk), .r (Fresh[65]), .c ({signal_1788, signal_1180}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_981 ( .a ({signal_1596, signal_1059}), .b ({signal_1602, signal_1062}), .clk (clk), .r (Fresh[66]), .c ({signal_1789, signal_1181}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_982 ( .a ({signal_1600, signal_1061}), .b ({ciphertext_s1[43], ciphertext_s0[43]}), .clk (clk), .r (Fresh[67]), .c ({signal_1790, signal_1182}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_983 ( .a ({ciphertext_s1[42], ciphertext_s0[42]}), .b ({signal_1602, signal_1062}), .clk (clk), .r (Fresh[68]), .c ({signal_1791, signal_1183}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_984 ( .a ({signal_1588, signal_1055}), .b ({signal_1594, signal_1058}), .clk (clk), .r (Fresh[69]), .c ({signal_1792, signal_1184}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_985 ( .a ({signal_1592, signal_1057}), .b ({ciphertext_s1[39], ciphertext_s0[39]}), .clk (clk), .r (Fresh[70]), .c ({signal_1793, signal_1185}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_986 ( .a ({ciphertext_s1[38], ciphertext_s0[38]}), .b ({signal_1594, signal_1058}), .clk (clk), .r (Fresh[71]), .c ({signal_1794, signal_1186}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_987 ( .a ({signal_1548, signal_1035}), .b ({signal_1554, signal_1038}), .clk (clk), .r (Fresh[72]), .c ({signal_1795, signal_1187}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_988 ( .a ({signal_1552, signal_1037}), .b ({ciphertext_s1[19], ciphertext_s0[19]}), .clk (clk), .r (Fresh[73]), .c ({signal_1796, signal_1188}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_989 ( .a ({ciphertext_s1[18], ciphertext_s0[18]}), .b ({signal_1554, signal_1038}), .clk (clk), .r (Fresh[74]), .c ({signal_1797, signal_1189}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_990 ( .a ({signal_1572, signal_1047}), .b ({signal_1578, signal_1050}), .clk (clk), .r (Fresh[75]), .c ({signal_1798, signal_1190}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_991 ( .a ({signal_1576, signal_1049}), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .clk (clk), .r (Fresh[76]), .c ({signal_1799, signal_1191}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_992 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({signal_1578, signal_1050}), .clk (clk), .r (Fresh[77]), .c ({signal_1800, signal_1192}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_993 ( .a ({signal_1564, signal_1043}), .b ({signal_1570, signal_1046}), .clk (clk), .r (Fresh[78]), .c ({signal_1801, signal_1193}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_994 ( .a ({signal_1568, signal_1045}), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .clk (clk), .r (Fresh[79]), .c ({signal_1802, signal_1194}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_995 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({signal_1570, signal_1046}), .clk (clk), .r (Fresh[80]), .c ({signal_1803, signal_1195}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_996 ( .a ({signal_1556, signal_1039}), .b ({signal_1562, signal_1042}), .clk (clk), .r (Fresh[81]), .c ({signal_1804, signal_1196}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_997 ( .a ({signal_1560, signal_1041}), .b ({ciphertext_s1[23], ciphertext_s0[23]}), .clk (clk), .r (Fresh[82]), .c ({signal_1805, signal_1197}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_998 ( .a ({ciphertext_s1[22], ciphertext_s0[22]}), .b ({signal_1562, signal_1042}), .clk (clk), .r (Fresh[83]), .c ({signal_1806, signal_1198}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_999 ( .a ({signal_1524, signal_1023}), .b ({signal_1530, signal_1026}), .clk (clk), .r (Fresh[84]), .c ({signal_1807, signal_1199}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1000 ( .a ({signal_1528, signal_1025}), .b ({ciphertext_s1[7], ciphertext_s0[7]}), .clk (clk), .r (Fresh[85]), .c ({signal_1808, signal_1200}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1001 ( .a ({ciphertext_s1[6], ciphertext_s0[6]}), .b ({signal_1530, signal_1026}), .clk (clk), .r (Fresh[86]), .c ({signal_1809, signal_1201}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1002 ( .a ({signal_1532, signal_1027}), .b ({signal_1538, signal_1030}), .clk (clk), .r (Fresh[87]), .c ({signal_1810, signal_1202}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1003 ( .a ({signal_1536, signal_1029}), .b ({ciphertext_s1[11], ciphertext_s0[11]}), .clk (clk), .r (Fresh[88]), .c ({signal_1811, signal_1203}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1004 ( .a ({ciphertext_s1[10], ciphertext_s0[10]}), .b ({signal_1538, signal_1030}), .clk (clk), .r (Fresh[89]), .c ({signal_1812, signal_1204}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1005 ( .a ({signal_1540, signal_1031}), .b ({signal_1546, signal_1034}), .clk (clk), .r (Fresh[90]), .c ({signal_1813, signal_1205}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1006 ( .a ({signal_1544, signal_1033}), .b ({ciphertext_s1[15], ciphertext_s0[15]}), .clk (clk), .r (Fresh[91]), .c ({signal_1814, signal_1206}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1007 ( .a ({ciphertext_s1[14], ciphertext_s0[14]}), .b ({signal_1546, signal_1034}), .clk (clk), .r (Fresh[92]), .c ({signal_1815, signal_1207}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1008 ( .a ({signal_1516, signal_1019}), .b ({signal_1522, signal_1022}), .clk (clk), .r (Fresh[93]), .c ({signal_1816, signal_1208}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1009 ( .a ({signal_1520, signal_1021}), .b ({ciphertext_s1[3], ciphertext_s0[3]}), .clk (clk), .r (Fresh[94]), .c ({signal_1817, signal_1209}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1010 ( .a ({ciphertext_s1[2], ciphertext_s0[2]}), .b ({signal_1522, signal_1022}), .clk (clk), .r (Fresh[95]), .c ({signal_1818, signal_1210}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1011 ( .a ({signal_1755, signal_1147}), .b ({signal_1819, signal_1211}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1012 ( .a ({signal_1756, signal_1148}), .b ({signal_1820, signal_1212}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1013 ( .a ({signal_1757, signal_1149}), .b ({signal_1821, signal_1213}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1014 ( .a ({signal_1758, signal_1150}), .b ({signal_1822, signal_1214}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1015 ( .a ({signal_1759, signal_1151}), .b ({signal_1823, signal_1215}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1016 ( .a ({signal_1760, signal_1152}), .b ({signal_1824, signal_1216}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1017 ( .a ({signal_1761, signal_1153}), .b ({signal_1825, signal_1217}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1018 ( .a ({signal_1762, signal_1154}), .b ({signal_1826, signal_1218}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1019 ( .a ({signal_1763, signal_1155}), .b ({signal_1827, signal_1219}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1020 ( .a ({signal_1764, signal_1156}), .b ({signal_1828, signal_1220}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1021 ( .a ({signal_1765, signal_1157}), .b ({signal_1829, signal_1221}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1022 ( .a ({signal_1766, signal_1158}), .b ({signal_1830, signal_1222}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1023 ( .a ({signal_1767, signal_1159}), .b ({signal_1831, signal_1223}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1024 ( .a ({signal_1768, signal_1160}), .b ({signal_1832, signal_1224}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1025 ( .a ({signal_1769, signal_1161}), .b ({signal_1833, signal_1225}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1026 ( .a ({signal_1770, signal_1162}), .b ({signal_1834, signal_1226}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1027 ( .a ({signal_1771, signal_1163}), .b ({signal_1835, signal_1227}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1028 ( .a ({signal_1772, signal_1164}), .b ({signal_1836, signal_1228}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1029 ( .a ({signal_1773, signal_1165}), .b ({signal_1837, signal_1229}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1030 ( .a ({signal_1774, signal_1166}), .b ({signal_1838, signal_1230}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1031 ( .a ({signal_1775, signal_1167}), .b ({signal_1839, signal_1231}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1032 ( .a ({signal_1776, signal_1168}), .b ({signal_1840, signal_1232}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1033 ( .a ({signal_1777, signal_1169}), .b ({signal_1841, signal_1233}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1034 ( .a ({signal_1778, signal_1170}), .b ({signal_1842, signal_1234}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1035 ( .a ({signal_1779, signal_1171}), .b ({signal_1843, signal_1235}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1036 ( .a ({signal_1780, signal_1172}), .b ({signal_1844, signal_1236}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1037 ( .a ({signal_1781, signal_1173}), .b ({signal_1845, signal_1237}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1038 ( .a ({signal_1782, signal_1174}), .b ({signal_1846, signal_1238}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1039 ( .a ({signal_1783, signal_1175}), .b ({signal_1847, signal_1239}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1040 ( .a ({signal_1784, signal_1176}), .b ({signal_1848, signal_1240}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1041 ( .a ({signal_1785, signal_1177}), .b ({signal_1849, signal_1241}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1042 ( .a ({signal_1786, signal_1178}), .b ({signal_1850, signal_1242}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1043 ( .a ({signal_1787, signal_1179}), .b ({signal_1851, signal_1243}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1044 ( .a ({signal_1788, signal_1180}), .b ({signal_1852, signal_1244}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1045 ( .a ({signal_1789, signal_1181}), .b ({signal_1853, signal_1245}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1046 ( .a ({signal_1790, signal_1182}), .b ({signal_1854, signal_1246}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1047 ( .a ({signal_1791, signal_1183}), .b ({signal_1855, signal_1247}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1048 ( .a ({signal_1792, signal_1184}), .b ({signal_1856, signal_1248}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1049 ( .a ({signal_1793, signal_1185}), .b ({signal_1857, signal_1249}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1050 ( .a ({signal_1794, signal_1186}), .b ({signal_1858, signal_1250}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1051 ( .a ({signal_1795, signal_1187}), .b ({signal_1859, signal_1251}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1052 ( .a ({signal_1796, signal_1188}), .b ({signal_1860, signal_1252}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1053 ( .a ({signal_1797, signal_1189}), .b ({signal_1861, signal_1253}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1054 ( .a ({signal_1798, signal_1190}), .b ({signal_1862, signal_1254}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1055 ( .a ({signal_1799, signal_1191}), .b ({signal_1863, signal_1255}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1056 ( .a ({signal_1800, signal_1192}), .b ({signal_1864, signal_1256}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1057 ( .a ({signal_1801, signal_1193}), .b ({signal_1865, signal_1257}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1058 ( .a ({signal_1802, signal_1194}), .b ({signal_1866, signal_1258}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1059 ( .a ({signal_1803, signal_1195}), .b ({signal_1867, signal_1259}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1060 ( .a ({signal_1804, signal_1196}), .b ({signal_1868, signal_1260}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1061 ( .a ({signal_1805, signal_1197}), .b ({signal_1869, signal_1261}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1062 ( .a ({signal_1806, signal_1198}), .b ({signal_1870, signal_1262}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1063 ( .a ({signal_1807, signal_1199}), .b ({signal_1871, signal_1263}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1064 ( .a ({signal_1808, signal_1200}), .b ({signal_1872, signal_1264}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1065 ( .a ({signal_1809, signal_1201}), .b ({signal_1873, signal_1265}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1066 ( .a ({signal_1810, signal_1202}), .b ({signal_1874, signal_1266}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1067 ( .a ({signal_1811, signal_1203}), .b ({signal_1875, signal_1267}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1068 ( .a ({signal_1812, signal_1204}), .b ({signal_1876, signal_1268}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1069 ( .a ({signal_1813, signal_1205}), .b ({signal_1877, signal_1269}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1070 ( .a ({signal_1814, signal_1206}), .b ({signal_1878, signal_1270}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1071 ( .a ({signal_1815, signal_1207}), .b ({signal_1879, signal_1271}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1072 ( .a ({signal_1816, signal_1208}), .b ({signal_1880, signal_1272}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1073 ( .a ({signal_1817, signal_1209}), .b ({signal_1881, signal_1273}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1074 ( .a ({signal_1818, signal_1210}), .b ({signal_1882, signal_1274}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1075 ( .a ({signal_1640, signal_1081}), .b ({signal_1723, signal_1115}), .clk (clk), .r (Fresh[96]), .c ({signal_1883, signal_1275}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1076 ( .a ({signal_1616, signal_1069}), .b ({signal_1724, signal_1116}), .clk (clk), .r (Fresh[97]), .c ({signal_1884, signal_1276}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1077 ( .a ({signal_1624, signal_1073}), .b ({signal_1725, signal_1117}), .clk (clk), .r (Fresh[98]), .c ({signal_1885, signal_1277}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1078 ( .a ({signal_1632, signal_1077}), .b ({signal_1726, signal_1118}), .clk (clk), .r (Fresh[99]), .c ({signal_1886, signal_1278}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1079 ( .a ({signal_1584, signal_1053}), .b ({signal_1727, signal_1119}), .clk (clk), .r (Fresh[100]), .c ({signal_1887, signal_1279}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1080 ( .a ({signal_1608, signal_1065}), .b ({signal_1728, signal_1120}), .clk (clk), .r (Fresh[101]), .c ({signal_1888, signal_1280}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1081 ( .a ({signal_1600, signal_1061}), .b ({signal_1729, signal_1121}), .clk (clk), .r (Fresh[102]), .c ({signal_1889, signal_1281}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1082 ( .a ({signal_1592, signal_1057}), .b ({signal_1730, signal_1122}), .clk (clk), .r (Fresh[103]), .c ({signal_1890, signal_1282}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1083 ( .a ({signal_1552, signal_1037}), .b ({signal_1731, signal_1123}), .clk (clk), .r (Fresh[104]), .c ({signal_1891, signal_1283}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1084 ( .a ({signal_1576, signal_1049}), .b ({signal_1732, signal_1124}), .clk (clk), .r (Fresh[105]), .c ({signal_1892, signal_1284}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1085 ( .a ({signal_1568, signal_1045}), .b ({signal_1733, signal_1125}), .clk (clk), .r (Fresh[106]), .c ({signal_1893, signal_1285}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1086 ( .a ({signal_1560, signal_1041}), .b ({signal_1734, signal_1126}), .clk (clk), .r (Fresh[107]), .c ({signal_1894, signal_1286}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1087 ( .a ({signal_1528, signal_1025}), .b ({signal_1735, signal_1127}), .clk (clk), .r (Fresh[108]), .c ({signal_1895, signal_1287}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1088 ( .a ({signal_1536, signal_1029}), .b ({signal_1736, signal_1128}), .clk (clk), .r (Fresh[109]), .c ({signal_1896, signal_1288}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1089 ( .a ({signal_1544, signal_1033}), .b ({signal_1737, signal_1129}), .clk (clk), .r (Fresh[110]), .c ({signal_1897, signal_1289}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1090 ( .a ({signal_1520, signal_1021}), .b ({signal_1738, signal_1130}), .clk (clk), .r (Fresh[111]), .c ({signal_1898, signal_1290}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1091 ( .a ({signal_1638, signal_1080}), .b ({signal_1739, signal_1131}), .clk (clk), .r (Fresh[112]), .c ({signal_1899, signal_1291}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1092 ( .a ({signal_1614, signal_1068}), .b ({signal_1740, signal_1132}), .clk (clk), .r (Fresh[113]), .c ({signal_1900, signal_1292}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1093 ( .a ({signal_1622, signal_1072}), .b ({signal_1741, signal_1133}), .clk (clk), .r (Fresh[114]), .c ({signal_1901, signal_1293}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1094 ( .a ({signal_1630, signal_1076}), .b ({signal_1742, signal_1134}), .clk (clk), .r (Fresh[115]), .c ({signal_1902, signal_1294}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1095 ( .a ({signal_1582, signal_1052}), .b ({signal_1743, signal_1135}), .clk (clk), .r (Fresh[116]), .c ({signal_1903, signal_1295}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1096 ( .a ({signal_1606, signal_1064}), .b ({signal_1744, signal_1136}), .clk (clk), .r (Fresh[117]), .c ({signal_1904, signal_1296}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1097 ( .a ({signal_1598, signal_1060}), .b ({signal_1745, signal_1137}), .clk (clk), .r (Fresh[118]), .c ({signal_1905, signal_1297}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1098 ( .a ({signal_1590, signal_1056}), .b ({signal_1746, signal_1138}), .clk (clk), .r (Fresh[119]), .c ({signal_1906, signal_1298}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1099 ( .a ({signal_1550, signal_1036}), .b ({signal_1747, signal_1139}), .clk (clk), .r (Fresh[120]), .c ({signal_1907, signal_1299}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1100 ( .a ({signal_1574, signal_1048}), .b ({signal_1748, signal_1140}), .clk (clk), .r (Fresh[121]), .c ({signal_1908, signal_1300}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1101 ( .a ({signal_1566, signal_1044}), .b ({signal_1749, signal_1141}), .clk (clk), .r (Fresh[122]), .c ({signal_1909, signal_1301}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1102 ( .a ({signal_1558, signal_1040}), .b ({signal_1750, signal_1142}), .clk (clk), .r (Fresh[123]), .c ({signal_1910, signal_1302}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1103 ( .a ({signal_1526, signal_1024}), .b ({signal_1751, signal_1143}), .clk (clk), .r (Fresh[124]), .c ({signal_1911, signal_1303}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1104 ( .a ({signal_1534, signal_1028}), .b ({signal_1752, signal_1144}), .clk (clk), .r (Fresh[125]), .c ({signal_1912, signal_1304}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1105 ( .a ({signal_1542, signal_1032}), .b ({signal_1753, signal_1145}), .clk (clk), .r (Fresh[126]), .c ({signal_1913, signal_1305}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1106 ( .a ({signal_1518, signal_1020}), .b ({signal_1754, signal_1146}), .clk (clk), .r (Fresh[127]), .c ({signal_1914, signal_1306}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1107 ( .a ({signal_1883, signal_1275}), .b ({signal_2059, signal_1307}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1108 ( .a ({signal_1884, signal_1276}), .b ({signal_2060, signal_1308}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1109 ( .a ({signal_1885, signal_1277}), .b ({signal_2061, signal_1309}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1110 ( .a ({signal_1886, signal_1278}), .b ({signal_2062, signal_1310}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1111 ( .a ({signal_1887, signal_1279}), .b ({signal_2063, signal_1311}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1112 ( .a ({signal_1888, signal_1280}), .b ({signal_2064, signal_1312}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1113 ( .a ({signal_1889, signal_1281}), .b ({signal_2065, signal_1313}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1114 ( .a ({signal_1890, signal_1282}), .b ({signal_2066, signal_1314}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1115 ( .a ({signal_1891, signal_1283}), .b ({signal_2067, signal_1315}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1116 ( .a ({signal_1892, signal_1284}), .b ({signal_2068, signal_1316}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1117 ( .a ({signal_1893, signal_1285}), .b ({signal_2069, signal_1317}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1118 ( .a ({signal_1894, signal_1286}), .b ({signal_2070, signal_1318}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1119 ( .a ({signal_1895, signal_1287}), .b ({signal_2071, signal_1319}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1120 ( .a ({signal_1896, signal_1288}), .b ({signal_2072, signal_1320}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1121 ( .a ({signal_1897, signal_1289}), .b ({signal_2073, signal_1321}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1122 ( .a ({signal_1898, signal_1290}), .b ({signal_2074, signal_1322}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1123 ( .a ({signal_1899, signal_1291}), .b ({signal_2075, signal_1323}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1124 ( .a ({signal_1900, signal_1292}), .b ({signal_2076, signal_1324}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1125 ( .a ({signal_1901, signal_1293}), .b ({signal_2077, signal_1325}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1126 ( .a ({signal_1902, signal_1294}), .b ({signal_2078, signal_1326}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1127 ( .a ({signal_1903, signal_1295}), .b ({signal_2079, signal_1327}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1128 ( .a ({signal_1904, signal_1296}), .b ({signal_2080, signal_1328}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1129 ( .a ({signal_1905, signal_1297}), .b ({signal_2081, signal_1329}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1130 ( .a ({signal_1906, signal_1298}), .b ({signal_2082, signal_1330}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1131 ( .a ({signal_1907, signal_1299}), .b ({signal_2083, signal_1331}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1132 ( .a ({signal_1908, signal_1300}), .b ({signal_2084, signal_1332}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1133 ( .a ({signal_1909, signal_1301}), .b ({signal_2085, signal_1333}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1134 ( .a ({signal_1910, signal_1302}), .b ({signal_2086, signal_1334}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1135 ( .a ({signal_1911, signal_1303}), .b ({signal_2087, signal_1335}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1136 ( .a ({signal_1912, signal_1304}), .b ({signal_2088, signal_1336}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1137 ( .a ({signal_1913, signal_1305}), .b ({signal_2089, signal_1337}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1138 ( .a ({signal_1914, signal_1306}), .b ({signal_2090, signal_1338}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1139 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({signal_1819, signal_1211}), .clk (clk), .r (Fresh[128]), .c ({signal_2091, signal_1339}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1140 ( .a ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({signal_1820, signal_1212}), .clk (clk), .r (Fresh[129]), .c ({signal_2092, signal_1340}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1141 ( .a ({ciphertext_s1[52], ciphertext_s0[52]}), .b ({signal_1821, signal_1213}), .clk (clk), .r (Fresh[130]), .c ({signal_2093, signal_1341}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1142 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({signal_1822, signal_1214}), .clk (clk), .r (Fresh[131]), .c ({signal_2094, signal_1342}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1143 ( .a ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({signal_1823, signal_1215}), .clk (clk), .r (Fresh[132]), .c ({signal_2095, signal_1343}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1144 ( .a ({ciphertext_s1[44], ciphertext_s0[44]}), .b ({signal_1824, signal_1216}), .clk (clk), .r (Fresh[133]), .c ({signal_2096, signal_1344}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1145 ( .a ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({signal_1825, signal_1217}), .clk (clk), .r (Fresh[134]), .c ({signal_2097, signal_1345}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1146 ( .a ({ciphertext_s1[36], ciphertext_s0[36]}), .b ({signal_1826, signal_1218}), .clk (clk), .r (Fresh[135]), .c ({signal_2098, signal_1346}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1147 ( .a ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({signal_1827, signal_1219}), .clk (clk), .r (Fresh[136]), .c ({signal_2099, signal_1347}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1148 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({signal_1828, signal_1220}), .clk (clk), .r (Fresh[137]), .c ({signal_2100, signal_1348}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1149 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({signal_1829, signal_1221}), .clk (clk), .r (Fresh[138]), .c ({signal_2101, signal_1349}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1150 ( .a ({ciphertext_s1[20], ciphertext_s0[20]}), .b ({signal_1830, signal_1222}), .clk (clk), .r (Fresh[139]), .c ({signal_2102, signal_1350}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1151 ( .a ({ciphertext_s1[4], ciphertext_s0[4]}), .b ({signal_1831, signal_1223}), .clk (clk), .r (Fresh[140]), .c ({signal_2103, signal_1351}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1152 ( .a ({ciphertext_s1[8], ciphertext_s0[8]}), .b ({signal_1832, signal_1224}), .clk (clk), .r (Fresh[141]), .c ({signal_2104, signal_1352}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1153 ( .a ({ciphertext_s1[12], ciphertext_s0[12]}), .b ({signal_1833, signal_1225}), .clk (clk), .r (Fresh[142]), .c ({signal_2105, signal_1353}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1154 ( .a ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({signal_1834, signal_1226}), .clk (clk), .r (Fresh[143]), .c ({signal_2106, signal_1354}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1155 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({signal_1836, signal_1228}), .clk (clk), .r (Fresh[144]), .c ({signal_2107, signal_1355}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1156 ( .a ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({signal_1839, signal_1231}), .clk (clk), .r (Fresh[145]), .c ({signal_2108, signal_1356}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1157 ( .a ({ciphertext_s1[52], ciphertext_s0[52]}), .b ({signal_1842, signal_1234}), .clk (clk), .r (Fresh[146]), .c ({signal_2109, signal_1357}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1158 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({signal_1845, signal_1237}), .clk (clk), .r (Fresh[147]), .c ({signal_2110, signal_1358}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1159 ( .a ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({signal_1848, signal_1240}), .clk (clk), .r (Fresh[148]), .c ({signal_2111, signal_1359}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1160 ( .a ({ciphertext_s1[44], ciphertext_s0[44]}), .b ({signal_1851, signal_1243}), .clk (clk), .r (Fresh[149]), .c ({signal_2112, signal_1360}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1161 ( .a ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({signal_1854, signal_1246}), .clk (clk), .r (Fresh[150]), .c ({signal_2113, signal_1361}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1162 ( .a ({ciphertext_s1[36], ciphertext_s0[36]}), .b ({signal_1857, signal_1249}), .clk (clk), .r (Fresh[151]), .c ({signal_2114, signal_1362}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1163 ( .a ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({signal_1860, signal_1252}), .clk (clk), .r (Fresh[152]), .c ({signal_2115, signal_1363}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1164 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({signal_1863, signal_1255}), .clk (clk), .r (Fresh[153]), .c ({signal_2116, signal_1364}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1165 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({signal_1866, signal_1258}), .clk (clk), .r (Fresh[154]), .c ({signal_2117, signal_1365}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1166 ( .a ({ciphertext_s1[20], ciphertext_s0[20]}), .b ({signal_1869, signal_1261}), .clk (clk), .r (Fresh[155]), .c ({signal_2118, signal_1366}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1167 ( .a ({ciphertext_s1[4], ciphertext_s0[4]}), .b ({signal_1872, signal_1264}), .clk (clk), .r (Fresh[156]), .c ({signal_2119, signal_1367}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1168 ( .a ({ciphertext_s1[8], ciphertext_s0[8]}), .b ({signal_1875, signal_1267}), .clk (clk), .r (Fresh[157]), .c ({signal_2120, signal_1368}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1169 ( .a ({ciphertext_s1[12], ciphertext_s0[12]}), .b ({signal_1878, signal_1270}), .clk (clk), .r (Fresh[158]), .c ({signal_2121, signal_1369}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1170 ( .a ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({signal_1881, signal_1273}), .clk (clk), .r (Fresh[159]), .c ({signal_2122, signal_1370}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1171 ( .a ({signal_2091, signal_1339}), .b ({signal_2131, signal_1371}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1172 ( .a ({signal_2092, signal_1340}), .b ({signal_2132, signal_1372}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1173 ( .a ({signal_2093, signal_1341}), .b ({signal_2133, signal_1373}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1174 ( .a ({signal_2094, signal_1342}), .b ({signal_2134, signal_1374}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1175 ( .a ({signal_2095, signal_1343}), .b ({signal_2135, signal_1375}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1176 ( .a ({signal_2096, signal_1344}), .b ({signal_2136, signal_1376}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1177 ( .a ({signal_2097, signal_1345}), .b ({signal_2137, signal_1377}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1178 ( .a ({signal_2098, signal_1346}), .b ({signal_2138, signal_1378}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1179 ( .a ({signal_2099, signal_1347}), .b ({signal_2139, signal_1379}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1180 ( .a ({signal_2100, signal_1348}), .b ({signal_2140, signal_1380}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1181 ( .a ({signal_2101, signal_1349}), .b ({signal_2141, signal_1381}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1182 ( .a ({signal_2102, signal_1350}), .b ({signal_2142, signal_1382}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1183 ( .a ({signal_2103, signal_1351}), .b ({signal_2143, signal_1383}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1184 ( .a ({signal_2104, signal_1352}), .b ({signal_2144, signal_1384}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1185 ( .a ({signal_2105, signal_1353}), .b ({signal_2145, signal_1385}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1186 ( .a ({signal_2106, signal_1354}), .b ({signal_2146, signal_1386}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1187 ( .a ({signal_2107, signal_1355}), .b ({signal_2147, signal_1387}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1188 ( .a ({signal_2108, signal_1356}), .b ({signal_2148, signal_1388}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1189 ( .a ({signal_2109, signal_1357}), .b ({signal_2149, signal_1389}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1190 ( .a ({signal_2110, signal_1358}), .b ({signal_2150, signal_1390}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1191 ( .a ({signal_2111, signal_1359}), .b ({signal_2151, signal_1391}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1192 ( .a ({signal_2112, signal_1360}), .b ({signal_2152, signal_1392}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1193 ( .a ({signal_2113, signal_1361}), .b ({signal_2153, signal_1393}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1194 ( .a ({signal_2114, signal_1362}), .b ({signal_2154, signal_1394}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1195 ( .a ({signal_2115, signal_1363}), .b ({signal_2155, signal_1395}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1196 ( .a ({signal_2116, signal_1364}), .b ({signal_2156, signal_1396}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1197 ( .a ({signal_2117, signal_1365}), .b ({signal_2157, signal_1397}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1198 ( .a ({signal_2118, signal_1366}), .b ({signal_2158, signal_1398}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1199 ( .a ({signal_2119, signal_1367}), .b ({signal_2159, signal_1399}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1200 ( .a ({signal_2120, signal_1368}), .b ({signal_2160, signal_1400}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1201 ( .a ({signal_2121, signal_1369}), .b ({signal_2161, signal_1401}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1202 ( .a ({signal_2122, signal_1370}), .b ({signal_2162, signal_1402}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1 ( .s (rst), .b ({signal_2307, signal_773}), .a ({plaintext_s1[1], plaintext_s0[1]}), .c ({signal_2340, signal_869}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3 ( .s (rst), .b ({signal_2211, signal_771}), .a ({plaintext_s1[3], plaintext_s0[3]}), .c ({signal_2260, signal_867}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_5 ( .s (rst), .b ({signal_2308, signal_769}), .a ({plaintext_s1[5], plaintext_s0[5]}), .c ({signal_2342, signal_865}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_7 ( .s (rst), .b ({signal_2212, signal_767}), .a ({plaintext_s1[7], plaintext_s0[7]}), .c ({signal_2262, signal_863}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_9 ( .s (rst), .b ({signal_2309, signal_765}), .a ({plaintext_s1[9], plaintext_s0[9]}), .c ({signal_2344, signal_861}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_11 ( .s (rst), .b ({signal_2213, signal_763}), .a ({plaintext_s1[11], plaintext_s0[11]}), .c ({signal_2264, signal_859}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_13 ( .s (rst), .b ({signal_2310, signal_761}), .a ({plaintext_s1[13], plaintext_s0[13]}), .c ({signal_2346, signal_857}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_15 ( .s (rst), .b ({signal_2214, signal_759}), .a ({plaintext_s1[15], plaintext_s0[15]}), .c ({signal_2266, signal_855}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_17 ( .s (rst), .b ({signal_2311, signal_757}), .a ({plaintext_s1[17], plaintext_s0[17]}), .c ({signal_2348, signal_853}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_19 ( .s (rst), .b ({signal_2215, signal_755}), .a ({plaintext_s1[19], plaintext_s0[19]}), .c ({signal_2268, signal_851}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_21 ( .s (rst), .b ({signal_2312, signal_753}), .a ({plaintext_s1[21], plaintext_s0[21]}), .c ({signal_2350, signal_849}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_23 ( .s (rst), .b ({signal_2216, signal_751}), .a ({plaintext_s1[23], plaintext_s0[23]}), .c ({signal_2270, signal_847}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_25 ( .s (rst), .b ({signal_2313, signal_749}), .a ({plaintext_s1[25], plaintext_s0[25]}), .c ({signal_2352, signal_845}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_27 ( .s (rst), .b ({signal_2217, signal_747}), .a ({plaintext_s1[27], plaintext_s0[27]}), .c ({signal_2272, signal_843}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_29 ( .s (rst), .b ({signal_2314, signal_745}), .a ({plaintext_s1[29], plaintext_s0[29]}), .c ({signal_2354, signal_841}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_31 ( .s (rst), .b ({signal_2218, signal_743}), .a ({plaintext_s1[31], plaintext_s0[31]}), .c ({signal_2274, signal_839}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_33 ( .s (rst), .b ({signal_2315, signal_741}), .a ({plaintext_s1[33], plaintext_s0[33]}), .c ({signal_2356, signal_805}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_35 ( .s (rst), .b ({signal_2219, signal_739}), .a ({plaintext_s1[35], plaintext_s0[35]}), .c ({signal_2276, signal_803}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_37 ( .s (rst), .b ({signal_2316, signal_737}), .a ({plaintext_s1[37], plaintext_s0[37]}), .c ({signal_2358, signal_801}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_39 ( .s (rst), .b ({signal_2220, signal_735}), .a ({plaintext_s1[39], plaintext_s0[39]}), .c ({signal_2278, signal_799}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_41 ( .s (rst), .b ({signal_2317, signal_733}), .a ({plaintext_s1[41], plaintext_s0[41]}), .c ({signal_2360, signal_797}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_43 ( .s (rst), .b ({signal_2221, signal_731}), .a ({plaintext_s1[43], plaintext_s0[43]}), .c ({signal_2280, signal_795}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_45 ( .s (rst), .b ({signal_2318, signal_729}), .a ({plaintext_s1[45], plaintext_s0[45]}), .c ({signal_2362, signal_793}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_47 ( .s (rst), .b ({signal_2222, signal_727}), .a ({plaintext_s1[47], plaintext_s0[47]}), .c ({signal_2282, signal_791}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_49 ( .s (rst), .b ({signal_2319, signal_725}), .a ({plaintext_s1[49], plaintext_s0[49]}), .c ({signal_2364, signal_789}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_51 ( .s (rst), .b ({signal_2223, signal_723}), .a ({plaintext_s1[51], plaintext_s0[51]}), .c ({signal_2284, signal_787}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_53 ( .s (rst), .b ({signal_2320, signal_721}), .a ({plaintext_s1[53], plaintext_s0[53]}), .c ({signal_2366, signal_785}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_55 ( .s (rst), .b ({signal_2224, signal_719}), .a ({plaintext_s1[55], plaintext_s0[55]}), .c ({signal_2286, signal_783}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_57 ( .s (rst), .b ({signal_2321, signal_717}), .a ({plaintext_s1[57], plaintext_s0[57]}), .c ({signal_2368, signal_781}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_59 ( .s (rst), .b ({signal_2225, signal_715}), .a ({plaintext_s1[59], plaintext_s0[59]}), .c ({signal_2288, signal_779}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_61 ( .s (rst), .b ({signal_2322, signal_713}), .a ({plaintext_s1[61], plaintext_s0[61]}), .c ({signal_2370, signal_777}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_63 ( .s (rst), .b ({signal_2226, signal_711}), .a ({plaintext_s1[63], plaintext_s0[63]}), .c ({signal_2290, signal_775}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_69 ( .a ({signal_2488, signal_271}), .b ({signal_2487, signal_272}), .c ({signal_2526, signal_821}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_70 ( .a ({signal_2348, signal_853}), .b ({signal_2340, signal_869}), .c ({signal_2487, signal_272}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_71 ( .a ({1'b0, 1'b0}), .b ({signal_2364, signal_789}), .c ({signal_2488, signal_271}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_72 ( .a ({signal_2489, signal_273}), .b ({signal_2340, signal_869}), .c ({signal_2527, signal_837}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_73 ( .a ({1'b0, 1'b0}), .b ({signal_2356, signal_805}), .c ({signal_2489, signal_273}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_79 ( .a ({signal_2372, signal_277}), .b ({signal_2371, signal_278}), .c ({signal_2490, signal_819}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_80 ( .a ({signal_2268, signal_851}), .b ({signal_2260, signal_867}), .c ({signal_2371, signal_278}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_81 ( .a ({1'b0, 1'b0}), .b ({signal_2284, signal_787}), .c ({signal_2372, signal_277}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_82 ( .a ({signal_2373, signal_279}), .b ({signal_2260, signal_867}), .c ({signal_2491, signal_835}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_83 ( .a ({1'b0, 1'b0}), .b ({signal_2276, signal_803}), .c ({signal_2373, signal_279}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_89 ( .a ({signal_2493, signal_283}), .b ({signal_2492, signal_284}), .c ({signal_2534, signal_817}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_90 ( .a ({signal_2350, signal_849}), .b ({signal_2342, signal_865}), .c ({signal_2492, signal_284}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_91 ( .a ({1'b0, 1'b0}), .b ({signal_2366, signal_785}), .c ({signal_2493, signal_283}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_92 ( .a ({signal_2494, signal_285}), .b ({signal_2342, signal_865}), .c ({signal_2535, signal_833}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_93 ( .a ({1'b0, 1'b0}), .b ({signal_2358, signal_801}), .c ({signal_2494, signal_285}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_99 ( .a ({signal_2375, signal_289}), .b ({signal_2374, signal_290}), .c ({signal_2495, signal_815}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_100 ( .a ({signal_2270, signal_847}), .b ({signal_2262, signal_863}), .c ({signal_2374, signal_290}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_101 ( .a ({1'b0, 1'b0}), .b ({signal_2286, signal_783}), .c ({signal_2375, signal_289}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_102 ( .a ({signal_2376, signal_291}), .b ({signal_2262, signal_863}), .c ({signal_2496, signal_831}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_103 ( .a ({1'b0, 1'b0}), .b ({signal_2278, signal_799}), .c ({signal_2376, signal_291}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_109 ( .a ({signal_2498, signal_295}), .b ({signal_2497, signal_296}), .c ({signal_2542, signal_813}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_110 ( .a ({signal_2352, signal_845}), .b ({signal_2344, signal_861}), .c ({signal_2497, signal_296}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_111 ( .a ({1'b0, 1'b0}), .b ({signal_2368, signal_781}), .c ({signal_2498, signal_295}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_112 ( .a ({signal_2499, signal_297}), .b ({signal_2344, signal_861}), .c ({signal_2543, signal_829}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_113 ( .a ({1'b0, 1'b0}), .b ({signal_2360, signal_797}), .c ({signal_2499, signal_297}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_119 ( .a ({signal_2378, signal_301}), .b ({signal_2377, signal_302}), .c ({signal_2500, signal_811}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_120 ( .a ({signal_2272, signal_843}), .b ({signal_2264, signal_859}), .c ({signal_2377, signal_302}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_121 ( .a ({1'b0, 1'b0}), .b ({signal_2288, signal_779}), .c ({signal_2378, signal_301}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_122 ( .a ({signal_2379, signal_303}), .b ({signal_2264, signal_859}), .c ({signal_2501, signal_827}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_123 ( .a ({1'b0, 1'b0}), .b ({signal_2280, signal_795}), .c ({signal_2379, signal_303}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_129 ( .a ({signal_2503, signal_307}), .b ({signal_2502, signal_308}), .c ({signal_2550, signal_809}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_130 ( .a ({signal_2354, signal_841}), .b ({signal_2346, signal_857}), .c ({signal_2502, signal_308}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_131 ( .a ({1'b0, 1'b0}), .b ({signal_2370, signal_777}), .c ({signal_2503, signal_307}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_132 ( .a ({signal_2504, signal_309}), .b ({signal_2346, signal_857}), .c ({signal_2551, signal_825}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_133 ( .a ({1'b0, 1'b0}), .b ({signal_2362, signal_793}), .c ({signal_2504, signal_309}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_139 ( .a ({signal_2381, signal_313}), .b ({signal_2380, signal_314}), .c ({signal_2505, signal_807}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_140 ( .a ({signal_2274, signal_839}), .b ({signal_2266, signal_855}), .c ({signal_2380, signal_314}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_141 ( .a ({1'b0, 1'b0}), .b ({signal_2290, signal_775}), .c ({signal_2381, signal_313}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_142 ( .a ({signal_2382, signal_315}), .b ({signal_2266, signal_855}), .c ({signal_2506, signal_823}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_143 ( .a ({1'b0, 1'b0}), .b ({signal_2282, signal_791}), .c ({signal_2382, signal_315}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_146 ( .a ({signal_2603, signal_317}), .b ({signal_2031, signal_885}), .c ({signal_2636, signal_949}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_147 ( .a ({1'b0, 1'b0}), .b ({signal_2526, signal_821}), .c ({signal_2603, signal_317}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_150 ( .a ({signal_2555, signal_319}), .b ({signal_2037, signal_883}), .c ({signal_2604, signal_947}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_151 ( .a ({1'b0, 1'b0}), .b ({signal_2490, signal_819}), .c ({signal_2555, signal_319}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_154 ( .a ({signal_2605, signal_321}), .b ({signal_1710, signal_881}), .c ({signal_2639, signal_945}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_155 ( .a ({1'b0, 1'b0}), .b ({signal_2534, signal_817}), .c ({signal_2605, signal_321}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_158 ( .a ({signal_2556, signal_323}), .b ({signal_2043, signal_879}), .c ({signal_2606, signal_943}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_159 ( .a ({1'b0, 1'b0}), .b ({signal_2495, signal_815}), .c ({signal_2556, signal_323}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_162 ( .a ({signal_2607, signal_325}), .b ({signal_2046, signal_877}), .c ({signal_2642, signal_941}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_163 ( .a ({1'b0, 1'b0}), .b ({signal_2542, signal_813}), .c ({signal_2607, signal_325}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_166 ( .a ({signal_2557, signal_327}), .b ({signal_1719, signal_875}), .c ({signal_2608, signal_939}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_167 ( .a ({1'b0, 1'b0}), .b ({signal_2500, signal_811}), .c ({signal_2557, signal_327}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_170 ( .a ({signal_2609, signal_329}), .b ({signal_2055, signal_873}), .c ({signal_2645, signal_937}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_171 ( .a ({1'b0, 1'b0}), .b ({signal_2550, signal_809}), .c ({signal_2609, signal_329}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_174 ( .a ({signal_2558, signal_331}), .b ({signal_2058, signal_871}), .c ({signal_2610, signal_935}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_175 ( .a ({1'b0, 1'b0}), .b ({signal_2505, signal_807}), .c ({signal_2558, signal_331}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_179 ( .a ({signal_2611, signal_334}), .b ({signal_2124, signal_335}), .c ({signal_2648, signal_957}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_181 ( .a ({1'b0, 1'b0}), .b ({signal_2543, signal_829}), .c ({signal_2611, signal_334}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_185 ( .a ({signal_2559, signal_338}), .b ({signal_2126, signal_339}), .c ({signal_2612, signal_955}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_187 ( .a ({1'b0, 1'b0}), .b ({signal_2501, signal_827}), .c ({signal_2559, signal_338}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_191 ( .a ({signal_2613, signal_342}), .b ({signal_2128, signal_343}), .c ({signal_2651, signal_953}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_193 ( .a ({1'b0, 1'b0}), .b ({signal_2551, signal_825}), .c ({signal_2613, signal_342}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_197 ( .a ({signal_2560, signal_346}), .b ({signal_2130, signal_347}), .c ({signal_2614, signal_951}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_199 ( .a ({1'b0, 1'b0}), .b ({signal_2506, signal_823}), .c ({signal_2560, signal_346}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_202 ( .a ({signal_2507, signal_349}), .b ({signal_1917, signal_933}), .c ({signal_2562, signal_997}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_203 ( .a ({1'b0, 1'b0}), .b ({signal_2340, signal_869}), .c ({signal_2507, signal_349}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_206 ( .a ({signal_2383, signal_351}), .b ({signal_1920, signal_931}), .c ({signal_2508, signal_995}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_207 ( .a ({1'b0, 1'b0}), .b ({signal_2260, signal_867}), .c ({signal_2383, signal_351}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_210 ( .a ({signal_2509, signal_353}), .b ({signal_1926, signal_929}), .c ({signal_2565, signal_993}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_211 ( .a ({1'b0, 1'b0}), .b ({signal_2342, signal_865}), .c ({signal_2509, signal_353}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_214 ( .a ({signal_2384, signal_355}), .b ({signal_1932, signal_927}), .c ({signal_2510, signal_991}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_215 ( .a ({1'b0, 1'b0}), .b ({signal_2262, signal_863}), .c ({signal_2384, signal_355}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_218 ( .a ({signal_2511, signal_357}), .b ({signal_1938, signal_925}), .c ({signal_2568, signal_989}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_219 ( .a ({1'b0, 1'b0}), .b ({signal_2344, signal_861}), .c ({signal_2511, signal_357}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_222 ( .a ({signal_2385, signal_359}), .b ({signal_1944, signal_923}), .c ({signal_2512, signal_987}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_223 ( .a ({1'b0, 1'b0}), .b ({signal_2264, signal_859}), .c ({signal_2385, signal_359}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_226 ( .a ({signal_2513, signal_361}), .b ({signal_1950, signal_921}), .c ({signal_2571, signal_985}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_227 ( .a ({1'b0, 1'b0}), .b ({signal_2346, signal_857}), .c ({signal_2513, signal_361}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_230 ( .a ({signal_2386, signal_363}), .b ({signal_1956, signal_919}), .c ({signal_2514, signal_983}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_231 ( .a ({1'b0, 1'b0}), .b ({signal_2266, signal_855}), .c ({signal_2386, signal_363}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_234 ( .a ({signal_2515, signal_365}), .b ({signal_1962, signal_917}), .c ({signal_2574, signal_981}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_235 ( .a ({1'b0, 1'b0}), .b ({signal_2348, signal_853}), .c ({signal_2515, signal_365}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_238 ( .a ({signal_2387, signal_367}), .b ({signal_1968, signal_915}), .c ({signal_2516, signal_979}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_239 ( .a ({1'b0, 1'b0}), .b ({signal_2268, signal_851}), .c ({signal_2387, signal_367}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_242 ( .a ({signal_2517, signal_369}), .b ({signal_1974, signal_913}), .c ({signal_2577, signal_977}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_243 ( .a ({1'b0, 1'b0}), .b ({signal_2350, signal_849}), .c ({signal_2517, signal_369}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_246 ( .a ({signal_2388, signal_371}), .b ({signal_1686, signal_911}), .c ({signal_2518, signal_975}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_247 ( .a ({1'b0, 1'b0}), .b ({signal_2270, signal_847}), .c ({signal_2388, signal_371}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_250 ( .a ({signal_2519, signal_373}), .b ({signal_1692, signal_909}), .c ({signal_2580, signal_973}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_251 ( .a ({1'b0, 1'b0}), .b ({signal_2352, signal_845}), .c ({signal_2519, signal_373}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_254 ( .a ({signal_2389, signal_375}), .b ({signal_1698, signal_907}), .c ({signal_2520, signal_971}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_255 ( .a ({1'b0, 1'b0}), .b ({signal_2272, signal_843}), .c ({signal_2389, signal_375}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_258 ( .a ({signal_2521, signal_377}), .b ({signal_1980, signal_905}), .c ({signal_2583, signal_969}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_259 ( .a ({1'b0, 1'b0}), .b ({signal_2354, signal_841}), .c ({signal_2521, signal_377}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_262 ( .a ({signal_2390, signal_379}), .b ({signal_1986, signal_903}), .c ({signal_2522, signal_967}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_263 ( .a ({1'b0, 1'b0}), .b ({signal_2274, signal_839}), .c ({signal_2390, signal_379}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_266 ( .a ({signal_2631, signal_381}), .b ({signal_1701, signal_901}), .c ({signal_2654, signal_965}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_267 ( .a ({1'b0, 1'b0}), .b ({signal_2527, signal_837}), .c ({signal_2631, signal_381}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_270 ( .a ({signal_2585, signal_383}), .b ({signal_1995, signal_899}), .c ({signal_2632, signal_963}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_271 ( .a ({1'b0, 1'b0}), .b ({signal_2491, signal_835}), .c ({signal_2585, signal_383}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_274 ( .a ({signal_2633, signal_385}), .b ({signal_1998, signal_897}), .c ({signal_2657, signal_961}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_275 ( .a ({1'b0, 1'b0}), .b ({signal_2535, signal_833}), .c ({signal_2633, signal_385}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_278 ( .a ({signal_2586, signal_387}), .b ({signal_1707, signal_895}), .c ({signal_2634, signal_959}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_279 ( .a ({1'b0, 1'b0}), .b ({signal_2496, signal_831}), .c ({signal_2586, signal_387}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1203 ( .a ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({signal_2059, signal_1307}), .clk (clk), .r (Fresh[160]), .c ({signal_2163, signal_1403}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1204 ( .a ({ciphertext_s1[49], ciphertext_s0[49]}), .b ({signal_2060, signal_1308}), .clk (clk), .r (Fresh[161]), .c ({signal_2164, signal_1404}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1205 ( .a ({ciphertext_s1[53], ciphertext_s0[53]}), .b ({signal_2061, signal_1309}), .clk (clk), .r (Fresh[162]), .c ({signal_2165, signal_1405}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1206 ( .a ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({signal_2062, signal_1310}), .clk (clk), .r (Fresh[163]), .c ({signal_2166, signal_1406}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1207 ( .a ({ciphertext_s1[33], ciphertext_s0[33]}), .b ({signal_2063, signal_1311}), .clk (clk), .r (Fresh[164]), .c ({signal_2167, signal_1407}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1208 ( .a ({ciphertext_s1[45], ciphertext_s0[45]}), .b ({signal_2064, signal_1312}), .clk (clk), .r (Fresh[165]), .c ({signal_2168, signal_1408}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1209 ( .a ({ciphertext_s1[41], ciphertext_s0[41]}), .b ({signal_2065, signal_1313}), .clk (clk), .r (Fresh[166]), .c ({signal_2169, signal_1409}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1210 ( .a ({ciphertext_s1[37], ciphertext_s0[37]}), .b ({signal_2066, signal_1314}), .clk (clk), .r (Fresh[167]), .c ({signal_2170, signal_1410}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1211 ( .a ({ciphertext_s1[17], ciphertext_s0[17]}), .b ({signal_2067, signal_1315}), .clk (clk), .r (Fresh[168]), .c ({signal_2171, signal_1411}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1212 ( .a ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({signal_2068, signal_1316}), .clk (clk), .r (Fresh[169]), .c ({signal_2172, signal_1412}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1213 ( .a ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({signal_2069, signal_1317}), .clk (clk), .r (Fresh[170]), .c ({signal_2173, signal_1413}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1214 ( .a ({ciphertext_s1[21], ciphertext_s0[21]}), .b ({signal_2070, signal_1318}), .clk (clk), .r (Fresh[171]), .c ({signal_2174, signal_1414}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1215 ( .a ({ciphertext_s1[5], ciphertext_s0[5]}), .b ({signal_2071, signal_1319}), .clk (clk), .r (Fresh[172]), .c ({signal_2175, signal_1415}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1216 ( .a ({ciphertext_s1[9], ciphertext_s0[9]}), .b ({signal_2072, signal_1320}), .clk (clk), .r (Fresh[173]), .c ({signal_2176, signal_1416}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1217 ( .a ({ciphertext_s1[13], ciphertext_s0[13]}), .b ({signal_2073, signal_1321}), .clk (clk), .r (Fresh[174]), .c ({signal_2177, signal_1417}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1218 ( .a ({ciphertext_s1[1], ciphertext_s0[1]}), .b ({signal_2074, signal_1322}), .clk (clk), .r (Fresh[175]), .c ({signal_2178, signal_1418}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1219 ( .a ({signal_1835, signal_1227}), .b ({signal_2075, signal_1323}), .clk (clk), .r (Fresh[176]), .c ({signal_2179, signal_1419}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1220 ( .a ({signal_1838, signal_1230}), .b ({signal_2076, signal_1324}), .clk (clk), .r (Fresh[177]), .c ({signal_2180, signal_1420}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1221 ( .a ({signal_1841, signal_1233}), .b ({signal_2077, signal_1325}), .clk (clk), .r (Fresh[178]), .c ({signal_2181, signal_1421}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1222 ( .a ({signal_1844, signal_1236}), .b ({signal_2078, signal_1326}), .clk (clk), .r (Fresh[179]), .c ({signal_2182, signal_1422}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1223 ( .a ({signal_1847, signal_1239}), .b ({signal_2079, signal_1327}), .clk (clk), .r (Fresh[180]), .c ({signal_2183, signal_1423}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1224 ( .a ({signal_1850, signal_1242}), .b ({signal_2080, signal_1328}), .clk (clk), .r (Fresh[181]), .c ({signal_2184, signal_1424}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1225 ( .a ({signal_1853, signal_1245}), .b ({signal_2081, signal_1329}), .clk (clk), .r (Fresh[182]), .c ({signal_2185, signal_1425}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1226 ( .a ({signal_1856, signal_1248}), .b ({signal_2082, signal_1330}), .clk (clk), .r (Fresh[183]), .c ({signal_2186, signal_1426}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1227 ( .a ({signal_1859, signal_1251}), .b ({signal_2083, signal_1331}), .clk (clk), .r (Fresh[184]), .c ({signal_2187, signal_1427}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1228 ( .a ({signal_1862, signal_1254}), .b ({signal_2084, signal_1332}), .clk (clk), .r (Fresh[185]), .c ({signal_2188, signal_1428}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1229 ( .a ({signal_1865, signal_1257}), .b ({signal_2085, signal_1333}), .clk (clk), .r (Fresh[186]), .c ({signal_2189, signal_1429}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1230 ( .a ({signal_1868, signal_1260}), .b ({signal_2086, signal_1334}), .clk (clk), .r (Fresh[187]), .c ({signal_2190, signal_1430}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1231 ( .a ({signal_1871, signal_1263}), .b ({signal_2087, signal_1335}), .clk (clk), .r (Fresh[188]), .c ({signal_2191, signal_1431}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1232 ( .a ({signal_1874, signal_1266}), .b ({signal_2088, signal_1336}), .clk (clk), .r (Fresh[189]), .c ({signal_2192, signal_1432}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1233 ( .a ({signal_1877, signal_1269}), .b ({signal_2089, signal_1337}), .clk (clk), .r (Fresh[190]), .c ({signal_2193, signal_1433}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1234 ( .a ({signal_1880, signal_1272}), .b ({signal_2090, signal_1338}), .clk (clk), .r (Fresh[191]), .c ({signal_2194, signal_1434}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1235 ( .a ({signal_2163, signal_1403}), .b ({signal_2195, signal_1435}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1236 ( .a ({signal_2164, signal_1404}), .b ({signal_2196, signal_1436}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1237 ( .a ({signal_2165, signal_1405}), .b ({signal_2197, signal_1437}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1238 ( .a ({signal_2166, signal_1406}), .b ({signal_2198, signal_1438}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1239 ( .a ({signal_2167, signal_1407}), .b ({signal_2199, signal_1439}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1240 ( .a ({signal_2168, signal_1408}), .b ({signal_2200, signal_1440}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1241 ( .a ({signal_2169, signal_1409}), .b ({signal_2201, signal_1441}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1242 ( .a ({signal_2170, signal_1410}), .b ({signal_2202, signal_1442}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1243 ( .a ({signal_2171, signal_1411}), .b ({signal_2203, signal_1443}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1244 ( .a ({signal_2172, signal_1412}), .b ({signal_2204, signal_1444}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1245 ( .a ({signal_2173, signal_1413}), .b ({signal_2205, signal_1445}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1246 ( .a ({signal_2174, signal_1414}), .b ({signal_2206, signal_1446}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1247 ( .a ({signal_2175, signal_1415}), .b ({signal_2207, signal_1447}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1248 ( .a ({signal_2176, signal_1416}), .b ({signal_2208, signal_1448}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1249 ( .a ({signal_2177, signal_1417}), .b ({signal_2209, signal_1449}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1250 ( .a ({signal_2178, signal_1418}), .b ({signal_2210, signal_1450}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1251 ( .a ({signal_2179, signal_1419}), .b ({signal_2211, signal_771}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1252 ( .a ({signal_2180, signal_1420}), .b ({signal_2212, signal_767}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1253 ( .a ({signal_2181, signal_1421}), .b ({signal_2213, signal_763}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1254 ( .a ({signal_2182, signal_1422}), .b ({signal_2214, signal_759}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1255 ( .a ({signal_2183, signal_1423}), .b ({signal_2215, signal_755}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1256 ( .a ({signal_2184, signal_1424}), .b ({signal_2216, signal_751}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1257 ( .a ({signal_2185, signal_1425}), .b ({signal_2217, signal_747}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1258 ( .a ({signal_2186, signal_1426}), .b ({signal_2218, signal_743}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1259 ( .a ({signal_2187, signal_1427}), .b ({signal_2219, signal_739}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1260 ( .a ({signal_2188, signal_1428}), .b ({signal_2220, signal_735}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1261 ( .a ({signal_2189, signal_1429}), .b ({signal_2221, signal_731}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1262 ( .a ({signal_2190, signal_1430}), .b ({signal_2222, signal_727}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1263 ( .a ({signal_2191, signal_1431}), .b ({signal_2223, signal_723}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1264 ( .a ({signal_2192, signal_1432}), .b ({signal_2224, signal_719}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1265 ( .a ({signal_2193, signal_1433}), .b ({signal_2225, signal_715}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1266 ( .a ({signal_2194, signal_1434}), .b ({signal_2226, signal_711}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1267 ( .a ({signal_1638, signal_1080}), .b ({signal_2131, signal_1371}), .clk (clk), .r (Fresh[192]), .c ({signal_2227, signal_1451}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1268 ( .a ({signal_1614, signal_1068}), .b ({signal_2132, signal_1372}), .clk (clk), .r (Fresh[193]), .c ({signal_2228, signal_1452}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1269 ( .a ({signal_1622, signal_1072}), .b ({signal_2133, signal_1373}), .clk (clk), .r (Fresh[194]), .c ({signal_2229, signal_1453}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1270 ( .a ({signal_1630, signal_1076}), .b ({signal_2134, signal_1374}), .clk (clk), .r (Fresh[195]), .c ({signal_2230, signal_1454}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1271 ( .a ({signal_1582, signal_1052}), .b ({signal_2135, signal_1375}), .clk (clk), .r (Fresh[196]), .c ({signal_2231, signal_1455}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1272 ( .a ({signal_1606, signal_1064}), .b ({signal_2136, signal_1376}), .clk (clk), .r (Fresh[197]), .c ({signal_2232, signal_1456}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1273 ( .a ({signal_1598, signal_1060}), .b ({signal_2137, signal_1377}), .clk (clk), .r (Fresh[198]), .c ({signal_2233, signal_1457}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1274 ( .a ({signal_1590, signal_1056}), .b ({signal_2138, signal_1378}), .clk (clk), .r (Fresh[199]), .c ({signal_2234, signal_1458}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1275 ( .a ({signal_1550, signal_1036}), .b ({signal_2139, signal_1379}), .clk (clk), .r (Fresh[200]), .c ({signal_2235, signal_1459}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1276 ( .a ({signal_1574, signal_1048}), .b ({signal_2140, signal_1380}), .clk (clk), .r (Fresh[201]), .c ({signal_2236, signal_1460}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1277 ( .a ({signal_1566, signal_1044}), .b ({signal_2141, signal_1381}), .clk (clk), .r (Fresh[202]), .c ({signal_2237, signal_1461}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1278 ( .a ({signal_1558, signal_1040}), .b ({signal_2142, signal_1382}), .clk (clk), .r (Fresh[203]), .c ({signal_2238, signal_1462}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1279 ( .a ({signal_1526, signal_1024}), .b ({signal_2143, signal_1383}), .clk (clk), .r (Fresh[204]), .c ({signal_2239, signal_1463}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1280 ( .a ({signal_1534, signal_1028}), .b ({signal_2144, signal_1384}), .clk (clk), .r (Fresh[205]), .c ({signal_2240, signal_1464}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1281 ( .a ({signal_1542, signal_1032}), .b ({signal_2145, signal_1385}), .clk (clk), .r (Fresh[206]), .c ({signal_2241, signal_1465}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1282 ( .a ({signal_1518, signal_1020}), .b ({signal_2146, signal_1386}), .clk (clk), .r (Fresh[207]), .c ({signal_2242, signal_1466}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1283 ( .a ({signal_1837, signal_1229}), .b ({signal_2147, signal_1387}), .clk (clk), .r (Fresh[208]), .c ({signal_2243, signal_1467}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1284 ( .a ({signal_1840, signal_1232}), .b ({signal_2148, signal_1388}), .clk (clk), .r (Fresh[209]), .c ({signal_2244, signal_1468}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1285 ( .a ({signal_1843, signal_1235}), .b ({signal_2149, signal_1389}), .clk (clk), .r (Fresh[210]), .c ({signal_2245, signal_1469}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1286 ( .a ({signal_1846, signal_1238}), .b ({signal_2150, signal_1390}), .clk (clk), .r (Fresh[211]), .c ({signal_2246, signal_1470}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1287 ( .a ({signal_1849, signal_1241}), .b ({signal_2151, signal_1391}), .clk (clk), .r (Fresh[212]), .c ({signal_2247, signal_1471}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1288 ( .a ({signal_1852, signal_1244}), .b ({signal_2152, signal_1392}), .clk (clk), .r (Fresh[213]), .c ({signal_2248, signal_1472}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1289 ( .a ({signal_1855, signal_1247}), .b ({signal_2153, signal_1393}), .clk (clk), .r (Fresh[214]), .c ({signal_2249, signal_1473}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1290 ( .a ({signal_1858, signal_1250}), .b ({signal_2154, signal_1394}), .clk (clk), .r (Fresh[215]), .c ({signal_2250, signal_1474}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1291 ( .a ({signal_1861, signal_1253}), .b ({signal_2155, signal_1395}), .clk (clk), .r (Fresh[216]), .c ({signal_2251, signal_1475}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1292 ( .a ({signal_1864, signal_1256}), .b ({signal_2156, signal_1396}), .clk (clk), .r (Fresh[217]), .c ({signal_2252, signal_1476}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1293 ( .a ({signal_1867, signal_1259}), .b ({signal_2157, signal_1397}), .clk (clk), .r (Fresh[218]), .c ({signal_2253, signal_1477}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1294 ( .a ({signal_1870, signal_1262}), .b ({signal_2158, signal_1398}), .clk (clk), .r (Fresh[219]), .c ({signal_2254, signal_1478}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1295 ( .a ({signal_1873, signal_1265}), .b ({signal_2159, signal_1399}), .clk (clk), .r (Fresh[220]), .c ({signal_2255, signal_1479}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1296 ( .a ({signal_1876, signal_1268}), .b ({signal_2160, signal_1400}), .clk (clk), .r (Fresh[221]), .c ({signal_2256, signal_1480}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1297 ( .a ({signal_1879, signal_1271}), .b ({signal_2161, signal_1401}), .clk (clk), .r (Fresh[222]), .c ({signal_2257, signal_1481}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1298 ( .a ({signal_1882, signal_1274}), .b ({signal_2162, signal_1402}), .clk (clk), .r (Fresh[223]), .c ({signal_2258, signal_1482}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1299 ( .a ({signal_2227, signal_1451}), .b ({signal_2291, signal_1483}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1300 ( .a ({signal_2228, signal_1452}), .b ({signal_2292, signal_1484}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1301 ( .a ({signal_2229, signal_1453}), .b ({signal_2293, signal_1485}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1302 ( .a ({signal_2230, signal_1454}), .b ({signal_2294, signal_1486}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1303 ( .a ({signal_2231, signal_1455}), .b ({signal_2295, signal_1487}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1304 ( .a ({signal_2232, signal_1456}), .b ({signal_2296, signal_1488}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1305 ( .a ({signal_2233, signal_1457}), .b ({signal_2297, signal_1489}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1306 ( .a ({signal_2234, signal_1458}), .b ({signal_2298, signal_1490}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1307 ( .a ({signal_2235, signal_1459}), .b ({signal_2299, signal_1491}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1308 ( .a ({signal_2236, signal_1460}), .b ({signal_2300, signal_1492}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1309 ( .a ({signal_2237, signal_1461}), .b ({signal_2301, signal_1493}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1310 ( .a ({signal_2238, signal_1462}), .b ({signal_2302, signal_1494}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1311 ( .a ({signal_2239, signal_1463}), .b ({signal_2303, signal_1495}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1312 ( .a ({signal_2240, signal_1464}), .b ({signal_2304, signal_1496}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1313 ( .a ({signal_2241, signal_1465}), .b ({signal_2305, signal_1497}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1314 ( .a ({signal_2242, signal_1466}), .b ({signal_2306, signal_1498}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1315 ( .a ({signal_2243, signal_1467}), .b ({signal_2307, signal_773}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1316 ( .a ({signal_2244, signal_1468}), .b ({signal_2308, signal_769}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1317 ( .a ({signal_2245, signal_1469}), .b ({signal_2309, signal_765}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1318 ( .a ({signal_2246, signal_1470}), .b ({signal_2310, signal_761}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1319 ( .a ({signal_2247, signal_1471}), .b ({signal_2311, signal_757}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1320 ( .a ({signal_2248, signal_1472}), .b ({signal_2312, signal_753}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1321 ( .a ({signal_2249, signal_1473}), .b ({signal_2313, signal_749}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1322 ( .a ({signal_2250, signal_1474}), .b ({signal_2314, signal_745}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1323 ( .a ({signal_2251, signal_1475}), .b ({signal_2315, signal_741}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1324 ( .a ({signal_2252, signal_1476}), .b ({signal_2316, signal_737}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1325 ( .a ({signal_2253, signal_1477}), .b ({signal_2317, signal_733}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1326 ( .a ({signal_2254, signal_1478}), .b ({signal_2318, signal_729}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1327 ( .a ({signal_2255, signal_1479}), .b ({signal_2319, signal_725}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1328 ( .a ({signal_2256, signal_1480}), .b ({signal_2320, signal_721}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1329 ( .a ({signal_2257, signal_1481}), .b ({signal_2321, signal_717}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1330 ( .a ({signal_2258, signal_1482}), .b ({signal_2322, signal_713}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    mux2_masked #(.security_order(1), .pipeline(0)) cell_0 ( .s (rst), .b ({signal_2407, signal_774}), .a ({plaintext_s1[0], plaintext_s0[0]}), .c ({signal_2424, signal_870}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_2 ( .s (rst), .b ({signal_2391, signal_772}), .a ({plaintext_s1[2], plaintext_s0[2]}), .c ({signal_2426, signal_868}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_4 ( .s (rst), .b ({signal_2408, signal_770}), .a ({plaintext_s1[4], plaintext_s0[4]}), .c ({signal_2428, signal_866}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_6 ( .s (rst), .b ({signal_2392, signal_768}), .a ({plaintext_s1[6], plaintext_s0[6]}), .c ({signal_2430, signal_864}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_8 ( .s (rst), .b ({signal_2409, signal_766}), .a ({plaintext_s1[8], plaintext_s0[8]}), .c ({signal_2432, signal_862}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_10 ( .s (rst), .b ({signal_2393, signal_764}), .a ({plaintext_s1[10], plaintext_s0[10]}), .c ({signal_2434, signal_860}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_12 ( .s (rst), .b ({signal_2410, signal_762}), .a ({plaintext_s1[12], plaintext_s0[12]}), .c ({signal_2436, signal_858}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_14 ( .s (rst), .b ({signal_2394, signal_760}), .a ({plaintext_s1[14], plaintext_s0[14]}), .c ({signal_2438, signal_856}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_16 ( .s (rst), .b ({signal_2411, signal_758}), .a ({plaintext_s1[16], plaintext_s0[16]}), .c ({signal_2440, signal_854}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_18 ( .s (rst), .b ({signal_2395, signal_756}), .a ({plaintext_s1[18], plaintext_s0[18]}), .c ({signal_2442, signal_852}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_20 ( .s (rst), .b ({signal_2412, signal_754}), .a ({plaintext_s1[20], plaintext_s0[20]}), .c ({signal_2444, signal_850}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_22 ( .s (rst), .b ({signal_2396, signal_752}), .a ({plaintext_s1[22], plaintext_s0[22]}), .c ({signal_2446, signal_848}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_24 ( .s (rst), .b ({signal_2413, signal_750}), .a ({plaintext_s1[24], plaintext_s0[24]}), .c ({signal_2448, signal_846}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_26 ( .s (rst), .b ({signal_2397, signal_748}), .a ({plaintext_s1[26], plaintext_s0[26]}), .c ({signal_2450, signal_844}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_28 ( .s (rst), .b ({signal_2414, signal_746}), .a ({plaintext_s1[28], plaintext_s0[28]}), .c ({signal_2452, signal_842}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_30 ( .s (rst), .b ({signal_2398, signal_744}), .a ({plaintext_s1[30], plaintext_s0[30]}), .c ({signal_2454, signal_840}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_32 ( .s (rst), .b ({signal_2415, signal_742}), .a ({plaintext_s1[32], plaintext_s0[32]}), .c ({signal_2456, signal_806}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_34 ( .s (rst), .b ({signal_2399, signal_740}), .a ({plaintext_s1[34], plaintext_s0[34]}), .c ({signal_2458, signal_804}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_36 ( .s (rst), .b ({signal_2416, signal_738}), .a ({plaintext_s1[36], plaintext_s0[36]}), .c ({signal_2460, signal_802}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_38 ( .s (rst), .b ({signal_2400, signal_736}), .a ({plaintext_s1[38], plaintext_s0[38]}), .c ({signal_2462, signal_800}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_40 ( .s (rst), .b ({signal_2417, signal_734}), .a ({plaintext_s1[40], plaintext_s0[40]}), .c ({signal_2464, signal_798}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_42 ( .s (rst), .b ({signal_2401, signal_732}), .a ({plaintext_s1[42], plaintext_s0[42]}), .c ({signal_2466, signal_796}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_44 ( .s (rst), .b ({signal_2418, signal_730}), .a ({plaintext_s1[44], plaintext_s0[44]}), .c ({signal_2468, signal_794}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_46 ( .s (rst), .b ({signal_2402, signal_728}), .a ({plaintext_s1[46], plaintext_s0[46]}), .c ({signal_2470, signal_792}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_48 ( .s (rst), .b ({signal_2419, signal_726}), .a ({plaintext_s1[48], plaintext_s0[48]}), .c ({signal_2472, signal_790}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_50 ( .s (rst), .b ({signal_2403, signal_724}), .a ({plaintext_s1[50], plaintext_s0[50]}), .c ({signal_2474, signal_788}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_52 ( .s (rst), .b ({signal_2420, signal_722}), .a ({plaintext_s1[52], plaintext_s0[52]}), .c ({signal_2476, signal_786}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_54 ( .s (rst), .b ({signal_2404, signal_720}), .a ({plaintext_s1[54], plaintext_s0[54]}), .c ({signal_2478, signal_784}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_56 ( .s (rst), .b ({signal_2421, signal_718}), .a ({plaintext_s1[56], plaintext_s0[56]}), .c ({signal_2480, signal_782}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_58 ( .s (rst), .b ({signal_2405, signal_716}), .a ({plaintext_s1[58], plaintext_s0[58]}), .c ({signal_2482, signal_780}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_60 ( .s (rst), .b ({signal_2422, signal_714}), .a ({plaintext_s1[60], plaintext_s0[60]}), .c ({signal_2484, signal_778}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_62 ( .s (rst), .b ({signal_2406, signal_712}), .a ({plaintext_s1[62], plaintext_s0[62]}), .c ({signal_2486, signal_776}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_64 ( .a ({signal_2524, signal_268}), .b ({signal_2523, signal_269}), .c ({signal_2587, signal_822}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_65 ( .a ({signal_2440, signal_854}), .b ({signal_2424, signal_870}), .c ({signal_2523, signal_269}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_66 ( .a ({1'b0, 1'b0}), .b ({signal_2472, signal_790}), .c ({signal_2524, signal_268}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_67 ( .a ({signal_2525, signal_270}), .b ({signal_2424, signal_870}), .c ({signal_2588, signal_838}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_68 ( .a ({1'b0, 1'b0}), .b ({signal_2456, signal_806}), .c ({signal_2525, signal_270}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_74 ( .a ({signal_2529, signal_274}), .b ({signal_2528, signal_275}), .c ({signal_2589, signal_820}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_75 ( .a ({signal_2442, signal_852}), .b ({signal_2426, signal_868}), .c ({signal_2528, signal_275}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_76 ( .a ({1'b0, 1'b0}), .b ({signal_2474, signal_788}), .c ({signal_2529, signal_274}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_77 ( .a ({signal_2530, signal_276}), .b ({signal_2426, signal_868}), .c ({signal_2590, signal_836}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_78 ( .a ({1'b0, 1'b0}), .b ({signal_2458, signal_804}), .c ({signal_2530, signal_276}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_84 ( .a ({signal_2532, signal_280}), .b ({signal_2531, signal_281}), .c ({signal_2591, signal_818}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_85 ( .a ({signal_2444, signal_850}), .b ({signal_2428, signal_866}), .c ({signal_2531, signal_281}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_86 ( .a ({1'b0, 1'b0}), .b ({signal_2476, signal_786}), .c ({signal_2532, signal_280}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_87 ( .a ({signal_2533, signal_282}), .b ({signal_2428, signal_866}), .c ({signal_2592, signal_834}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_88 ( .a ({1'b0, 1'b0}), .b ({signal_2460, signal_802}), .c ({signal_2533, signal_282}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_94 ( .a ({signal_2537, signal_286}), .b ({signal_2536, signal_287}), .c ({signal_2593, signal_816}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_95 ( .a ({signal_2446, signal_848}), .b ({signal_2430, signal_864}), .c ({signal_2536, signal_287}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_96 ( .a ({1'b0, 1'b0}), .b ({signal_2478, signal_784}), .c ({signal_2537, signal_286}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_97 ( .a ({signal_2538, signal_288}), .b ({signal_2430, signal_864}), .c ({signal_2594, signal_832}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_98 ( .a ({1'b0, 1'b0}), .b ({signal_2462, signal_800}), .c ({signal_2538, signal_288}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_104 ( .a ({signal_2540, signal_292}), .b ({signal_2539, signal_293}), .c ({signal_2595, signal_814}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_105 ( .a ({signal_2448, signal_846}), .b ({signal_2432, signal_862}), .c ({signal_2539, signal_293}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_106 ( .a ({1'b0, 1'b0}), .b ({signal_2480, signal_782}), .c ({signal_2540, signal_292}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_107 ( .a ({signal_2541, signal_294}), .b ({signal_2432, signal_862}), .c ({signal_2596, signal_830}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_108 ( .a ({1'b0, 1'b0}), .b ({signal_2464, signal_798}), .c ({signal_2541, signal_294}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_114 ( .a ({signal_2545, signal_298}), .b ({signal_2544, signal_299}), .c ({signal_2597, signal_812}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_115 ( .a ({signal_2450, signal_844}), .b ({signal_2434, signal_860}), .c ({signal_2544, signal_299}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_116 ( .a ({1'b0, 1'b0}), .b ({signal_2482, signal_780}), .c ({signal_2545, signal_298}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_117 ( .a ({signal_2546, signal_300}), .b ({signal_2434, signal_860}), .c ({signal_2598, signal_828}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_118 ( .a ({1'b0, 1'b0}), .b ({signal_2466, signal_796}), .c ({signal_2546, signal_300}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_124 ( .a ({signal_2548, signal_304}), .b ({signal_2547, signal_305}), .c ({signal_2599, signal_810}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_125 ( .a ({signal_2452, signal_842}), .b ({signal_2436, signal_858}), .c ({signal_2547, signal_305}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_126 ( .a ({1'b0, 1'b0}), .b ({signal_2484, signal_778}), .c ({signal_2548, signal_304}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_127 ( .a ({signal_2549, signal_306}), .b ({signal_2436, signal_858}), .c ({signal_2600, signal_826}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_128 ( .a ({1'b0, 1'b0}), .b ({signal_2468, signal_794}), .c ({signal_2549, signal_306}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_134 ( .a ({signal_2553, signal_310}), .b ({signal_2552, signal_311}), .c ({signal_2601, signal_808}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_135 ( .a ({signal_2454, signal_840}), .b ({signal_2438, signal_856}), .c ({signal_2552, signal_311}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_136 ( .a ({1'b0, 1'b0}), .b ({signal_2486, signal_776}), .c ({signal_2553, signal_310}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_137 ( .a ({signal_2554, signal_312}), .b ({signal_2438, signal_856}), .c ({signal_2602, signal_824}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_138 ( .a ({1'b0, 1'b0}), .b ({signal_2470, signal_792}), .c ({signal_2554, signal_312}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_144 ( .a ({signal_2635, signal_316}), .b ({signal_2028, signal_886}), .c ({signal_2659, signal_950}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_145 ( .a ({1'b0, 1'b0}), .b ({signal_2587, signal_822}), .c ({signal_2635, signal_316}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_148 ( .a ({signal_2637, signal_318}), .b ({signal_2034, signal_884}), .c ({signal_2660, signal_948}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_149 ( .a ({1'b0, 1'b0}), .b ({signal_2589, signal_820}), .c ({signal_2637, signal_318}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_152 ( .a ({signal_2638, signal_320}), .b ({signal_2040, signal_882}), .c ({signal_2661, signal_946}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_153 ( .a ({1'b0, 1'b0}), .b ({signal_2591, signal_818}), .c ({signal_2638, signal_320}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_156 ( .a ({signal_2640, signal_322}), .b ({signal_1713, signal_880}), .c ({signal_2662, signal_944}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_157 ( .a ({1'b0, 1'b0}), .b ({signal_2593, signal_816}), .c ({signal_2640, signal_322}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_160 ( .a ({signal_2641, signal_324}), .b ({signal_1716, signal_878}), .c ({signal_2663, signal_942}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_161 ( .a ({1'b0, 1'b0}), .b ({signal_2595, signal_814}), .c ({signal_2641, signal_324}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_164 ( .a ({signal_2643, signal_326}), .b ({signal_2049, signal_876}), .c ({signal_2664, signal_940}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_165 ( .a ({1'b0, 1'b0}), .b ({signal_2597, signal_812}), .c ({signal_2643, signal_326}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_168 ( .a ({signal_2644, signal_328}), .b ({signal_2052, signal_874}), .c ({signal_2665, signal_938}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_169 ( .a ({1'b0, 1'b0}), .b ({signal_2599, signal_810}), .c ({signal_2644, signal_328}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_172 ( .a ({signal_2646, signal_330}), .b ({signal_1722, signal_872}), .c ({signal_2666, signal_936}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_173 ( .a ({1'b0, 1'b0}), .b ({signal_2601, signal_808}), .c ({signal_2646, signal_330}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_176 ( .a ({signal_2647, signal_332}), .b ({signal_2123, signal_333}), .c ({signal_2667, signal_958}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_178 ( .a ({1'b0, 1'b0}), .b ({signal_2596, signal_830}), .c ({signal_2647, signal_332}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_182 ( .a ({signal_2649, signal_336}), .b ({signal_2125, signal_337}), .c ({signal_2668, signal_956}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_184 ( .a ({1'b0, 1'b0}), .b ({signal_2598, signal_828}), .c ({signal_2649, signal_336}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_188 ( .a ({signal_2650, signal_340}), .b ({signal_2127, signal_341}), .c ({signal_2669, signal_954}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_190 ( .a ({1'b0, 1'b0}), .b ({signal_2600, signal_826}), .c ({signal_2650, signal_340}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_194 ( .a ({signal_2652, signal_344}), .b ({signal_2129, signal_345}), .c ({signal_2670, signal_952}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_196 ( .a ({1'b0, 1'b0}), .b ({signal_2602, signal_824}), .c ({signal_2652, signal_344}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_200 ( .a ({signal_2561, signal_348}), .b ({signal_1677, signal_934}), .c ({signal_2615, signal_998}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_201 ( .a ({1'b0, 1'b0}), .b ({signal_2424, signal_870}), .c ({signal_2561, signal_348}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_204 ( .a ({signal_2563, signal_350}), .b ({signal_1680, signal_932}), .c ({signal_2616, signal_996}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_205 ( .a ({1'b0, 1'b0}), .b ({signal_2426, signal_868}), .c ({signal_2563, signal_350}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_208 ( .a ({signal_2564, signal_352}), .b ({signal_1923, signal_930}), .c ({signal_2617, signal_994}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_209 ( .a ({1'b0, 1'b0}), .b ({signal_2428, signal_866}), .c ({signal_2564, signal_352}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_212 ( .a ({signal_2566, signal_354}), .b ({signal_1929, signal_928}), .c ({signal_2618, signal_992}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_213 ( .a ({1'b0, 1'b0}), .b ({signal_2430, signal_864}), .c ({signal_2566, signal_354}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_216 ( .a ({signal_2567, signal_356}), .b ({signal_1935, signal_926}), .c ({signal_2619, signal_990}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_217 ( .a ({1'b0, 1'b0}), .b ({signal_2432, signal_862}), .c ({signal_2567, signal_356}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_220 ( .a ({signal_2569, signal_358}), .b ({signal_1941, signal_924}), .c ({signal_2620, signal_988}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_221 ( .a ({1'b0, 1'b0}), .b ({signal_2434, signal_860}), .c ({signal_2569, signal_358}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_224 ( .a ({signal_2570, signal_360}), .b ({signal_1947, signal_922}), .c ({signal_2621, signal_986}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_225 ( .a ({1'b0, 1'b0}), .b ({signal_2436, signal_858}), .c ({signal_2570, signal_360}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_228 ( .a ({signal_2572, signal_362}), .b ({signal_1953, signal_920}), .c ({signal_2622, signal_984}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_229 ( .a ({1'b0, 1'b0}), .b ({signal_2438, signal_856}), .c ({signal_2572, signal_362}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_232 ( .a ({signal_2573, signal_364}), .b ({signal_1959, signal_918}), .c ({signal_2623, signal_982}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_233 ( .a ({1'b0, 1'b0}), .b ({signal_2440, signal_854}), .c ({signal_2573, signal_364}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_236 ( .a ({signal_2575, signal_366}), .b ({signal_1965, signal_916}), .c ({signal_2624, signal_980}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_237 ( .a ({1'b0, 1'b0}), .b ({signal_2442, signal_852}), .c ({signal_2575, signal_366}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_240 ( .a ({signal_2576, signal_368}), .b ({signal_1971, signal_914}), .c ({signal_2625, signal_978}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_241 ( .a ({1'b0, 1'b0}), .b ({signal_2444, signal_850}), .c ({signal_2576, signal_368}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_244 ( .a ({signal_2578, signal_370}), .b ({signal_1683, signal_912}), .c ({signal_2626, signal_976}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_245 ( .a ({1'b0, 1'b0}), .b ({signal_2446, signal_848}), .c ({signal_2578, signal_370}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_248 ( .a ({signal_2579, signal_372}), .b ({signal_1689, signal_910}), .c ({signal_2627, signal_974}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_249 ( .a ({1'b0, 1'b0}), .b ({signal_2448, signal_846}), .c ({signal_2579, signal_372}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_252 ( .a ({signal_2581, signal_374}), .b ({signal_1695, signal_908}), .c ({signal_2628, signal_972}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_253 ( .a ({1'b0, 1'b0}), .b ({signal_2450, signal_844}), .c ({signal_2581, signal_374}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_256 ( .a ({signal_2582, signal_376}), .b ({signal_1977, signal_906}), .c ({signal_2629, signal_970}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_257 ( .a ({1'b0, 1'b0}), .b ({signal_2452, signal_842}), .c ({signal_2582, signal_376}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_260 ( .a ({signal_2584, signal_378}), .b ({signal_1983, signal_904}), .c ({signal_2630, signal_968}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_261 ( .a ({1'b0, 1'b0}), .b ({signal_2454, signal_840}), .c ({signal_2584, signal_378}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_264 ( .a ({signal_2653, signal_380}), .b ({signal_1989, signal_902}), .c ({signal_2671, signal_966}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_265 ( .a ({1'b0, 1'b0}), .b ({signal_2588, signal_838}), .c ({signal_2653, signal_380}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_268 ( .a ({signal_2655, signal_382}), .b ({signal_1992, signal_900}), .c ({signal_2672, signal_964}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_269 ( .a ({1'b0, 1'b0}), .b ({signal_2590, signal_836}), .c ({signal_2655, signal_382}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_272 ( .a ({signal_2656, signal_384}), .b ({signal_1704, signal_898}), .c ({signal_2673, signal_962}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_273 ( .a ({1'b0, 1'b0}), .b ({signal_2592, signal_834}), .c ({signal_2656, signal_384}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_276 ( .a ({signal_2658, signal_386}), .b ({signal_2001, signal_896}), .c ({signal_2674, signal_960}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) cell_277 ( .a ({1'b0, 1'b0}), .b ({signal_2594, signal_832}), .c ({signal_2658, signal_386}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1331 ( .a ({signal_1835, signal_1227}), .b ({signal_2195, signal_1435}), .clk (clk), .r (Fresh[224]), .c ({signal_2323, signal_1499}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1332 ( .a ({signal_1838, signal_1230}), .b ({signal_2196, signal_1436}), .clk (clk), .r (Fresh[225]), .c ({signal_2324, signal_1500}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1333 ( .a ({signal_1841, signal_1233}), .b ({signal_2197, signal_1437}), .clk (clk), .r (Fresh[226]), .c ({signal_2325, signal_1501}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1334 ( .a ({signal_1844, signal_1236}), .b ({signal_2198, signal_1438}), .clk (clk), .r (Fresh[227]), .c ({signal_2326, signal_1502}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1335 ( .a ({signal_1847, signal_1239}), .b ({signal_2199, signal_1439}), .clk (clk), .r (Fresh[228]), .c ({signal_2327, signal_1503}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1336 ( .a ({signal_1850, signal_1242}), .b ({signal_2200, signal_1440}), .clk (clk), .r (Fresh[229]), .c ({signal_2328, signal_1504}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1337 ( .a ({signal_1853, signal_1245}), .b ({signal_2201, signal_1441}), .clk (clk), .r (Fresh[230]), .c ({signal_2329, signal_1505}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1338 ( .a ({signal_1856, signal_1248}), .b ({signal_2202, signal_1442}), .clk (clk), .r (Fresh[231]), .c ({signal_2330, signal_1506}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1339 ( .a ({signal_1859, signal_1251}), .b ({signal_2203, signal_1443}), .clk (clk), .r (Fresh[232]), .c ({signal_2331, signal_1507}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1340 ( .a ({signal_1862, signal_1254}), .b ({signal_2204, signal_1444}), .clk (clk), .r (Fresh[233]), .c ({signal_2332, signal_1508}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1341 ( .a ({signal_1865, signal_1257}), .b ({signal_2205, signal_1445}), .clk (clk), .r (Fresh[234]), .c ({signal_2333, signal_1509}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1342 ( .a ({signal_1868, signal_1260}), .b ({signal_2206, signal_1446}), .clk (clk), .r (Fresh[235]), .c ({signal_2334, signal_1510}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1343 ( .a ({signal_1871, signal_1263}), .b ({signal_2207, signal_1447}), .clk (clk), .r (Fresh[236]), .c ({signal_2335, signal_1511}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1344 ( .a ({signal_1874, signal_1266}), .b ({signal_2208, signal_1448}), .clk (clk), .r (Fresh[237]), .c ({signal_2336, signal_1512}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1345 ( .a ({signal_1877, signal_1269}), .b ({signal_2209, signal_1449}), .clk (clk), .r (Fresh[238]), .c ({signal_2337, signal_1513}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1346 ( .a ({signal_1880, signal_1272}), .b ({signal_2210, signal_1450}), .clk (clk), .r (Fresh[239]), .c ({signal_2338, signal_1514}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1347 ( .a ({signal_2323, signal_1499}), .b ({signal_2391, signal_772}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1348 ( .a ({signal_2324, signal_1500}), .b ({signal_2392, signal_768}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1349 ( .a ({signal_2325, signal_1501}), .b ({signal_2393, signal_764}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1350 ( .a ({signal_2326, signal_1502}), .b ({signal_2394, signal_760}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1351 ( .a ({signal_2327, signal_1503}), .b ({signal_2395, signal_756}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1352 ( .a ({signal_2328, signal_1504}), .b ({signal_2396, signal_752}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1353 ( .a ({signal_2329, signal_1505}), .b ({signal_2397, signal_748}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1354 ( .a ({signal_2330, signal_1506}), .b ({signal_2398, signal_744}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1355 ( .a ({signal_2331, signal_1507}), .b ({signal_2399, signal_740}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1356 ( .a ({signal_2332, signal_1508}), .b ({signal_2400, signal_736}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1357 ( .a ({signal_2333, signal_1509}), .b ({signal_2401, signal_732}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1358 ( .a ({signal_2334, signal_1510}), .b ({signal_2402, signal_728}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1359 ( .a ({signal_2335, signal_1511}), .b ({signal_2403, signal_724}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1360 ( .a ({signal_2336, signal_1512}), .b ({signal_2404, signal_720}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1361 ( .a ({signal_2337, signal_1513}), .b ({signal_2405, signal_716}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1362 ( .a ({signal_2338, signal_1514}), .b ({signal_2406, signal_712}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1363 ( .a ({signal_1739, signal_1131}), .b ({signal_2291, signal_1483}), .clk (clk), .r (Fresh[240]), .c ({signal_2407, signal_774}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1364 ( .a ({signal_1740, signal_1132}), .b ({signal_2292, signal_1484}), .clk (clk), .r (Fresh[241]), .c ({signal_2408, signal_770}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1365 ( .a ({signal_1741, signal_1133}), .b ({signal_2293, signal_1485}), .clk (clk), .r (Fresh[242]), .c ({signal_2409, signal_766}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1366 ( .a ({signal_1742, signal_1134}), .b ({signal_2294, signal_1486}), .clk (clk), .r (Fresh[243]), .c ({signal_2410, signal_762}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1367 ( .a ({signal_1743, signal_1135}), .b ({signal_2295, signal_1487}), .clk (clk), .r (Fresh[244]), .c ({signal_2411, signal_758}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1368 ( .a ({signal_1744, signal_1136}), .b ({signal_2296, signal_1488}), .clk (clk), .r (Fresh[245]), .c ({signal_2412, signal_754}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1369 ( .a ({signal_1745, signal_1137}), .b ({signal_2297, signal_1489}), .clk (clk), .r (Fresh[246]), .c ({signal_2413, signal_750}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1370 ( .a ({signal_1746, signal_1138}), .b ({signal_2298, signal_1490}), .clk (clk), .r (Fresh[247]), .c ({signal_2414, signal_746}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1371 ( .a ({signal_1747, signal_1139}), .b ({signal_2299, signal_1491}), .clk (clk), .r (Fresh[248]), .c ({signal_2415, signal_742}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1372 ( .a ({signal_1748, signal_1140}), .b ({signal_2300, signal_1492}), .clk (clk), .r (Fresh[249]), .c ({signal_2416, signal_738}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1373 ( .a ({signal_1749, signal_1141}), .b ({signal_2301, signal_1493}), .clk (clk), .r (Fresh[250]), .c ({signal_2417, signal_734}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1374 ( .a ({signal_1750, signal_1142}), .b ({signal_2302, signal_1494}), .clk (clk), .r (Fresh[251]), .c ({signal_2418, signal_730}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1375 ( .a ({signal_1751, signal_1143}), .b ({signal_2303, signal_1495}), .clk (clk), .r (Fresh[252]), .c ({signal_2419, signal_726}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1376 ( .a ({signal_1752, signal_1144}), .b ({signal_2304, signal_1496}), .clk (clk), .r (Fresh[253]), .c ({signal_2420, signal_722}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1377 ( .a ({signal_1753, signal_1145}), .b ({signal_2305, signal_1497}), .clk (clk), .r (Fresh[254]), .c ({signal_2421, signal_718}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1378 ( .a ({signal_1754, signal_1146}), .b ({signal_2306, signal_1498}), .clk (clk), .r (Fresh[255]), .c ({signal_2422, signal_714}) ) ;

    /* register cells */
    reg_masked #(.security_order(1), .pipeline(0)) cell_281 ( .clk (signal_2931), .D ({signal_2610, signal_935}), .Q ({ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_283 ( .clk (signal_2931), .D ({signal_2666, signal_936}), .Q ({ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_285 ( .clk (signal_2931), .D ({signal_2645, signal_937}), .Q ({ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_287 ( .clk (signal_2931), .D ({signal_2665, signal_938}), .Q ({ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_289 ( .clk (signal_2931), .D ({signal_2608, signal_939}), .Q ({ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_291 ( .clk (signal_2931), .D ({signal_2664, signal_940}), .Q ({ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_293 ( .clk (signal_2931), .D ({signal_2642, signal_941}), .Q ({ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_295 ( .clk (signal_2931), .D ({signal_2663, signal_942}), .Q ({ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_297 ( .clk (signal_2931), .D ({signal_2606, signal_943}), .Q ({ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_299 ( .clk (signal_2931), .D ({signal_2662, signal_944}), .Q ({ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_301 ( .clk (signal_2931), .D ({signal_2639, signal_945}), .Q ({ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_303 ( .clk (signal_2931), .D ({signal_2661, signal_946}), .Q ({ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_305 ( .clk (signal_2931), .D ({signal_2604, signal_947}), .Q ({ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_307 ( .clk (signal_2931), .D ({signal_2660, signal_948}), .Q ({ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_309 ( .clk (signal_2931), .D ({signal_2636, signal_949}), .Q ({ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_311 ( .clk (signal_2931), .D ({signal_2659, signal_950}), .Q ({ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_313 ( .clk (signal_2931), .D ({signal_2614, signal_951}), .Q ({ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_315 ( .clk (signal_2931), .D ({signal_2670, signal_952}), .Q ({ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_317 ( .clk (signal_2931), .D ({signal_2651, signal_953}), .Q ({ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_319 ( .clk (signal_2931), .D ({signal_2669, signal_954}), .Q ({ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_321 ( .clk (signal_2931), .D ({signal_2612, signal_955}), .Q ({ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_323 ( .clk (signal_2931), .D ({signal_2668, signal_956}), .Q ({ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_325 ( .clk (signal_2931), .D ({signal_2648, signal_957}), .Q ({ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_327 ( .clk (signal_2931), .D ({signal_2667, signal_958}), .Q ({ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_329 ( .clk (signal_2931), .D ({signal_2634, signal_959}), .Q ({ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_331 ( .clk (signal_2931), .D ({signal_2674, signal_960}), .Q ({ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_333 ( .clk (signal_2931), .D ({signal_2657, signal_961}), .Q ({ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_335 ( .clk (signal_2931), .D ({signal_2673, signal_962}), .Q ({ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_337 ( .clk (signal_2931), .D ({signal_2632, signal_963}), .Q ({ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_339 ( .clk (signal_2931), .D ({signal_2672, signal_964}), .Q ({ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_341 ( .clk (signal_2931), .D ({signal_2654, signal_965}), .Q ({ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_343 ( .clk (signal_2931), .D ({signal_2671, signal_966}), .Q ({ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_345 ( .clk (signal_2931), .D ({signal_2522, signal_967}), .Q ({ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_347 ( .clk (signal_2931), .D ({signal_2630, signal_968}), .Q ({ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_349 ( .clk (signal_2931), .D ({signal_2583, signal_969}), .Q ({ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_351 ( .clk (signal_2931), .D ({signal_2629, signal_970}), .Q ({ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_353 ( .clk (signal_2931), .D ({signal_2520, signal_971}), .Q ({ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_355 ( .clk (signal_2931), .D ({signal_2628, signal_972}), .Q ({ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_357 ( .clk (signal_2931), .D ({signal_2580, signal_973}), .Q ({ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_359 ( .clk (signal_2931), .D ({signal_2627, signal_974}), .Q ({ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_361 ( .clk (signal_2931), .D ({signal_2518, signal_975}), .Q ({ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_363 ( .clk (signal_2931), .D ({signal_2626, signal_976}), .Q ({ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_365 ( .clk (signal_2931), .D ({signal_2577, signal_977}), .Q ({ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_367 ( .clk (signal_2931), .D ({signal_2625, signal_978}), .Q ({ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_369 ( .clk (signal_2931), .D ({signal_2516, signal_979}), .Q ({ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_371 ( .clk (signal_2931), .D ({signal_2624, signal_980}), .Q ({ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_373 ( .clk (signal_2931), .D ({signal_2574, signal_981}), .Q ({ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_375 ( .clk (signal_2931), .D ({signal_2623, signal_982}), .Q ({ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_377 ( .clk (signal_2931), .D ({signal_2514, signal_983}), .Q ({ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_379 ( .clk (signal_2931), .D ({signal_2622, signal_984}), .Q ({ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_381 ( .clk (signal_2931), .D ({signal_2571, signal_985}), .Q ({ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_383 ( .clk (signal_2931), .D ({signal_2621, signal_986}), .Q ({ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_385 ( .clk (signal_2931), .D ({signal_2512, signal_987}), .Q ({ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_387 ( .clk (signal_2931), .D ({signal_2620, signal_988}), .Q ({ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_389 ( .clk (signal_2931), .D ({signal_2568, signal_989}), .Q ({ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_391 ( .clk (signal_2931), .D ({signal_2619, signal_990}), .Q ({ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_393 ( .clk (signal_2931), .D ({signal_2510, signal_991}), .Q ({ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_395 ( .clk (signal_2931), .D ({signal_2618, signal_992}), .Q ({ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_397 ( .clk (signal_2931), .D ({signal_2565, signal_993}), .Q ({ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_399 ( .clk (signal_2931), .D ({signal_2617, signal_994}), .Q ({ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_401 ( .clk (signal_2931), .D ({signal_2508, signal_995}), .Q ({ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_403 ( .clk (signal_2931), .D ({signal_2616, signal_996}), .Q ({ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_405 ( .clk (signal_2931), .D ({signal_2562, signal_997}), .Q ({ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_407 ( .clk (signal_2931), .D ({signal_2615, signal_998}), .Q ({ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    DFF_X1 cell_789 ( .CK (signal_2931), .D (signal_1008), .Q (signal_1001), .QN () ) ;
    DFF_X1 cell_791 ( .CK (signal_2931), .D (signal_1009), .Q (signal_1002), .QN () ) ;
    DFF_X1 cell_793 ( .CK (signal_2931), .D (signal_1010), .Q (signal_1003), .QN () ) ;
    DFF_X1 cell_795 ( .CK (signal_2931), .D (signal_1011), .Q (signal_1004), .QN () ) ;
    DFF_X1 cell_797 ( .CK (signal_2931), .D (signal_1012), .Q (signal_1005), .QN () ) ;
    DFF_X1 cell_799 ( .CK (signal_2931), .D (signal_1013), .Q (signal_1006), .QN () ) ;
    DFF_X1 cell_801 ( .CK (signal_2931), .D (signal_1014), .Q (signal_1007), .QN () ) ;
    DFF_X1 cell_814 ( .CK (signal_2931), .D (signal_1017), .Q (signal_1015), .QN () ) ;
    DFF_X1 cell_816 ( .CK (signal_2931), .D (signal_1018), .Q (signal_1016), .QN () ) ;
    DFF_X1 cell_818 ( .CK (signal_2931), .D (signal_267), .Q (done), .QN () ) ;
endmodule
