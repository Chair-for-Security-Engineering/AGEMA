
module AES_GHPCLL_ClockGating_d1 ( plaintext_s0, key_s0, clk, start, 
        plaintext_s1, key_s1, Fresh, ciphertext_s0, done, ciphertext_s1, Synch
 );
  input [127:0] plaintext_s0;
  input [127:0] key_s0;
  input [127:0] plaintext_s1;
  input [127:0] key_s1;
  input [135:0] Fresh;
  output [127:0] ciphertext_s0;
  output [127:0] ciphertext_s1;
  input clk, start;
  output done, Synch;
  wire   new_AGEMA_signal_1984, new_AGEMA_signal_1983, new_AGEMA_signal_1987,
         new_AGEMA_signal_1986, new_AGEMA_signal_1990, new_AGEMA_signal_1989,
         new_AGEMA_signal_1993, new_AGEMA_signal_1992, new_AGEMA_signal_1996,
         new_AGEMA_signal_1995, new_AGEMA_signal_1999, new_AGEMA_signal_1998,
         new_AGEMA_signal_2002, new_AGEMA_signal_2001, new_AGEMA_signal_2005,
         new_AGEMA_signal_2004, intselXOR, ctrl_N14, nReset,
         ctrl_seq6_SFF_0_QD, ctrl_seq6_SFF_1_QD, ctrl_seq6_SFF_2_QD,
         ctrl_seq6_SFF_3_QD, ctrl_seq6_SFF_4_QD, ctrl_seq4_SFF_0_QD,
         ctrl_seq4_SFF_1_QD, new_AGEMA_signal_3126,
         stateArray_S00reg_gff_1_SFF_0_QD, new_AGEMA_signal_2156,
         new_AGEMA_signal_3127, stateArray_S00reg_gff_1_SFF_1_QD,
         new_AGEMA_signal_2159, new_AGEMA_signal_3128,
         stateArray_S00reg_gff_1_SFF_2_QD, new_AGEMA_signal_2162,
         new_AGEMA_signal_3129, stateArray_S00reg_gff_1_SFF_3_QD,
         new_AGEMA_signal_2165, new_AGEMA_signal_3130,
         stateArray_S00reg_gff_1_SFF_4_QD, new_AGEMA_signal_2168,
         new_AGEMA_signal_3131, stateArray_S00reg_gff_1_SFF_5_QD,
         new_AGEMA_signal_2171, new_AGEMA_signal_3132,
         stateArray_S00reg_gff_1_SFF_6_QD, new_AGEMA_signal_2174,
         new_AGEMA_signal_3133, stateArray_S00reg_gff_1_SFF_7_QD,
         new_AGEMA_signal_2177, new_AGEMA_signal_3134,
         stateArray_S01reg_gff_1_SFF_0_QD, new_AGEMA_signal_2180,
         new_AGEMA_signal_3135, stateArray_S01reg_gff_1_SFF_1_QD,
         new_AGEMA_signal_2183, new_AGEMA_signal_3136,
         stateArray_S01reg_gff_1_SFF_2_QD, new_AGEMA_signal_2186,
         new_AGEMA_signal_3137, stateArray_S01reg_gff_1_SFF_3_QD,
         new_AGEMA_signal_2189, new_AGEMA_signal_3138,
         stateArray_S01reg_gff_1_SFF_4_QD, new_AGEMA_signal_2192,
         new_AGEMA_signal_3139, stateArray_S01reg_gff_1_SFF_5_QD,
         new_AGEMA_signal_2195, new_AGEMA_signal_3140,
         stateArray_S01reg_gff_1_SFF_6_QD, new_AGEMA_signal_2198,
         new_AGEMA_signal_3141, stateArray_S01reg_gff_1_SFF_7_QD,
         new_AGEMA_signal_2201, new_AGEMA_signal_3142,
         stateArray_S02reg_gff_1_SFF_0_QD, new_AGEMA_signal_2204,
         new_AGEMA_signal_3143, stateArray_S02reg_gff_1_SFF_1_QD,
         new_AGEMA_signal_2207, new_AGEMA_signal_3144,
         stateArray_S02reg_gff_1_SFF_2_QD, new_AGEMA_signal_2210,
         new_AGEMA_signal_3145, stateArray_S02reg_gff_1_SFF_3_QD,
         new_AGEMA_signal_2213, new_AGEMA_signal_3146,
         stateArray_S02reg_gff_1_SFF_4_QD, new_AGEMA_signal_2216,
         new_AGEMA_signal_3147, stateArray_S02reg_gff_1_SFF_5_QD,
         new_AGEMA_signal_2219, new_AGEMA_signal_3148,
         stateArray_S02reg_gff_1_SFF_6_QD, new_AGEMA_signal_2222,
         new_AGEMA_signal_3149, stateArray_S02reg_gff_1_SFF_7_QD,
         new_AGEMA_signal_2225, new_AGEMA_signal_3150,
         stateArray_S03reg_gff_1_SFF_0_QD, new_AGEMA_signal_3046,
         new_AGEMA_signal_3151, stateArray_S03reg_gff_1_SFF_1_QD,
         new_AGEMA_signal_3048, new_AGEMA_signal_3152,
         stateArray_S03reg_gff_1_SFF_2_QD, new_AGEMA_signal_3050,
         new_AGEMA_signal_3153, stateArray_S03reg_gff_1_SFF_3_QD,
         new_AGEMA_signal_3052, new_AGEMA_signal_3154,
         stateArray_S03reg_gff_1_SFF_4_QD, new_AGEMA_signal_3054,
         new_AGEMA_signal_3155, stateArray_S03reg_gff_1_SFF_5_QD,
         new_AGEMA_signal_3056, new_AGEMA_signal_3156,
         stateArray_S03reg_gff_1_SFF_6_QD, new_AGEMA_signal_3058,
         new_AGEMA_signal_3157, stateArray_S03reg_gff_1_SFF_7_QD,
         new_AGEMA_signal_3060, new_AGEMA_signal_3158,
         stateArray_S10reg_gff_1_SFF_0_QD, new_AGEMA_signal_2228,
         new_AGEMA_signal_3159, stateArray_S10reg_gff_1_SFF_1_QD,
         new_AGEMA_signal_2231, new_AGEMA_signal_3160,
         stateArray_S10reg_gff_1_SFF_2_QD, new_AGEMA_signal_2234,
         new_AGEMA_signal_3161, stateArray_S10reg_gff_1_SFF_3_QD,
         new_AGEMA_signal_2237, new_AGEMA_signal_3162,
         stateArray_S10reg_gff_1_SFF_4_QD, new_AGEMA_signal_2240,
         new_AGEMA_signal_3163, stateArray_S10reg_gff_1_SFF_5_QD,
         new_AGEMA_signal_2243, new_AGEMA_signal_3164,
         stateArray_S10reg_gff_1_SFF_6_QD, new_AGEMA_signal_2246,
         new_AGEMA_signal_3165, stateArray_S10reg_gff_1_SFF_7_QD,
         new_AGEMA_signal_2249, new_AGEMA_signal_3166,
         stateArray_S11reg_gff_1_SFF_0_QD, new_AGEMA_signal_2252,
         new_AGEMA_signal_3167, stateArray_S11reg_gff_1_SFF_1_QD,
         new_AGEMA_signal_2255, new_AGEMA_signal_3168,
         stateArray_S11reg_gff_1_SFF_2_QD, new_AGEMA_signal_2258,
         new_AGEMA_signal_3169, stateArray_S11reg_gff_1_SFF_3_QD,
         new_AGEMA_signal_2261, new_AGEMA_signal_3170,
         stateArray_S11reg_gff_1_SFF_4_QD, new_AGEMA_signal_2264,
         new_AGEMA_signal_3171, stateArray_S11reg_gff_1_SFF_5_QD,
         new_AGEMA_signal_2267, new_AGEMA_signal_3172,
         stateArray_S11reg_gff_1_SFF_6_QD, new_AGEMA_signal_2270,
         new_AGEMA_signal_3173, stateArray_S11reg_gff_1_SFF_7_QD,
         new_AGEMA_signal_2273, new_AGEMA_signal_3174,
         stateArray_S12reg_gff_1_SFF_0_QD, new_AGEMA_signal_2276,
         new_AGEMA_signal_3175, stateArray_S12reg_gff_1_SFF_1_QD,
         new_AGEMA_signal_2279, new_AGEMA_signal_3176,
         stateArray_S12reg_gff_1_SFF_2_QD, new_AGEMA_signal_2282,
         new_AGEMA_signal_3177, stateArray_S12reg_gff_1_SFF_3_QD,
         new_AGEMA_signal_2285, new_AGEMA_signal_3178,
         stateArray_S12reg_gff_1_SFF_4_QD, new_AGEMA_signal_2288,
         new_AGEMA_signal_3179, stateArray_S12reg_gff_1_SFF_5_QD,
         new_AGEMA_signal_2291, new_AGEMA_signal_3180,
         stateArray_S12reg_gff_1_SFF_6_QD, new_AGEMA_signal_2294,
         new_AGEMA_signal_3181, stateArray_S12reg_gff_1_SFF_7_QD,
         new_AGEMA_signal_2297, new_AGEMA_signal_3182,
         stateArray_S13reg_gff_1_SFF_0_QD, new_AGEMA_signal_3062,
         new_AGEMA_signal_3183, stateArray_S13reg_gff_1_SFF_1_QD,
         new_AGEMA_signal_3064, new_AGEMA_signal_3184,
         stateArray_S13reg_gff_1_SFF_2_QD, new_AGEMA_signal_3066,
         new_AGEMA_signal_3185, stateArray_S13reg_gff_1_SFF_3_QD,
         new_AGEMA_signal_3068, new_AGEMA_signal_3186,
         stateArray_S13reg_gff_1_SFF_4_QD, new_AGEMA_signal_3070,
         new_AGEMA_signal_3187, stateArray_S13reg_gff_1_SFF_5_QD,
         new_AGEMA_signal_3072, new_AGEMA_signal_3188,
         stateArray_S13reg_gff_1_SFF_6_QD, new_AGEMA_signal_3074,
         new_AGEMA_signal_3189, stateArray_S13reg_gff_1_SFF_7_QD,
         new_AGEMA_signal_3076, new_AGEMA_signal_3190,
         stateArray_S20reg_gff_1_SFF_0_QD, new_AGEMA_signal_2300,
         new_AGEMA_signal_3191, stateArray_S20reg_gff_1_SFF_1_QD,
         new_AGEMA_signal_2303, new_AGEMA_signal_3192,
         stateArray_S20reg_gff_1_SFF_2_QD, new_AGEMA_signal_2306,
         new_AGEMA_signal_3193, stateArray_S20reg_gff_1_SFF_3_QD,
         new_AGEMA_signal_2309, new_AGEMA_signal_3194,
         stateArray_S20reg_gff_1_SFF_4_QD, new_AGEMA_signal_2312,
         new_AGEMA_signal_3195, stateArray_S20reg_gff_1_SFF_5_QD,
         new_AGEMA_signal_2315, new_AGEMA_signal_3196,
         stateArray_S20reg_gff_1_SFF_6_QD, new_AGEMA_signal_2318,
         new_AGEMA_signal_3197, stateArray_S20reg_gff_1_SFF_7_QD,
         new_AGEMA_signal_2321, new_AGEMA_signal_3198,
         stateArray_S21reg_gff_1_SFF_0_QD, new_AGEMA_signal_2324,
         new_AGEMA_signal_3199, stateArray_S21reg_gff_1_SFF_1_QD,
         new_AGEMA_signal_2327, new_AGEMA_signal_3200,
         stateArray_S21reg_gff_1_SFF_2_QD, new_AGEMA_signal_2330,
         new_AGEMA_signal_3201, stateArray_S21reg_gff_1_SFF_3_QD,
         new_AGEMA_signal_2333, new_AGEMA_signal_3202,
         stateArray_S21reg_gff_1_SFF_4_QD, new_AGEMA_signal_2336,
         new_AGEMA_signal_3203, stateArray_S21reg_gff_1_SFF_5_QD,
         new_AGEMA_signal_2339, new_AGEMA_signal_3204,
         stateArray_S21reg_gff_1_SFF_6_QD, new_AGEMA_signal_2342,
         new_AGEMA_signal_3205, stateArray_S21reg_gff_1_SFF_7_QD,
         new_AGEMA_signal_2345, new_AGEMA_signal_3206,
         stateArray_S22reg_gff_1_SFF_0_QD, new_AGEMA_signal_2348,
         new_AGEMA_signal_3207, stateArray_S22reg_gff_1_SFF_1_QD,
         new_AGEMA_signal_2351, new_AGEMA_signal_3208,
         stateArray_S22reg_gff_1_SFF_2_QD, new_AGEMA_signal_2354,
         new_AGEMA_signal_3209, stateArray_S22reg_gff_1_SFF_3_QD,
         new_AGEMA_signal_2357, new_AGEMA_signal_3210,
         stateArray_S22reg_gff_1_SFF_4_QD, new_AGEMA_signal_2360,
         new_AGEMA_signal_3211, stateArray_S22reg_gff_1_SFF_5_QD,
         new_AGEMA_signal_2363, new_AGEMA_signal_3212,
         stateArray_S22reg_gff_1_SFF_6_QD, new_AGEMA_signal_2366,
         new_AGEMA_signal_3213, stateArray_S22reg_gff_1_SFF_7_QD,
         new_AGEMA_signal_2369, new_AGEMA_signal_3214,
         stateArray_S23reg_gff_1_SFF_0_QD, new_AGEMA_signal_3078,
         new_AGEMA_signal_3215, stateArray_S23reg_gff_1_SFF_1_QD,
         new_AGEMA_signal_3080, new_AGEMA_signal_3216,
         stateArray_S23reg_gff_1_SFF_2_QD, new_AGEMA_signal_3082,
         new_AGEMA_signal_3217, stateArray_S23reg_gff_1_SFF_3_QD,
         new_AGEMA_signal_3084, new_AGEMA_signal_3218,
         stateArray_S23reg_gff_1_SFF_4_QD, new_AGEMA_signal_3086,
         new_AGEMA_signal_3219, stateArray_S23reg_gff_1_SFF_5_QD,
         new_AGEMA_signal_3088, new_AGEMA_signal_3220,
         stateArray_S23reg_gff_1_SFF_6_QD, new_AGEMA_signal_3090,
         new_AGEMA_signal_3221, stateArray_S23reg_gff_1_SFF_7_QD,
         new_AGEMA_signal_3092, new_AGEMA_signal_3222,
         stateArray_S30reg_gff_1_SFF_0_QD, new_AGEMA_signal_2372,
         new_AGEMA_signal_3223, stateArray_S30reg_gff_1_SFF_1_QD,
         new_AGEMA_signal_2375, new_AGEMA_signal_3224,
         stateArray_S30reg_gff_1_SFF_2_QD, new_AGEMA_signal_2378,
         new_AGEMA_signal_3225, stateArray_S30reg_gff_1_SFF_3_QD,
         new_AGEMA_signal_2381, new_AGEMA_signal_3226,
         stateArray_S30reg_gff_1_SFF_4_QD, new_AGEMA_signal_2384,
         new_AGEMA_signal_3227, stateArray_S30reg_gff_1_SFF_5_QD,
         new_AGEMA_signal_2387, new_AGEMA_signal_3228,
         stateArray_S30reg_gff_1_SFF_6_QD, new_AGEMA_signal_2390,
         new_AGEMA_signal_3229, stateArray_S30reg_gff_1_SFF_7_QD,
         new_AGEMA_signal_2393, new_AGEMA_signal_3230,
         stateArray_S31reg_gff_1_SFF_0_QD, new_AGEMA_signal_2396,
         new_AGEMA_signal_3231, stateArray_S31reg_gff_1_SFF_1_QD,
         new_AGEMA_signal_2399, new_AGEMA_signal_3232,
         stateArray_S31reg_gff_1_SFF_2_QD, new_AGEMA_signal_2402,
         new_AGEMA_signal_3233, stateArray_S31reg_gff_1_SFF_3_QD,
         new_AGEMA_signal_2405, new_AGEMA_signal_3234,
         stateArray_S31reg_gff_1_SFF_4_QD, new_AGEMA_signal_2408,
         new_AGEMA_signal_3235, stateArray_S31reg_gff_1_SFF_5_QD,
         new_AGEMA_signal_2411, new_AGEMA_signal_3236,
         stateArray_S31reg_gff_1_SFF_6_QD, new_AGEMA_signal_2414,
         new_AGEMA_signal_3237, stateArray_S31reg_gff_1_SFF_7_QD,
         new_AGEMA_signal_2417, new_AGEMA_signal_3238,
         stateArray_S32reg_gff_1_SFF_0_QD, new_AGEMA_signal_2420,
         new_AGEMA_signal_3239, stateArray_S32reg_gff_1_SFF_1_QD,
         new_AGEMA_signal_2423, new_AGEMA_signal_3240,
         stateArray_S32reg_gff_1_SFF_2_QD, new_AGEMA_signal_2426,
         new_AGEMA_signal_3241, stateArray_S32reg_gff_1_SFF_3_QD,
         new_AGEMA_signal_2429, new_AGEMA_signal_3242,
         stateArray_S32reg_gff_1_SFF_4_QD, new_AGEMA_signal_2432,
         new_AGEMA_signal_3243, stateArray_S32reg_gff_1_SFF_5_QD,
         new_AGEMA_signal_2435, new_AGEMA_signal_3244,
         stateArray_S32reg_gff_1_SFF_6_QD, new_AGEMA_signal_2438,
         new_AGEMA_signal_3245, stateArray_S32reg_gff_1_SFF_7_QD,
         new_AGEMA_signal_2441, new_AGEMA_signal_3008, new_AGEMA_signal_2880,
         new_AGEMA_signal_3009, new_AGEMA_signal_2881, new_AGEMA_signal_3010,
         new_AGEMA_signal_2882, new_AGEMA_signal_3011, new_AGEMA_signal_2883,
         new_AGEMA_signal_3012, new_AGEMA_signal_2884, new_AGEMA_signal_3013,
         new_AGEMA_signal_2885, new_AGEMA_signal_3014, new_AGEMA_signal_2886,
         new_AGEMA_signal_3015, new_AGEMA_signal_2887, new_AGEMA_signal_3016,
         new_AGEMA_signal_2872, new_AGEMA_signal_3017, new_AGEMA_signal_2873,
         new_AGEMA_signal_3018, new_AGEMA_signal_2874, new_AGEMA_signal_3019,
         new_AGEMA_signal_2875, new_AGEMA_signal_3020, new_AGEMA_signal_2876,
         new_AGEMA_signal_3021, new_AGEMA_signal_2877, new_AGEMA_signal_3022,
         new_AGEMA_signal_2878, new_AGEMA_signal_3023, new_AGEMA_signal_2879,
         new_AGEMA_signal_3024, new_AGEMA_signal_2864, new_AGEMA_signal_3025,
         new_AGEMA_signal_2865, new_AGEMA_signal_3026, new_AGEMA_signal_2866,
         new_AGEMA_signal_3027, new_AGEMA_signal_2867, new_AGEMA_signal_3028,
         new_AGEMA_signal_2868, new_AGEMA_signal_3029, new_AGEMA_signal_2869,
         new_AGEMA_signal_3030, new_AGEMA_signal_2870, new_AGEMA_signal_3031,
         new_AGEMA_signal_2871, new_AGEMA_signal_2860, new_AGEMA_signal_2825,
         new_AGEMA_signal_2861, new_AGEMA_signal_2849, new_AGEMA_signal_2834,
         new_AGEMA_signal_2823, new_AGEMA_signal_2862, new_AGEMA_signal_2848,
         new_AGEMA_signal_2863, new_AGEMA_signal_2847, new_AGEMA_signal_2835,
         new_AGEMA_signal_2820, new_AGEMA_signal_2836, new_AGEMA_signal_2819,
         new_AGEMA_signal_2837, new_AGEMA_signal_2818, new_AGEMA_signal_2817,
         new_AGEMA_signal_2846, new_AGEMA_signal_2815, new_AGEMA_signal_2845,
         new_AGEMA_signal_2844, new_AGEMA_signal_2812, new_AGEMA_signal_2811,
         new_AGEMA_signal_2810, new_AGEMA_signal_2809, new_AGEMA_signal_2843,
         new_AGEMA_signal_2807, new_AGEMA_signal_2842, new_AGEMA_signal_2841,
         new_AGEMA_signal_2804, new_AGEMA_signal_2803, new_AGEMA_signal_2802,
         new_AGEMA_signal_2801, new_AGEMA_signal_2840, new_AGEMA_signal_2799,
         new_AGEMA_signal_2839, new_AGEMA_signal_2838, new_AGEMA_signal_2796,
         new_AGEMA_signal_2795, new_AGEMA_signal_2794, new_AGEMA_signal_2007,
         new_AGEMA_signal_2006, KeyArray_outS01ser_7_, new_AGEMA_signal_2009,
         new_AGEMA_signal_2008, KeyArray_outS01ser_6_, new_AGEMA_signal_2011,
         new_AGEMA_signal_2010, KeyArray_outS01ser_5_, new_AGEMA_signal_2013,
         new_AGEMA_signal_2012, KeyArray_outS01ser_4_, new_AGEMA_signal_2015,
         new_AGEMA_signal_2014, KeyArray_outS01ser_3_, new_AGEMA_signal_2017,
         new_AGEMA_signal_2016, KeyArray_outS01ser_2_, new_AGEMA_signal_2019,
         new_AGEMA_signal_2018, KeyArray_outS01ser_1_, new_AGEMA_signal_2021,
         new_AGEMA_signal_2020, KeyArray_outS01ser_0_, new_AGEMA_signal_3375,
         KeyArray_S00reg_gff_1_SFF_0_n5, new_AGEMA_signal_3267,
         KeyArray_S00reg_gff_1_SFF_0_QD, new_AGEMA_signal_2491,
         new_AGEMA_signal_3247, new_AGEMA_signal_3376,
         KeyArray_S00reg_gff_1_SFF_1_n6, new_AGEMA_signal_3268,
         KeyArray_S00reg_gff_1_SFF_1_QD, new_AGEMA_signal_2494,
         new_AGEMA_signal_3249, new_AGEMA_signal_3377,
         KeyArray_S00reg_gff_1_SFF_2_n6, new_AGEMA_signal_3269,
         KeyArray_S00reg_gff_1_SFF_2_QD, new_AGEMA_signal_2497,
         new_AGEMA_signal_3251, new_AGEMA_signal_3378,
         KeyArray_S00reg_gff_1_SFF_3_n6, new_AGEMA_signal_3270,
         KeyArray_S00reg_gff_1_SFF_3_QD, new_AGEMA_signal_2500,
         new_AGEMA_signal_3253, new_AGEMA_signal_3379,
         KeyArray_S00reg_gff_1_SFF_4_n6, new_AGEMA_signal_3271,
         KeyArray_S00reg_gff_1_SFF_4_QD, new_AGEMA_signal_2503,
         new_AGEMA_signal_3255, new_AGEMA_signal_3380,
         KeyArray_S00reg_gff_1_SFF_5_n6, new_AGEMA_signal_3272,
         KeyArray_S00reg_gff_1_SFF_5_QD, new_AGEMA_signal_2506,
         new_AGEMA_signal_3257, new_AGEMA_signal_3381,
         KeyArray_S00reg_gff_1_SFF_6_n6, new_AGEMA_signal_3273,
         KeyArray_S00reg_gff_1_SFF_6_QD, new_AGEMA_signal_2509,
         new_AGEMA_signal_3259, new_AGEMA_signal_3382,
         KeyArray_S00reg_gff_1_SFF_7_n6, new_AGEMA_signal_3274,
         KeyArray_S00reg_gff_1_SFF_7_QD, new_AGEMA_signal_2512,
         new_AGEMA_signal_3261, new_AGEMA_signal_3275,
         KeyArray_S01reg_gff_1_SFF_0_n6, new_AGEMA_signal_2888,
         KeyArray_S01reg_gff_1_SFF_0_QD, new_AGEMA_signal_2515,
         new_AGEMA_signal_2444, new_AGEMA_signal_3276,
         KeyArray_S01reg_gff_1_SFF_1_n6, new_AGEMA_signal_2889,
         KeyArray_S01reg_gff_1_SFF_1_QD, new_AGEMA_signal_2518,
         new_AGEMA_signal_2447, new_AGEMA_signal_3277,
         KeyArray_S01reg_gff_1_SFF_2_n6, new_AGEMA_signal_2890,
         KeyArray_S01reg_gff_1_SFF_2_QD, new_AGEMA_signal_2521,
         new_AGEMA_signal_2450, new_AGEMA_signal_3278,
         KeyArray_S01reg_gff_1_SFF_3_n6, new_AGEMA_signal_2891,
         KeyArray_S01reg_gff_1_SFF_3_QD, new_AGEMA_signal_2524,
         new_AGEMA_signal_2453, new_AGEMA_signal_3279,
         KeyArray_S01reg_gff_1_SFF_4_n6, new_AGEMA_signal_2892,
         KeyArray_S01reg_gff_1_SFF_4_QD, new_AGEMA_signal_2527,
         new_AGEMA_signal_2456, new_AGEMA_signal_3280,
         KeyArray_S01reg_gff_1_SFF_5_n6, new_AGEMA_signal_2893,
         KeyArray_S01reg_gff_1_SFF_5_QD, new_AGEMA_signal_2530,
         new_AGEMA_signal_2459, new_AGEMA_signal_3281,
         KeyArray_S01reg_gff_1_SFF_6_n6, new_AGEMA_signal_2894,
         KeyArray_S01reg_gff_1_SFF_6_QD, new_AGEMA_signal_2533,
         new_AGEMA_signal_2462, new_AGEMA_signal_3282,
         KeyArray_S01reg_gff_1_SFF_7_n6, new_AGEMA_signal_2895,
         KeyArray_S01reg_gff_1_SFF_7_QD, new_AGEMA_signal_2536,
         new_AGEMA_signal_2465, new_AGEMA_signal_3283,
         KeyArray_S02reg_gff_1_SFF_0_n6, new_AGEMA_signal_2896,
         KeyArray_S02reg_gff_1_SFF_0_QD, new_AGEMA_signal_2443,
         new_AGEMA_signal_2539, new_AGEMA_signal_2468, new_AGEMA_signal_3284,
         KeyArray_S02reg_gff_1_SFF_1_n6, new_AGEMA_signal_2897,
         KeyArray_S02reg_gff_1_SFF_1_QD, new_AGEMA_signal_2446,
         new_AGEMA_signal_2542, new_AGEMA_signal_2471, new_AGEMA_signal_3285,
         KeyArray_S02reg_gff_1_SFF_2_n6, new_AGEMA_signal_2898,
         KeyArray_S02reg_gff_1_SFF_2_QD, new_AGEMA_signal_2449,
         new_AGEMA_signal_2545, new_AGEMA_signal_2474, new_AGEMA_signal_3286,
         KeyArray_S02reg_gff_1_SFF_3_n6, new_AGEMA_signal_2899,
         KeyArray_S02reg_gff_1_SFF_3_QD, new_AGEMA_signal_2452,
         new_AGEMA_signal_2548, new_AGEMA_signal_2477, new_AGEMA_signal_3287,
         KeyArray_S02reg_gff_1_SFF_4_n6, new_AGEMA_signal_2900,
         KeyArray_S02reg_gff_1_SFF_4_QD, new_AGEMA_signal_2455,
         new_AGEMA_signal_2551, new_AGEMA_signal_2480, new_AGEMA_signal_3288,
         KeyArray_S02reg_gff_1_SFF_5_n6, new_AGEMA_signal_2901,
         KeyArray_S02reg_gff_1_SFF_5_QD, new_AGEMA_signal_2458,
         new_AGEMA_signal_2554, new_AGEMA_signal_2483, new_AGEMA_signal_3289,
         KeyArray_S02reg_gff_1_SFF_6_n6, new_AGEMA_signal_2902,
         KeyArray_S02reg_gff_1_SFF_6_QD, new_AGEMA_signal_2461,
         new_AGEMA_signal_2557, new_AGEMA_signal_2486, new_AGEMA_signal_3290,
         KeyArray_S02reg_gff_1_SFF_7_n6, new_AGEMA_signal_2903,
         KeyArray_S02reg_gff_1_SFF_7_QD, new_AGEMA_signal_2464,
         new_AGEMA_signal_2560, new_AGEMA_signal_2489, new_AGEMA_signal_3291,
         KeyArray_S03reg_gff_1_SFF_0_n6, new_AGEMA_signal_2904,
         KeyArray_S03reg_gff_1_SFF_0_QD, new_AGEMA_signal_2467,
         new_AGEMA_signal_2563, new_AGEMA_signal_2492, new_AGEMA_signal_3292,
         KeyArray_S03reg_gff_1_SFF_1_n6, new_AGEMA_signal_2905,
         KeyArray_S03reg_gff_1_SFF_1_QD, new_AGEMA_signal_2470,
         new_AGEMA_signal_2566, new_AGEMA_signal_2495, new_AGEMA_signal_3293,
         KeyArray_S03reg_gff_1_SFF_2_n6, new_AGEMA_signal_2906,
         KeyArray_S03reg_gff_1_SFF_2_QD, new_AGEMA_signal_2473,
         new_AGEMA_signal_2569, new_AGEMA_signal_2498, new_AGEMA_signal_3294,
         KeyArray_S03reg_gff_1_SFF_3_n6, new_AGEMA_signal_2907,
         KeyArray_S03reg_gff_1_SFF_3_QD, new_AGEMA_signal_2476,
         new_AGEMA_signal_2572, new_AGEMA_signal_2501, new_AGEMA_signal_3295,
         KeyArray_S03reg_gff_1_SFF_4_n6, new_AGEMA_signal_2908,
         KeyArray_S03reg_gff_1_SFF_4_QD, new_AGEMA_signal_2479,
         new_AGEMA_signal_2575, new_AGEMA_signal_2504, new_AGEMA_signal_3296,
         KeyArray_S03reg_gff_1_SFF_5_n5, new_AGEMA_signal_2909,
         KeyArray_S03reg_gff_1_SFF_5_QD, new_AGEMA_signal_2482,
         new_AGEMA_signal_2578, new_AGEMA_signal_2507, new_AGEMA_signal_3297,
         KeyArray_S03reg_gff_1_SFF_6_n5, new_AGEMA_signal_2910,
         KeyArray_S03reg_gff_1_SFF_6_QD, new_AGEMA_signal_2485,
         new_AGEMA_signal_2581, new_AGEMA_signal_2510, new_AGEMA_signal_3298,
         KeyArray_S03reg_gff_1_SFF_7_n5, new_AGEMA_signal_2911,
         KeyArray_S03reg_gff_1_SFF_7_QD, new_AGEMA_signal_2488,
         new_AGEMA_signal_2584, new_AGEMA_signal_2513, new_AGEMA_signal_3299,
         KeyArray_S10reg_gff_1_SFF_0_n5, new_AGEMA_signal_2912,
         KeyArray_S10reg_gff_1_SFF_0_QD, new_AGEMA_signal_2587,
         new_AGEMA_signal_2516, new_AGEMA_signal_3300,
         KeyArray_S10reg_gff_1_SFF_1_n5, new_AGEMA_signal_2913,
         KeyArray_S10reg_gff_1_SFF_1_QD, new_AGEMA_signal_2590,
         new_AGEMA_signal_2519, new_AGEMA_signal_3301,
         KeyArray_S10reg_gff_1_SFF_2_n5, new_AGEMA_signal_2914,
         KeyArray_S10reg_gff_1_SFF_2_QD, new_AGEMA_signal_2593,
         new_AGEMA_signal_2522, new_AGEMA_signal_3302,
         KeyArray_S10reg_gff_1_SFF_3_n5, new_AGEMA_signal_2915,
         KeyArray_S10reg_gff_1_SFF_3_QD, new_AGEMA_signal_2596,
         new_AGEMA_signal_2525, new_AGEMA_signal_3303,
         KeyArray_S10reg_gff_1_SFF_4_n5, new_AGEMA_signal_2916,
         KeyArray_S10reg_gff_1_SFF_4_QD, new_AGEMA_signal_2599,
         new_AGEMA_signal_2528, new_AGEMA_signal_3304,
         KeyArray_S10reg_gff_1_SFF_5_n5, new_AGEMA_signal_2917,
         KeyArray_S10reg_gff_1_SFF_5_QD, new_AGEMA_signal_2602,
         new_AGEMA_signal_2531, new_AGEMA_signal_3305,
         KeyArray_S10reg_gff_1_SFF_6_n5, new_AGEMA_signal_2918,
         KeyArray_S10reg_gff_1_SFF_6_QD, new_AGEMA_signal_2605,
         new_AGEMA_signal_2534, new_AGEMA_signal_3306,
         KeyArray_S10reg_gff_1_SFF_7_n5, new_AGEMA_signal_2919,
         KeyArray_S10reg_gff_1_SFF_7_QD, new_AGEMA_signal_2608,
         new_AGEMA_signal_2537, new_AGEMA_signal_3307,
         KeyArray_S11reg_gff_1_SFF_0_n6, new_AGEMA_signal_2920,
         KeyArray_S11reg_gff_1_SFF_0_QD, new_AGEMA_signal_2611,
         new_AGEMA_signal_2540, new_AGEMA_signal_3308,
         KeyArray_S11reg_gff_1_SFF_1_n6, new_AGEMA_signal_2921,
         KeyArray_S11reg_gff_1_SFF_1_QD, new_AGEMA_signal_2614,
         new_AGEMA_signal_2543, new_AGEMA_signal_3309,
         KeyArray_S11reg_gff_1_SFF_2_n6, new_AGEMA_signal_2922,
         KeyArray_S11reg_gff_1_SFF_2_QD, new_AGEMA_signal_2617,
         new_AGEMA_signal_2546, new_AGEMA_signal_3310,
         KeyArray_S11reg_gff_1_SFF_3_n6, new_AGEMA_signal_2923,
         KeyArray_S11reg_gff_1_SFF_3_QD, new_AGEMA_signal_2620,
         new_AGEMA_signal_2549, new_AGEMA_signal_3311,
         KeyArray_S11reg_gff_1_SFF_4_n6, new_AGEMA_signal_2924,
         KeyArray_S11reg_gff_1_SFF_4_QD, new_AGEMA_signal_2623,
         new_AGEMA_signal_2552, new_AGEMA_signal_3312,
         KeyArray_S11reg_gff_1_SFF_5_n6, new_AGEMA_signal_2925,
         KeyArray_S11reg_gff_1_SFF_5_QD, new_AGEMA_signal_2626,
         new_AGEMA_signal_2555, new_AGEMA_signal_3313,
         KeyArray_S11reg_gff_1_SFF_6_n6, new_AGEMA_signal_2926,
         KeyArray_S11reg_gff_1_SFF_6_QD, new_AGEMA_signal_2629,
         new_AGEMA_signal_2558, new_AGEMA_signal_3314,
         KeyArray_S11reg_gff_1_SFF_7_n6, new_AGEMA_signal_2927,
         KeyArray_S11reg_gff_1_SFF_7_QD, new_AGEMA_signal_2632,
         new_AGEMA_signal_2561, new_AGEMA_signal_3093,
         KeyArray_S12reg_gff_1_SFF_0_n6, new_AGEMA_signal_2928,
         KeyArray_S12reg_gff_1_SFF_0_QD, new_AGEMA_signal_2635,
         new_AGEMA_signal_2564, new_AGEMA_signal_3094,
         KeyArray_S12reg_gff_1_SFF_1_n6, new_AGEMA_signal_2929,
         KeyArray_S12reg_gff_1_SFF_1_QD, new_AGEMA_signal_2638,
         new_AGEMA_signal_2567, new_AGEMA_signal_3095,
         KeyArray_S12reg_gff_1_SFF_2_n6, new_AGEMA_signal_2930,
         KeyArray_S12reg_gff_1_SFF_2_QD, new_AGEMA_signal_2641,
         new_AGEMA_signal_2570, new_AGEMA_signal_3096,
         KeyArray_S12reg_gff_1_SFF_3_n6, new_AGEMA_signal_2931,
         KeyArray_S12reg_gff_1_SFF_3_QD, new_AGEMA_signal_2644,
         new_AGEMA_signal_2573, new_AGEMA_signal_3097,
         KeyArray_S12reg_gff_1_SFF_4_n6, new_AGEMA_signal_2932,
         KeyArray_S12reg_gff_1_SFF_4_QD, new_AGEMA_signal_2647,
         new_AGEMA_signal_2576, new_AGEMA_signal_3098,
         KeyArray_S12reg_gff_1_SFF_5_n6, new_AGEMA_signal_2933,
         KeyArray_S12reg_gff_1_SFF_5_QD, new_AGEMA_signal_2650,
         new_AGEMA_signal_2579, new_AGEMA_signal_3099,
         KeyArray_S12reg_gff_1_SFF_6_n6, new_AGEMA_signal_2934,
         KeyArray_S12reg_gff_1_SFF_6_QD, new_AGEMA_signal_2653,
         new_AGEMA_signal_2582, new_AGEMA_signal_3100,
         KeyArray_S12reg_gff_1_SFF_7_n6, new_AGEMA_signal_2935,
         KeyArray_S12reg_gff_1_SFF_7_QD, new_AGEMA_signal_2656,
         new_AGEMA_signal_2585, new_AGEMA_signal_3101,
         KeyArray_S13reg_gff_1_SFF_0_n6, new_AGEMA_signal_2936,
         KeyArray_S13reg_gff_1_SFF_0_QD, new_AGEMA_signal_2659,
         new_AGEMA_signal_2588, new_AGEMA_signal_3102,
         KeyArray_S13reg_gff_1_SFF_1_n6, new_AGEMA_signal_2937,
         KeyArray_S13reg_gff_1_SFF_1_QD, new_AGEMA_signal_2662,
         new_AGEMA_signal_2591, new_AGEMA_signal_3103,
         KeyArray_S13reg_gff_1_SFF_2_n6, new_AGEMA_signal_2938,
         KeyArray_S13reg_gff_1_SFF_2_QD, new_AGEMA_signal_2665,
         new_AGEMA_signal_2594, new_AGEMA_signal_3104,
         KeyArray_S13reg_gff_1_SFF_3_n6, new_AGEMA_signal_2939,
         KeyArray_S13reg_gff_1_SFF_3_QD, new_AGEMA_signal_2668,
         new_AGEMA_signal_2597, new_AGEMA_signal_3105,
         KeyArray_S13reg_gff_1_SFF_4_n6, new_AGEMA_signal_2940,
         KeyArray_S13reg_gff_1_SFF_4_QD, new_AGEMA_signal_2671,
         new_AGEMA_signal_2600, new_AGEMA_signal_3106,
         KeyArray_S13reg_gff_1_SFF_5_n5, new_AGEMA_signal_2941,
         KeyArray_S13reg_gff_1_SFF_5_QD, new_AGEMA_signal_2674,
         new_AGEMA_signal_2603, new_AGEMA_signal_3107,
         KeyArray_S13reg_gff_1_SFF_6_n5, new_AGEMA_signal_2942,
         KeyArray_S13reg_gff_1_SFF_6_QD, new_AGEMA_signal_2677,
         new_AGEMA_signal_2606, new_AGEMA_signal_3108,
         KeyArray_S13reg_gff_1_SFF_7_n5, new_AGEMA_signal_2943,
         KeyArray_S13reg_gff_1_SFF_7_QD, new_AGEMA_signal_2680,
         new_AGEMA_signal_2609, new_AGEMA_signal_3315,
         KeyArray_S20reg_gff_1_SFF_0_n5, new_AGEMA_signal_2944,
         KeyArray_S20reg_gff_1_SFF_0_QD, new_AGEMA_signal_2683,
         new_AGEMA_signal_2612, new_AGEMA_signal_3316,
         KeyArray_S20reg_gff_1_SFF_1_n5, new_AGEMA_signal_2945,
         KeyArray_S20reg_gff_1_SFF_1_QD, new_AGEMA_signal_2686,
         new_AGEMA_signal_2615, new_AGEMA_signal_3317,
         KeyArray_S20reg_gff_1_SFF_2_n5, new_AGEMA_signal_2946,
         KeyArray_S20reg_gff_1_SFF_2_QD, new_AGEMA_signal_2689,
         new_AGEMA_signal_2618, new_AGEMA_signal_3318,
         KeyArray_S20reg_gff_1_SFF_3_n5, new_AGEMA_signal_2947,
         KeyArray_S20reg_gff_1_SFF_3_QD, new_AGEMA_signal_2692,
         new_AGEMA_signal_2621, new_AGEMA_signal_3319,
         KeyArray_S20reg_gff_1_SFF_4_n5, new_AGEMA_signal_2948,
         KeyArray_S20reg_gff_1_SFF_4_QD, new_AGEMA_signal_2695,
         new_AGEMA_signal_2624, new_AGEMA_signal_3320,
         KeyArray_S20reg_gff_1_SFF_5_n5, new_AGEMA_signal_2949,
         KeyArray_S20reg_gff_1_SFF_5_QD, new_AGEMA_signal_2698,
         new_AGEMA_signal_2627, new_AGEMA_signal_3321,
         KeyArray_S20reg_gff_1_SFF_6_n5, new_AGEMA_signal_2950,
         KeyArray_S20reg_gff_1_SFF_6_QD, new_AGEMA_signal_2701,
         new_AGEMA_signal_2630, new_AGEMA_signal_3322,
         KeyArray_S20reg_gff_1_SFF_7_n5, new_AGEMA_signal_2951,
         KeyArray_S20reg_gff_1_SFF_7_QD, new_AGEMA_signal_2704,
         new_AGEMA_signal_2633, new_AGEMA_signal_3323,
         KeyArray_S21reg_gff_1_SFF_0_n6, new_AGEMA_signal_2952,
         KeyArray_S21reg_gff_1_SFF_0_QD, new_AGEMA_signal_2707,
         new_AGEMA_signal_2636, new_AGEMA_signal_3324,
         KeyArray_S21reg_gff_1_SFF_1_n6, new_AGEMA_signal_2953,
         KeyArray_S21reg_gff_1_SFF_1_QD, new_AGEMA_signal_2710,
         new_AGEMA_signal_2639, new_AGEMA_signal_3325,
         KeyArray_S21reg_gff_1_SFF_2_n6, new_AGEMA_signal_2954,
         KeyArray_S21reg_gff_1_SFF_2_QD, new_AGEMA_signal_2713,
         new_AGEMA_signal_2642, new_AGEMA_signal_3326,
         KeyArray_S21reg_gff_1_SFF_3_n6, new_AGEMA_signal_2955,
         KeyArray_S21reg_gff_1_SFF_3_QD, new_AGEMA_signal_2716,
         new_AGEMA_signal_2645, new_AGEMA_signal_3327,
         KeyArray_S21reg_gff_1_SFF_4_n6, new_AGEMA_signal_2956,
         KeyArray_S21reg_gff_1_SFF_4_QD, new_AGEMA_signal_2719,
         new_AGEMA_signal_2648, new_AGEMA_signal_3328,
         KeyArray_S21reg_gff_1_SFF_5_n6, new_AGEMA_signal_2957,
         KeyArray_S21reg_gff_1_SFF_5_QD, new_AGEMA_signal_2722,
         new_AGEMA_signal_2651, new_AGEMA_signal_3329,
         KeyArray_S21reg_gff_1_SFF_6_n6, new_AGEMA_signal_2958,
         KeyArray_S21reg_gff_1_SFF_6_QD, new_AGEMA_signal_2725,
         new_AGEMA_signal_2654, new_AGEMA_signal_3330,
         KeyArray_S21reg_gff_1_SFF_7_n6, new_AGEMA_signal_2959,
         KeyArray_S21reg_gff_1_SFF_7_QD, new_AGEMA_signal_2728,
         new_AGEMA_signal_2657, new_AGEMA_signal_3331,
         KeyArray_S22reg_gff_1_SFF_0_n6, new_AGEMA_signal_2960,
         KeyArray_S22reg_gff_1_SFF_0_QD, new_AGEMA_signal_2731,
         new_AGEMA_signal_2660, new_AGEMA_signal_3332,
         KeyArray_S22reg_gff_1_SFF_1_n6, new_AGEMA_signal_2961,
         KeyArray_S22reg_gff_1_SFF_1_QD, new_AGEMA_signal_2734,
         new_AGEMA_signal_2663, new_AGEMA_signal_3333,
         KeyArray_S22reg_gff_1_SFF_2_n6, new_AGEMA_signal_2962,
         KeyArray_S22reg_gff_1_SFF_2_QD, new_AGEMA_signal_2737,
         new_AGEMA_signal_2666, new_AGEMA_signal_3334,
         KeyArray_S22reg_gff_1_SFF_3_n6, new_AGEMA_signal_2963,
         KeyArray_S22reg_gff_1_SFF_3_QD, new_AGEMA_signal_2740,
         new_AGEMA_signal_2669, new_AGEMA_signal_3335,
         KeyArray_S22reg_gff_1_SFF_4_n6, new_AGEMA_signal_2964,
         KeyArray_S22reg_gff_1_SFF_4_QD, new_AGEMA_signal_2743,
         new_AGEMA_signal_2672, new_AGEMA_signal_3336,
         KeyArray_S22reg_gff_1_SFF_5_n6, new_AGEMA_signal_2965,
         KeyArray_S22reg_gff_1_SFF_5_QD, new_AGEMA_signal_2746,
         new_AGEMA_signal_2675, new_AGEMA_signal_3337,
         KeyArray_S22reg_gff_1_SFF_6_n6, new_AGEMA_signal_2966,
         KeyArray_S22reg_gff_1_SFF_6_QD, new_AGEMA_signal_2749,
         new_AGEMA_signal_2678, new_AGEMA_signal_3338,
         KeyArray_S22reg_gff_1_SFF_7_n6, new_AGEMA_signal_2967,
         KeyArray_S22reg_gff_1_SFF_7_QD, new_AGEMA_signal_2752,
         new_AGEMA_signal_2681, new_AGEMA_signal_3339,
         KeyArray_S23reg_gff_1_SFF_0_n6, new_AGEMA_signal_2968,
         KeyArray_S23reg_gff_1_SFF_0_QD, new_AGEMA_signal_2755,
         new_AGEMA_signal_2684, new_AGEMA_signal_3340,
         KeyArray_S23reg_gff_1_SFF_1_n6, new_AGEMA_signal_2969,
         KeyArray_S23reg_gff_1_SFF_1_QD, new_AGEMA_signal_2758,
         new_AGEMA_signal_2687, new_AGEMA_signal_3341,
         KeyArray_S23reg_gff_1_SFF_2_n6, new_AGEMA_signal_2970,
         KeyArray_S23reg_gff_1_SFF_2_QD, new_AGEMA_signal_2761,
         new_AGEMA_signal_2690, new_AGEMA_signal_3342,
         KeyArray_S23reg_gff_1_SFF_3_n6, new_AGEMA_signal_2971,
         KeyArray_S23reg_gff_1_SFF_3_QD, new_AGEMA_signal_2764,
         new_AGEMA_signal_2693, new_AGEMA_signal_3343,
         KeyArray_S23reg_gff_1_SFF_4_n6, new_AGEMA_signal_2972,
         KeyArray_S23reg_gff_1_SFF_4_QD, new_AGEMA_signal_2767,
         new_AGEMA_signal_2696, new_AGEMA_signal_3344,
         KeyArray_S23reg_gff_1_SFF_5_n5, new_AGEMA_signal_2973,
         KeyArray_S23reg_gff_1_SFF_5_QD, new_AGEMA_signal_2770,
         new_AGEMA_signal_2699, new_AGEMA_signal_3345,
         KeyArray_S23reg_gff_1_SFF_6_n5, new_AGEMA_signal_2974,
         KeyArray_S23reg_gff_1_SFF_6_QD, new_AGEMA_signal_2773,
         new_AGEMA_signal_2702, new_AGEMA_signal_3346,
         KeyArray_S23reg_gff_1_SFF_7_n5, new_AGEMA_signal_2975,
         KeyArray_S23reg_gff_1_SFF_7_QD, new_AGEMA_signal_2776,
         new_AGEMA_signal_2705, new_AGEMA_signal_3347,
         KeyArray_S31reg_gff_1_SFF_0_n6, new_AGEMA_signal_2976,
         KeyArray_S31reg_gff_1_SFF_0_QD, new_AGEMA_signal_2732,
         new_AGEMA_signal_3348, KeyArray_S31reg_gff_1_SFF_1_n6,
         new_AGEMA_signal_2977, KeyArray_S31reg_gff_1_SFF_1_QD,
         new_AGEMA_signal_2735, new_AGEMA_signal_3349,
         KeyArray_S31reg_gff_1_SFF_2_n6, new_AGEMA_signal_2978,
         KeyArray_S31reg_gff_1_SFF_2_QD, new_AGEMA_signal_2738,
         new_AGEMA_signal_3350, KeyArray_S31reg_gff_1_SFF_3_n6,
         new_AGEMA_signal_2979, KeyArray_S31reg_gff_1_SFF_3_QD,
         new_AGEMA_signal_2741, new_AGEMA_signal_3351,
         KeyArray_S31reg_gff_1_SFF_4_n6, new_AGEMA_signal_2980,
         KeyArray_S31reg_gff_1_SFF_4_QD, new_AGEMA_signal_2744,
         new_AGEMA_signal_3352, KeyArray_S31reg_gff_1_SFF_5_n6,
         new_AGEMA_signal_2981, KeyArray_S31reg_gff_1_SFF_5_QD,
         new_AGEMA_signal_2747, new_AGEMA_signal_3353,
         KeyArray_S31reg_gff_1_SFF_6_n6, new_AGEMA_signal_2982,
         KeyArray_S31reg_gff_1_SFF_6_QD, new_AGEMA_signal_2750,
         new_AGEMA_signal_3354, KeyArray_S31reg_gff_1_SFF_7_n6,
         new_AGEMA_signal_2983, KeyArray_S31reg_gff_1_SFF_7_QD,
         new_AGEMA_signal_2753, new_AGEMA_signal_3355,
         KeyArray_S32reg_gff_1_SFF_0_n6, new_AGEMA_signal_2984,
         KeyArray_S32reg_gff_1_SFF_0_QD, new_AGEMA_signal_2756,
         new_AGEMA_signal_3356, KeyArray_S32reg_gff_1_SFF_1_n6,
         new_AGEMA_signal_2985, KeyArray_S32reg_gff_1_SFF_1_QD,
         new_AGEMA_signal_2759, new_AGEMA_signal_3357,
         KeyArray_S32reg_gff_1_SFF_2_n6, new_AGEMA_signal_2986,
         KeyArray_S32reg_gff_1_SFF_2_QD, new_AGEMA_signal_2762,
         new_AGEMA_signal_3358, KeyArray_S32reg_gff_1_SFF_3_n6,
         new_AGEMA_signal_2987, KeyArray_S32reg_gff_1_SFF_3_QD,
         new_AGEMA_signal_2765, new_AGEMA_signal_3359,
         KeyArray_S32reg_gff_1_SFF_4_n6, new_AGEMA_signal_2988,
         KeyArray_S32reg_gff_1_SFF_4_QD, new_AGEMA_signal_2768,
         new_AGEMA_signal_3360, KeyArray_S32reg_gff_1_SFF_5_n6,
         new_AGEMA_signal_2989, KeyArray_S32reg_gff_1_SFF_5_QD,
         new_AGEMA_signal_2771, new_AGEMA_signal_3361,
         KeyArray_S32reg_gff_1_SFF_6_n5, new_AGEMA_signal_2990,
         KeyArray_S32reg_gff_1_SFF_6_QD, new_AGEMA_signal_2774,
         new_AGEMA_signal_3362, KeyArray_S32reg_gff_1_SFF_7_n5,
         new_AGEMA_signal_2991, KeyArray_S32reg_gff_1_SFF_7_QD,
         new_AGEMA_signal_2777, new_AGEMA_signal_3363,
         KeyArray_S33reg_gff_1_SFF_0_n5, new_AGEMA_signal_2992,
         KeyArray_S33reg_gff_1_SFF_0_QD, new_AGEMA_signal_2779,
         new_AGEMA_signal_3364, KeyArray_S33reg_gff_1_SFF_1_n5,
         new_AGEMA_signal_2993, KeyArray_S33reg_gff_1_SFF_1_QD,
         new_AGEMA_signal_2781, new_AGEMA_signal_3365,
         KeyArray_S33reg_gff_1_SFF_2_n5, new_AGEMA_signal_2994,
         KeyArray_S33reg_gff_1_SFF_2_QD, new_AGEMA_signal_2783,
         new_AGEMA_signal_3366, KeyArray_S33reg_gff_1_SFF_3_n5,
         new_AGEMA_signal_2995, KeyArray_S33reg_gff_1_SFF_3_QD,
         new_AGEMA_signal_2785, new_AGEMA_signal_3367,
         KeyArray_S33reg_gff_1_SFF_4_n5, new_AGEMA_signal_2996,
         KeyArray_S33reg_gff_1_SFF_4_QD, new_AGEMA_signal_2787,
         new_AGEMA_signal_3368, KeyArray_S33reg_gff_1_SFF_5_n5,
         new_AGEMA_signal_2997, KeyArray_S33reg_gff_1_SFF_5_QD,
         new_AGEMA_signal_2789, new_AGEMA_signal_3369,
         KeyArray_S33reg_gff_1_SFF_6_n5, new_AGEMA_signal_2998,
         KeyArray_S33reg_gff_1_SFF_6_QD, new_AGEMA_signal_2791,
         new_AGEMA_signal_3370, KeyArray_S33reg_gff_1_SFF_7_n5,
         new_AGEMA_signal_2999, KeyArray_S33reg_gff_1_SFF_7_QD,
         new_AGEMA_signal_2793, new_AGEMA_signal_3109, new_AGEMA_signal_3110,
         new_AGEMA_signal_3111, new_AGEMA_signal_3112, new_AGEMA_signal_3113,
         new_AGEMA_signal_3114, new_AGEMA_signal_3115, new_AGEMA_signal_3116,
         new_AGEMA_signal_2708, new_AGEMA_signal_2711, new_AGEMA_signal_2714,
         new_AGEMA_signal_2717, new_AGEMA_signal_2720, new_AGEMA_signal_2723,
         new_AGEMA_signal_2726, new_AGEMA_signal_2729, new_AGEMA_signal_2024,
         MixColumns_line0_n15, new_AGEMA_signal_2122, MixColumns_line0_n16,
         new_AGEMA_signal_2051, new_AGEMA_signal_2027, MixColumns_line0_n13,
         new_AGEMA_signal_2123, MixColumns_line0_n14, new_AGEMA_signal_2053,
         new_AGEMA_signal_2030, MixColumns_line0_n11, new_AGEMA_signal_2124,
         MixColumns_line0_n12, new_AGEMA_signal_2055, new_AGEMA_signal_2033,
         MixColumns_line0_n9, new_AGEMA_signal_2797, MixColumns_line0_n10,
         new_AGEMA_signal_2127, MixColumns_line0_S02_1, new_AGEMA_signal_2046,
         new_AGEMA_signal_2036, MixColumns_line0_n7, new_AGEMA_signal_2798,
         MixColumns_line0_n8, new_AGEMA_signal_2128, new_AGEMA_signal_2047,
         new_AGEMA_signal_2039, MixColumns_line0_n5, new_AGEMA_signal_2125,
         MixColumns_line0_n6, new_AGEMA_signal_2058, new_AGEMA_signal_2042,
         MixColumns_line0_n3, new_AGEMA_signal_2800, MixColumns_line0_n4,
         new_AGEMA_signal_2129, new_AGEMA_signal_2048, new_AGEMA_signal_2045,
         MixColumns_line0_n1, new_AGEMA_signal_2126, MixColumns_line0_n2,
         new_AGEMA_signal_2060, MixColumns_line0_timesTHREE_input2_1,
         new_AGEMA_signal_2062, new_AGEMA_signal_2063, new_AGEMA_signal_2064,
         new_AGEMA_signal_2065, MixColumns_line1_n15, new_AGEMA_signal_2130,
         MixColumns_line1_n16, new_AGEMA_signal_2076, new_AGEMA_signal_2066,
         MixColumns_line1_n13, new_AGEMA_signal_2131, MixColumns_line1_n14,
         new_AGEMA_signal_2077, new_AGEMA_signal_2067, MixColumns_line1_n11,
         new_AGEMA_signal_2132, MixColumns_line1_n12, new_AGEMA_signal_2078,
         new_AGEMA_signal_2068, MixColumns_line1_n9, new_AGEMA_signal_2805,
         MixColumns_line1_n10, new_AGEMA_signal_2135, new_AGEMA_signal_2073,
         MixColumns_line1_S02_4_, new_AGEMA_signal_2069, MixColumns_line1_n7,
         new_AGEMA_signal_2806, MixColumns_line1_n8, new_AGEMA_signal_2136,
         new_AGEMA_signal_2074, MixColumns_line1_S02_3_, new_AGEMA_signal_2070,
         MixColumns_line1_n5, new_AGEMA_signal_2133, MixColumns_line1_n6,
         new_AGEMA_signal_2079, new_AGEMA_signal_2071, MixColumns_line1_n3,
         new_AGEMA_signal_2808, MixColumns_line1_n4, new_AGEMA_signal_2137,
         new_AGEMA_signal_2075, MixColumns_line1_S02_1_, new_AGEMA_signal_2072,
         MixColumns_line1_n1, new_AGEMA_signal_2134, MixColumns_line1_n2,
         new_AGEMA_signal_2080, MixColumns_line1_timesTHREE_input2_1,
         new_AGEMA_signal_2081, new_AGEMA_signal_2082, new_AGEMA_signal_2083,
         new_AGEMA_signal_2084, MixColumns_line2_n15, new_AGEMA_signal_2138,
         MixColumns_line2_n16, new_AGEMA_signal_2095, new_AGEMA_signal_2085,
         MixColumns_line2_n13, new_AGEMA_signal_2139, MixColumns_line2_n14,
         new_AGEMA_signal_2096, new_AGEMA_signal_2086, MixColumns_line2_n11,
         new_AGEMA_signal_2140, MixColumns_line2_n12, new_AGEMA_signal_2097,
         new_AGEMA_signal_2087, MixColumns_line2_n9, new_AGEMA_signal_2813,
         MixColumns_line2_n10, new_AGEMA_signal_2143, new_AGEMA_signal_2092,
         MixColumns_line2_S02_4_, new_AGEMA_signal_2088, MixColumns_line2_n7,
         new_AGEMA_signal_2814, MixColumns_line2_n8, new_AGEMA_signal_2144,
         new_AGEMA_signal_2093, MixColumns_line2_S02_3_, new_AGEMA_signal_2089,
         MixColumns_line2_n5, new_AGEMA_signal_2141, MixColumns_line2_n6,
         new_AGEMA_signal_2098, new_AGEMA_signal_2090, MixColumns_line2_n3,
         new_AGEMA_signal_2816, MixColumns_line2_n4, new_AGEMA_signal_2145,
         new_AGEMA_signal_2094, MixColumns_line2_S02_1_, new_AGEMA_signal_2091,
         MixColumns_line2_n1, new_AGEMA_signal_2142, MixColumns_line2_n2,
         new_AGEMA_signal_2099, MixColumns_line2_timesTHREE_input2_1,
         new_AGEMA_signal_2100, new_AGEMA_signal_2101, new_AGEMA_signal_2102,
         new_AGEMA_signal_2103, MixColumns_line3_n15, new_AGEMA_signal_2146,
         MixColumns_line3_n16, new_AGEMA_signal_2114, new_AGEMA_signal_2104,
         MixColumns_line3_n13, new_AGEMA_signal_2147, MixColumns_line3_n14,
         new_AGEMA_signal_2115, new_AGEMA_signal_2105, MixColumns_line3_n11,
         new_AGEMA_signal_2148, MixColumns_line3_n12, new_AGEMA_signal_2116,
         new_AGEMA_signal_2106, MixColumns_line3_n9, new_AGEMA_signal_2821,
         MixColumns_line3_n10, new_AGEMA_signal_2151, new_AGEMA_signal_2111,
         MixColumns_line3_S02_4_, new_AGEMA_signal_2107, MixColumns_line3_n7,
         new_AGEMA_signal_2822, MixColumns_line3_n8, new_AGEMA_signal_2152,
         new_AGEMA_signal_2112, MixColumns_line3_S02_3_, new_AGEMA_signal_2108,
         MixColumns_line3_n5, new_AGEMA_signal_2149, MixColumns_line3_n6,
         new_AGEMA_signal_2117, new_AGEMA_signal_2109, MixColumns_line3_n3,
         new_AGEMA_signal_2824, MixColumns_line3_n4, new_AGEMA_signal_2153,
         new_AGEMA_signal_2113, MixColumns_line3_S02_1_, new_AGEMA_signal_2110,
         MixColumns_line3_n1, new_AGEMA_signal_2150, MixColumns_line3_n2,
         new_AGEMA_signal_2118, new_AGEMA_signal_2119,
         MixColumns_line3_timesTHREE_input2_4_, new_AGEMA_signal_2120,
         MixColumns_line3_timesTHREE_input2_3_, new_AGEMA_signal_2121,
         MixColumns_line3_timesTHREE_input2_1_, calcRCon_n51, calcRCon_n50,
         calcRCon_n49, calcRCon_n48, calcRCon_n47, calcRCon_n46, calcRCon_n45,
         calcRCon_n44, new_AGEMA_signal_2826, new_AGEMA_signal_2827,
         new_AGEMA_signal_2828, new_AGEMA_signal_2829, new_AGEMA_signal_2830,
         new_AGEMA_signal_2831, new_AGEMA_signal_2832, new_AGEMA_signal_2833,
         new_AGEMA_signal_2850, Inst_bSbox_T1, new_AGEMA_signal_2851,
         Inst_bSbox_T2, new_AGEMA_signal_2852, Inst_bSbox_T3,
         new_AGEMA_signal_2853, Inst_bSbox_T4, new_AGEMA_signal_2854,
         Inst_bSbox_T5, new_AGEMA_signal_3000, Inst_bSbox_T6,
         new_AGEMA_signal_2855, Inst_bSbox_T7, new_AGEMA_signal_3032,
         Inst_bSbox_T8, new_AGEMA_signal_3001, Inst_bSbox_T9,
         new_AGEMA_signal_3033, Inst_bSbox_T10, new_AGEMA_signal_2856,
         Inst_bSbox_T11, new_AGEMA_signal_2857, Inst_bSbox_T12,
         new_AGEMA_signal_3002, Inst_bSbox_T13, new_AGEMA_signal_3034,
         Inst_bSbox_T14, new_AGEMA_signal_3003, Inst_bSbox_T15,
         new_AGEMA_signal_3004, Inst_bSbox_T16, new_AGEMA_signal_3035,
         Inst_bSbox_T17, new_AGEMA_signal_2858, Inst_bSbox_T18,
         new_AGEMA_signal_3005, Inst_bSbox_T19, new_AGEMA_signal_3036,
         Inst_bSbox_T20, new_AGEMA_signal_2859, Inst_bSbox_T21,
         new_AGEMA_signal_3006, Inst_bSbox_T22, new_AGEMA_signal_3037,
         Inst_bSbox_T23, new_AGEMA_signal_3117, Inst_bSbox_T24,
         new_AGEMA_signal_3118, Inst_bSbox_T25, new_AGEMA_signal_3038,
         Inst_bSbox_T26, new_AGEMA_signal_3007, Inst_bSbox_T27, clk_gated,
         new_AGEMA_signal_3039, Inst_bSbox_M1, new_AGEMA_signal_3119,
         Inst_bSbox_M2, new_AGEMA_signal_3120, Inst_bSbox_M3,
         new_AGEMA_signal_3040, Inst_bSbox_M4, new_AGEMA_signal_3121,
         Inst_bSbox_M5, new_AGEMA_signal_3041, Inst_bSbox_M6,
         new_AGEMA_signal_3042, Inst_bSbox_M7, new_AGEMA_signal_3122,
         Inst_bSbox_M8, new_AGEMA_signal_3123, Inst_bSbox_M9,
         new_AGEMA_signal_3262, Inst_bSbox_M10, new_AGEMA_signal_3043,
         Inst_bSbox_M11, new_AGEMA_signal_3044, Inst_bSbox_M12,
         new_AGEMA_signal_3124, Inst_bSbox_M13, new_AGEMA_signal_3125,
         Inst_bSbox_M14, new_AGEMA_signal_3263, Inst_bSbox_M15,
         new_AGEMA_signal_3264, Inst_bSbox_M16, new_AGEMA_signal_3265,
         Inst_bSbox_M17, new_AGEMA_signal_3266, Inst_bSbox_M18,
         new_AGEMA_signal_3371, Inst_bSbox_M19, new_AGEMA_signal_3372,
         Inst_bSbox_M20, new_AGEMA_signal_3373, Inst_bSbox_M21,
         new_AGEMA_signal_3374, Inst_bSbox_M22, new_AGEMA_signal_3383,
         Inst_bSbox_M23, new_AGEMA_signal_3387, Inst_bSbox_M24,
         new_AGEMA_signal_3385, Inst_bSbox_M27, new_AGEMA_signal_3384,
         Inst_bSbox_M25, new_AGEMA_signal_3388, Inst_bSbox_M26,
         new_AGEMA_signal_3389, Inst_bSbox_M28, new_AGEMA_signal_3390,
         Inst_bSbox_M31, new_AGEMA_signal_3391, Inst_bSbox_M33,
         new_AGEMA_signal_3386, Inst_bSbox_M34, new_AGEMA_signal_3396,
         Inst_bSbox_M36, new_AGEMA_signal_3392, Inst_bSbox_M29,
         new_AGEMA_signal_3393, Inst_bSbox_M30, new_AGEMA_signal_3394,
         Inst_bSbox_M32, new_AGEMA_signal_3395, Inst_bSbox_M35,
         new_AGEMA_signal_3397, Inst_bSbox_M37, new_AGEMA_signal_3398,
         Inst_bSbox_M38, new_AGEMA_signal_3399, Inst_bSbox_M39,
         new_AGEMA_signal_3400, Inst_bSbox_M40, new_AGEMA_signal_3401,
         Inst_bSbox_M41, new_AGEMA_signal_3402, Inst_bSbox_M42,
         new_AGEMA_signal_3403, Inst_bSbox_M43, new_AGEMA_signal_3404,
         Inst_bSbox_M44, new_AGEMA_signal_3413, Inst_bSbox_M45,
         new_AGEMA_signal_3455, new_AGEMA_signal_3454, new_AGEMA_signal_3464,
         new_AGEMA_signal_3463, new_AGEMA_signal_3465, new_AGEMA_signal_3462,
         new_AGEMA_signal_3466, new_AGEMA_signal_3461, new_AGEMA_signal_3467,
         new_AGEMA_signal_3460, new_AGEMA_signal_3468, new_AGEMA_signal_3459,
         new_AGEMA_signal_3469, new_AGEMA_signal_3458, new_AGEMA_signal_3470,
         new_AGEMA_signal_3457, new_AGEMA_signal_3497,
         stateArray_S33reg_gff_1_SFF_0_QD, new_AGEMA_signal_3488,
         new_AGEMA_signal_3520, stateArray_S33reg_gff_1_SFF_1_QD,
         new_AGEMA_signal_3499, new_AGEMA_signal_3521,
         stateArray_S33reg_gff_1_SFF_2_QD, new_AGEMA_signal_3501,
         new_AGEMA_signal_3522, stateArray_S33reg_gff_1_SFF_3_QD,
         new_AGEMA_signal_3503, new_AGEMA_signal_3523,
         stateArray_S33reg_gff_1_SFF_4_QD, new_AGEMA_signal_3505,
         new_AGEMA_signal_3524, stateArray_S33reg_gff_1_SFF_5_QD,
         new_AGEMA_signal_3507, new_AGEMA_signal_3525,
         stateArray_S33reg_gff_1_SFF_6_QD, new_AGEMA_signal_3509,
         new_AGEMA_signal_3526, stateArray_S33reg_gff_1_SFF_7_QD,
         new_AGEMA_signal_3511, new_AGEMA_signal_3471, new_AGEMA_signal_3480,
         new_AGEMA_signal_3481, new_AGEMA_signal_3482, new_AGEMA_signal_3483,
         new_AGEMA_signal_3484, new_AGEMA_signal_3485, new_AGEMA_signal_3486,
         new_AGEMA_signal_3489, new_AGEMA_signal_3472, KeyArray_n55,
         new_AGEMA_signal_3490, new_AGEMA_signal_3473, KeyArray_n54,
         new_AGEMA_signal_3491, new_AGEMA_signal_3474, KeyArray_n53,
         new_AGEMA_signal_3492, new_AGEMA_signal_3475, KeyArray_n52,
         new_AGEMA_signal_3493, new_AGEMA_signal_3476, KeyArray_n51,
         new_AGEMA_signal_3494, new_AGEMA_signal_3477, KeyArray_n50,
         new_AGEMA_signal_3495, new_AGEMA_signal_3478, KeyArray_n49,
         new_AGEMA_signal_3479, new_AGEMA_signal_3456, KeyArray_n48,
         new_AGEMA_signal_3512, KeyArray_S30reg_gff_1_SFF_0_n5,
         new_AGEMA_signal_3496, KeyArray_S30reg_gff_1_SFF_0_QD,
         new_AGEMA_signal_3527, KeyArray_S30reg_gff_1_SFF_1_n5,
         new_AGEMA_signal_3513, KeyArray_S30reg_gff_1_SFF_1_QD,
         new_AGEMA_signal_3528, KeyArray_S30reg_gff_1_SFF_2_n5,
         new_AGEMA_signal_3514, KeyArray_S30reg_gff_1_SFF_2_QD,
         new_AGEMA_signal_3529, KeyArray_S30reg_gff_1_SFF_3_n5,
         new_AGEMA_signal_3515, KeyArray_S30reg_gff_1_SFF_3_QD,
         new_AGEMA_signal_3530, KeyArray_S30reg_gff_1_SFF_4_n5,
         new_AGEMA_signal_3516, KeyArray_S30reg_gff_1_SFF_4_QD,
         new_AGEMA_signal_3531, KeyArray_S30reg_gff_1_SFF_5_n5,
         new_AGEMA_signal_3517, KeyArray_S30reg_gff_1_SFF_5_QD,
         new_AGEMA_signal_3532, KeyArray_S30reg_gff_1_SFF_6_n5,
         new_AGEMA_signal_3518, KeyArray_S30reg_gff_1_SFF_6_QD,
         new_AGEMA_signal_3533, KeyArray_S30reg_gff_1_SFF_7_n5,
         new_AGEMA_signal_3519, KeyArray_S30reg_gff_1_SFF_7_QD,
         new_AGEMA_signal_3414, Inst_bSbox_M46, new_AGEMA_signal_3405,
         Inst_bSbox_M47, new_AGEMA_signal_3406, Inst_bSbox_M48,
         new_AGEMA_signal_3415, Inst_bSbox_M49, new_AGEMA_signal_3407,
         Inst_bSbox_M50, new_AGEMA_signal_3408, Inst_bSbox_M51,
         new_AGEMA_signal_3416, Inst_bSbox_M52, new_AGEMA_signal_3425,
         Inst_bSbox_M53, new_AGEMA_signal_3417, Inst_bSbox_M54,
         new_AGEMA_signal_3418, Inst_bSbox_M55, new_AGEMA_signal_3409,
         Inst_bSbox_M56, new_AGEMA_signal_3410, Inst_bSbox_M57,
         new_AGEMA_signal_3419, Inst_bSbox_M58, new_AGEMA_signal_3411,
         Inst_bSbox_M59, new_AGEMA_signal_3412, Inst_bSbox_M60,
         new_AGEMA_signal_3420, Inst_bSbox_M61, new_AGEMA_signal_3426,
         Inst_bSbox_M62, new_AGEMA_signal_3421, Inst_bSbox_M63,
         new_AGEMA_signal_3435, Inst_bSbox_L0, new_AGEMA_signal_3422,
         Inst_bSbox_L1, new_AGEMA_signal_3427, Inst_bSbox_L2,
         new_AGEMA_signal_3428, Inst_bSbox_L3, new_AGEMA_signal_3429,
         Inst_bSbox_L4, new_AGEMA_signal_3430, Inst_bSbox_L5,
         new_AGEMA_signal_3436, Inst_bSbox_L6, new_AGEMA_signal_3437,
         Inst_bSbox_L7, new_AGEMA_signal_3423, Inst_bSbox_L8,
         new_AGEMA_signal_3438, Inst_bSbox_L9, new_AGEMA_signal_3439,
         Inst_bSbox_L10, new_AGEMA_signal_3440, Inst_bSbox_L11,
         new_AGEMA_signal_3424, Inst_bSbox_L12, new_AGEMA_signal_3444,
         Inst_bSbox_L13, new_AGEMA_signal_3431, Inst_bSbox_L14,
         new_AGEMA_signal_3432, Inst_bSbox_L15, new_AGEMA_signal_3445,
         Inst_bSbox_L16, new_AGEMA_signal_3433, Inst_bSbox_L17,
         new_AGEMA_signal_3434, Inst_bSbox_L18, new_AGEMA_signal_3441,
         Inst_bSbox_L19, new_AGEMA_signal_3446, Inst_bSbox_L20,
         new_AGEMA_signal_3447, Inst_bSbox_L21, new_AGEMA_signal_3442,
         Inst_bSbox_L22, new_AGEMA_signal_3443, Inst_bSbox_L23,
         new_AGEMA_signal_3448, Inst_bSbox_L24, new_AGEMA_signal_3449,
         Inst_bSbox_L25, new_AGEMA_signal_3450, Inst_bSbox_L26,
         new_AGEMA_signal_3451, Inst_bSbox_L27, new_AGEMA_signal_3452,
         Inst_bSbox_L28, new_AGEMA_signal_3453, Inst_bSbox_L29, n3, n36, n114,
         n124, n125, n126, n128, n129, n130, n131, n133, n135, n136, n137,
         n138, n139, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244,
         Inst_bSbox_XOR_T6_U1_Ins_1_n2, ClockGatingInst_n5,
         ClockGatingInst_n10, ClockGatingInst_n9, ClockGatingInst_n8,
         ClockGatingInst_n7, ClockGatingInst_n6, ClockGatingInst_n4,
         ClockGatingInst_n3, ClockGatingInst_n2, ClockGatingInst_n1,
         ClockGatingInst_LatchedEnable, ClockGatingInst_N7,
         ClockGatingInst_ShiftRegister_5_, Inst_bSbox_AND_M1_U1_n3,
         Inst_bSbox_AND_M1_U1_n2, Inst_bSbox_AND_M1_U1_n1,
         Inst_bSbox_AND_M1_U1_out0_mid_0_, Inst_bSbox_AND_M1_U1_Step1_ins_n17,
         Inst_bSbox_AND_M1_U1_Step1_ins_n16,
         Inst_bSbox_AND_M1_U1_Step1_ins_n15,
         Inst_bSbox_AND_M1_U1_Step1_ins_n14,
         Inst_bSbox_AND_M1_U1_Step1_ins_n13,
         Inst_bSbox_AND_M1_U1_Step2_inst_n11,
         Inst_bSbox_AND_M1_U1_Step2_inst_n10,
         Inst_bSbox_AND_M1_U1_Step2_inst_n9, Inst_bSbox_AND_M2_U1_n11,
         Inst_bSbox_AND_M2_U1_n10, Inst_bSbox_AND_M2_U1_n9,
         Inst_bSbox_AND_M2_U1_out0_mid_0_, Inst_bSbox_AND_M2_U1_Step1_ins_n17,
         Inst_bSbox_AND_M2_U1_Step1_ins_n16,
         Inst_bSbox_AND_M2_U1_Step1_ins_n15,
         Inst_bSbox_AND_M2_U1_Step1_ins_n14,
         Inst_bSbox_AND_M2_U1_Step1_ins_n13,
         Inst_bSbox_AND_M2_U1_Step2_inst_n11,
         Inst_bSbox_AND_M2_U1_Step2_inst_n10,
         Inst_bSbox_AND_M2_U1_Step2_inst_n9, Inst_bSbox_AND_M4_U1_n11,
         Inst_bSbox_AND_M4_U1_n10, Inst_bSbox_AND_M4_U1_n9,
         Inst_bSbox_AND_M4_U1_out0_mid_0_, Inst_bSbox_AND_M4_U1_Step1_ins_n17,
         Inst_bSbox_AND_M4_U1_Step1_ins_n16,
         Inst_bSbox_AND_M4_U1_Step1_ins_n15,
         Inst_bSbox_AND_M4_U1_Step1_ins_n14,
         Inst_bSbox_AND_M4_U1_Step1_ins_n13,
         Inst_bSbox_AND_M4_U1_Step2_inst_n11,
         Inst_bSbox_AND_M4_U1_Step2_inst_n10,
         Inst_bSbox_AND_M4_U1_Step2_inst_n9, Inst_bSbox_AND_M6_U1_n11,
         Inst_bSbox_AND_M6_U1_n10, Inst_bSbox_AND_M6_U1_n9,
         Inst_bSbox_AND_M6_U1_out0_mid_0_, Inst_bSbox_AND_M6_U1_Step1_ins_n17,
         Inst_bSbox_AND_M6_U1_Step1_ins_n16,
         Inst_bSbox_AND_M6_U1_Step1_ins_n15,
         Inst_bSbox_AND_M6_U1_Step1_ins_n14,
         Inst_bSbox_AND_M6_U1_Step1_ins_n13,
         Inst_bSbox_AND_M6_U1_Step2_inst_n11,
         Inst_bSbox_AND_M6_U1_Step2_inst_n10,
         Inst_bSbox_AND_M6_U1_Step2_inst_n9, Inst_bSbox_AND_M7_U1_n11,
         Inst_bSbox_AND_M7_U1_n10, Inst_bSbox_AND_M7_U1_n9,
         Inst_bSbox_AND_M7_U1_out0_mid_0_, Inst_bSbox_AND_M7_U1_Step1_ins_n17,
         Inst_bSbox_AND_M7_U1_Step1_ins_n16,
         Inst_bSbox_AND_M7_U1_Step1_ins_n15,
         Inst_bSbox_AND_M7_U1_Step1_ins_n14,
         Inst_bSbox_AND_M7_U1_Step1_ins_n13,
         Inst_bSbox_AND_M7_U1_Step2_inst_n11,
         Inst_bSbox_AND_M7_U1_Step2_inst_n10,
         Inst_bSbox_AND_M7_U1_Step2_inst_n9, Inst_bSbox_AND_M9_U1_n11,
         Inst_bSbox_AND_M9_U1_n10, Inst_bSbox_AND_M9_U1_n9,
         Inst_bSbox_AND_M9_U1_out0_mid_0_, Inst_bSbox_AND_M9_U1_Step1_ins_n17,
         Inst_bSbox_AND_M9_U1_Step1_ins_n16,
         Inst_bSbox_AND_M9_U1_Step1_ins_n15,
         Inst_bSbox_AND_M9_U1_Step1_ins_n14,
         Inst_bSbox_AND_M9_U1_Step1_ins_n13,
         Inst_bSbox_AND_M9_U1_Step2_inst_n11,
         Inst_bSbox_AND_M9_U1_Step2_inst_n10,
         Inst_bSbox_AND_M9_U1_Step2_inst_n9, Inst_bSbox_AND_M11_U1_n11,
         Inst_bSbox_AND_M11_U1_n10, Inst_bSbox_AND_M11_U1_n9,
         Inst_bSbox_AND_M11_U1_out0_mid_0_,
         Inst_bSbox_AND_M11_U1_Step1_ins_n17,
         Inst_bSbox_AND_M11_U1_Step1_ins_n16,
         Inst_bSbox_AND_M11_U1_Step1_ins_n15,
         Inst_bSbox_AND_M11_U1_Step1_ins_n14,
         Inst_bSbox_AND_M11_U1_Step1_ins_n13,
         Inst_bSbox_AND_M11_U1_Step2_inst_n11,
         Inst_bSbox_AND_M11_U1_Step2_inst_n10,
         Inst_bSbox_AND_M11_U1_Step2_inst_n9, Inst_bSbox_AND_M12_U1_n11,
         Inst_bSbox_AND_M12_U1_n10, Inst_bSbox_AND_M12_U1_n9,
         Inst_bSbox_AND_M12_U1_out0_mid_0_,
         Inst_bSbox_AND_M12_U1_Step1_ins_n17,
         Inst_bSbox_AND_M12_U1_Step1_ins_n16,
         Inst_bSbox_AND_M12_U1_Step1_ins_n15,
         Inst_bSbox_AND_M12_U1_Step1_ins_n14,
         Inst_bSbox_AND_M12_U1_Step1_ins_n13,
         Inst_bSbox_AND_M12_U1_Step2_inst_n11,
         Inst_bSbox_AND_M12_U1_Step2_inst_n10,
         Inst_bSbox_AND_M12_U1_Step2_inst_n9, Inst_bSbox_AND_M14_U1_n11,
         Inst_bSbox_AND_M14_U1_n10, Inst_bSbox_AND_M14_U1_n9,
         Inst_bSbox_AND_M14_U1_out0_mid_0_,
         Inst_bSbox_AND_M14_U1_Step1_ins_n17,
         Inst_bSbox_AND_M14_U1_Step1_ins_n16,
         Inst_bSbox_AND_M14_U1_Step1_ins_n15,
         Inst_bSbox_AND_M14_U1_Step1_ins_n14,
         Inst_bSbox_AND_M14_U1_Step1_ins_n13,
         Inst_bSbox_AND_M14_U1_Step2_inst_n11,
         Inst_bSbox_AND_M14_U1_Step2_inst_n10,
         Inst_bSbox_AND_M14_U1_Step2_inst_n9, Inst_bSbox_AND_M25_U1_n11,
         Inst_bSbox_AND_M25_U1_n10, Inst_bSbox_AND_M25_U1_n9,
         Inst_bSbox_AND_M25_U1_out0_mid_0_,
         Inst_bSbox_AND_M25_U1_Step1_ins_n17,
         Inst_bSbox_AND_M25_U1_Step1_ins_n16,
         Inst_bSbox_AND_M25_U1_Step1_ins_n15,
         Inst_bSbox_AND_M25_U1_Step1_ins_n14,
         Inst_bSbox_AND_M25_U1_Step1_ins_n13,
         Inst_bSbox_AND_M25_U1_Step2_inst_n11,
         Inst_bSbox_AND_M25_U1_Step2_inst_n10,
         Inst_bSbox_AND_M25_U1_Step2_inst_n9, Inst_bSbox_AND_M31_U1_n11,
         Inst_bSbox_AND_M31_U1_n10, Inst_bSbox_AND_M31_U1_n9,
         Inst_bSbox_AND_M31_U1_out0_mid_0_,
         Inst_bSbox_AND_M31_U1_Step1_ins_n17,
         Inst_bSbox_AND_M31_U1_Step1_ins_n16,
         Inst_bSbox_AND_M31_U1_Step1_ins_n15,
         Inst_bSbox_AND_M31_U1_Step1_ins_n14,
         Inst_bSbox_AND_M31_U1_Step1_ins_n13,
         Inst_bSbox_AND_M31_U1_Step2_inst_n11,
         Inst_bSbox_AND_M31_U1_Step2_inst_n10,
         Inst_bSbox_AND_M31_U1_Step2_inst_n9, Inst_bSbox_AND_M34_U1_n11,
         Inst_bSbox_AND_M34_U1_n10, Inst_bSbox_AND_M34_U1_n9,
         Inst_bSbox_AND_M34_U1_out0_mid_0_,
         Inst_bSbox_AND_M34_U1_Step1_ins_n17,
         Inst_bSbox_AND_M34_U1_Step1_ins_n16,
         Inst_bSbox_AND_M34_U1_Step1_ins_n15,
         Inst_bSbox_AND_M34_U1_Step1_ins_n14,
         Inst_bSbox_AND_M34_U1_Step1_ins_n13,
         Inst_bSbox_AND_M34_U1_Step2_inst_n11,
         Inst_bSbox_AND_M34_U1_Step2_inst_n10,
         Inst_bSbox_AND_M34_U1_Step2_inst_n9, Inst_bSbox_AND_M29_U1_n11,
         Inst_bSbox_AND_M29_U1_n10, Inst_bSbox_AND_M29_U1_n9,
         Inst_bSbox_AND_M29_U1_out0_mid_0_,
         Inst_bSbox_AND_M29_U1_Step1_ins_n17,
         Inst_bSbox_AND_M29_U1_Step1_ins_n16,
         Inst_bSbox_AND_M29_U1_Step1_ins_n15,
         Inst_bSbox_AND_M29_U1_Step1_ins_n14,
         Inst_bSbox_AND_M29_U1_Step1_ins_n13,
         Inst_bSbox_AND_M29_U1_Step2_inst_n11,
         Inst_bSbox_AND_M29_U1_Step2_inst_n10,
         Inst_bSbox_AND_M29_U1_Step2_inst_n9, Inst_bSbox_AND_M30_U1_n11,
         Inst_bSbox_AND_M30_U1_n10, Inst_bSbox_AND_M30_U1_n9,
         Inst_bSbox_AND_M30_U1_out0_mid_0_,
         Inst_bSbox_AND_M30_U1_Step1_ins_n17,
         Inst_bSbox_AND_M30_U1_Step1_ins_n16,
         Inst_bSbox_AND_M30_U1_Step1_ins_n15,
         Inst_bSbox_AND_M30_U1_Step1_ins_n14,
         Inst_bSbox_AND_M30_U1_Step1_ins_n13,
         Inst_bSbox_AND_M30_U1_Step2_inst_n11,
         Inst_bSbox_AND_M30_U1_Step2_inst_n10,
         Inst_bSbox_AND_M30_U1_Step2_inst_n9, Inst_bSbox_AND_M32_U1_n11,
         Inst_bSbox_AND_M32_U1_n10, Inst_bSbox_AND_M32_U1_n9,
         Inst_bSbox_AND_M32_U1_out0_mid_0_,
         Inst_bSbox_AND_M32_U1_Step1_ins_n17,
         Inst_bSbox_AND_M32_U1_Step1_ins_n16,
         Inst_bSbox_AND_M32_U1_Step1_ins_n15,
         Inst_bSbox_AND_M32_U1_Step1_ins_n14,
         Inst_bSbox_AND_M32_U1_Step1_ins_n13,
         Inst_bSbox_AND_M32_U1_Step2_inst_n11,
         Inst_bSbox_AND_M32_U1_Step2_inst_n10,
         Inst_bSbox_AND_M32_U1_Step2_inst_n9, Inst_bSbox_AND_M35_U1_n11,
         Inst_bSbox_AND_M35_U1_n10, Inst_bSbox_AND_M35_U1_n9,
         Inst_bSbox_AND_M35_U1_out0_mid_0_,
         Inst_bSbox_AND_M35_U1_Step1_ins_n17,
         Inst_bSbox_AND_M35_U1_Step1_ins_n16,
         Inst_bSbox_AND_M35_U1_Step1_ins_n15,
         Inst_bSbox_AND_M35_U1_Step1_ins_n14,
         Inst_bSbox_AND_M35_U1_Step1_ins_n13,
         Inst_bSbox_AND_M35_U1_Step2_inst_n11,
         Inst_bSbox_AND_M35_U1_Step2_inst_n10,
         Inst_bSbox_AND_M35_U1_Step2_inst_n9, Inst_bSbox_AND_M46_U1_n11,
         Inst_bSbox_AND_M46_U1_n10, Inst_bSbox_AND_M46_U1_n9,
         Inst_bSbox_AND_M46_U1_out0_mid_0_,
         Inst_bSbox_AND_M46_U1_Step1_ins_n17,
         Inst_bSbox_AND_M46_U1_Step1_ins_n16,
         Inst_bSbox_AND_M46_U1_Step1_ins_n15,
         Inst_bSbox_AND_M46_U1_Step1_ins_n14,
         Inst_bSbox_AND_M46_U1_Step1_ins_n13,
         Inst_bSbox_AND_M46_U1_Step2_inst_n11,
         Inst_bSbox_AND_M46_U1_Step2_inst_n10,
         Inst_bSbox_AND_M46_U1_Step2_inst_n9, Inst_bSbox_AND_M47_U1_n11,
         Inst_bSbox_AND_M47_U1_n10, Inst_bSbox_AND_M47_U1_n9,
         Inst_bSbox_AND_M47_U1_out0_mid_0_,
         Inst_bSbox_AND_M47_U1_Step1_ins_n17,
         Inst_bSbox_AND_M47_U1_Step1_ins_n16,
         Inst_bSbox_AND_M47_U1_Step1_ins_n15,
         Inst_bSbox_AND_M47_U1_Step1_ins_n14,
         Inst_bSbox_AND_M47_U1_Step1_ins_n13,
         Inst_bSbox_AND_M47_U1_Step2_inst_n11,
         Inst_bSbox_AND_M47_U1_Step2_inst_n10,
         Inst_bSbox_AND_M47_U1_Step2_inst_n9, Inst_bSbox_AND_M48_U1_n11,
         Inst_bSbox_AND_M48_U1_n10, Inst_bSbox_AND_M48_U1_n9,
         Inst_bSbox_AND_M48_U1_out0_mid_0_,
         Inst_bSbox_AND_M48_U1_Step1_ins_n17,
         Inst_bSbox_AND_M48_U1_Step1_ins_n16,
         Inst_bSbox_AND_M48_U1_Step1_ins_n15,
         Inst_bSbox_AND_M48_U1_Step1_ins_n14,
         Inst_bSbox_AND_M48_U1_Step1_ins_n13,
         Inst_bSbox_AND_M48_U1_Step2_inst_n11,
         Inst_bSbox_AND_M48_U1_Step2_inst_n10,
         Inst_bSbox_AND_M48_U1_Step2_inst_n9, Inst_bSbox_AND_M49_U1_n11,
         Inst_bSbox_AND_M49_U1_n10, Inst_bSbox_AND_M49_U1_n9,
         Inst_bSbox_AND_M49_U1_out0_mid_0_,
         Inst_bSbox_AND_M49_U1_Step1_ins_n17,
         Inst_bSbox_AND_M49_U1_Step1_ins_n16,
         Inst_bSbox_AND_M49_U1_Step1_ins_n15,
         Inst_bSbox_AND_M49_U1_Step1_ins_n14,
         Inst_bSbox_AND_M49_U1_Step1_ins_n13,
         Inst_bSbox_AND_M49_U1_Step2_inst_n11,
         Inst_bSbox_AND_M49_U1_Step2_inst_n10,
         Inst_bSbox_AND_M49_U1_Step2_inst_n9, Inst_bSbox_AND_M50_U1_n11,
         Inst_bSbox_AND_M50_U1_n10, Inst_bSbox_AND_M50_U1_n9,
         Inst_bSbox_AND_M50_U1_out0_mid_0_,
         Inst_bSbox_AND_M50_U1_Step1_ins_n17,
         Inst_bSbox_AND_M50_U1_Step1_ins_n16,
         Inst_bSbox_AND_M50_U1_Step1_ins_n15,
         Inst_bSbox_AND_M50_U1_Step1_ins_n14,
         Inst_bSbox_AND_M50_U1_Step1_ins_n13,
         Inst_bSbox_AND_M50_U1_Step2_inst_n11,
         Inst_bSbox_AND_M50_U1_Step2_inst_n10,
         Inst_bSbox_AND_M50_U1_Step2_inst_n9, Inst_bSbox_AND_M51_U1_n11,
         Inst_bSbox_AND_M51_U1_n10, Inst_bSbox_AND_M51_U1_n9,
         Inst_bSbox_AND_M51_U1_out0_mid_0_,
         Inst_bSbox_AND_M51_U1_Step1_ins_n17,
         Inst_bSbox_AND_M51_U1_Step1_ins_n16,
         Inst_bSbox_AND_M51_U1_Step1_ins_n15,
         Inst_bSbox_AND_M51_U1_Step1_ins_n14,
         Inst_bSbox_AND_M51_U1_Step1_ins_n13,
         Inst_bSbox_AND_M51_U1_Step2_inst_n11,
         Inst_bSbox_AND_M51_U1_Step2_inst_n10,
         Inst_bSbox_AND_M51_U1_Step2_inst_n9, Inst_bSbox_AND_M52_U1_n11,
         Inst_bSbox_AND_M52_U1_n10, Inst_bSbox_AND_M52_U1_n9,
         Inst_bSbox_AND_M52_U1_out0_mid_0_,
         Inst_bSbox_AND_M52_U1_Step1_ins_n17,
         Inst_bSbox_AND_M52_U1_Step1_ins_n16,
         Inst_bSbox_AND_M52_U1_Step1_ins_n15,
         Inst_bSbox_AND_M52_U1_Step1_ins_n14,
         Inst_bSbox_AND_M52_U1_Step1_ins_n13,
         Inst_bSbox_AND_M52_U1_Step2_inst_n11,
         Inst_bSbox_AND_M52_U1_Step2_inst_n10,
         Inst_bSbox_AND_M52_U1_Step2_inst_n9, Inst_bSbox_AND_M53_U1_n11,
         Inst_bSbox_AND_M53_U1_n10, Inst_bSbox_AND_M53_U1_n9,
         Inst_bSbox_AND_M53_U1_out0_mid_0_,
         Inst_bSbox_AND_M53_U1_Step1_ins_n17,
         Inst_bSbox_AND_M53_U1_Step1_ins_n16,
         Inst_bSbox_AND_M53_U1_Step1_ins_n15,
         Inst_bSbox_AND_M53_U1_Step1_ins_n14,
         Inst_bSbox_AND_M53_U1_Step1_ins_n13,
         Inst_bSbox_AND_M53_U1_Step2_inst_n11,
         Inst_bSbox_AND_M53_U1_Step2_inst_n10,
         Inst_bSbox_AND_M53_U1_Step2_inst_n9, Inst_bSbox_AND_M54_U1_n11,
         Inst_bSbox_AND_M54_U1_n10, Inst_bSbox_AND_M54_U1_n9,
         Inst_bSbox_AND_M54_U1_out0_mid_0_,
         Inst_bSbox_AND_M54_U1_Step1_ins_n17,
         Inst_bSbox_AND_M54_U1_Step1_ins_n16,
         Inst_bSbox_AND_M54_U1_Step1_ins_n15,
         Inst_bSbox_AND_M54_U1_Step1_ins_n14,
         Inst_bSbox_AND_M54_U1_Step1_ins_n13,
         Inst_bSbox_AND_M54_U1_Step2_inst_n11,
         Inst_bSbox_AND_M54_U1_Step2_inst_n10,
         Inst_bSbox_AND_M54_U1_Step2_inst_n9, Inst_bSbox_AND_M55_U1_n11,
         Inst_bSbox_AND_M55_U1_n10, Inst_bSbox_AND_M55_U1_n9,
         Inst_bSbox_AND_M55_U1_out0_mid_0_,
         Inst_bSbox_AND_M55_U1_Step1_ins_n17,
         Inst_bSbox_AND_M55_U1_Step1_ins_n16,
         Inst_bSbox_AND_M55_U1_Step1_ins_n15,
         Inst_bSbox_AND_M55_U1_Step1_ins_n14,
         Inst_bSbox_AND_M55_U1_Step1_ins_n13,
         Inst_bSbox_AND_M55_U1_Step2_inst_n11,
         Inst_bSbox_AND_M55_U1_Step2_inst_n10,
         Inst_bSbox_AND_M55_U1_Step2_inst_n9, Inst_bSbox_AND_M56_U1_n11,
         Inst_bSbox_AND_M56_U1_n10, Inst_bSbox_AND_M56_U1_n9,
         Inst_bSbox_AND_M56_U1_out0_mid_0_,
         Inst_bSbox_AND_M56_U1_Step1_ins_n17,
         Inst_bSbox_AND_M56_U1_Step1_ins_n16,
         Inst_bSbox_AND_M56_U1_Step1_ins_n15,
         Inst_bSbox_AND_M56_U1_Step1_ins_n14,
         Inst_bSbox_AND_M56_U1_Step1_ins_n13,
         Inst_bSbox_AND_M56_U1_Step2_inst_n11,
         Inst_bSbox_AND_M56_U1_Step2_inst_n10,
         Inst_bSbox_AND_M56_U1_Step2_inst_n9, Inst_bSbox_AND_M57_U1_n11,
         Inst_bSbox_AND_M57_U1_n10, Inst_bSbox_AND_M57_U1_n9,
         Inst_bSbox_AND_M57_U1_out0_mid_0_,
         Inst_bSbox_AND_M57_U1_Step1_ins_n17,
         Inst_bSbox_AND_M57_U1_Step1_ins_n16,
         Inst_bSbox_AND_M57_U1_Step1_ins_n15,
         Inst_bSbox_AND_M57_U1_Step1_ins_n14,
         Inst_bSbox_AND_M57_U1_Step1_ins_n13,
         Inst_bSbox_AND_M57_U1_Step2_inst_n11,
         Inst_bSbox_AND_M57_U1_Step2_inst_n10,
         Inst_bSbox_AND_M57_U1_Step2_inst_n9, Inst_bSbox_AND_M58_U1_n11,
         Inst_bSbox_AND_M58_U1_n10, Inst_bSbox_AND_M58_U1_n9,
         Inst_bSbox_AND_M58_U1_out0_mid_0_,
         Inst_bSbox_AND_M58_U1_Step1_ins_n17,
         Inst_bSbox_AND_M58_U1_Step1_ins_n16,
         Inst_bSbox_AND_M58_U1_Step1_ins_n15,
         Inst_bSbox_AND_M58_U1_Step1_ins_n14,
         Inst_bSbox_AND_M58_U1_Step1_ins_n13,
         Inst_bSbox_AND_M58_U1_Step2_inst_n11,
         Inst_bSbox_AND_M58_U1_Step2_inst_n10,
         Inst_bSbox_AND_M58_U1_Step2_inst_n9, Inst_bSbox_AND_M59_U1_n11,
         Inst_bSbox_AND_M59_U1_n10, Inst_bSbox_AND_M59_U1_n9,
         Inst_bSbox_AND_M59_U1_out0_mid_0_,
         Inst_bSbox_AND_M59_U1_Step1_ins_n17,
         Inst_bSbox_AND_M59_U1_Step1_ins_n16,
         Inst_bSbox_AND_M59_U1_Step1_ins_n15,
         Inst_bSbox_AND_M59_U1_Step1_ins_n14,
         Inst_bSbox_AND_M59_U1_Step1_ins_n13,
         Inst_bSbox_AND_M59_U1_Step2_inst_n11,
         Inst_bSbox_AND_M59_U1_Step2_inst_n10,
         Inst_bSbox_AND_M59_U1_Step2_inst_n9, Inst_bSbox_AND_M60_U1_n11,
         Inst_bSbox_AND_M60_U1_n10, Inst_bSbox_AND_M60_U1_n9,
         Inst_bSbox_AND_M60_U1_out0_mid_0_,
         Inst_bSbox_AND_M60_U1_Step1_ins_n17,
         Inst_bSbox_AND_M60_U1_Step1_ins_n16,
         Inst_bSbox_AND_M60_U1_Step1_ins_n15,
         Inst_bSbox_AND_M60_U1_Step1_ins_n14,
         Inst_bSbox_AND_M60_U1_Step1_ins_n13,
         Inst_bSbox_AND_M60_U1_Step2_inst_n11,
         Inst_bSbox_AND_M60_U1_Step2_inst_n10,
         Inst_bSbox_AND_M60_U1_Step2_inst_n9, Inst_bSbox_AND_M61_U1_n11,
         Inst_bSbox_AND_M61_U1_n10, Inst_bSbox_AND_M61_U1_n9,
         Inst_bSbox_AND_M61_U1_out0_mid_0_,
         Inst_bSbox_AND_M61_U1_Step1_ins_n17,
         Inst_bSbox_AND_M61_U1_Step1_ins_n16,
         Inst_bSbox_AND_M61_U1_Step1_ins_n15,
         Inst_bSbox_AND_M61_U1_Step1_ins_n14,
         Inst_bSbox_AND_M61_U1_Step1_ins_n13,
         Inst_bSbox_AND_M61_U1_Step2_inst_n11,
         Inst_bSbox_AND_M61_U1_Step2_inst_n10,
         Inst_bSbox_AND_M61_U1_Step2_inst_n9, Inst_bSbox_AND_M62_U1_n11,
         Inst_bSbox_AND_M62_U1_n10, Inst_bSbox_AND_M62_U1_n9,
         Inst_bSbox_AND_M62_U1_out0_mid_0_,
         Inst_bSbox_AND_M62_U1_Step1_ins_n17,
         Inst_bSbox_AND_M62_U1_Step1_ins_n16,
         Inst_bSbox_AND_M62_U1_Step1_ins_n15,
         Inst_bSbox_AND_M62_U1_Step1_ins_n14,
         Inst_bSbox_AND_M62_U1_Step1_ins_n13,
         Inst_bSbox_AND_M62_U1_Step2_inst_n11,
         Inst_bSbox_AND_M62_U1_Step2_inst_n10,
         Inst_bSbox_AND_M62_U1_Step2_inst_n9, Inst_bSbox_AND_M63_U1_n11,
         Inst_bSbox_AND_M63_U1_n10, Inst_bSbox_AND_M63_U1_n9,
         Inst_bSbox_AND_M63_U1_out0_mid_0_,
         Inst_bSbox_AND_M63_U1_Step1_ins_n17,
         Inst_bSbox_AND_M63_U1_Step1_ins_n16,
         Inst_bSbox_AND_M63_U1_Step1_ins_n15,
         Inst_bSbox_AND_M63_U1_Step1_ins_n14,
         Inst_bSbox_AND_M63_U1_Step1_ins_n13,
         Inst_bSbox_AND_M63_U1_Step2_inst_n11,
         Inst_bSbox_AND_M63_U1_Step2_inst_n10,
         Inst_bSbox_AND_M63_U1_Step2_inst_n9;
  wire   [7:0] StateOutXORroundKey;
  wire   [7:0] keyStateIn;
  wire   [7:0] stateArray_inS00ser;
  wire   [7:0] stateArray_inS01ser;
  wire   [7:0] stateArray_inS02ser;
  wire   [7:0] stateArray_inS03ser;
  wire   [7:0] stateArray_inS10ser;
  wire   [7:0] stateArray_inS11ser;
  wire   [7:0] stateArray_inS12ser;
  wire   [7:0] stateArray_inS13ser;
  wire   [7:0] stateArray_inS20ser;
  wire   [7:0] stateArray_inS21ser;
  wire   [7:0] stateArray_inS22ser;
  wire   [7:0] stateArray_inS23ser;
  wire   [7:0] stateArray_inS30ser;
  wire   [7:0] stateArray_inS31ser;
  wire   [7:0] stateArray_inS32ser;
  wire   [7:0] stateArray_outS10ser_MC;
  wire   [31:0] StateInMC;
  wire   [7:0] stateArray_outS20ser_MC;
  wire   [7:0] stateArray_outS30ser_MC;
  wire   [31:0] MCout;
  wire   [7:0] KeyArray_outS01ser_XOR_00;
  wire   [7:0] KeyArray_outS10ser;
  wire   [7:0] KeyArray_inS00ser;
  wire   [7:0] KeyArray_outS11ser;
  wire   [7:0] KeyArray_inS01ser;
  wire   [7:0] KeyArray_outS02ser;
  wire   [7:0] KeyArray_outS12ser;
  wire   [7:0] KeyArray_inS02ser;
  wire   [7:0] KeyArray_outS03ser;
  wire   [7:0] keySBIn;
  wire   [7:0] KeyArray_inS03ser;
  wire   [7:0] KeyArray_outS20ser;
  wire   [7:0] KeyArray_inS10ser;
  wire   [7:0] KeyArray_outS21ser;
  wire   [7:0] KeyArray_inS11ser;
  wire   [7:0] KeyArray_outS22ser;
  wire   [7:0] KeyArray_inS12ser;
  wire   [7:0] KeyArray_outS23ser;
  wire   [7:0] KeyArray_inS13ser;
  wire   [7:0] KeyArray_outS30ser;
  wire   [7:0] KeyArray_inS20ser;
  wire   [7:0] KeyArray_outS31ser;
  wire   [7:0] KeyArray_inS21ser;
  wire   [7:0] KeyArray_outS32ser;
  wire   [7:0] KeyArray_inS22ser;
  wire   [7:0] KeyArray_outS33ser;
  wire   [7:0] KeyArray_inS23ser;
  wire   [7:0] KeyArray_inS31ser;
  wire   [7:0] KeyArray_inS32ser;
  wire   [7:0] KeyArray_inS33ser;
  wire   [7:0] KeyArray_outS01ser_p;
  wire   [7:0] KeyArray_inS30ser;
  wire   [7:0] MixColumns_line0_S13;
  wire   [4:3] MixColumns_line0_S02;
  wire   [4:3] MixColumns_line0_timesTHREE_input2;
  wire   [7:0] MixColumns_line1_S13;
  wire   [4:3] MixColumns_line1_timesTHREE_input2;
  wire   [7:0] MixColumns_line2_S13;
  wire   [4:3] MixColumns_line2_timesTHREE_input2;
  wire   [7:0] MixColumns_line3_S13;
  wire   [7:0] roundConstant;
  wire   [7:0] SboxIn;
  wire   [7:0] StateIn;
  wire   [7:0] SboxOut;
  wire   [7:0] stateArray_inS33ser;
  wire   [7:0] stateArray_input_MC;
  wire   [7:0] KeyArray_inS30par;
  wire   [3:0] Inst_bSbox_AND_M1_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M1_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M1_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M2_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M2_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M2_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M4_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M4_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M4_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M6_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M6_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M6_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M7_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M7_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M7_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M9_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M9_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M9_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M11_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M11_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M11_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M12_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M12_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M12_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M14_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M14_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M14_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M25_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M25_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M25_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M31_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M31_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M31_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M34_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M34_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M34_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M29_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M29_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M29_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M30_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M30_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M30_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M32_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M32_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M32_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M35_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M35_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M35_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M46_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M46_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M46_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M47_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M47_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M47_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M48_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M48_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M48_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M49_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M49_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M49_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M50_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M50_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M50_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M51_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M51_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M51_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M52_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M52_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M52_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M53_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M53_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M53_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M54_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M54_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M54_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M55_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M55_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M55_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M56_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M56_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M56_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M57_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M57_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M57_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M58_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M58_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M58_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M59_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M59_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M59_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M60_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M60_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M60_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M61_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M61_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M61_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M62_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M62_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M62_U1_Step1_ins_Step1;
  wire   [3:0] Inst_bSbox_AND_M63_U1_Step1_reg;
  wire   [1:0] Inst_bSbox_AND_M63_U1_in1_reg;
  wire   [3:0] Inst_bSbox_AND_M63_U1_Step1_ins_Step1;

  DFF_X1 ctrl_CSselMC_reg_FF_FF ( .D(ctrl_N14), .CK(clk_gated), .Q(), .QN(n124) );
  DFF_X1 nReset_reg_FF_FF ( .D(n114), .CK(clk_gated), .Q(nReset), .QN(n149) );
  DFF_X1 ctrl_seq6_SFF_3_Q_reg_FF_FF ( .D(ctrl_seq6_SFF_3_QD), .CK(clk_gated), 
        .Q(n126), .QN() );
  DFF_X1 ctrl_seq6_SFF_1_Q_reg_FF_FF ( .D(ctrl_seq6_SFF_1_QD), .CK(clk_gated), 
        .Q(n125), .QN() );
  DFF_X1 ctrl_seq6_SFF_4_Q_reg_FF_FF ( .D(ctrl_seq6_SFF_4_QD), .CK(clk_gated), 
        .Q(), .QN(n155) );
  DFF_X1 ctrl_seq6_SFF_2_Q_reg_FF_FF ( .D(ctrl_seq6_SFF_2_QD), .CK(clk_gated), 
        .Q(n133), .QN() );
  DFF_X1 ctrl_seq6_SFF_0_Q_reg_FF_FF ( .D(ctrl_seq6_SFF_0_QD), .CK(clk_gated), 
        .Q(), .QN(n148) );
  DFF_X1 ctrl_seq4_SFF_0_Q_reg_FF_FF ( .D(ctrl_seq4_SFF_0_QD), .CK(clk_gated), 
        .Q(n139), .QN(n154) );
  DFF_X1 ctrl_seq4_SFF_1_Q_reg_FF_FF ( .D(ctrl_seq4_SFF_1_QD), .CK(clk_gated), 
        .Q(n3), .QN() );
  DFF_X1 ctrl_CSenRC_reg_FF_FF ( .D(n193), .CK(clk_gated), .Q(), .QN(n143) );
  DFF_X1 calcRCon_s_current_state_reg_7__FF_FF ( .D(calcRCon_n44), .CK(
        clk_gated), .Q(n129), .QN(n146) );
  DFF_X1 calcRCon_s_current_state_reg_2__FF_FF ( .D(calcRCon_n49), .CK(
        clk_gated), .Q(n137), .QN(n144) );
  DFF_X1 calcRCon_s_current_state_reg_0__FF_FF ( .D(calcRCon_n51), .CK(
        clk_gated), .Q(n128), .QN(n147) );
  DFF_X1 calcRCon_s_current_state_reg_3__FF_FF ( .D(calcRCon_n48), .CK(
        clk_gated), .Q(n131), .QN(n153) );
  DFF_X1 calcRCon_s_current_state_reg_4__FF_FF ( .D(calcRCon_n47), .CK(
        clk_gated), .Q(n135), .QN(n151) );
  DFF_X1 calcRCon_s_current_state_reg_1__FF_FF ( .D(calcRCon_n50), .CK(
        clk_gated), .Q(n138), .QN(n152) );
  DFF_X1 calcRCon_s_current_state_reg_6__FF_FF ( .D(calcRCon_n45), .CK(
        clk_gated), .Q(n130), .QN(n150) );
  DFF_X1 calcRCon_s_current_state_reg_5__FF_FF ( .D(calcRCon_n46), .CK(
        clk_gated), .Q(n136), .QN(n145) );
  BUF_X1 U111 ( .A(n36), .Z(n199) );
  BUF_X1 U112 ( .A(n36), .Z(n193) );
  BUF_X1 U113 ( .A(n36), .Z(n195) );
  BUF_X1 U114 ( .A(n36), .Z(n196) );
  BUF_X1 U115 ( .A(n36), .Z(n192) );
  BUF_X1 U116 ( .A(n204), .Z(n203) );
  BUF_X1 U117 ( .A(n36), .Z(n201) );
  BUF_X1 U118 ( .A(n36), .Z(n200) );
  BUF_X1 U119 ( .A(n204), .Z(n202) );
  BUF_X1 U120 ( .A(n36), .Z(n204) );
  NOR2_X1 U121 ( .A1(n231), .A2(n232), .ZN(n36) );
  INV_X1 U122 ( .A(n142), .ZN(n173) );
  INV_X1 U123 ( .A(n142), .ZN(n174) );
  OR2_X1 U124 ( .A1(n124), .A2(n231), .ZN(n142) );
  BUF_X1 U125 ( .A(n196), .Z(n194) );
  INV_X1 U126 ( .A(n201), .ZN(n188) );
  INV_X1 U127 ( .A(n201), .ZN(n181) );
  INV_X1 U128 ( .A(n196), .ZN(n178) );
  INV_X1 U129 ( .A(n199), .ZN(n179) );
  INV_X1 U130 ( .A(n193), .ZN(n182) );
  INV_X1 U131 ( .A(n193), .ZN(n187) );
  INV_X1 U132 ( .A(n142), .ZN(n165) );
  INV_X1 U133 ( .A(n142), .ZN(n167) );
  INV_X1 U134 ( .A(n142), .ZN(n171) );
  INV_X1 U135 ( .A(n193), .ZN(n186) );
  INV_X1 U136 ( .A(n199), .ZN(n183) );
  INV_X1 U137 ( .A(n199), .ZN(n177) );
  INV_X1 U138 ( .A(n196), .ZN(n185) );
  INV_X1 U139 ( .A(n142), .ZN(n176) );
  INV_X1 U140 ( .A(n142), .ZN(n166) );
  INV_X1 U141 ( .A(n195), .ZN(n184) );
  INV_X1 U142 ( .A(n142), .ZN(n164) );
  INV_X1 U143 ( .A(n195), .ZN(n180) );
  INV_X1 U144 ( .A(n142), .ZN(n170) );
  INV_X1 U145 ( .A(n142), .ZN(n168) );
  INV_X1 U146 ( .A(n142), .ZN(n172) );
  INV_X1 U147 ( .A(n142), .ZN(n169) );
  BUF_X1 U148 ( .A(n193), .Z(n191) );
  BUF_X1 U149 ( .A(n195), .Z(n197) );
  INV_X1 U150 ( .A(n142), .ZN(n162) );
  BUF_X1 U151 ( .A(n141), .Z(n158) );
  INV_X1 U152 ( .A(n198), .ZN(n190) );
  INV_X1 U153 ( .A(n142), .ZN(n161) );
  INV_X1 U154 ( .A(n201), .ZN(n189) );
  INV_X1 U155 ( .A(n142), .ZN(n160) );
  INV_X1 U156 ( .A(n142), .ZN(n163) );
  INV_X1 U157 ( .A(n142), .ZN(n175) );
  BUF_X1 U158 ( .A(n141), .Z(n157) );
  BUF_X1 U159 ( .A(n141), .Z(n156) );
  BUF_X1 U160 ( .A(n141), .Z(n159) );
  INV_X1 U161 ( .A(n241), .ZN(n141) );
  OR4_X1 U162 ( .A1(n125), .A2(n133), .A3(n126), .A4(n240), .ZN(n232) );
  INV_X1 U163 ( .A(nReset), .ZN(n231) );
  INV_X1 U164 ( .A(n149), .ZN(n225) );
  INV_X1 U165 ( .A(n149), .ZN(n224) );
  INV_X1 U166 ( .A(n149), .ZN(n229) );
  INV_X1 U167 ( .A(n149), .ZN(n223) );
  INV_X1 U168 ( .A(n149), .ZN(n226) );
  INV_X1 U169 ( .A(n149), .ZN(n222) );
  INV_X1 U170 ( .A(n149), .ZN(n221) );
  INV_X1 U171 ( .A(n149), .ZN(n220) );
  INV_X1 U172 ( .A(n149), .ZN(n219) );
  INV_X1 U173 ( .A(n149), .ZN(n227) );
  AOI211_X4 U174 ( .C1(n244), .C2(n243), .A(n242), .B(n231), .ZN(intselXOR) );
  INV_X1 U175 ( .A(n149), .ZN(n230) );
  NAND2_X1 U176 ( .A1(n148), .A2(n155), .ZN(n240) );
  INV_X1 U177 ( .A(n149), .ZN(n228) );
  BUF_X1 U178 ( .A(n36), .Z(n198) );
  INV_X1 U179 ( .A(n231), .ZN(n205) );
  INV_X1 U180 ( .A(n149), .ZN(n206) );
  INV_X1 U181 ( .A(n149), .ZN(n207) );
  INV_X1 U182 ( .A(n149), .ZN(n208) );
  INV_X1 U183 ( .A(n149), .ZN(n209) );
  INV_X1 U184 ( .A(n149), .ZN(n210) );
  INV_X1 U185 ( .A(n149), .ZN(n211) );
  INV_X1 U186 ( .A(n149), .ZN(n212) );
  INV_X1 U187 ( .A(n149), .ZN(n213) );
  INV_X1 U188 ( .A(n149), .ZN(n214) );
  INV_X1 U189 ( .A(n231), .ZN(n215) );
  INV_X1 U190 ( .A(n231), .ZN(n216) );
  INV_X1 U191 ( .A(n231), .ZN(n217) );
  INV_X1 U192 ( .A(n231), .ZN(n218) );
  OAI221_X1 U193 ( .B1(n192), .B2(n146), .C1(n190), .C2(n150), .A(n225), .ZN(
        calcRCon_n44) );
  NAND2_X1 U194 ( .A1(n214), .A2(n232), .ZN(n239) );
  OAI22_X1 U195 ( .A1(n190), .A2(n145), .B1(n239), .B2(n150), .ZN(calcRCon_n45) );
  OAI22_X1 U196 ( .A1(n190), .A2(n151), .B1(n239), .B2(n145), .ZN(calcRCon_n46) );
  NAND2_X1 U197 ( .A1(n129), .A2(n199), .ZN(n237) );
  NOR2_X1 U198 ( .A1(n129), .A2(n190), .ZN(n235) );
  INV_X1 U199 ( .A(n239), .ZN(n238) );
  AOI22_X1 U200 ( .A1(n131), .A2(n235), .B1(n135), .B2(n238), .ZN(n233) );
  OAI21_X1 U201 ( .B1(n131), .B2(n237), .A(n233), .ZN(calcRCon_n47) );
  AOI22_X1 U202 ( .A1(n131), .A2(n190), .B1(n235), .B2(n137), .ZN(n234) );
  OAI211_X1 U203 ( .C1(n137), .C2(n237), .A(n224), .B(n234), .ZN(calcRCon_n48)
         );
  OAI221_X1 U204 ( .B1(n195), .B2(n144), .C1(n190), .C2(n152), .A(n227), .ZN(
        calcRCon_n49) );
  AOI22_X1 U205 ( .A1(n235), .A2(n128), .B1(n238), .B2(n138), .ZN(n236) );
  OAI21_X1 U206 ( .B1(n128), .B2(n237), .A(n236), .ZN(calcRCon_n50) );
  OAI211_X1 U207 ( .C1(n199), .C2(n147), .A(n230), .B(n237), .ZN(calcRCon_n51)
         );
  NOR2_X1 U208 ( .A1(n3), .A2(n139), .ZN(n242) );
  OAI21_X1 U209 ( .B1(n242), .B2(n142), .A(n190), .ZN(ctrl_N14) );
  NAND2_X1 U210 ( .A1(n238), .A2(n3), .ZN(ctrl_seq4_SFF_0_QD) );
  NOR2_X1 U211 ( .A1(n239), .A2(n154), .ZN(ctrl_seq4_SFF_1_QD) );
  OAI211_X1 U212 ( .C1(n148), .C2(n155), .A(n226), .B(n240), .ZN(
        ctrl_seq6_SFF_0_QD) );
  NOR2_X1 U213 ( .A1(n231), .A2(n148), .ZN(ctrl_seq6_SFF_1_QD) );
  OR2_X1 U214 ( .A1(n125), .A2(n231), .ZN(ctrl_seq6_SFF_2_QD) );
  AND2_X1 U215 ( .A1(n229), .A2(n133), .ZN(ctrl_seq6_SFF_3_QD) );
  OR2_X1 U216 ( .A1(n126), .A2(n231), .ZN(ctrl_seq6_SFF_4_QD) );
  NAND4_X1 U217 ( .A1(n135), .A2(n137), .A3(n138), .A4(n136), .ZN(n241) );
  NOR4_X1 U218 ( .A1(n3), .A2(n190), .A3(n154), .A4(n241), .ZN(done) );
  NOR4_X1 U219 ( .A1(n138), .A2(n144), .A3(n153), .A4(n147), .ZN(n244) );
  NOR4_X1 U220 ( .A1(n130), .A2(n135), .A3(n136), .A4(n146), .ZN(n243) );
  NOR2_X1 U221 ( .A1(n147), .A2(n143), .ZN(roundConstant[0]) );
  NOR2_X1 U222 ( .A1(n152), .A2(n143), .ZN(roundConstant[1]) );
  NOR2_X1 U223 ( .A1(n144), .A2(n143), .ZN(roundConstant[2]) );
  NOR2_X1 U224 ( .A1(n153), .A2(n143), .ZN(roundConstant[3]) );
  NOR2_X1 U225 ( .A1(n151), .A2(n143), .ZN(roundConstant[4]) );
  NOR2_X1 U226 ( .A1(n145), .A2(n143), .ZN(roundConstant[5]) );
  NOR2_X1 U227 ( .A1(n150), .A2(n143), .ZN(roundConstant[6]) );
  NOR2_X1 U228 ( .A1(n146), .A2(n143), .ZN(roundConstant[7]) );
  INV_X1 U229 ( .A(start), .ZN(n114) );
  XOR2_X1 U29_Ins_0_U1 ( .A(ciphertext_s0[120]), .B(keyStateIn[0]), .Z(
        StateOutXORroundKey[0]) );
  XOR2_X1 U29_Ins_1_U1 ( .A(ciphertext_s1[120]), .B(new_AGEMA_signal_1983), 
        .Z(new_AGEMA_signal_1984) );
  XOR2_X1 U30_Ins_0_U1 ( .A(ciphertext_s0[121]), .B(keyStateIn[1]), .Z(
        StateOutXORroundKey[1]) );
  XOR2_X1 U30_Ins_1_U1 ( .A(ciphertext_s1[121]), .B(new_AGEMA_signal_1986), 
        .Z(new_AGEMA_signal_1987) );
  XOR2_X1 U31_Ins_0_U1 ( .A(ciphertext_s0[122]), .B(keyStateIn[2]), .Z(
        StateOutXORroundKey[2]) );
  XOR2_X1 U31_Ins_1_U1 ( .A(ciphertext_s1[122]), .B(new_AGEMA_signal_1989), 
        .Z(new_AGEMA_signal_1990) );
  XOR2_X1 U32_Ins_0_U1 ( .A(ciphertext_s0[123]), .B(keyStateIn[3]), .Z(
        StateOutXORroundKey[3]) );
  XOR2_X1 U32_Ins_1_U1 ( .A(ciphertext_s1[123]), .B(new_AGEMA_signal_1992), 
        .Z(new_AGEMA_signal_1993) );
  XOR2_X1 U33_Ins_0_U1 ( .A(ciphertext_s0[124]), .B(keyStateIn[4]), .Z(
        StateOutXORroundKey[4]) );
  XOR2_X1 U33_Ins_1_U1 ( .A(ciphertext_s1[124]), .B(new_AGEMA_signal_1995), 
        .Z(new_AGEMA_signal_1996) );
  XOR2_X1 U34_Ins_0_U1 ( .A(ciphertext_s0[125]), .B(keyStateIn[5]), .Z(
        StateOutXORroundKey[5]) );
  XOR2_X1 U34_Ins_1_U1 ( .A(ciphertext_s1[125]), .B(new_AGEMA_signal_1998), 
        .Z(new_AGEMA_signal_1999) );
  XOR2_X1 U35_Ins_0_U1 ( .A(ciphertext_s0[126]), .B(keyStateIn[6]), .Z(
        StateOutXORroundKey[6]) );
  XOR2_X1 U35_Ins_1_U1 ( .A(ciphertext_s1[126]), .B(new_AGEMA_signal_2001), 
        .Z(new_AGEMA_signal_2002) );
  XOR2_X1 U36_Ins_0_U1 ( .A(ciphertext_s0[127]), .B(keyStateIn[7]), .Z(
        StateOutXORroundKey[7]) );
  XOR2_X1 U36_Ins_1_U1 ( .A(ciphertext_s1[127]), .B(new_AGEMA_signal_2004), 
        .Z(new_AGEMA_signal_2005) );
  MUX2_X1 stateArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS00ser[0]), .B(ciphertext_s0[120]), .S(n191), .Z(
        stateArray_S00reg_gff_1_SFF_0_QD) );
  MUX2_X1 stateArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2156), .B(ciphertext_s1[120]), .S(n191), .Z(
        new_AGEMA_signal_3126) );
  MUX2_X1 stateArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS00ser[1]), .B(ciphertext_s0[121]), .S(n201), .Z(
        stateArray_S00reg_gff_1_SFF_1_QD) );
  MUX2_X1 stateArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2159), .B(ciphertext_s1[121]), .S(n201), .Z(
        new_AGEMA_signal_3127) );
  MUX2_X1 stateArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS00ser[2]), .B(ciphertext_s0[122]), .S(n193), .Z(
        stateArray_S00reg_gff_1_SFF_2_QD) );
  MUX2_X1 stateArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2162), .B(ciphertext_s1[122]), .S(n193), .Z(
        new_AGEMA_signal_3128) );
  MUX2_X1 stateArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS00ser[3]), .B(ciphertext_s0[123]), .S(n192), .Z(
        stateArray_S00reg_gff_1_SFF_3_QD) );
  MUX2_X1 stateArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2165), .B(ciphertext_s1[123]), .S(n192), .Z(
        new_AGEMA_signal_3129) );
  MUX2_X1 stateArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS00ser[4]), .B(ciphertext_s0[124]), .S(n196), .Z(
        stateArray_S00reg_gff_1_SFF_4_QD) );
  MUX2_X1 stateArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2168), .B(ciphertext_s1[124]), .S(n196), .Z(
        new_AGEMA_signal_3130) );
  MUX2_X1 stateArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS00ser[5]), .B(ciphertext_s0[125]), .S(n199), .Z(
        stateArray_S00reg_gff_1_SFF_5_QD) );
  MUX2_X1 stateArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2171), .B(ciphertext_s1[125]), .S(n199), .Z(
        new_AGEMA_signal_3131) );
  MUX2_X1 stateArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS00ser[6]), .B(ciphertext_s0[126]), .S(n200), .Z(
        stateArray_S00reg_gff_1_SFF_6_QD) );
  MUX2_X1 stateArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2174), .B(ciphertext_s1[126]), .S(n200), .Z(
        new_AGEMA_signal_3132) );
  MUX2_X1 stateArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS00ser[7]), .B(ciphertext_s0[127]), .S(n195), .Z(
        stateArray_S00reg_gff_1_SFF_7_QD) );
  MUX2_X1 stateArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2177), .B(ciphertext_s1[127]), .S(n195), .Z(
        new_AGEMA_signal_3133) );
  MUX2_X1 stateArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS01ser[0]), .B(ciphertext_s0[112]), .S(n199), .Z(
        stateArray_S01reg_gff_1_SFF_0_QD) );
  MUX2_X1 stateArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2180), .B(ciphertext_s1[112]), .S(n199), .Z(
        new_AGEMA_signal_3134) );
  MUX2_X1 stateArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS01ser[1]), .B(ciphertext_s0[113]), .S(n195), .Z(
        stateArray_S01reg_gff_1_SFF_1_QD) );
  MUX2_X1 stateArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2183), .B(ciphertext_s1[113]), .S(n195), .Z(
        new_AGEMA_signal_3135) );
  MUX2_X1 stateArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS01ser[2]), .B(ciphertext_s0[114]), .S(n192), .Z(
        stateArray_S01reg_gff_1_SFF_2_QD) );
  MUX2_X1 stateArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2186), .B(ciphertext_s1[114]), .S(n192), .Z(
        new_AGEMA_signal_3136) );
  MUX2_X1 stateArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS01ser[3]), .B(ciphertext_s0[115]), .S(n195), .Z(
        stateArray_S01reg_gff_1_SFF_3_QD) );
  MUX2_X1 stateArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2189), .B(ciphertext_s1[115]), .S(n195), .Z(
        new_AGEMA_signal_3137) );
  MUX2_X1 stateArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS01ser[4]), .B(ciphertext_s0[116]), .S(n200), .Z(
        stateArray_S01reg_gff_1_SFF_4_QD) );
  MUX2_X1 stateArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2192), .B(ciphertext_s1[116]), .S(n200), .Z(
        new_AGEMA_signal_3138) );
  MUX2_X1 stateArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS01ser[5]), .B(ciphertext_s0[117]), .S(n201), .Z(
        stateArray_S01reg_gff_1_SFF_5_QD) );
  MUX2_X1 stateArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2195), .B(ciphertext_s1[117]), .S(n201), .Z(
        new_AGEMA_signal_3139) );
  MUX2_X1 stateArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS01ser[6]), .B(ciphertext_s0[118]), .S(n193), .Z(
        stateArray_S01reg_gff_1_SFF_6_QD) );
  MUX2_X1 stateArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2198), .B(ciphertext_s1[118]), .S(n193), .Z(
        new_AGEMA_signal_3140) );
  MUX2_X1 stateArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS01ser[7]), .B(ciphertext_s0[119]), .S(n196), .Z(
        stateArray_S01reg_gff_1_SFF_7_QD) );
  MUX2_X1 stateArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2201), .B(ciphertext_s1[119]), .S(n196), .Z(
        new_AGEMA_signal_3141) );
  MUX2_X1 stateArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS02ser[0]), .B(ciphertext_s0[104]), .S(n192), .Z(
        stateArray_S02reg_gff_1_SFF_0_QD) );
  MUX2_X1 stateArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2204), .B(ciphertext_s1[104]), .S(n192), .Z(
        new_AGEMA_signal_3142) );
  MUX2_X1 stateArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS02ser[1]), .B(ciphertext_s0[105]), .S(n195), .Z(
        stateArray_S02reg_gff_1_SFF_1_QD) );
  MUX2_X1 stateArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2207), .B(ciphertext_s1[105]), .S(n195), .Z(
        new_AGEMA_signal_3143) );
  MUX2_X1 stateArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS02ser[2]), .B(ciphertext_s0[106]), .S(n200), .Z(
        stateArray_S02reg_gff_1_SFF_2_QD) );
  MUX2_X1 stateArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2210), .B(ciphertext_s1[106]), .S(n200), .Z(
        new_AGEMA_signal_3144) );
  MUX2_X1 stateArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS02ser[3]), .B(ciphertext_s0[107]), .S(n196), .Z(
        stateArray_S02reg_gff_1_SFF_3_QD) );
  MUX2_X1 stateArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2213), .B(ciphertext_s1[107]), .S(n196), .Z(
        new_AGEMA_signal_3145) );
  MUX2_X1 stateArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS02ser[4]), .B(ciphertext_s0[108]), .S(n199), .Z(
        stateArray_S02reg_gff_1_SFF_4_QD) );
  MUX2_X1 stateArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2216), .B(ciphertext_s1[108]), .S(n199), .Z(
        new_AGEMA_signal_3146) );
  MUX2_X1 stateArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS02ser[5]), .B(ciphertext_s0[109]), .S(n192), .Z(
        stateArray_S02reg_gff_1_SFF_5_QD) );
  MUX2_X1 stateArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2219), .B(ciphertext_s1[109]), .S(n192), .Z(
        new_AGEMA_signal_3147) );
  MUX2_X1 stateArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS02ser[6]), .B(ciphertext_s0[110]), .S(n193), .Z(
        stateArray_S02reg_gff_1_SFF_6_QD) );
  MUX2_X1 stateArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2222), .B(ciphertext_s1[110]), .S(n193), .Z(
        new_AGEMA_signal_3148) );
  MUX2_X1 stateArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS02ser[7]), .B(ciphertext_s0[111]), .S(n201), .Z(
        stateArray_S02reg_gff_1_SFF_7_QD) );
  MUX2_X1 stateArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2225), .B(ciphertext_s1[111]), .S(n201), .Z(
        new_AGEMA_signal_3149) );
  MUX2_X1 stateArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS03ser[0]), .B(ciphertext_s0[96]), .S(n196), .Z(
        stateArray_S03reg_gff_1_SFF_0_QD) );
  MUX2_X1 stateArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3046), .B(ciphertext_s1[96]), .S(n196), .Z(
        new_AGEMA_signal_3150) );
  MUX2_X1 stateArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS03ser[1]), .B(ciphertext_s0[97]), .S(n203), .Z(
        stateArray_S03reg_gff_1_SFF_1_QD) );
  MUX2_X1 stateArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3048), .B(ciphertext_s1[97]), .S(n203), .Z(
        new_AGEMA_signal_3151) );
  MUX2_X1 stateArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS03ser[2]), .B(ciphertext_s0[98]), .S(n202), .Z(
        stateArray_S03reg_gff_1_SFF_2_QD) );
  MUX2_X1 stateArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3050), .B(ciphertext_s1[98]), .S(n202), .Z(
        new_AGEMA_signal_3152) );
  MUX2_X1 stateArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS03ser[3]), .B(ciphertext_s0[99]), .S(n203), .Z(
        stateArray_S03reg_gff_1_SFF_3_QD) );
  MUX2_X1 stateArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3052), .B(ciphertext_s1[99]), .S(n203), .Z(
        new_AGEMA_signal_3153) );
  MUX2_X1 stateArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS03ser[4]), .B(ciphertext_s0[100]), .S(n204), .Z(
        stateArray_S03reg_gff_1_SFF_4_QD) );
  MUX2_X1 stateArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3054), .B(ciphertext_s1[100]), .S(n204), .Z(
        new_AGEMA_signal_3154) );
  MUX2_X1 stateArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS03ser[5]), .B(ciphertext_s0[101]), .S(n203), .Z(
        stateArray_S03reg_gff_1_SFF_5_QD) );
  MUX2_X1 stateArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3056), .B(ciphertext_s1[101]), .S(n203), .Z(
        new_AGEMA_signal_3155) );
  MUX2_X1 stateArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS03ser[6]), .B(ciphertext_s0[102]), .S(n204), .Z(
        stateArray_S03reg_gff_1_SFF_6_QD) );
  MUX2_X1 stateArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3058), .B(ciphertext_s1[102]), .S(n204), .Z(
        new_AGEMA_signal_3156) );
  MUX2_X1 stateArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS03ser[7]), .B(ciphertext_s0[103]), .S(n198), .Z(
        stateArray_S03reg_gff_1_SFF_7_QD) );
  MUX2_X1 stateArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3060), .B(ciphertext_s1[103]), .S(n198), .Z(
        new_AGEMA_signal_3157) );
  MUX2_X1 stateArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS10ser[0]), .B(ciphertext_s0[80]), .S(n204), .Z(
        stateArray_S10reg_gff_1_SFF_0_QD) );
  MUX2_X1 stateArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2228), .B(ciphertext_s1[80]), .S(n204), .Z(
        new_AGEMA_signal_3158) );
  MUX2_X1 stateArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS10ser[1]), .B(ciphertext_s0[81]), .S(n203), .Z(
        stateArray_S10reg_gff_1_SFF_1_QD) );
  MUX2_X1 stateArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2231), .B(ciphertext_s1[81]), .S(n203), .Z(
        new_AGEMA_signal_3159) );
  MUX2_X1 stateArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS10ser[2]), .B(ciphertext_s0[82]), .S(n204), .Z(
        stateArray_S10reg_gff_1_SFF_2_QD) );
  MUX2_X1 stateArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2234), .B(ciphertext_s1[82]), .S(n204), .Z(
        new_AGEMA_signal_3160) );
  MUX2_X1 stateArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS10ser[3]), .B(ciphertext_s0[83]), .S(n194), .Z(
        stateArray_S10reg_gff_1_SFF_3_QD) );
  MUX2_X1 stateArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2237), .B(ciphertext_s1[83]), .S(n194), .Z(
        new_AGEMA_signal_3161) );
  MUX2_X1 stateArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS10ser[4]), .B(ciphertext_s0[84]), .S(n193), .Z(
        stateArray_S10reg_gff_1_SFF_4_QD) );
  MUX2_X1 stateArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2240), .B(ciphertext_s1[84]), .S(n193), .Z(
        new_AGEMA_signal_3162) );
  MUX2_X1 stateArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS10ser[5]), .B(ciphertext_s0[85]), .S(n203), .Z(
        stateArray_S10reg_gff_1_SFF_5_QD) );
  MUX2_X1 stateArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2243), .B(ciphertext_s1[85]), .S(n203), .Z(
        new_AGEMA_signal_3163) );
  MUX2_X1 stateArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS10ser[6]), .B(ciphertext_s0[86]), .S(n198), .Z(
        stateArray_S10reg_gff_1_SFF_6_QD) );
  MUX2_X1 stateArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2246), .B(ciphertext_s1[86]), .S(n198), .Z(
        new_AGEMA_signal_3164) );
  MUX2_X1 stateArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS10ser[7]), .B(ciphertext_s0[87]), .S(n198), .Z(
        stateArray_S10reg_gff_1_SFF_7_QD) );
  MUX2_X1 stateArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2249), .B(ciphertext_s1[87]), .S(n198), .Z(
        new_AGEMA_signal_3165) );
  MUX2_X1 stateArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS11ser[0]), .B(ciphertext_s0[72]), .S(n203), .Z(
        stateArray_S11reg_gff_1_SFF_0_QD) );
  MUX2_X1 stateArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2252), .B(ciphertext_s1[72]), .S(n203), .Z(
        new_AGEMA_signal_3166) );
  MUX2_X1 stateArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS11ser[1]), .B(ciphertext_s0[73]), .S(n203), .Z(
        stateArray_S11reg_gff_1_SFF_1_QD) );
  MUX2_X1 stateArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2255), .B(ciphertext_s1[73]), .S(n203), .Z(
        new_AGEMA_signal_3167) );
  MUX2_X1 stateArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS11ser[2]), .B(ciphertext_s0[74]), .S(n204), .Z(
        stateArray_S11reg_gff_1_SFF_2_QD) );
  MUX2_X1 stateArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2258), .B(ciphertext_s1[74]), .S(n204), .Z(
        new_AGEMA_signal_3168) );
  MUX2_X1 stateArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS11ser[3]), .B(ciphertext_s0[75]), .S(n204), .Z(
        stateArray_S11reg_gff_1_SFF_3_QD) );
  MUX2_X1 stateArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2261), .B(ciphertext_s1[75]), .S(n204), .Z(
        new_AGEMA_signal_3169) );
  MUX2_X1 stateArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS11ser[4]), .B(ciphertext_s0[76]), .S(n195), .Z(
        stateArray_S11reg_gff_1_SFF_4_QD) );
  MUX2_X1 stateArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2264), .B(ciphertext_s1[76]), .S(n195), .Z(
        new_AGEMA_signal_3170) );
  MUX2_X1 stateArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS11ser[5]), .B(ciphertext_s0[77]), .S(n202), .Z(
        stateArray_S11reg_gff_1_SFF_5_QD) );
  MUX2_X1 stateArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2267), .B(ciphertext_s1[77]), .S(n202), .Z(
        new_AGEMA_signal_3171) );
  MUX2_X1 stateArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS11ser[6]), .B(ciphertext_s0[78]), .S(n204), .Z(
        stateArray_S11reg_gff_1_SFF_6_QD) );
  MUX2_X1 stateArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2270), .B(ciphertext_s1[78]), .S(n204), .Z(
        new_AGEMA_signal_3172) );
  MUX2_X1 stateArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS11ser[7]), .B(ciphertext_s0[79]), .S(n202), .Z(
        stateArray_S11reg_gff_1_SFF_7_QD) );
  MUX2_X1 stateArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2273), .B(ciphertext_s1[79]), .S(n202), .Z(
        new_AGEMA_signal_3173) );
  MUX2_X1 stateArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS12ser[0]), .B(ciphertext_s0[64]), .S(n204), .Z(
        stateArray_S12reg_gff_1_SFF_0_QD) );
  MUX2_X1 stateArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2276), .B(ciphertext_s1[64]), .S(n204), .Z(
        new_AGEMA_signal_3174) );
  MUX2_X1 stateArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS12ser[1]), .B(ciphertext_s0[65]), .S(n204), .Z(
        stateArray_S12reg_gff_1_SFF_1_QD) );
  MUX2_X1 stateArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2279), .B(ciphertext_s1[65]), .S(n204), .Z(
        new_AGEMA_signal_3175) );
  MUX2_X1 stateArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS12ser[2]), .B(ciphertext_s0[66]), .S(n202), .Z(
        stateArray_S12reg_gff_1_SFF_2_QD) );
  MUX2_X1 stateArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2282), .B(ciphertext_s1[66]), .S(n202), .Z(
        new_AGEMA_signal_3176) );
  MUX2_X1 stateArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS12ser[3]), .B(ciphertext_s0[67]), .S(n203), .Z(
        stateArray_S12reg_gff_1_SFF_3_QD) );
  MUX2_X1 stateArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2285), .B(ciphertext_s1[67]), .S(n203), .Z(
        new_AGEMA_signal_3177) );
  MUX2_X1 stateArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS12ser[4]), .B(ciphertext_s0[68]), .S(n203), .Z(
        stateArray_S12reg_gff_1_SFF_4_QD) );
  MUX2_X1 stateArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2288), .B(ciphertext_s1[68]), .S(n203), .Z(
        new_AGEMA_signal_3178) );
  MUX2_X1 stateArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS12ser[5]), .B(ciphertext_s0[69]), .S(n203), .Z(
        stateArray_S12reg_gff_1_SFF_5_QD) );
  MUX2_X1 stateArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2291), .B(ciphertext_s1[69]), .S(n203), .Z(
        new_AGEMA_signal_3179) );
  MUX2_X1 stateArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS12ser[6]), .B(ciphertext_s0[70]), .S(n194), .Z(
        stateArray_S12reg_gff_1_SFF_6_QD) );
  MUX2_X1 stateArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2294), .B(ciphertext_s1[70]), .S(n194), .Z(
        new_AGEMA_signal_3180) );
  MUX2_X1 stateArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS12ser[7]), .B(ciphertext_s0[71]), .S(n202), .Z(
        stateArray_S12reg_gff_1_SFF_7_QD) );
  MUX2_X1 stateArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2297), .B(ciphertext_s1[71]), .S(n202), .Z(
        new_AGEMA_signal_3181) );
  MUX2_X1 stateArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS13ser[0]), .B(ciphertext_s0[88]), .S(n202), .Z(
        stateArray_S13reg_gff_1_SFF_0_QD) );
  MUX2_X1 stateArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3062), .B(ciphertext_s1[88]), .S(n202), .Z(
        new_AGEMA_signal_3182) );
  MUX2_X1 stateArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS13ser[1]), .B(ciphertext_s0[89]), .S(n202), .Z(
        stateArray_S13reg_gff_1_SFF_1_QD) );
  MUX2_X1 stateArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3064), .B(ciphertext_s1[89]), .S(n202), .Z(
        new_AGEMA_signal_3183) );
  MUX2_X1 stateArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS13ser[2]), .B(ciphertext_s0[90]), .S(n202), .Z(
        stateArray_S13reg_gff_1_SFF_2_QD) );
  MUX2_X1 stateArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3066), .B(ciphertext_s1[90]), .S(n202), .Z(
        new_AGEMA_signal_3184) );
  MUX2_X1 stateArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS13ser[3]), .B(ciphertext_s0[91]), .S(n197), .Z(
        stateArray_S13reg_gff_1_SFF_3_QD) );
  MUX2_X1 stateArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3068), .B(ciphertext_s1[91]), .S(n197), .Z(
        new_AGEMA_signal_3185) );
  MUX2_X1 stateArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS13ser[4]), .B(ciphertext_s0[92]), .S(n201), .Z(
        stateArray_S13reg_gff_1_SFF_4_QD) );
  MUX2_X1 stateArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3070), .B(ciphertext_s1[92]), .S(n201), .Z(
        new_AGEMA_signal_3186) );
  MUX2_X1 stateArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS13ser[5]), .B(ciphertext_s0[93]), .S(n191), .Z(
        stateArray_S13reg_gff_1_SFF_5_QD) );
  MUX2_X1 stateArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3072), .B(ciphertext_s1[93]), .S(n191), .Z(
        new_AGEMA_signal_3187) );
  MUX2_X1 stateArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS13ser[6]), .B(ciphertext_s0[94]), .S(n197), .Z(
        stateArray_S13reg_gff_1_SFF_6_QD) );
  MUX2_X1 stateArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3074), .B(ciphertext_s1[94]), .S(n197), .Z(
        new_AGEMA_signal_3188) );
  MUX2_X1 stateArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS13ser[7]), .B(ciphertext_s0[95]), .S(n191), .Z(
        stateArray_S13reg_gff_1_SFF_7_QD) );
  MUX2_X1 stateArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3076), .B(ciphertext_s1[95]), .S(n191), .Z(
        new_AGEMA_signal_3189) );
  MUX2_X1 stateArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS20ser[0]), .B(ciphertext_s0[40]), .S(n196), .Z(
        stateArray_S20reg_gff_1_SFF_0_QD) );
  MUX2_X1 stateArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2300), .B(ciphertext_s1[40]), .S(n196), .Z(
        new_AGEMA_signal_3190) );
  MUX2_X1 stateArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS20ser[1]), .B(ciphertext_s0[41]), .S(n202), .Z(
        stateArray_S20reg_gff_1_SFF_1_QD) );
  MUX2_X1 stateArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2303), .B(ciphertext_s1[41]), .S(n202), .Z(
        new_AGEMA_signal_3191) );
  MUX2_X1 stateArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS20ser[2]), .B(ciphertext_s0[42]), .S(n201), .Z(
        stateArray_S20reg_gff_1_SFF_2_QD) );
  MUX2_X1 stateArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2306), .B(ciphertext_s1[42]), .S(n201), .Z(
        new_AGEMA_signal_3192) );
  MUX2_X1 stateArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS20ser[3]), .B(ciphertext_s0[43]), .S(n193), .Z(
        stateArray_S20reg_gff_1_SFF_3_QD) );
  MUX2_X1 stateArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2309), .B(ciphertext_s1[43]), .S(n193), .Z(
        new_AGEMA_signal_3193) );
  MUX2_X1 stateArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS20ser[4]), .B(ciphertext_s0[44]), .S(n194), .Z(
        stateArray_S20reg_gff_1_SFF_4_QD) );
  MUX2_X1 stateArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2312), .B(ciphertext_s1[44]), .S(n194), .Z(
        new_AGEMA_signal_3194) );
  MUX2_X1 stateArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS20ser[5]), .B(ciphertext_s0[45]), .S(n194), .Z(
        stateArray_S20reg_gff_1_SFF_5_QD) );
  MUX2_X1 stateArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2315), .B(ciphertext_s1[45]), .S(n194), .Z(
        new_AGEMA_signal_3195) );
  MUX2_X1 stateArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS20ser[6]), .B(ciphertext_s0[46]), .S(n194), .Z(
        stateArray_S20reg_gff_1_SFF_6_QD) );
  MUX2_X1 stateArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2318), .B(ciphertext_s1[46]), .S(n194), .Z(
        new_AGEMA_signal_3196) );
  MUX2_X1 stateArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS20ser[7]), .B(ciphertext_s0[47]), .S(n201), .Z(
        stateArray_S20reg_gff_1_SFF_7_QD) );
  MUX2_X1 stateArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2321), .B(ciphertext_s1[47]), .S(n201), .Z(
        new_AGEMA_signal_3197) );
  MUX2_X1 stateArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS21ser[0]), .B(ciphertext_s0[32]), .S(n201), .Z(
        stateArray_S21reg_gff_1_SFF_0_QD) );
  MUX2_X1 stateArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2324), .B(ciphertext_s1[32]), .S(n201), .Z(
        new_AGEMA_signal_3198) );
  MUX2_X1 stateArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS21ser[1]), .B(ciphertext_s0[33]), .S(n201), .Z(
        stateArray_S21reg_gff_1_SFF_1_QD) );
  MUX2_X1 stateArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2327), .B(ciphertext_s1[33]), .S(n201), .Z(
        new_AGEMA_signal_3199) );
  MUX2_X1 stateArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS21ser[2]), .B(ciphertext_s0[34]), .S(n200), .Z(
        stateArray_S21reg_gff_1_SFF_2_QD) );
  MUX2_X1 stateArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2330), .B(ciphertext_s1[34]), .S(n200), .Z(
        new_AGEMA_signal_3200) );
  MUX2_X1 stateArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS21ser[3]), .B(ciphertext_s0[35]), .S(n200), .Z(
        stateArray_S21reg_gff_1_SFF_3_QD) );
  MUX2_X1 stateArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2333), .B(ciphertext_s1[35]), .S(n200), .Z(
        new_AGEMA_signal_3201) );
  MUX2_X1 stateArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS21ser[4]), .B(ciphertext_s0[36]), .S(n200), .Z(
        stateArray_S21reg_gff_1_SFF_4_QD) );
  MUX2_X1 stateArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2336), .B(ciphertext_s1[36]), .S(n200), .Z(
        new_AGEMA_signal_3202) );
  MUX2_X1 stateArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS21ser[5]), .B(ciphertext_s0[37]), .S(n199), .Z(
        stateArray_S21reg_gff_1_SFF_5_QD) );
  MUX2_X1 stateArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2339), .B(ciphertext_s1[37]), .S(n199), .Z(
        new_AGEMA_signal_3203) );
  MUX2_X1 stateArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS21ser[6]), .B(ciphertext_s0[38]), .S(n199), .Z(
        stateArray_S21reg_gff_1_SFF_6_QD) );
  MUX2_X1 stateArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2342), .B(ciphertext_s1[38]), .S(n199), .Z(
        new_AGEMA_signal_3204) );
  MUX2_X1 stateArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS21ser[7]), .B(ciphertext_s0[39]), .S(n199), .Z(
        stateArray_S21reg_gff_1_SFF_7_QD) );
  MUX2_X1 stateArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2345), .B(ciphertext_s1[39]), .S(n199), .Z(
        new_AGEMA_signal_3205) );
  MUX2_X1 stateArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS22ser[0]), .B(ciphertext_s0[56]), .S(n191), .Z(
        stateArray_S22reg_gff_1_SFF_0_QD) );
  MUX2_X1 stateArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2348), .B(ciphertext_s1[56]), .S(n191), .Z(
        new_AGEMA_signal_3206) );
  MUX2_X1 stateArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS22ser[1]), .B(ciphertext_s0[57]), .S(n197), .Z(
        stateArray_S22reg_gff_1_SFF_1_QD) );
  MUX2_X1 stateArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2351), .B(ciphertext_s1[57]), .S(n197), .Z(
        new_AGEMA_signal_3207) );
  MUX2_X1 stateArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS22ser[2]), .B(ciphertext_s0[58]), .S(n191), .Z(
        stateArray_S22reg_gff_1_SFF_2_QD) );
  MUX2_X1 stateArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2354), .B(ciphertext_s1[58]), .S(n191), .Z(
        new_AGEMA_signal_3208) );
  MUX2_X1 stateArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS22ser[3]), .B(ciphertext_s0[59]), .S(n198), .Z(
        stateArray_S22reg_gff_1_SFF_3_QD) );
  MUX2_X1 stateArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2357), .B(ciphertext_s1[59]), .S(n198), .Z(
        new_AGEMA_signal_3209) );
  MUX2_X1 stateArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS22ser[4]), .B(ciphertext_s0[60]), .S(n198), .Z(
        stateArray_S22reg_gff_1_SFF_4_QD) );
  MUX2_X1 stateArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2360), .B(ciphertext_s1[60]), .S(n198), .Z(
        new_AGEMA_signal_3210) );
  MUX2_X1 stateArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS22ser[5]), .B(ciphertext_s0[61]), .S(n198), .Z(
        stateArray_S22reg_gff_1_SFF_5_QD) );
  MUX2_X1 stateArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2363), .B(ciphertext_s1[61]), .S(n198), .Z(
        new_AGEMA_signal_3211) );
  MUX2_X1 stateArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS22ser[6]), .B(ciphertext_s0[62]), .S(n197), .Z(
        stateArray_S22reg_gff_1_SFF_6_QD) );
  MUX2_X1 stateArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2366), .B(ciphertext_s1[62]), .S(n197), .Z(
        new_AGEMA_signal_3212) );
  MUX2_X1 stateArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS22ser[7]), .B(ciphertext_s0[63]), .S(n197), .Z(
        stateArray_S22reg_gff_1_SFF_7_QD) );
  MUX2_X1 stateArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2369), .B(ciphertext_s1[63]), .S(n197), .Z(
        new_AGEMA_signal_3213) );
  MUX2_X1 stateArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS23ser[0]), .B(ciphertext_s0[48]), .S(n197), .Z(
        stateArray_S23reg_gff_1_SFF_0_QD) );
  MUX2_X1 stateArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3078), .B(ciphertext_s1[48]), .S(n197), .Z(
        new_AGEMA_signal_3214) );
  MUX2_X1 stateArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS23ser[1]), .B(ciphertext_s0[49]), .S(n196), .Z(
        stateArray_S23reg_gff_1_SFF_1_QD) );
  MUX2_X1 stateArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3080), .B(ciphertext_s1[49]), .S(n196), .Z(
        new_AGEMA_signal_3215) );
  MUX2_X1 stateArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS23ser[2]), .B(ciphertext_s0[50]), .S(n196), .Z(
        stateArray_S23reg_gff_1_SFF_2_QD) );
  MUX2_X1 stateArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3082), .B(ciphertext_s1[50]), .S(n196), .Z(
        new_AGEMA_signal_3216) );
  MUX2_X1 stateArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS23ser[3]), .B(ciphertext_s0[51]), .S(n196), .Z(
        stateArray_S23reg_gff_1_SFF_3_QD) );
  MUX2_X1 stateArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3084), .B(ciphertext_s1[51]), .S(n196), .Z(
        new_AGEMA_signal_3217) );
  MUX2_X1 stateArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS23ser[4]), .B(ciphertext_s0[52]), .S(n195), .Z(
        stateArray_S23reg_gff_1_SFF_4_QD) );
  MUX2_X1 stateArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3086), .B(ciphertext_s1[52]), .S(n195), .Z(
        new_AGEMA_signal_3218) );
  MUX2_X1 stateArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS23ser[5]), .B(ciphertext_s0[53]), .S(n195), .Z(
        stateArray_S23reg_gff_1_SFF_5_QD) );
  MUX2_X1 stateArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3088), .B(ciphertext_s1[53]), .S(n195), .Z(
        new_AGEMA_signal_3219) );
  MUX2_X1 stateArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS23ser[6]), .B(ciphertext_s0[54]), .S(n195), .Z(
        stateArray_S23reg_gff_1_SFF_6_QD) );
  MUX2_X1 stateArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3090), .B(ciphertext_s1[54]), .S(n195), .Z(
        new_AGEMA_signal_3220) );
  MUX2_X1 stateArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS23ser[7]), .B(ciphertext_s0[55]), .S(n198), .Z(
        stateArray_S23reg_gff_1_SFF_7_QD) );
  MUX2_X1 stateArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3092), .B(ciphertext_s1[55]), .S(n198), .Z(
        new_AGEMA_signal_3221) );
  MUX2_X1 stateArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS30ser[0]), .B(ciphertext_s0[0]), .S(n200), .Z(
        stateArray_S30reg_gff_1_SFF_0_QD) );
  MUX2_X1 stateArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2372), .B(ciphertext_s1[0]), .S(n200), .Z(
        new_AGEMA_signal_3222) );
  MUX2_X1 stateArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS30ser[1]), .B(ciphertext_s0[1]), .S(n200), .Z(
        stateArray_S30reg_gff_1_SFF_1_QD) );
  MUX2_X1 stateArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2375), .B(ciphertext_s1[1]), .S(n200), .Z(
        new_AGEMA_signal_3223) );
  MUX2_X1 stateArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS30ser[2]), .B(ciphertext_s0[2]), .S(n200), .Z(
        stateArray_S30reg_gff_1_SFF_2_QD) );
  MUX2_X1 stateArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2378), .B(ciphertext_s1[2]), .S(n200), .Z(
        new_AGEMA_signal_3224) );
  MUX2_X1 stateArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS30ser[3]), .B(ciphertext_s0[3]), .S(n192), .Z(
        stateArray_S30reg_gff_1_SFF_3_QD) );
  MUX2_X1 stateArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2381), .B(ciphertext_s1[3]), .S(n192), .Z(
        new_AGEMA_signal_3225) );
  MUX2_X1 stateArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS30ser[4]), .B(ciphertext_s0[4]), .S(n197), .Z(
        stateArray_S30reg_gff_1_SFF_4_QD) );
  MUX2_X1 stateArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2384), .B(ciphertext_s1[4]), .S(n197), .Z(
        new_AGEMA_signal_3226) );
  MUX2_X1 stateArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS30ser[5]), .B(ciphertext_s0[5]), .S(n192), .Z(
        stateArray_S30reg_gff_1_SFF_5_QD) );
  MUX2_X1 stateArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2387), .B(ciphertext_s1[5]), .S(n192), .Z(
        new_AGEMA_signal_3227) );
  MUX2_X1 stateArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS30ser[6]), .B(ciphertext_s0[6]), .S(n36), .Z(
        stateArray_S30reg_gff_1_SFF_6_QD) );
  MUX2_X1 stateArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2390), .B(ciphertext_s1[6]), .S(n36), .Z(
        new_AGEMA_signal_3228) );
  MUX2_X1 stateArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS30ser[7]), .B(ciphertext_s0[7]), .S(n198), .Z(
        stateArray_S30reg_gff_1_SFF_7_QD) );
  MUX2_X1 stateArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2393), .B(ciphertext_s1[7]), .S(n198), .Z(
        new_AGEMA_signal_3229) );
  MUX2_X1 stateArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS31ser[0]), .B(ciphertext_s0[24]), .S(n36), .Z(
        stateArray_S31reg_gff_1_SFF_0_QD) );
  MUX2_X1 stateArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2396), .B(ciphertext_s1[24]), .S(n36), .Z(
        new_AGEMA_signal_3230) );
  MUX2_X1 stateArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS31ser[1]), .B(ciphertext_s0[25]), .S(n194), .Z(
        stateArray_S31reg_gff_1_SFF_1_QD) );
  MUX2_X1 stateArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2399), .B(ciphertext_s1[25]), .S(n194), .Z(
        new_AGEMA_signal_3231) );
  MUX2_X1 stateArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS31ser[2]), .B(ciphertext_s0[26]), .S(n194), .Z(
        stateArray_S31reg_gff_1_SFF_2_QD) );
  MUX2_X1 stateArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2402), .B(ciphertext_s1[26]), .S(n194), .Z(
        new_AGEMA_signal_3232) );
  MUX2_X1 stateArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS31ser[3]), .B(ciphertext_s0[27]), .S(n194), .Z(
        stateArray_S31reg_gff_1_SFF_3_QD) );
  MUX2_X1 stateArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2405), .B(ciphertext_s1[27]), .S(n194), .Z(
        new_AGEMA_signal_3233) );
  MUX2_X1 stateArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS31ser[4]), .B(ciphertext_s0[28]), .S(n193), .Z(
        stateArray_S31reg_gff_1_SFF_4_QD) );
  MUX2_X1 stateArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2408), .B(ciphertext_s1[28]), .S(n193), .Z(
        new_AGEMA_signal_3234) );
  MUX2_X1 stateArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS31ser[5]), .B(ciphertext_s0[29]), .S(n193), .Z(
        stateArray_S31reg_gff_1_SFF_5_QD) );
  MUX2_X1 stateArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2411), .B(ciphertext_s1[29]), .S(n193), .Z(
        new_AGEMA_signal_3235) );
  MUX2_X1 stateArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS31ser[6]), .B(ciphertext_s0[30]), .S(n193), .Z(
        stateArray_S31reg_gff_1_SFF_6_QD) );
  MUX2_X1 stateArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2414), .B(ciphertext_s1[30]), .S(n193), .Z(
        new_AGEMA_signal_3236) );
  MUX2_X1 stateArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS31ser[7]), .B(ciphertext_s0[31]), .S(n194), .Z(
        stateArray_S31reg_gff_1_SFF_7_QD) );
  MUX2_X1 stateArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2417), .B(ciphertext_s1[31]), .S(n194), .Z(
        new_AGEMA_signal_3237) );
  MUX2_X1 stateArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS32ser[0]), .B(ciphertext_s0[16]), .S(n198), .Z(
        stateArray_S32reg_gff_1_SFF_0_QD) );
  MUX2_X1 stateArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2420), .B(ciphertext_s1[16]), .S(n198), .Z(
        new_AGEMA_signal_3238) );
  MUX2_X1 stateArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS32ser[1]), .B(ciphertext_s0[17]), .S(n194), .Z(
        stateArray_S32reg_gff_1_SFF_1_QD) );
  MUX2_X1 stateArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2423), .B(ciphertext_s1[17]), .S(n194), .Z(
        new_AGEMA_signal_3239) );
  MUX2_X1 stateArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS32ser[2]), .B(ciphertext_s0[18]), .S(n191), .Z(
        stateArray_S32reg_gff_1_SFF_2_QD) );
  MUX2_X1 stateArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2426), .B(ciphertext_s1[18]), .S(n191), .Z(
        new_AGEMA_signal_3240) );
  MUX2_X1 stateArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS32ser[3]), .B(ciphertext_s0[19]), .S(n197), .Z(
        stateArray_S32reg_gff_1_SFF_3_QD) );
  MUX2_X1 stateArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2429), .B(ciphertext_s1[19]), .S(n197), .Z(
        new_AGEMA_signal_3241) );
  MUX2_X1 stateArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS32ser[4]), .B(ciphertext_s0[20]), .S(n199), .Z(
        stateArray_S32reg_gff_1_SFF_4_QD) );
  MUX2_X1 stateArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2432), .B(ciphertext_s1[20]), .S(n199), .Z(
        new_AGEMA_signal_3242) );
  MUX2_X1 stateArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS32ser[5]), .B(ciphertext_s0[21]), .S(n200), .Z(
        stateArray_S32reg_gff_1_SFF_5_QD) );
  MUX2_X1 stateArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2435), .B(ciphertext_s1[21]), .S(n200), .Z(
        new_AGEMA_signal_3243) );
  MUX2_X1 stateArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS32ser[6]), .B(ciphertext_s0[22]), .S(n202), .Z(
        stateArray_S32reg_gff_1_SFF_6_QD) );
  MUX2_X1 stateArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2438), .B(ciphertext_s1[22]), .S(n202), .Z(
        new_AGEMA_signal_3244) );
  MUX2_X1 stateArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS32ser[7]), .B(ciphertext_s0[23]), .S(n191), .Z(
        stateArray_S32reg_gff_1_SFF_7_QD) );
  MUX2_X1 stateArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2441), .B(ciphertext_s1[23]), .S(n191), .Z(
        new_AGEMA_signal_3245) );
  MUX2_X1 stateArray_MUX_inS00ser_mux_inst_0_U1_Ins_0_U1 ( .A(
        plaintext_s0[120]), .B(ciphertext_s0[112]), .S(n205), .Z(
        stateArray_inS00ser[0]) );
  MUX2_X1 stateArray_MUX_inS00ser_mux_inst_0_U1_Ins_1_U1 ( .A(
        plaintext_s1[120]), .B(ciphertext_s1[112]), .S(n205), .Z(
        new_AGEMA_signal_2156) );
  MUX2_X1 stateArray_MUX_inS00ser_mux_inst_1_U1_Ins_0_U1 ( .A(
        plaintext_s0[121]), .B(ciphertext_s0[113]), .S(n223), .Z(
        stateArray_inS00ser[1]) );
  MUX2_X1 stateArray_MUX_inS00ser_mux_inst_1_U1_Ins_1_U1 ( .A(
        plaintext_s1[121]), .B(ciphertext_s1[113]), .S(n223), .Z(
        new_AGEMA_signal_2159) );
  MUX2_X1 stateArray_MUX_inS00ser_mux_inst_2_U1_Ins_0_U1 ( .A(
        plaintext_s0[122]), .B(ciphertext_s0[114]), .S(n222), .Z(
        stateArray_inS00ser[2]) );
  MUX2_X1 stateArray_MUX_inS00ser_mux_inst_2_U1_Ins_1_U1 ( .A(
        plaintext_s1[122]), .B(ciphertext_s1[114]), .S(n222), .Z(
        new_AGEMA_signal_2162) );
  MUX2_X1 stateArray_MUX_inS00ser_mux_inst_3_U1_Ins_0_U1 ( .A(
        plaintext_s0[123]), .B(ciphertext_s0[115]), .S(n218), .Z(
        stateArray_inS00ser[3]) );
  MUX2_X1 stateArray_MUX_inS00ser_mux_inst_3_U1_Ins_1_U1 ( .A(
        plaintext_s1[123]), .B(ciphertext_s1[115]), .S(n218), .Z(
        new_AGEMA_signal_2165) );
  MUX2_X1 stateArray_MUX_inS00ser_mux_inst_4_U1_Ins_0_U1 ( .A(
        plaintext_s0[124]), .B(ciphertext_s0[116]), .S(n221), .Z(
        stateArray_inS00ser[4]) );
  MUX2_X1 stateArray_MUX_inS00ser_mux_inst_4_U1_Ins_1_U1 ( .A(
        plaintext_s1[124]), .B(ciphertext_s1[116]), .S(n221), .Z(
        new_AGEMA_signal_2168) );
  MUX2_X1 stateArray_MUX_inS00ser_mux_inst_5_U1_Ins_0_U1 ( .A(
        plaintext_s0[125]), .B(ciphertext_s0[117]), .S(n205), .Z(
        stateArray_inS00ser[5]) );
  MUX2_X1 stateArray_MUX_inS00ser_mux_inst_5_U1_Ins_1_U1 ( .A(
        plaintext_s1[125]), .B(ciphertext_s1[117]), .S(n205), .Z(
        new_AGEMA_signal_2171) );
  MUX2_X1 stateArray_MUX_inS00ser_mux_inst_6_U1_Ins_0_U1 ( .A(
        plaintext_s0[126]), .B(ciphertext_s0[118]), .S(n224), .Z(
        stateArray_inS00ser[6]) );
  MUX2_X1 stateArray_MUX_inS00ser_mux_inst_6_U1_Ins_1_U1 ( .A(
        plaintext_s1[126]), .B(ciphertext_s1[118]), .S(n224), .Z(
        new_AGEMA_signal_2174) );
  MUX2_X1 stateArray_MUX_inS00ser_mux_inst_7_U1_Ins_0_U1 ( .A(
        plaintext_s0[127]), .B(ciphertext_s0[119]), .S(n229), .Z(
        stateArray_inS00ser[7]) );
  MUX2_X1 stateArray_MUX_inS00ser_mux_inst_7_U1_Ins_1_U1 ( .A(
        plaintext_s1[127]), .B(ciphertext_s1[119]), .S(n229), .Z(
        new_AGEMA_signal_2177) );
  MUX2_X1 stateArray_MUX_inS01ser_mux_inst_0_U1_Ins_0_U1 ( .A(
        plaintext_s0[112]), .B(ciphertext_s0[104]), .S(n226), .Z(
        stateArray_inS01ser[0]) );
  MUX2_X1 stateArray_MUX_inS01ser_mux_inst_0_U1_Ins_1_U1 ( .A(
        plaintext_s1[112]), .B(ciphertext_s1[104]), .S(n226), .Z(
        new_AGEMA_signal_2180) );
  MUX2_X1 stateArray_MUX_inS01ser_mux_inst_1_U1_Ins_0_U1 ( .A(
        plaintext_s0[113]), .B(ciphertext_s0[105]), .S(n228), .Z(
        stateArray_inS01ser[1]) );
  MUX2_X1 stateArray_MUX_inS01ser_mux_inst_1_U1_Ins_1_U1 ( .A(
        plaintext_s1[113]), .B(ciphertext_s1[105]), .S(n228), .Z(
        new_AGEMA_signal_2183) );
  MUX2_X1 stateArray_MUX_inS01ser_mux_inst_2_U1_Ins_0_U1 ( .A(
        plaintext_s0[114]), .B(ciphertext_s0[106]), .S(n223), .Z(
        stateArray_inS01ser[2]) );
  MUX2_X1 stateArray_MUX_inS01ser_mux_inst_2_U1_Ins_1_U1 ( .A(
        plaintext_s1[114]), .B(ciphertext_s1[106]), .S(n223), .Z(
        new_AGEMA_signal_2186) );
  MUX2_X1 stateArray_MUX_inS01ser_mux_inst_3_U1_Ins_0_U1 ( .A(
        plaintext_s0[115]), .B(ciphertext_s0[107]), .S(n225), .Z(
        stateArray_inS01ser[3]) );
  MUX2_X1 stateArray_MUX_inS01ser_mux_inst_3_U1_Ins_1_U1 ( .A(
        plaintext_s1[115]), .B(ciphertext_s1[107]), .S(n225), .Z(
        new_AGEMA_signal_2189) );
  MUX2_X1 stateArray_MUX_inS01ser_mux_inst_4_U1_Ins_0_U1 ( .A(
        plaintext_s0[116]), .B(ciphertext_s0[108]), .S(n230), .Z(
        stateArray_inS01ser[4]) );
  MUX2_X1 stateArray_MUX_inS01ser_mux_inst_4_U1_Ins_1_U1 ( .A(
        plaintext_s1[116]), .B(ciphertext_s1[108]), .S(n230), .Z(
        new_AGEMA_signal_2192) );
  MUX2_X1 stateArray_MUX_inS01ser_mux_inst_5_U1_Ins_0_U1 ( .A(
        plaintext_s0[117]), .B(ciphertext_s0[109]), .S(n227), .Z(
        stateArray_inS01ser[5]) );
  MUX2_X1 stateArray_MUX_inS01ser_mux_inst_5_U1_Ins_1_U1 ( .A(
        plaintext_s1[117]), .B(ciphertext_s1[109]), .S(n227), .Z(
        new_AGEMA_signal_2195) );
  MUX2_X1 stateArray_MUX_inS01ser_mux_inst_6_U1_Ins_0_U1 ( .A(
        plaintext_s0[118]), .B(ciphertext_s0[110]), .S(n229), .Z(
        stateArray_inS01ser[6]) );
  MUX2_X1 stateArray_MUX_inS01ser_mux_inst_6_U1_Ins_1_U1 ( .A(
        plaintext_s1[118]), .B(ciphertext_s1[110]), .S(n229), .Z(
        new_AGEMA_signal_2198) );
  MUX2_X1 stateArray_MUX_inS01ser_mux_inst_7_U1_Ins_0_U1 ( .A(
        plaintext_s0[119]), .B(ciphertext_s0[111]), .S(n226), .Z(
        stateArray_inS01ser[7]) );
  MUX2_X1 stateArray_MUX_inS01ser_mux_inst_7_U1_Ins_1_U1 ( .A(
        plaintext_s1[119]), .B(ciphertext_s1[111]), .S(n226), .Z(
        new_AGEMA_signal_2201) );
  MUX2_X1 stateArray_MUX_inS02ser_mux_inst_0_U1_Ins_0_U1 ( .A(
        plaintext_s0[104]), .B(ciphertext_s0[96]), .S(n228), .Z(
        stateArray_inS02ser[0]) );
  MUX2_X1 stateArray_MUX_inS02ser_mux_inst_0_U1_Ins_1_U1 ( .A(
        plaintext_s1[104]), .B(ciphertext_s1[96]), .S(n228), .Z(
        new_AGEMA_signal_2204) );
  MUX2_X1 stateArray_MUX_inS02ser_mux_inst_1_U1_Ins_0_U1 ( .A(
        plaintext_s0[105]), .B(ciphertext_s0[97]), .S(n223), .Z(
        stateArray_inS02ser[1]) );
  MUX2_X1 stateArray_MUX_inS02ser_mux_inst_1_U1_Ins_1_U1 ( .A(
        plaintext_s1[105]), .B(ciphertext_s1[97]), .S(n223), .Z(
        new_AGEMA_signal_2207) );
  MUX2_X1 stateArray_MUX_inS02ser_mux_inst_2_U1_Ins_0_U1 ( .A(
        plaintext_s0[106]), .B(ciphertext_s0[98]), .S(n224), .Z(
        stateArray_inS02ser[2]) );
  MUX2_X1 stateArray_MUX_inS02ser_mux_inst_2_U1_Ins_1_U1 ( .A(
        plaintext_s1[106]), .B(ciphertext_s1[98]), .S(n224), .Z(
        new_AGEMA_signal_2210) );
  MUX2_X1 stateArray_MUX_inS02ser_mux_inst_3_U1_Ins_0_U1 ( .A(
        plaintext_s0[107]), .B(ciphertext_s0[99]), .S(n230), .Z(
        stateArray_inS02ser[3]) );
  MUX2_X1 stateArray_MUX_inS02ser_mux_inst_3_U1_Ins_1_U1 ( .A(
        plaintext_s1[107]), .B(ciphertext_s1[99]), .S(n230), .Z(
        new_AGEMA_signal_2213) );
  MUX2_X1 stateArray_MUX_inS02ser_mux_inst_4_U1_Ins_0_U1 ( .A(
        plaintext_s0[108]), .B(ciphertext_s0[100]), .S(n208), .Z(
        stateArray_inS02ser[4]) );
  MUX2_X1 stateArray_MUX_inS02ser_mux_inst_4_U1_Ins_1_U1 ( .A(
        plaintext_s1[108]), .B(ciphertext_s1[100]), .S(n208), .Z(
        new_AGEMA_signal_2216) );
  MUX2_X1 stateArray_MUX_inS02ser_mux_inst_5_U1_Ins_0_U1 ( .A(
        plaintext_s0[109]), .B(ciphertext_s0[101]), .S(n211), .Z(
        stateArray_inS02ser[5]) );
  MUX2_X1 stateArray_MUX_inS02ser_mux_inst_5_U1_Ins_1_U1 ( .A(
        plaintext_s1[109]), .B(ciphertext_s1[101]), .S(n211), .Z(
        new_AGEMA_signal_2219) );
  MUX2_X1 stateArray_MUX_inS02ser_mux_inst_6_U1_Ins_0_U1 ( .A(
        plaintext_s0[110]), .B(ciphertext_s0[102]), .S(n210), .Z(
        stateArray_inS02ser[6]) );
  MUX2_X1 stateArray_MUX_inS02ser_mux_inst_6_U1_Ins_1_U1 ( .A(
        plaintext_s1[110]), .B(ciphertext_s1[102]), .S(n210), .Z(
        new_AGEMA_signal_2222) );
  MUX2_X1 stateArray_MUX_inS02ser_mux_inst_7_U1_Ins_0_U1 ( .A(
        plaintext_s0[111]), .B(ciphertext_s0[103]), .S(n209), .Z(
        stateArray_inS02ser[7]) );
  MUX2_X1 stateArray_MUX_inS02ser_mux_inst_7_U1_Ins_1_U1 ( .A(
        plaintext_s1[111]), .B(ciphertext_s1[103]), .S(n209), .Z(
        new_AGEMA_signal_2225) );
  MUX2_X1 stateArray_MUX_outS10_MC_mux_inst_0_U1_Ins_0_U1 ( .A(
        ciphertext_s0[88]), .B(StateInMC[24]), .S(n160), .Z(
        stateArray_outS10ser_MC[0]) );
  MUX2_X1 stateArray_MUX_outS10_MC_mux_inst_0_U1_Ins_1_U1 ( .A(
        ciphertext_s1[88]), .B(new_AGEMA_signal_2880), .S(n160), .Z(
        new_AGEMA_signal_3008) );
  MUX2_X1 stateArray_MUX_outS10_MC_mux_inst_1_U1_Ins_0_U1 ( .A(
        ciphertext_s0[89]), .B(StateInMC[25]), .S(n160), .Z(
        stateArray_outS10ser_MC[1]) );
  MUX2_X1 stateArray_MUX_outS10_MC_mux_inst_1_U1_Ins_1_U1 ( .A(
        ciphertext_s1[89]), .B(new_AGEMA_signal_2881), .S(n160), .Z(
        new_AGEMA_signal_3009) );
  MUX2_X1 stateArray_MUX_outS10_MC_mux_inst_2_U1_Ins_0_U1 ( .A(
        ciphertext_s0[90]), .B(StateInMC[26]), .S(n160), .Z(
        stateArray_outS10ser_MC[2]) );
  MUX2_X1 stateArray_MUX_outS10_MC_mux_inst_2_U1_Ins_1_U1 ( .A(
        ciphertext_s1[90]), .B(new_AGEMA_signal_2882), .S(n160), .Z(
        new_AGEMA_signal_3010) );
  MUX2_X1 stateArray_MUX_outS10_MC_mux_inst_3_U1_Ins_0_U1 ( .A(
        ciphertext_s0[91]), .B(StateInMC[27]), .S(n160), .Z(
        stateArray_outS10ser_MC[3]) );
  MUX2_X1 stateArray_MUX_outS10_MC_mux_inst_3_U1_Ins_1_U1 ( .A(
        ciphertext_s1[91]), .B(new_AGEMA_signal_2883), .S(n160), .Z(
        new_AGEMA_signal_3011) );
  MUX2_X1 stateArray_MUX_outS10_MC_mux_inst_4_U1_Ins_0_U1 ( .A(
        ciphertext_s0[92]), .B(StateInMC[28]), .S(n160), .Z(
        stateArray_outS10ser_MC[4]) );
  MUX2_X1 stateArray_MUX_outS10_MC_mux_inst_4_U1_Ins_1_U1 ( .A(
        ciphertext_s1[92]), .B(new_AGEMA_signal_2884), .S(n160), .Z(
        new_AGEMA_signal_3012) );
  MUX2_X1 stateArray_MUX_outS10_MC_mux_inst_5_U1_Ins_0_U1 ( .A(
        ciphertext_s0[93]), .B(StateInMC[29]), .S(n160), .Z(
        stateArray_outS10ser_MC[5]) );
  MUX2_X1 stateArray_MUX_outS10_MC_mux_inst_5_U1_Ins_1_U1 ( .A(
        ciphertext_s1[93]), .B(new_AGEMA_signal_2885), .S(n160), .Z(
        new_AGEMA_signal_3013) );
  MUX2_X1 stateArray_MUX_outS10_MC_mux_inst_6_U1_Ins_0_U1 ( .A(
        ciphertext_s0[94]), .B(StateInMC[30]), .S(n160), .Z(
        stateArray_outS10ser_MC[6]) );
  MUX2_X1 stateArray_MUX_outS10_MC_mux_inst_6_U1_Ins_1_U1 ( .A(
        ciphertext_s1[94]), .B(new_AGEMA_signal_2886), .S(n160), .Z(
        new_AGEMA_signal_3014) );
  MUX2_X1 stateArray_MUX_outS10_MC_mux_inst_7_U1_Ins_0_U1 ( .A(
        ciphertext_s0[95]), .B(StateInMC[31]), .S(n161), .Z(
        stateArray_outS10ser_MC[7]) );
  MUX2_X1 stateArray_MUX_outS10_MC_mux_inst_7_U1_Ins_1_U1 ( .A(
        ciphertext_s1[95]), .B(new_AGEMA_signal_2887), .S(n161), .Z(
        new_AGEMA_signal_3015) );
  MUX2_X1 stateArray_MUX_inS03ser_mux_inst_0_U1_Ins_0_U1 ( .A(plaintext_s0[96]), .B(stateArray_outS10ser_MC[0]), .S(n212), .Z(stateArray_inS03ser[0]) );
  MUX2_X1 stateArray_MUX_inS03ser_mux_inst_0_U1_Ins_1_U1 ( .A(plaintext_s1[96]), .B(new_AGEMA_signal_3008), .S(n212), .Z(new_AGEMA_signal_3046) );
  MUX2_X1 stateArray_MUX_inS03ser_mux_inst_1_U1_Ins_0_U1 ( .A(plaintext_s0[97]), .B(stateArray_outS10ser_MC[1]), .S(n206), .Z(stateArray_inS03ser[1]) );
  MUX2_X1 stateArray_MUX_inS03ser_mux_inst_1_U1_Ins_1_U1 ( .A(plaintext_s1[97]), .B(new_AGEMA_signal_3009), .S(n206), .Z(new_AGEMA_signal_3048) );
  MUX2_X1 stateArray_MUX_inS03ser_mux_inst_2_U1_Ins_0_U1 ( .A(plaintext_s0[98]), .B(stateArray_outS10ser_MC[2]), .S(n213), .Z(stateArray_inS03ser[2]) );
  MUX2_X1 stateArray_MUX_inS03ser_mux_inst_2_U1_Ins_1_U1 ( .A(plaintext_s1[98]), .B(new_AGEMA_signal_3010), .S(n213), .Z(new_AGEMA_signal_3050) );
  MUX2_X1 stateArray_MUX_inS03ser_mux_inst_3_U1_Ins_0_U1 ( .A(plaintext_s0[99]), .B(stateArray_outS10ser_MC[3]), .S(n228), .Z(stateArray_inS03ser[3]) );
  MUX2_X1 stateArray_MUX_inS03ser_mux_inst_3_U1_Ins_1_U1 ( .A(plaintext_s1[99]), .B(new_AGEMA_signal_3011), .S(n228), .Z(new_AGEMA_signal_3052) );
  MUX2_X1 stateArray_MUX_inS03ser_mux_inst_4_U1_Ins_0_U1 ( .A(
        plaintext_s0[100]), .B(stateArray_outS10ser_MC[4]), .S(n207), .Z(
        stateArray_inS03ser[4]) );
  MUX2_X1 stateArray_MUX_inS03ser_mux_inst_4_U1_Ins_1_U1 ( .A(
        plaintext_s1[100]), .B(new_AGEMA_signal_3012), .S(n207), .Z(
        new_AGEMA_signal_3054) );
  MUX2_X1 stateArray_MUX_inS03ser_mux_inst_5_U1_Ins_0_U1 ( .A(
        plaintext_s0[101]), .B(stateArray_outS10ser_MC[5]), .S(n223), .Z(
        stateArray_inS03ser[5]) );
  MUX2_X1 stateArray_MUX_inS03ser_mux_inst_5_U1_Ins_1_U1 ( .A(
        plaintext_s1[101]), .B(new_AGEMA_signal_3013), .S(n223), .Z(
        new_AGEMA_signal_3056) );
  MUX2_X1 stateArray_MUX_inS03ser_mux_inst_6_U1_Ins_0_U1 ( .A(
        plaintext_s0[102]), .B(stateArray_outS10ser_MC[6]), .S(n209), .Z(
        stateArray_inS03ser[6]) );
  MUX2_X1 stateArray_MUX_inS03ser_mux_inst_6_U1_Ins_1_U1 ( .A(
        plaintext_s1[102]), .B(new_AGEMA_signal_3014), .S(n209), .Z(
        new_AGEMA_signal_3058) );
  MUX2_X1 stateArray_MUX_inS03ser_mux_inst_7_U1_Ins_0_U1 ( .A(
        plaintext_s0[103]), .B(stateArray_outS10ser_MC[7]), .S(n227), .Z(
        stateArray_inS03ser[7]) );
  MUX2_X1 stateArray_MUX_inS03ser_mux_inst_7_U1_Ins_1_U1 ( .A(
        plaintext_s1[103]), .B(new_AGEMA_signal_3015), .S(n227), .Z(
        new_AGEMA_signal_3060) );
  MUX2_X1 stateArray_MUX_inS10ser_mux_inst_0_U1_Ins_0_U1 ( .A(plaintext_s0[88]), .B(ciphertext_s0[80]), .S(n210), .Z(stateArray_inS10ser[0]) );
  MUX2_X1 stateArray_MUX_inS10ser_mux_inst_0_U1_Ins_1_U1 ( .A(plaintext_s1[88]), .B(ciphertext_s1[80]), .S(n210), .Z(new_AGEMA_signal_2228) );
  MUX2_X1 stateArray_MUX_inS10ser_mux_inst_1_U1_Ins_0_U1 ( .A(plaintext_s0[89]), .B(ciphertext_s0[81]), .S(n225), .Z(stateArray_inS10ser[1]) );
  MUX2_X1 stateArray_MUX_inS10ser_mux_inst_1_U1_Ins_1_U1 ( .A(plaintext_s1[89]), .B(ciphertext_s1[81]), .S(n225), .Z(new_AGEMA_signal_2231) );
  MUX2_X1 stateArray_MUX_inS10ser_mux_inst_2_U1_Ins_0_U1 ( .A(plaintext_s0[90]), .B(ciphertext_s0[82]), .S(n219), .Z(stateArray_inS10ser[2]) );
  MUX2_X1 stateArray_MUX_inS10ser_mux_inst_2_U1_Ins_1_U1 ( .A(plaintext_s1[90]), .B(ciphertext_s1[82]), .S(n219), .Z(new_AGEMA_signal_2234) );
  MUX2_X1 stateArray_MUX_inS10ser_mux_inst_3_U1_Ins_0_U1 ( .A(plaintext_s0[91]), .B(ciphertext_s0[83]), .S(n219), .Z(stateArray_inS10ser[3]) );
  MUX2_X1 stateArray_MUX_inS10ser_mux_inst_3_U1_Ins_1_U1 ( .A(plaintext_s1[91]), .B(ciphertext_s1[83]), .S(n219), .Z(new_AGEMA_signal_2237) );
  MUX2_X1 stateArray_MUX_inS10ser_mux_inst_4_U1_Ins_0_U1 ( .A(plaintext_s0[92]), .B(ciphertext_s0[84]), .S(n219), .Z(stateArray_inS10ser[4]) );
  MUX2_X1 stateArray_MUX_inS10ser_mux_inst_4_U1_Ins_1_U1 ( .A(plaintext_s1[92]), .B(ciphertext_s1[84]), .S(n219), .Z(new_AGEMA_signal_2240) );
  MUX2_X1 stateArray_MUX_inS10ser_mux_inst_5_U1_Ins_0_U1 ( .A(plaintext_s0[93]), .B(ciphertext_s0[85]), .S(n219), .Z(stateArray_inS10ser[5]) );
  MUX2_X1 stateArray_MUX_inS10ser_mux_inst_5_U1_Ins_1_U1 ( .A(plaintext_s1[93]), .B(ciphertext_s1[85]), .S(n219), .Z(new_AGEMA_signal_2243) );
  MUX2_X1 stateArray_MUX_inS10ser_mux_inst_6_U1_Ins_0_U1 ( .A(plaintext_s0[94]), .B(ciphertext_s0[86]), .S(n219), .Z(stateArray_inS10ser[6]) );
  MUX2_X1 stateArray_MUX_inS10ser_mux_inst_6_U1_Ins_1_U1 ( .A(plaintext_s1[94]), .B(ciphertext_s1[86]), .S(n219), .Z(new_AGEMA_signal_2246) );
  MUX2_X1 stateArray_MUX_inS10ser_mux_inst_7_U1_Ins_0_U1 ( .A(plaintext_s0[95]), .B(ciphertext_s0[87]), .S(n219), .Z(stateArray_inS10ser[7]) );
  MUX2_X1 stateArray_MUX_inS10ser_mux_inst_7_U1_Ins_1_U1 ( .A(plaintext_s1[95]), .B(ciphertext_s1[87]), .S(n219), .Z(new_AGEMA_signal_2249) );
  MUX2_X1 stateArray_MUX_inS11ser_mux_inst_0_U1_Ins_0_U1 ( .A(plaintext_s0[80]), .B(ciphertext_s0[72]), .S(n219), .Z(stateArray_inS11ser[0]) );
  MUX2_X1 stateArray_MUX_inS11ser_mux_inst_0_U1_Ins_1_U1 ( .A(plaintext_s1[80]), .B(ciphertext_s1[72]), .S(n219), .Z(new_AGEMA_signal_2252) );
  MUX2_X1 stateArray_MUX_inS11ser_mux_inst_1_U1_Ins_0_U1 ( .A(plaintext_s0[81]), .B(ciphertext_s0[73]), .S(n220), .Z(stateArray_inS11ser[1]) );
  MUX2_X1 stateArray_MUX_inS11ser_mux_inst_1_U1_Ins_1_U1 ( .A(plaintext_s1[81]), .B(ciphertext_s1[73]), .S(n220), .Z(new_AGEMA_signal_2255) );
  MUX2_X1 stateArray_MUX_inS11ser_mux_inst_2_U1_Ins_0_U1 ( .A(plaintext_s0[82]), .B(ciphertext_s0[74]), .S(n220), .Z(stateArray_inS11ser[2]) );
  MUX2_X1 stateArray_MUX_inS11ser_mux_inst_2_U1_Ins_1_U1 ( .A(plaintext_s1[82]), .B(ciphertext_s1[74]), .S(n220), .Z(new_AGEMA_signal_2258) );
  MUX2_X1 stateArray_MUX_inS11ser_mux_inst_3_U1_Ins_0_U1 ( .A(plaintext_s0[83]), .B(ciphertext_s0[75]), .S(n220), .Z(stateArray_inS11ser[3]) );
  MUX2_X1 stateArray_MUX_inS11ser_mux_inst_3_U1_Ins_1_U1 ( .A(plaintext_s1[83]), .B(ciphertext_s1[75]), .S(n220), .Z(new_AGEMA_signal_2261) );
  MUX2_X1 stateArray_MUX_inS11ser_mux_inst_4_U1_Ins_0_U1 ( .A(plaintext_s0[84]), .B(ciphertext_s0[76]), .S(n220), .Z(stateArray_inS11ser[4]) );
  MUX2_X1 stateArray_MUX_inS11ser_mux_inst_4_U1_Ins_1_U1 ( .A(plaintext_s1[84]), .B(ciphertext_s1[76]), .S(n220), .Z(new_AGEMA_signal_2264) );
  MUX2_X1 stateArray_MUX_inS11ser_mux_inst_5_U1_Ins_0_U1 ( .A(plaintext_s0[85]), .B(ciphertext_s0[77]), .S(n220), .Z(stateArray_inS11ser[5]) );
  MUX2_X1 stateArray_MUX_inS11ser_mux_inst_5_U1_Ins_1_U1 ( .A(plaintext_s1[85]), .B(ciphertext_s1[77]), .S(n220), .Z(new_AGEMA_signal_2267) );
  MUX2_X1 stateArray_MUX_inS11ser_mux_inst_6_U1_Ins_0_U1 ( .A(plaintext_s0[86]), .B(ciphertext_s0[78]), .S(n220), .Z(stateArray_inS11ser[6]) );
  MUX2_X1 stateArray_MUX_inS11ser_mux_inst_6_U1_Ins_1_U1 ( .A(plaintext_s1[86]), .B(ciphertext_s1[78]), .S(n220), .Z(new_AGEMA_signal_2270) );
  MUX2_X1 stateArray_MUX_inS11ser_mux_inst_7_U1_Ins_0_U1 ( .A(plaintext_s0[87]), .B(ciphertext_s0[79]), .S(n220), .Z(stateArray_inS11ser[7]) );
  MUX2_X1 stateArray_MUX_inS11ser_mux_inst_7_U1_Ins_1_U1 ( .A(plaintext_s1[87]), .B(ciphertext_s1[79]), .S(n220), .Z(new_AGEMA_signal_2273) );
  MUX2_X1 stateArray_MUX_inS12ser_mux_inst_0_U1_Ins_0_U1 ( .A(plaintext_s0[72]), .B(ciphertext_s0[64]), .S(n221), .Z(stateArray_inS12ser[0]) );
  MUX2_X1 stateArray_MUX_inS12ser_mux_inst_0_U1_Ins_1_U1 ( .A(plaintext_s1[72]), .B(ciphertext_s1[64]), .S(n221), .Z(new_AGEMA_signal_2276) );
  MUX2_X1 stateArray_MUX_inS12ser_mux_inst_1_U1_Ins_0_U1 ( .A(plaintext_s0[73]), .B(ciphertext_s0[65]), .S(n221), .Z(stateArray_inS12ser[1]) );
  MUX2_X1 stateArray_MUX_inS12ser_mux_inst_1_U1_Ins_1_U1 ( .A(plaintext_s1[73]), .B(ciphertext_s1[65]), .S(n221), .Z(new_AGEMA_signal_2279) );
  MUX2_X1 stateArray_MUX_inS12ser_mux_inst_2_U1_Ins_0_U1 ( .A(plaintext_s0[74]), .B(ciphertext_s0[66]), .S(n221), .Z(stateArray_inS12ser[2]) );
  MUX2_X1 stateArray_MUX_inS12ser_mux_inst_2_U1_Ins_1_U1 ( .A(plaintext_s1[74]), .B(ciphertext_s1[66]), .S(n221), .Z(new_AGEMA_signal_2282) );
  MUX2_X1 stateArray_MUX_inS12ser_mux_inst_3_U1_Ins_0_U1 ( .A(plaintext_s0[75]), .B(ciphertext_s0[67]), .S(n221), .Z(stateArray_inS12ser[3]) );
  MUX2_X1 stateArray_MUX_inS12ser_mux_inst_3_U1_Ins_1_U1 ( .A(plaintext_s1[75]), .B(ciphertext_s1[67]), .S(n221), .Z(new_AGEMA_signal_2285) );
  MUX2_X1 stateArray_MUX_inS12ser_mux_inst_4_U1_Ins_0_U1 ( .A(plaintext_s0[76]), .B(ciphertext_s0[68]), .S(n221), .Z(stateArray_inS12ser[4]) );
  MUX2_X1 stateArray_MUX_inS12ser_mux_inst_4_U1_Ins_1_U1 ( .A(plaintext_s1[76]), .B(ciphertext_s1[68]), .S(n221), .Z(new_AGEMA_signal_2288) );
  MUX2_X1 stateArray_MUX_inS12ser_mux_inst_5_U1_Ins_0_U1 ( .A(plaintext_s0[77]), .B(ciphertext_s0[69]), .S(n221), .Z(stateArray_inS12ser[5]) );
  MUX2_X1 stateArray_MUX_inS12ser_mux_inst_5_U1_Ins_1_U1 ( .A(plaintext_s1[77]), .B(ciphertext_s1[69]), .S(n221), .Z(new_AGEMA_signal_2291) );
  MUX2_X1 stateArray_MUX_inS12ser_mux_inst_6_U1_Ins_0_U1 ( .A(plaintext_s0[78]), .B(ciphertext_s0[70]), .S(n221), .Z(stateArray_inS12ser[6]) );
  MUX2_X1 stateArray_MUX_inS12ser_mux_inst_6_U1_Ins_1_U1 ( .A(plaintext_s1[78]), .B(ciphertext_s1[70]), .S(n221), .Z(new_AGEMA_signal_2294) );
  MUX2_X1 stateArray_MUX_inS12ser_mux_inst_7_U1_Ins_0_U1 ( .A(plaintext_s0[79]), .B(ciphertext_s0[71]), .S(n222), .Z(stateArray_inS12ser[7]) );
  MUX2_X1 stateArray_MUX_inS12ser_mux_inst_7_U1_Ins_1_U1 ( .A(plaintext_s1[79]), .B(ciphertext_s1[71]), .S(n222), .Z(new_AGEMA_signal_2297) );
  MUX2_X1 stateArray_MUX_outS20_MC_mux_inst_0_U1_Ins_0_U1 ( .A(
        ciphertext_s0[56]), .B(StateInMC[16]), .S(n161), .Z(
        stateArray_outS20ser_MC[0]) );
  MUX2_X1 stateArray_MUX_outS20_MC_mux_inst_0_U1_Ins_1_U1 ( .A(
        ciphertext_s1[56]), .B(new_AGEMA_signal_2872), .S(n161), .Z(
        new_AGEMA_signal_3016) );
  MUX2_X1 stateArray_MUX_outS20_MC_mux_inst_1_U1_Ins_0_U1 ( .A(
        ciphertext_s0[57]), .B(StateInMC[17]), .S(n161), .Z(
        stateArray_outS20ser_MC[1]) );
  MUX2_X1 stateArray_MUX_outS20_MC_mux_inst_1_U1_Ins_1_U1 ( .A(
        ciphertext_s1[57]), .B(new_AGEMA_signal_2873), .S(n161), .Z(
        new_AGEMA_signal_3017) );
  MUX2_X1 stateArray_MUX_outS20_MC_mux_inst_2_U1_Ins_0_U1 ( .A(
        ciphertext_s0[58]), .B(StateInMC[18]), .S(n161), .Z(
        stateArray_outS20ser_MC[2]) );
  MUX2_X1 stateArray_MUX_outS20_MC_mux_inst_2_U1_Ins_1_U1 ( .A(
        ciphertext_s1[58]), .B(new_AGEMA_signal_2874), .S(n161), .Z(
        new_AGEMA_signal_3018) );
  MUX2_X1 stateArray_MUX_outS20_MC_mux_inst_3_U1_Ins_0_U1 ( .A(
        ciphertext_s0[59]), .B(StateInMC[19]), .S(n161), .Z(
        stateArray_outS20ser_MC[3]) );
  MUX2_X1 stateArray_MUX_outS20_MC_mux_inst_3_U1_Ins_1_U1 ( .A(
        ciphertext_s1[59]), .B(new_AGEMA_signal_2875), .S(n161), .Z(
        new_AGEMA_signal_3019) );
  MUX2_X1 stateArray_MUX_outS20_MC_mux_inst_4_U1_Ins_0_U1 ( .A(
        ciphertext_s0[60]), .B(StateInMC[20]), .S(n161), .Z(
        stateArray_outS20ser_MC[4]) );
  MUX2_X1 stateArray_MUX_outS20_MC_mux_inst_4_U1_Ins_1_U1 ( .A(
        ciphertext_s1[60]), .B(new_AGEMA_signal_2876), .S(n161), .Z(
        new_AGEMA_signal_3020) );
  MUX2_X1 stateArray_MUX_outS20_MC_mux_inst_5_U1_Ins_0_U1 ( .A(
        ciphertext_s0[61]), .B(StateInMC[21]), .S(n161), .Z(
        stateArray_outS20ser_MC[5]) );
  MUX2_X1 stateArray_MUX_outS20_MC_mux_inst_5_U1_Ins_1_U1 ( .A(
        ciphertext_s1[61]), .B(new_AGEMA_signal_2877), .S(n161), .Z(
        new_AGEMA_signal_3021) );
  MUX2_X1 stateArray_MUX_outS20_MC_mux_inst_6_U1_Ins_0_U1 ( .A(
        ciphertext_s0[62]), .B(StateInMC[22]), .S(n162), .Z(
        stateArray_outS20ser_MC[6]) );
  MUX2_X1 stateArray_MUX_outS20_MC_mux_inst_6_U1_Ins_1_U1 ( .A(
        ciphertext_s1[62]), .B(new_AGEMA_signal_2878), .S(n162), .Z(
        new_AGEMA_signal_3022) );
  MUX2_X1 stateArray_MUX_outS20_MC_mux_inst_7_U1_Ins_0_U1 ( .A(
        ciphertext_s0[63]), .B(StateInMC[23]), .S(n162), .Z(
        stateArray_outS20ser_MC[7]) );
  MUX2_X1 stateArray_MUX_outS20_MC_mux_inst_7_U1_Ins_1_U1 ( .A(
        ciphertext_s1[63]), .B(new_AGEMA_signal_2879), .S(n162), .Z(
        new_AGEMA_signal_3023) );
  MUX2_X1 stateArray_MUX_inS13ser_mux_inst_0_U1_Ins_0_U1 ( .A(plaintext_s0[64]), .B(stateArray_outS20ser_MC[0]), .S(n222), .Z(stateArray_inS13ser[0]) );
  MUX2_X1 stateArray_MUX_inS13ser_mux_inst_0_U1_Ins_1_U1 ( .A(plaintext_s1[64]), .B(new_AGEMA_signal_3016), .S(n222), .Z(new_AGEMA_signal_3062) );
  MUX2_X1 stateArray_MUX_inS13ser_mux_inst_1_U1_Ins_0_U1 ( .A(plaintext_s0[65]), .B(stateArray_outS20ser_MC[1]), .S(n222), .Z(stateArray_inS13ser[1]) );
  MUX2_X1 stateArray_MUX_inS13ser_mux_inst_1_U1_Ins_1_U1 ( .A(plaintext_s1[65]), .B(new_AGEMA_signal_3017), .S(n222), .Z(new_AGEMA_signal_3064) );
  MUX2_X1 stateArray_MUX_inS13ser_mux_inst_2_U1_Ins_0_U1 ( .A(plaintext_s0[66]), .B(stateArray_outS20ser_MC[2]), .S(n222), .Z(stateArray_inS13ser[2]) );
  MUX2_X1 stateArray_MUX_inS13ser_mux_inst_2_U1_Ins_1_U1 ( .A(plaintext_s1[66]), .B(new_AGEMA_signal_3018), .S(n222), .Z(new_AGEMA_signal_3066) );
  MUX2_X1 stateArray_MUX_inS13ser_mux_inst_3_U1_Ins_0_U1 ( .A(plaintext_s0[67]), .B(stateArray_outS20ser_MC[3]), .S(n222), .Z(stateArray_inS13ser[3]) );
  MUX2_X1 stateArray_MUX_inS13ser_mux_inst_3_U1_Ins_1_U1 ( .A(plaintext_s1[67]), .B(new_AGEMA_signal_3019), .S(n222), .Z(new_AGEMA_signal_3068) );
  MUX2_X1 stateArray_MUX_inS13ser_mux_inst_4_U1_Ins_0_U1 ( .A(plaintext_s0[68]), .B(stateArray_outS20ser_MC[4]), .S(n222), .Z(stateArray_inS13ser[4]) );
  MUX2_X1 stateArray_MUX_inS13ser_mux_inst_4_U1_Ins_1_U1 ( .A(plaintext_s1[68]), .B(new_AGEMA_signal_3020), .S(n222), .Z(new_AGEMA_signal_3070) );
  MUX2_X1 stateArray_MUX_inS13ser_mux_inst_5_U1_Ins_0_U1 ( .A(plaintext_s0[69]), .B(stateArray_outS20ser_MC[5]), .S(n222), .Z(stateArray_inS13ser[5]) );
  MUX2_X1 stateArray_MUX_inS13ser_mux_inst_5_U1_Ins_1_U1 ( .A(plaintext_s1[69]), .B(new_AGEMA_signal_3021), .S(n222), .Z(new_AGEMA_signal_3072) );
  MUX2_X1 stateArray_MUX_inS13ser_mux_inst_6_U1_Ins_0_U1 ( .A(plaintext_s0[70]), .B(stateArray_outS20ser_MC[6]), .S(n223), .Z(stateArray_inS13ser[6]) );
  MUX2_X1 stateArray_MUX_inS13ser_mux_inst_6_U1_Ins_1_U1 ( .A(plaintext_s1[70]), .B(new_AGEMA_signal_3022), .S(n223), .Z(new_AGEMA_signal_3074) );
  MUX2_X1 stateArray_MUX_inS13ser_mux_inst_7_U1_Ins_0_U1 ( .A(plaintext_s0[71]), .B(stateArray_outS20ser_MC[7]), .S(n223), .Z(stateArray_inS13ser[7]) );
  MUX2_X1 stateArray_MUX_inS13ser_mux_inst_7_U1_Ins_1_U1 ( .A(plaintext_s1[71]), .B(new_AGEMA_signal_3023), .S(n223), .Z(new_AGEMA_signal_3076) );
  MUX2_X1 stateArray_MUX_inS20ser_mux_inst_0_U1_Ins_0_U1 ( .A(plaintext_s0[56]), .B(ciphertext_s0[48]), .S(n223), .Z(stateArray_inS20ser[0]) );
  MUX2_X1 stateArray_MUX_inS20ser_mux_inst_0_U1_Ins_1_U1 ( .A(plaintext_s1[56]), .B(ciphertext_s1[48]), .S(n223), .Z(new_AGEMA_signal_2300) );
  MUX2_X1 stateArray_MUX_inS20ser_mux_inst_1_U1_Ins_0_U1 ( .A(plaintext_s0[57]), .B(ciphertext_s0[49]), .S(n223), .Z(stateArray_inS20ser[1]) );
  MUX2_X1 stateArray_MUX_inS20ser_mux_inst_1_U1_Ins_1_U1 ( .A(plaintext_s1[57]), .B(ciphertext_s1[49]), .S(n223), .Z(new_AGEMA_signal_2303) );
  MUX2_X1 stateArray_MUX_inS20ser_mux_inst_2_U1_Ins_0_U1 ( .A(plaintext_s0[58]), .B(ciphertext_s0[50]), .S(n223), .Z(stateArray_inS20ser[2]) );
  MUX2_X1 stateArray_MUX_inS20ser_mux_inst_2_U1_Ins_1_U1 ( .A(plaintext_s1[58]), .B(ciphertext_s1[50]), .S(n223), .Z(new_AGEMA_signal_2306) );
  MUX2_X1 stateArray_MUX_inS20ser_mux_inst_3_U1_Ins_0_U1 ( .A(plaintext_s0[59]), .B(ciphertext_s0[51]), .S(n223), .Z(stateArray_inS20ser[3]) );
  MUX2_X1 stateArray_MUX_inS20ser_mux_inst_3_U1_Ins_1_U1 ( .A(plaintext_s1[59]), .B(ciphertext_s1[51]), .S(n223), .Z(new_AGEMA_signal_2309) );
  MUX2_X1 stateArray_MUX_inS20ser_mux_inst_4_U1_Ins_0_U1 ( .A(plaintext_s0[60]), .B(ciphertext_s0[52]), .S(n224), .Z(stateArray_inS20ser[4]) );
  MUX2_X1 stateArray_MUX_inS20ser_mux_inst_4_U1_Ins_1_U1 ( .A(plaintext_s1[60]), .B(ciphertext_s1[52]), .S(n224), .Z(new_AGEMA_signal_2312) );
  MUX2_X1 stateArray_MUX_inS20ser_mux_inst_5_U1_Ins_0_U1 ( .A(plaintext_s0[61]), .B(ciphertext_s0[53]), .S(n224), .Z(stateArray_inS20ser[5]) );
  MUX2_X1 stateArray_MUX_inS20ser_mux_inst_5_U1_Ins_1_U1 ( .A(plaintext_s1[61]), .B(ciphertext_s1[53]), .S(n224), .Z(new_AGEMA_signal_2315) );
  MUX2_X1 stateArray_MUX_inS20ser_mux_inst_6_U1_Ins_0_U1 ( .A(plaintext_s0[62]), .B(ciphertext_s0[54]), .S(n224), .Z(stateArray_inS20ser[6]) );
  MUX2_X1 stateArray_MUX_inS20ser_mux_inst_6_U1_Ins_1_U1 ( .A(plaintext_s1[62]), .B(ciphertext_s1[54]), .S(n224), .Z(new_AGEMA_signal_2318) );
  MUX2_X1 stateArray_MUX_inS20ser_mux_inst_7_U1_Ins_0_U1 ( .A(plaintext_s0[63]), .B(ciphertext_s0[55]), .S(n224), .Z(stateArray_inS20ser[7]) );
  MUX2_X1 stateArray_MUX_inS20ser_mux_inst_7_U1_Ins_1_U1 ( .A(plaintext_s1[63]), .B(ciphertext_s1[55]), .S(n224), .Z(new_AGEMA_signal_2321) );
  MUX2_X1 stateArray_MUX_inS21ser_mux_inst_0_U1_Ins_0_U1 ( .A(plaintext_s0[48]), .B(ciphertext_s0[40]), .S(n224), .Z(stateArray_inS21ser[0]) );
  MUX2_X1 stateArray_MUX_inS21ser_mux_inst_0_U1_Ins_1_U1 ( .A(plaintext_s1[48]), .B(ciphertext_s1[40]), .S(n224), .Z(new_AGEMA_signal_2324) );
  MUX2_X1 stateArray_MUX_inS21ser_mux_inst_1_U1_Ins_0_U1 ( .A(plaintext_s0[49]), .B(ciphertext_s0[41]), .S(n224), .Z(stateArray_inS21ser[1]) );
  MUX2_X1 stateArray_MUX_inS21ser_mux_inst_1_U1_Ins_1_U1 ( .A(plaintext_s1[49]), .B(ciphertext_s1[41]), .S(n224), .Z(new_AGEMA_signal_2327) );
  MUX2_X1 stateArray_MUX_inS21ser_mux_inst_2_U1_Ins_0_U1 ( .A(plaintext_s0[50]), .B(ciphertext_s0[42]), .S(n225), .Z(stateArray_inS21ser[2]) );
  MUX2_X1 stateArray_MUX_inS21ser_mux_inst_2_U1_Ins_1_U1 ( .A(plaintext_s1[50]), .B(ciphertext_s1[42]), .S(n225), .Z(new_AGEMA_signal_2330) );
  MUX2_X1 stateArray_MUX_inS21ser_mux_inst_3_U1_Ins_0_U1 ( .A(plaintext_s0[51]), .B(ciphertext_s0[43]), .S(n224), .Z(stateArray_inS21ser[3]) );
  MUX2_X1 stateArray_MUX_inS21ser_mux_inst_3_U1_Ins_1_U1 ( .A(plaintext_s1[51]), .B(ciphertext_s1[43]), .S(n224), .Z(new_AGEMA_signal_2333) );
  MUX2_X1 stateArray_MUX_inS21ser_mux_inst_4_U1_Ins_0_U1 ( .A(plaintext_s0[52]), .B(ciphertext_s0[44]), .S(n225), .Z(stateArray_inS21ser[4]) );
  MUX2_X1 stateArray_MUX_inS21ser_mux_inst_4_U1_Ins_1_U1 ( .A(plaintext_s1[52]), .B(ciphertext_s1[44]), .S(n225), .Z(new_AGEMA_signal_2336) );
  MUX2_X1 stateArray_MUX_inS21ser_mux_inst_5_U1_Ins_0_U1 ( .A(plaintext_s0[53]), .B(ciphertext_s0[45]), .S(n225), .Z(stateArray_inS21ser[5]) );
  MUX2_X1 stateArray_MUX_inS21ser_mux_inst_5_U1_Ins_1_U1 ( .A(plaintext_s1[53]), .B(ciphertext_s1[45]), .S(n225), .Z(new_AGEMA_signal_2339) );
  MUX2_X1 stateArray_MUX_inS21ser_mux_inst_6_U1_Ins_0_U1 ( .A(plaintext_s0[54]), .B(ciphertext_s0[46]), .S(n225), .Z(stateArray_inS21ser[6]) );
  MUX2_X1 stateArray_MUX_inS21ser_mux_inst_6_U1_Ins_1_U1 ( .A(plaintext_s1[54]), .B(ciphertext_s1[46]), .S(n225), .Z(new_AGEMA_signal_2342) );
  MUX2_X1 stateArray_MUX_inS21ser_mux_inst_7_U1_Ins_0_U1 ( .A(plaintext_s0[55]), .B(ciphertext_s0[47]), .S(n225), .Z(stateArray_inS21ser[7]) );
  MUX2_X1 stateArray_MUX_inS21ser_mux_inst_7_U1_Ins_1_U1 ( .A(plaintext_s1[55]), .B(ciphertext_s1[47]), .S(n225), .Z(new_AGEMA_signal_2345) );
  MUX2_X1 stateArray_MUX_inS22ser_mux_inst_0_U1_Ins_0_U1 ( .A(plaintext_s0[40]), .B(ciphertext_s0[32]), .S(n225), .Z(stateArray_inS22ser[0]) );
  MUX2_X1 stateArray_MUX_inS22ser_mux_inst_0_U1_Ins_1_U1 ( .A(plaintext_s1[40]), .B(ciphertext_s1[32]), .S(n225), .Z(new_AGEMA_signal_2348) );
  MUX2_X1 stateArray_MUX_inS22ser_mux_inst_1_U1_Ins_0_U1 ( .A(plaintext_s0[41]), .B(ciphertext_s0[33]), .S(n225), .Z(stateArray_inS22ser[1]) );
  MUX2_X1 stateArray_MUX_inS22ser_mux_inst_1_U1_Ins_1_U1 ( .A(plaintext_s1[41]), .B(ciphertext_s1[33]), .S(n225), .Z(new_AGEMA_signal_2351) );
  MUX2_X1 stateArray_MUX_inS22ser_mux_inst_2_U1_Ins_0_U1 ( .A(plaintext_s0[42]), .B(ciphertext_s0[34]), .S(n226), .Z(stateArray_inS22ser[2]) );
  MUX2_X1 stateArray_MUX_inS22ser_mux_inst_2_U1_Ins_1_U1 ( .A(plaintext_s1[42]), .B(ciphertext_s1[34]), .S(n226), .Z(new_AGEMA_signal_2354) );
  MUX2_X1 stateArray_MUX_inS22ser_mux_inst_3_U1_Ins_0_U1 ( .A(plaintext_s0[43]), .B(ciphertext_s0[35]), .S(n226), .Z(stateArray_inS22ser[3]) );
  MUX2_X1 stateArray_MUX_inS22ser_mux_inst_3_U1_Ins_1_U1 ( .A(plaintext_s1[43]), .B(ciphertext_s1[35]), .S(n226), .Z(new_AGEMA_signal_2357) );
  MUX2_X1 stateArray_MUX_inS22ser_mux_inst_4_U1_Ins_0_U1 ( .A(plaintext_s0[44]), .B(ciphertext_s0[36]), .S(n226), .Z(stateArray_inS22ser[4]) );
  MUX2_X1 stateArray_MUX_inS22ser_mux_inst_4_U1_Ins_1_U1 ( .A(plaintext_s1[44]), .B(ciphertext_s1[36]), .S(n226), .Z(new_AGEMA_signal_2360) );
  MUX2_X1 stateArray_MUX_inS22ser_mux_inst_5_U1_Ins_0_U1 ( .A(plaintext_s0[45]), .B(ciphertext_s0[37]), .S(n226), .Z(stateArray_inS22ser[5]) );
  MUX2_X1 stateArray_MUX_inS22ser_mux_inst_5_U1_Ins_1_U1 ( .A(plaintext_s1[45]), .B(ciphertext_s1[37]), .S(n226), .Z(new_AGEMA_signal_2363) );
  MUX2_X1 stateArray_MUX_inS22ser_mux_inst_6_U1_Ins_0_U1 ( .A(plaintext_s0[46]), .B(ciphertext_s0[38]), .S(n226), .Z(stateArray_inS22ser[6]) );
  MUX2_X1 stateArray_MUX_inS22ser_mux_inst_6_U1_Ins_1_U1 ( .A(plaintext_s1[46]), .B(ciphertext_s1[38]), .S(n226), .Z(new_AGEMA_signal_2366) );
  MUX2_X1 stateArray_MUX_inS22ser_mux_inst_7_U1_Ins_0_U1 ( .A(plaintext_s0[47]), .B(ciphertext_s0[39]), .S(n226), .Z(stateArray_inS22ser[7]) );
  MUX2_X1 stateArray_MUX_inS22ser_mux_inst_7_U1_Ins_1_U1 ( .A(plaintext_s1[47]), .B(ciphertext_s1[39]), .S(n226), .Z(new_AGEMA_signal_2369) );
  MUX2_X1 stateArray_MUX_outS30_MC_mux_inst_0_U1_Ins_0_U1 ( .A(
        ciphertext_s0[24]), .B(StateInMC[8]), .S(n162), .Z(
        stateArray_outS30ser_MC[0]) );
  MUX2_X1 stateArray_MUX_outS30_MC_mux_inst_0_U1_Ins_1_U1 ( .A(
        ciphertext_s1[24]), .B(new_AGEMA_signal_2864), .S(n162), .Z(
        new_AGEMA_signal_3024) );
  MUX2_X1 stateArray_MUX_outS30_MC_mux_inst_1_U1_Ins_0_U1 ( .A(
        ciphertext_s0[25]), .B(StateInMC[9]), .S(n162), .Z(
        stateArray_outS30ser_MC[1]) );
  MUX2_X1 stateArray_MUX_outS30_MC_mux_inst_1_U1_Ins_1_U1 ( .A(
        ciphertext_s1[25]), .B(new_AGEMA_signal_2865), .S(n162), .Z(
        new_AGEMA_signal_3025) );
  MUX2_X1 stateArray_MUX_outS30_MC_mux_inst_2_U1_Ins_0_U1 ( .A(
        ciphertext_s0[26]), .B(StateInMC[10]), .S(n162), .Z(
        stateArray_outS30ser_MC[2]) );
  MUX2_X1 stateArray_MUX_outS30_MC_mux_inst_2_U1_Ins_1_U1 ( .A(
        ciphertext_s1[26]), .B(new_AGEMA_signal_2866), .S(n162), .Z(
        new_AGEMA_signal_3026) );
  MUX2_X1 stateArray_MUX_outS30_MC_mux_inst_3_U1_Ins_0_U1 ( .A(
        ciphertext_s0[27]), .B(StateInMC[11]), .S(n162), .Z(
        stateArray_outS30ser_MC[3]) );
  MUX2_X1 stateArray_MUX_outS30_MC_mux_inst_3_U1_Ins_1_U1 ( .A(
        ciphertext_s1[27]), .B(new_AGEMA_signal_2867), .S(n162), .Z(
        new_AGEMA_signal_3027) );
  MUX2_X1 stateArray_MUX_outS30_MC_mux_inst_4_U1_Ins_0_U1 ( .A(
        ciphertext_s0[28]), .B(StateInMC[12]), .S(n162), .Z(
        stateArray_outS30ser_MC[4]) );
  MUX2_X1 stateArray_MUX_outS30_MC_mux_inst_4_U1_Ins_1_U1 ( .A(
        ciphertext_s1[28]), .B(new_AGEMA_signal_2868), .S(n162), .Z(
        new_AGEMA_signal_3028) );
  MUX2_X1 stateArray_MUX_outS30_MC_mux_inst_5_U1_Ins_0_U1 ( .A(
        ciphertext_s0[29]), .B(StateInMC[13]), .S(n163), .Z(
        stateArray_outS30ser_MC[5]) );
  MUX2_X1 stateArray_MUX_outS30_MC_mux_inst_5_U1_Ins_1_U1 ( .A(
        ciphertext_s1[29]), .B(new_AGEMA_signal_2869), .S(n163), .Z(
        new_AGEMA_signal_3029) );
  MUX2_X1 stateArray_MUX_outS30_MC_mux_inst_6_U1_Ins_0_U1 ( .A(
        ciphertext_s0[30]), .B(StateInMC[14]), .S(n163), .Z(
        stateArray_outS30ser_MC[6]) );
  MUX2_X1 stateArray_MUX_outS30_MC_mux_inst_6_U1_Ins_1_U1 ( .A(
        ciphertext_s1[30]), .B(new_AGEMA_signal_2870), .S(n163), .Z(
        new_AGEMA_signal_3030) );
  MUX2_X1 stateArray_MUX_outS30_MC_mux_inst_7_U1_Ins_0_U1 ( .A(
        ciphertext_s0[31]), .B(StateInMC[15]), .S(n163), .Z(
        stateArray_outS30ser_MC[7]) );
  MUX2_X1 stateArray_MUX_outS30_MC_mux_inst_7_U1_Ins_1_U1 ( .A(
        ciphertext_s1[31]), .B(new_AGEMA_signal_2871), .S(n163), .Z(
        new_AGEMA_signal_3031) );
  MUX2_X1 stateArray_MUX_inS23ser_mux_inst_0_U1_Ins_0_U1 ( .A(plaintext_s0[32]), .B(stateArray_outS30ser_MC[0]), .S(n227), .Z(stateArray_inS23ser[0]) );
  MUX2_X1 stateArray_MUX_inS23ser_mux_inst_0_U1_Ins_1_U1 ( .A(plaintext_s1[32]), .B(new_AGEMA_signal_3024), .S(n227), .Z(new_AGEMA_signal_3078) );
  MUX2_X1 stateArray_MUX_inS23ser_mux_inst_1_U1_Ins_0_U1 ( .A(plaintext_s0[33]), .B(stateArray_outS30ser_MC[1]), .S(n226), .Z(stateArray_inS23ser[1]) );
  MUX2_X1 stateArray_MUX_inS23ser_mux_inst_1_U1_Ins_1_U1 ( .A(plaintext_s1[33]), .B(new_AGEMA_signal_3025), .S(n226), .Z(new_AGEMA_signal_3080) );
  MUX2_X1 stateArray_MUX_inS23ser_mux_inst_2_U1_Ins_0_U1 ( .A(plaintext_s0[34]), .B(stateArray_outS30ser_MC[2]), .S(n227), .Z(stateArray_inS23ser[2]) );
  MUX2_X1 stateArray_MUX_inS23ser_mux_inst_2_U1_Ins_1_U1 ( .A(plaintext_s1[34]), .B(new_AGEMA_signal_3026), .S(n227), .Z(new_AGEMA_signal_3082) );
  MUX2_X1 stateArray_MUX_inS23ser_mux_inst_3_U1_Ins_0_U1 ( .A(plaintext_s0[35]), .B(stateArray_outS30ser_MC[3]), .S(n227), .Z(stateArray_inS23ser[3]) );
  MUX2_X1 stateArray_MUX_inS23ser_mux_inst_3_U1_Ins_1_U1 ( .A(plaintext_s1[35]), .B(new_AGEMA_signal_3027), .S(n227), .Z(new_AGEMA_signal_3084) );
  MUX2_X1 stateArray_MUX_inS23ser_mux_inst_4_U1_Ins_0_U1 ( .A(plaintext_s0[36]), .B(stateArray_outS30ser_MC[4]), .S(n227), .Z(stateArray_inS23ser[4]) );
  MUX2_X1 stateArray_MUX_inS23ser_mux_inst_4_U1_Ins_1_U1 ( .A(plaintext_s1[36]), .B(new_AGEMA_signal_3028), .S(n227), .Z(new_AGEMA_signal_3086) );
  MUX2_X1 stateArray_MUX_inS23ser_mux_inst_5_U1_Ins_0_U1 ( .A(plaintext_s0[37]), .B(stateArray_outS30ser_MC[5]), .S(n227), .Z(stateArray_inS23ser[5]) );
  MUX2_X1 stateArray_MUX_inS23ser_mux_inst_5_U1_Ins_1_U1 ( .A(plaintext_s1[37]), .B(new_AGEMA_signal_3029), .S(n227), .Z(new_AGEMA_signal_3088) );
  MUX2_X1 stateArray_MUX_inS23ser_mux_inst_6_U1_Ins_0_U1 ( .A(plaintext_s0[38]), .B(stateArray_outS30ser_MC[6]), .S(n227), .Z(stateArray_inS23ser[6]) );
  MUX2_X1 stateArray_MUX_inS23ser_mux_inst_6_U1_Ins_1_U1 ( .A(plaintext_s1[38]), .B(new_AGEMA_signal_3030), .S(n227), .Z(new_AGEMA_signal_3090) );
  MUX2_X1 stateArray_MUX_inS23ser_mux_inst_7_U1_Ins_0_U1 ( .A(plaintext_s0[39]), .B(stateArray_outS30ser_MC[7]), .S(n227), .Z(stateArray_inS23ser[7]) );
  MUX2_X1 stateArray_MUX_inS23ser_mux_inst_7_U1_Ins_1_U1 ( .A(plaintext_s1[39]), .B(new_AGEMA_signal_3031), .S(n227), .Z(new_AGEMA_signal_3092) );
  MUX2_X1 stateArray_MUX_inS30ser_mux_inst_0_U1_Ins_0_U1 ( .A(plaintext_s0[24]), .B(ciphertext_s0[16]), .S(n228), .Z(stateArray_inS30ser[0]) );
  MUX2_X1 stateArray_MUX_inS30ser_mux_inst_0_U1_Ins_1_U1 ( .A(plaintext_s1[24]), .B(ciphertext_s1[16]), .S(n228), .Z(new_AGEMA_signal_2372) );
  MUX2_X1 stateArray_MUX_inS30ser_mux_inst_1_U1_Ins_0_U1 ( .A(plaintext_s0[25]), .B(ciphertext_s0[17]), .S(n228), .Z(stateArray_inS30ser[1]) );
  MUX2_X1 stateArray_MUX_inS30ser_mux_inst_1_U1_Ins_1_U1 ( .A(plaintext_s1[25]), .B(ciphertext_s1[17]), .S(n228), .Z(new_AGEMA_signal_2375) );
  MUX2_X1 stateArray_MUX_inS30ser_mux_inst_2_U1_Ins_0_U1 ( .A(plaintext_s0[26]), .B(ciphertext_s0[18]), .S(n228), .Z(stateArray_inS30ser[2]) );
  MUX2_X1 stateArray_MUX_inS30ser_mux_inst_2_U1_Ins_1_U1 ( .A(plaintext_s1[26]), .B(ciphertext_s1[18]), .S(n228), .Z(new_AGEMA_signal_2378) );
  MUX2_X1 stateArray_MUX_inS30ser_mux_inst_3_U1_Ins_0_U1 ( .A(plaintext_s0[27]), .B(ciphertext_s0[19]), .S(n228), .Z(stateArray_inS30ser[3]) );
  MUX2_X1 stateArray_MUX_inS30ser_mux_inst_3_U1_Ins_1_U1 ( .A(plaintext_s1[27]), .B(ciphertext_s1[19]), .S(n228), .Z(new_AGEMA_signal_2381) );
  MUX2_X1 stateArray_MUX_inS30ser_mux_inst_4_U1_Ins_0_U1 ( .A(plaintext_s0[28]), .B(ciphertext_s0[20]), .S(n228), .Z(stateArray_inS30ser[4]) );
  MUX2_X1 stateArray_MUX_inS30ser_mux_inst_4_U1_Ins_1_U1 ( .A(plaintext_s1[28]), .B(ciphertext_s1[20]), .S(n228), .Z(new_AGEMA_signal_2384) );
  MUX2_X1 stateArray_MUX_inS30ser_mux_inst_5_U1_Ins_0_U1 ( .A(plaintext_s0[29]), .B(ciphertext_s0[21]), .S(n228), .Z(stateArray_inS30ser[5]) );
  MUX2_X1 stateArray_MUX_inS30ser_mux_inst_5_U1_Ins_1_U1 ( .A(plaintext_s1[29]), .B(ciphertext_s1[21]), .S(n228), .Z(new_AGEMA_signal_2387) );
  MUX2_X1 stateArray_MUX_inS30ser_mux_inst_6_U1_Ins_0_U1 ( .A(plaintext_s0[30]), .B(ciphertext_s0[22]), .S(n229), .Z(stateArray_inS30ser[6]) );
  MUX2_X1 stateArray_MUX_inS30ser_mux_inst_6_U1_Ins_1_U1 ( .A(plaintext_s1[30]), .B(ciphertext_s1[22]), .S(n229), .Z(new_AGEMA_signal_2390) );
  MUX2_X1 stateArray_MUX_inS30ser_mux_inst_7_U1_Ins_0_U1 ( .A(plaintext_s0[31]), .B(ciphertext_s0[23]), .S(n228), .Z(stateArray_inS30ser[7]) );
  MUX2_X1 stateArray_MUX_inS30ser_mux_inst_7_U1_Ins_1_U1 ( .A(plaintext_s1[31]), .B(ciphertext_s1[23]), .S(n228), .Z(new_AGEMA_signal_2393) );
  MUX2_X1 stateArray_MUX_inS31ser_mux_inst_0_U1_Ins_0_U1 ( .A(plaintext_s0[16]), .B(ciphertext_s0[8]), .S(n229), .Z(stateArray_inS31ser[0]) );
  MUX2_X1 stateArray_MUX_inS31ser_mux_inst_0_U1_Ins_1_U1 ( .A(plaintext_s1[16]), .B(ciphertext_s1[8]), .S(n229), .Z(new_AGEMA_signal_2396) );
  MUX2_X1 stateArray_MUX_inS31ser_mux_inst_1_U1_Ins_0_U1 ( .A(plaintext_s0[17]), .B(ciphertext_s0[9]), .S(n229), .Z(stateArray_inS31ser[1]) );
  MUX2_X1 stateArray_MUX_inS31ser_mux_inst_1_U1_Ins_1_U1 ( .A(plaintext_s1[17]), .B(ciphertext_s1[9]), .S(n229), .Z(new_AGEMA_signal_2399) );
  MUX2_X1 stateArray_MUX_inS31ser_mux_inst_2_U1_Ins_0_U1 ( .A(plaintext_s0[18]), .B(ciphertext_s0[10]), .S(n229), .Z(stateArray_inS31ser[2]) );
  MUX2_X1 stateArray_MUX_inS31ser_mux_inst_2_U1_Ins_1_U1 ( .A(plaintext_s1[18]), .B(ciphertext_s1[10]), .S(n229), .Z(new_AGEMA_signal_2402) );
  MUX2_X1 stateArray_MUX_inS31ser_mux_inst_3_U1_Ins_0_U1 ( .A(plaintext_s0[19]), .B(ciphertext_s0[11]), .S(n229), .Z(stateArray_inS31ser[3]) );
  MUX2_X1 stateArray_MUX_inS31ser_mux_inst_3_U1_Ins_1_U1 ( .A(plaintext_s1[19]), .B(ciphertext_s1[11]), .S(n229), .Z(new_AGEMA_signal_2405) );
  MUX2_X1 stateArray_MUX_inS31ser_mux_inst_4_U1_Ins_0_U1 ( .A(plaintext_s0[20]), .B(ciphertext_s0[12]), .S(n229), .Z(stateArray_inS31ser[4]) );
  MUX2_X1 stateArray_MUX_inS31ser_mux_inst_4_U1_Ins_1_U1 ( .A(plaintext_s1[20]), .B(ciphertext_s1[12]), .S(n229), .Z(new_AGEMA_signal_2408) );
  MUX2_X1 stateArray_MUX_inS31ser_mux_inst_5_U1_Ins_0_U1 ( .A(plaintext_s0[21]), .B(ciphertext_s0[13]), .S(n229), .Z(stateArray_inS31ser[5]) );
  MUX2_X1 stateArray_MUX_inS31ser_mux_inst_5_U1_Ins_1_U1 ( .A(plaintext_s1[21]), .B(ciphertext_s1[13]), .S(n229), .Z(new_AGEMA_signal_2411) );
  MUX2_X1 stateArray_MUX_inS31ser_mux_inst_6_U1_Ins_0_U1 ( .A(plaintext_s0[22]), .B(ciphertext_s0[14]), .S(n230), .Z(stateArray_inS31ser[6]) );
  MUX2_X1 stateArray_MUX_inS31ser_mux_inst_6_U1_Ins_1_U1 ( .A(plaintext_s1[22]), .B(ciphertext_s1[14]), .S(n230), .Z(new_AGEMA_signal_2414) );
  MUX2_X1 stateArray_MUX_inS31ser_mux_inst_7_U1_Ins_0_U1 ( .A(plaintext_s0[23]), .B(ciphertext_s0[15]), .S(n230), .Z(stateArray_inS31ser[7]) );
  MUX2_X1 stateArray_MUX_inS31ser_mux_inst_7_U1_Ins_1_U1 ( .A(plaintext_s1[23]), .B(ciphertext_s1[15]), .S(n230), .Z(new_AGEMA_signal_2417) );
  MUX2_X1 stateArray_MUX_inS32ser_mux_inst_0_U1_Ins_0_U1 ( .A(plaintext_s0[8]), 
        .B(ciphertext_s0[0]), .S(n230), .Z(stateArray_inS32ser[0]) );
  MUX2_X1 stateArray_MUX_inS32ser_mux_inst_0_U1_Ins_1_U1 ( .A(plaintext_s1[8]), 
        .B(ciphertext_s1[0]), .S(n230), .Z(new_AGEMA_signal_2420) );
  MUX2_X1 stateArray_MUX_inS32ser_mux_inst_1_U1_Ins_0_U1 ( .A(plaintext_s0[9]), 
        .B(ciphertext_s0[1]), .S(n230), .Z(stateArray_inS32ser[1]) );
  MUX2_X1 stateArray_MUX_inS32ser_mux_inst_1_U1_Ins_1_U1 ( .A(plaintext_s1[9]), 
        .B(ciphertext_s1[1]), .S(n230), .Z(new_AGEMA_signal_2423) );
  MUX2_X1 stateArray_MUX_inS32ser_mux_inst_2_U1_Ins_0_U1 ( .A(plaintext_s0[10]), .B(ciphertext_s0[2]), .S(n230), .Z(stateArray_inS32ser[2]) );
  MUX2_X1 stateArray_MUX_inS32ser_mux_inst_2_U1_Ins_1_U1 ( .A(plaintext_s1[10]), .B(ciphertext_s1[2]), .S(n230), .Z(new_AGEMA_signal_2426) );
  MUX2_X1 stateArray_MUX_inS32ser_mux_inst_3_U1_Ins_0_U1 ( .A(plaintext_s0[11]), .B(ciphertext_s0[3]), .S(n230), .Z(stateArray_inS32ser[3]) );
  MUX2_X1 stateArray_MUX_inS32ser_mux_inst_3_U1_Ins_1_U1 ( .A(plaintext_s1[11]), .B(ciphertext_s1[3]), .S(n230), .Z(new_AGEMA_signal_2429) );
  MUX2_X1 stateArray_MUX_inS32ser_mux_inst_4_U1_Ins_0_U1 ( .A(plaintext_s0[12]), .B(ciphertext_s0[4]), .S(n214), .Z(stateArray_inS32ser[4]) );
  MUX2_X1 stateArray_MUX_inS32ser_mux_inst_4_U1_Ins_1_U1 ( .A(plaintext_s1[12]), .B(ciphertext_s1[4]), .S(n214), .Z(new_AGEMA_signal_2432) );
  MUX2_X1 stateArray_MUX_inS32ser_mux_inst_5_U1_Ins_0_U1 ( .A(plaintext_s0[13]), .B(ciphertext_s0[5]), .S(n230), .Z(stateArray_inS32ser[5]) );
  MUX2_X1 stateArray_MUX_inS32ser_mux_inst_5_U1_Ins_1_U1 ( .A(plaintext_s1[13]), .B(ciphertext_s1[5]), .S(n230), .Z(new_AGEMA_signal_2435) );
  MUX2_X1 stateArray_MUX_inS32ser_mux_inst_6_U1_Ins_0_U1 ( .A(plaintext_s0[14]), .B(ciphertext_s0[6]), .S(n213), .Z(stateArray_inS32ser[6]) );
  MUX2_X1 stateArray_MUX_inS32ser_mux_inst_6_U1_Ins_1_U1 ( .A(plaintext_s1[14]), .B(ciphertext_s1[6]), .S(n213), .Z(new_AGEMA_signal_2438) );
  MUX2_X1 stateArray_MUX_inS32ser_mux_inst_7_U1_Ins_0_U1 ( .A(plaintext_s0[15]), .B(ciphertext_s0[7]), .S(n208), .Z(stateArray_inS32ser[7]) );
  MUX2_X1 stateArray_MUX_inS32ser_mux_inst_7_U1_Ins_1_U1 ( .A(plaintext_s1[15]), .B(ciphertext_s1[7]), .S(n208), .Z(new_AGEMA_signal_2441) );
  MUX2_X1 MUX_StateInMC_mux_inst_0_U1_Ins_0_U1 ( .A(MCout[0]), .B(
        ciphertext_s0[24]), .S(n156), .Z(StateInMC[0]) );
  MUX2_X1 MUX_StateInMC_mux_inst_0_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2825), 
        .B(ciphertext_s1[24]), .S(n156), .Z(new_AGEMA_signal_2860) );
  MUX2_X1 MUX_StateInMC_mux_inst_1_U1_Ins_0_U1 ( .A(MCout[1]), .B(
        ciphertext_s0[25]), .S(n159), .Z(StateInMC[1]) );
  MUX2_X1 MUX_StateInMC_mux_inst_1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2849), 
        .B(ciphertext_s1[25]), .S(n159), .Z(new_AGEMA_signal_2861) );
  MUX2_X1 MUX_StateInMC_mux_inst_2_U1_Ins_0_U1 ( .A(MCout[2]), .B(
        ciphertext_s0[26]), .S(n157), .Z(StateInMC[2]) );
  MUX2_X1 MUX_StateInMC_mux_inst_2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2823), 
        .B(ciphertext_s1[26]), .S(n157), .Z(new_AGEMA_signal_2834) );
  MUX2_X1 MUX_StateInMC_mux_inst_3_U1_Ins_0_U1 ( .A(MCout[3]), .B(
        ciphertext_s0[27]), .S(n158), .Z(StateInMC[3]) );
  MUX2_X1 MUX_StateInMC_mux_inst_3_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2848), 
        .B(ciphertext_s1[27]), .S(n158), .Z(new_AGEMA_signal_2862) );
  MUX2_X1 MUX_StateInMC_mux_inst_4_U1_Ins_0_U1 ( .A(MCout[4]), .B(
        ciphertext_s0[28]), .S(n141), .Z(StateInMC[4]) );
  MUX2_X1 MUX_StateInMC_mux_inst_4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2847), 
        .B(ciphertext_s1[28]), .S(n141), .Z(new_AGEMA_signal_2863) );
  MUX2_X1 MUX_StateInMC_mux_inst_5_U1_Ins_0_U1 ( .A(MCout[5]), .B(
        ciphertext_s0[29]), .S(n141), .Z(StateInMC[5]) );
  MUX2_X1 MUX_StateInMC_mux_inst_5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2820), 
        .B(ciphertext_s1[29]), .S(n141), .Z(new_AGEMA_signal_2835) );
  MUX2_X1 MUX_StateInMC_mux_inst_6_U1_Ins_0_U1 ( .A(MCout[6]), .B(
        ciphertext_s0[30]), .S(n141), .Z(StateInMC[6]) );
  MUX2_X1 MUX_StateInMC_mux_inst_6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2819), 
        .B(ciphertext_s1[30]), .S(n141), .Z(new_AGEMA_signal_2836) );
  MUX2_X1 MUX_StateInMC_mux_inst_7_U1_Ins_0_U1 ( .A(MCout[7]), .B(
        ciphertext_s0[31]), .S(n156), .Z(StateInMC[7]) );
  MUX2_X1 MUX_StateInMC_mux_inst_7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2818), 
        .B(ciphertext_s1[31]), .S(n156), .Z(new_AGEMA_signal_2837) );
  MUX2_X1 MUX_StateInMC_mux_inst_8_U1_Ins_0_U1 ( .A(MCout[8]), .B(
        ciphertext_s0[56]), .S(n156), .Z(StateInMC[8]) );
  MUX2_X1 MUX_StateInMC_mux_inst_8_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2817), 
        .B(ciphertext_s1[56]), .S(n156), .Z(new_AGEMA_signal_2864) );
  MUX2_X1 MUX_StateInMC_mux_inst_9_U1_Ins_0_U1 ( .A(MCout[9]), .B(
        ciphertext_s0[57]), .S(n156), .Z(StateInMC[9]) );
  MUX2_X1 MUX_StateInMC_mux_inst_9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2846), 
        .B(ciphertext_s1[57]), .S(n156), .Z(new_AGEMA_signal_2865) );
  MUX2_X1 MUX_StateInMC_mux_inst_10_U1_Ins_0_U1 ( .A(MCout[10]), .B(
        ciphertext_s0[58]), .S(n156), .Z(StateInMC[10]) );
  MUX2_X1 MUX_StateInMC_mux_inst_10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2815), 
        .B(ciphertext_s1[58]), .S(n156), .Z(new_AGEMA_signal_2866) );
  MUX2_X1 MUX_StateInMC_mux_inst_11_U1_Ins_0_U1 ( .A(MCout[11]), .B(
        ciphertext_s0[59]), .S(n156), .Z(StateInMC[11]) );
  MUX2_X1 MUX_StateInMC_mux_inst_11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2845), 
        .B(ciphertext_s1[59]), .S(n156), .Z(new_AGEMA_signal_2867) );
  MUX2_X1 MUX_StateInMC_mux_inst_12_U1_Ins_0_U1 ( .A(MCout[12]), .B(
        ciphertext_s0[60]), .S(n156), .Z(StateInMC[12]) );
  MUX2_X1 MUX_StateInMC_mux_inst_12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2844), 
        .B(ciphertext_s1[60]), .S(n156), .Z(new_AGEMA_signal_2868) );
  MUX2_X1 MUX_StateInMC_mux_inst_13_U1_Ins_0_U1 ( .A(MCout[13]), .B(
        ciphertext_s0[61]), .S(n156), .Z(StateInMC[13]) );
  MUX2_X1 MUX_StateInMC_mux_inst_13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2812), 
        .B(ciphertext_s1[61]), .S(n156), .Z(new_AGEMA_signal_2869) );
  MUX2_X1 MUX_StateInMC_mux_inst_14_U1_Ins_0_U1 ( .A(MCout[14]), .B(
        ciphertext_s0[62]), .S(n157), .Z(StateInMC[14]) );
  MUX2_X1 MUX_StateInMC_mux_inst_14_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2811), 
        .B(ciphertext_s1[62]), .S(n157), .Z(new_AGEMA_signal_2870) );
  MUX2_X1 MUX_StateInMC_mux_inst_15_U1_Ins_0_U1 ( .A(MCout[15]), .B(
        ciphertext_s0[63]), .S(n157), .Z(StateInMC[15]) );
  MUX2_X1 MUX_StateInMC_mux_inst_15_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2810), 
        .B(ciphertext_s1[63]), .S(n157), .Z(new_AGEMA_signal_2871) );
  MUX2_X1 MUX_StateInMC_mux_inst_16_U1_Ins_0_U1 ( .A(MCout[16]), .B(
        ciphertext_s0[88]), .S(n157), .Z(StateInMC[16]) );
  MUX2_X1 MUX_StateInMC_mux_inst_16_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2809), 
        .B(ciphertext_s1[88]), .S(n157), .Z(new_AGEMA_signal_2872) );
  MUX2_X1 MUX_StateInMC_mux_inst_17_U1_Ins_0_U1 ( .A(MCout[17]), .B(
        ciphertext_s0[89]), .S(n157), .Z(StateInMC[17]) );
  MUX2_X1 MUX_StateInMC_mux_inst_17_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2843), 
        .B(ciphertext_s1[89]), .S(n157), .Z(new_AGEMA_signal_2873) );
  MUX2_X1 MUX_StateInMC_mux_inst_18_U1_Ins_0_U1 ( .A(MCout[18]), .B(
        ciphertext_s0[90]), .S(n157), .Z(StateInMC[18]) );
  MUX2_X1 MUX_StateInMC_mux_inst_18_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2807), 
        .B(ciphertext_s1[90]), .S(n157), .Z(new_AGEMA_signal_2874) );
  MUX2_X1 MUX_StateInMC_mux_inst_19_U1_Ins_0_U1 ( .A(MCout[19]), .B(
        ciphertext_s0[91]), .S(n157), .Z(StateInMC[19]) );
  MUX2_X1 MUX_StateInMC_mux_inst_19_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2842), 
        .B(ciphertext_s1[91]), .S(n157), .Z(new_AGEMA_signal_2875) );
  MUX2_X1 MUX_StateInMC_mux_inst_20_U1_Ins_0_U1 ( .A(MCout[20]), .B(
        ciphertext_s0[92]), .S(n157), .Z(StateInMC[20]) );
  MUX2_X1 MUX_StateInMC_mux_inst_20_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2841), 
        .B(ciphertext_s1[92]), .S(n157), .Z(new_AGEMA_signal_2876) );
  MUX2_X1 MUX_StateInMC_mux_inst_21_U1_Ins_0_U1 ( .A(MCout[21]), .B(
        ciphertext_s0[93]), .S(n158), .Z(StateInMC[21]) );
  MUX2_X1 MUX_StateInMC_mux_inst_21_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2804), 
        .B(ciphertext_s1[93]), .S(n158), .Z(new_AGEMA_signal_2877) );
  MUX2_X1 MUX_StateInMC_mux_inst_22_U1_Ins_0_U1 ( .A(MCout[22]), .B(
        ciphertext_s0[94]), .S(n158), .Z(StateInMC[22]) );
  MUX2_X1 MUX_StateInMC_mux_inst_22_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2803), 
        .B(ciphertext_s1[94]), .S(n158), .Z(new_AGEMA_signal_2878) );
  MUX2_X1 MUX_StateInMC_mux_inst_23_U1_Ins_0_U1 ( .A(MCout[23]), .B(
        ciphertext_s0[95]), .S(n158), .Z(StateInMC[23]) );
  MUX2_X1 MUX_StateInMC_mux_inst_23_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2802), 
        .B(ciphertext_s1[95]), .S(n158), .Z(new_AGEMA_signal_2879) );
  MUX2_X1 MUX_StateInMC_mux_inst_24_U1_Ins_0_U1 ( .A(MCout[24]), .B(
        ciphertext_s0[120]), .S(n158), .Z(StateInMC[24]) );
  MUX2_X1 MUX_StateInMC_mux_inst_24_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2801), 
        .B(ciphertext_s1[120]), .S(n158), .Z(new_AGEMA_signal_2880) );
  MUX2_X1 MUX_StateInMC_mux_inst_25_U1_Ins_0_U1 ( .A(MCout[25]), .B(
        ciphertext_s0[121]), .S(n158), .Z(StateInMC[25]) );
  MUX2_X1 MUX_StateInMC_mux_inst_25_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2840), 
        .B(ciphertext_s1[121]), .S(n158), .Z(new_AGEMA_signal_2881) );
  MUX2_X1 MUX_StateInMC_mux_inst_26_U1_Ins_0_U1 ( .A(MCout[26]), .B(
        ciphertext_s0[122]), .S(n158), .Z(StateInMC[26]) );
  MUX2_X1 MUX_StateInMC_mux_inst_26_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2799), 
        .B(ciphertext_s1[122]), .S(n158), .Z(new_AGEMA_signal_2882) );
  MUX2_X1 MUX_StateInMC_mux_inst_27_U1_Ins_0_U1 ( .A(MCout[27]), .B(
        ciphertext_s0[123]), .S(n158), .Z(StateInMC[27]) );
  MUX2_X1 MUX_StateInMC_mux_inst_27_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2839), 
        .B(ciphertext_s1[123]), .S(n158), .Z(new_AGEMA_signal_2883) );
  MUX2_X1 MUX_StateInMC_mux_inst_28_U1_Ins_0_U1 ( .A(MCout[28]), .B(
        ciphertext_s0[124]), .S(n159), .Z(StateInMC[28]) );
  MUX2_X1 MUX_StateInMC_mux_inst_28_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2838), 
        .B(ciphertext_s1[124]), .S(n159), .Z(new_AGEMA_signal_2884) );
  MUX2_X1 MUX_StateInMC_mux_inst_29_U1_Ins_0_U1 ( .A(MCout[29]), .B(
        ciphertext_s0[125]), .S(n159), .Z(StateInMC[29]) );
  MUX2_X1 MUX_StateInMC_mux_inst_29_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2796), 
        .B(ciphertext_s1[125]), .S(n159), .Z(new_AGEMA_signal_2885) );
  MUX2_X1 MUX_StateInMC_mux_inst_30_U1_Ins_0_U1 ( .A(MCout[30]), .B(
        ciphertext_s0[126]), .S(n159), .Z(StateInMC[30]) );
  MUX2_X1 MUX_StateInMC_mux_inst_30_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2795), 
        .B(ciphertext_s1[126]), .S(n159), .Z(new_AGEMA_signal_2886) );
  MUX2_X1 MUX_StateInMC_mux_inst_31_U1_Ins_0_U1 ( .A(MCout[31]), .B(
        ciphertext_s0[127]), .S(n159), .Z(StateInMC[31]) );
  MUX2_X1 MUX_StateInMC_mux_inst_31_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2794), 
        .B(ciphertext_s1[127]), .S(n159), .Z(new_AGEMA_signal_2887) );
  XOR2_X1 KeyArray_U50_Ins_0_U1 ( .A(KeyArray_outS01ser_7_), .B(keyStateIn[7]), 
        .Z(KeyArray_outS01ser_XOR_00[7]) );
  XOR2_X1 KeyArray_U50_Ins_1_U1 ( .A(new_AGEMA_signal_2006), .B(
        new_AGEMA_signal_2004), .Z(new_AGEMA_signal_2007) );
  XOR2_X1 KeyArray_U49_Ins_0_U1 ( .A(KeyArray_outS01ser_6_), .B(keyStateIn[6]), 
        .Z(KeyArray_outS01ser_XOR_00[6]) );
  XOR2_X1 KeyArray_U49_Ins_1_U1 ( .A(new_AGEMA_signal_2008), .B(
        new_AGEMA_signal_2001), .Z(new_AGEMA_signal_2009) );
  XOR2_X1 KeyArray_U48_Ins_0_U1 ( .A(KeyArray_outS01ser_5_), .B(keyStateIn[5]), 
        .Z(KeyArray_outS01ser_XOR_00[5]) );
  XOR2_X1 KeyArray_U48_Ins_1_U1 ( .A(new_AGEMA_signal_2010), .B(
        new_AGEMA_signal_1998), .Z(new_AGEMA_signal_2011) );
  XOR2_X1 KeyArray_U47_Ins_0_U1 ( .A(KeyArray_outS01ser_4_), .B(keyStateIn[4]), 
        .Z(KeyArray_outS01ser_XOR_00[4]) );
  XOR2_X1 KeyArray_U47_Ins_1_U1 ( .A(new_AGEMA_signal_2012), .B(
        new_AGEMA_signal_1995), .Z(new_AGEMA_signal_2013) );
  XOR2_X1 KeyArray_U46_Ins_0_U1 ( .A(KeyArray_outS01ser_3_), .B(keyStateIn[3]), 
        .Z(KeyArray_outS01ser_XOR_00[3]) );
  XOR2_X1 KeyArray_U46_Ins_1_U1 ( .A(new_AGEMA_signal_2014), .B(
        new_AGEMA_signal_1992), .Z(new_AGEMA_signal_2015) );
  XOR2_X1 KeyArray_U45_Ins_0_U1 ( .A(KeyArray_outS01ser_2_), .B(keyStateIn[2]), 
        .Z(KeyArray_outS01ser_XOR_00[2]) );
  XOR2_X1 KeyArray_U45_Ins_1_U1 ( .A(new_AGEMA_signal_2016), .B(
        new_AGEMA_signal_1989), .Z(new_AGEMA_signal_2017) );
  XOR2_X1 KeyArray_U44_Ins_0_U1 ( .A(KeyArray_outS01ser_1_), .B(keyStateIn[1]), 
        .Z(KeyArray_outS01ser_XOR_00[1]) );
  XOR2_X1 KeyArray_U44_Ins_1_U1 ( .A(new_AGEMA_signal_2018), .B(
        new_AGEMA_signal_1986), .Z(new_AGEMA_signal_2019) );
  XOR2_X1 KeyArray_U43_Ins_0_U1 ( .A(KeyArray_outS01ser_0_), .B(keyStateIn[0]), 
        .Z(KeyArray_outS01ser_XOR_00[0]) );
  XOR2_X1 KeyArray_U43_Ins_1_U1 ( .A(new_AGEMA_signal_2020), .B(
        new_AGEMA_signal_1983), .Z(new_AGEMA_signal_2021) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_0_U1_Ins_0_U1 ( .A(keyStateIn[0]), .B(
        KeyArray_S00reg_gff_1_SFF_0_QD), .S(n177), .Z(
        KeyArray_S00reg_gff_1_SFF_0_n5) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_0_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1983), 
        .B(new_AGEMA_signal_3267), .S(n177), .Z(new_AGEMA_signal_3375) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS00ser[0]), .B(KeyArray_outS10ser[0]), .S(n163), .Z(
        KeyArray_S00reg_gff_1_SFF_0_QD) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3247), .B(new_AGEMA_signal_2491), .S(n163), .Z(
        new_AGEMA_signal_3267) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_1_U1_Ins_0_U1 ( .A(keyStateIn[1]), .B(
        KeyArray_S00reg_gff_1_SFF_1_QD), .S(n190), .Z(
        KeyArray_S00reg_gff_1_SFF_1_n6) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1986), 
        .B(new_AGEMA_signal_3268), .S(n190), .Z(new_AGEMA_signal_3376) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS00ser[1]), .B(KeyArray_outS10ser[1]), .S(n163), .Z(
        KeyArray_S00reg_gff_1_SFF_1_QD) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3249), .B(new_AGEMA_signal_2494), .S(n163), .Z(
        new_AGEMA_signal_3268) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_2_U1_Ins_0_U1 ( .A(keyStateIn[2]), .B(
        KeyArray_S00reg_gff_1_SFF_2_QD), .S(n189), .Z(
        KeyArray_S00reg_gff_1_SFF_2_n6) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1989), 
        .B(new_AGEMA_signal_3269), .S(n189), .Z(new_AGEMA_signal_3377) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS00ser[2]), .B(KeyArray_outS10ser[2]), .S(n163), .Z(
        KeyArray_S00reg_gff_1_SFF_2_QD) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3251), .B(new_AGEMA_signal_2497), .S(n163), .Z(
        new_AGEMA_signal_3269) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_3_U1_Ins_0_U1 ( .A(keyStateIn[3]), .B(
        KeyArray_S00reg_gff_1_SFF_3_QD), .S(n190), .Z(
        KeyArray_S00reg_gff_1_SFF_3_n6) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_3_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1992), 
        .B(new_AGEMA_signal_3270), .S(n190), .Z(new_AGEMA_signal_3378) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS00ser[3]), .B(KeyArray_outS10ser[3]), .S(n163), .Z(
        KeyArray_S00reg_gff_1_SFF_3_QD) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3253), .B(new_AGEMA_signal_2500), .S(n163), .Z(
        new_AGEMA_signal_3270) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_4_U1_Ins_0_U1 ( .A(keyStateIn[4]), .B(
        KeyArray_S00reg_gff_1_SFF_4_QD), .S(n189), .Z(
        KeyArray_S00reg_gff_1_SFF_4_n6) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1995), 
        .B(new_AGEMA_signal_3271), .S(n189), .Z(new_AGEMA_signal_3379) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS00ser[4]), .B(KeyArray_outS10ser[4]), .S(n161), .Z(
        KeyArray_S00reg_gff_1_SFF_4_QD) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3255), .B(new_AGEMA_signal_2503), .S(n161), .Z(
        new_AGEMA_signal_3271) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_5_U1_Ins_0_U1 ( .A(keyStateIn[5]), .B(
        KeyArray_S00reg_gff_1_SFF_5_QD), .S(n189), .Z(
        KeyArray_S00reg_gff_1_SFF_5_n6) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1998), 
        .B(new_AGEMA_signal_3272), .S(n189), .Z(new_AGEMA_signal_3380) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS00ser[5]), .B(KeyArray_outS10ser[5]), .S(n163), .Z(
        KeyArray_S00reg_gff_1_SFF_5_QD) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3257), .B(new_AGEMA_signal_2506), .S(n163), .Z(
        new_AGEMA_signal_3272) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_6_U1_Ins_0_U1 ( .A(keyStateIn[6]), .B(
        KeyArray_S00reg_gff_1_SFF_6_QD), .S(n189), .Z(
        KeyArray_S00reg_gff_1_SFF_6_n6) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2001), 
        .B(new_AGEMA_signal_3273), .S(n189), .Z(new_AGEMA_signal_3381) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS00ser[6]), .B(KeyArray_outS10ser[6]), .S(n160), .Z(
        KeyArray_S00reg_gff_1_SFF_6_QD) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3259), .B(new_AGEMA_signal_2509), .S(n160), .Z(
        new_AGEMA_signal_3273) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_7_U1_Ins_0_U1 ( .A(keyStateIn[7]), .B(
        KeyArray_S00reg_gff_1_SFF_7_QD), .S(n189), .Z(
        KeyArray_S00reg_gff_1_SFF_7_n6) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2004), 
        .B(new_AGEMA_signal_3274), .S(n189), .Z(new_AGEMA_signal_3382) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS00ser[7]), .B(KeyArray_outS10ser[7]), .S(n161), .Z(
        KeyArray_S00reg_gff_1_SFF_7_QD) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3261), .B(new_AGEMA_signal_2512), .S(n161), .Z(
        new_AGEMA_signal_3274) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_0_U1_Ins_0_U1 ( .A(KeyArray_outS01ser_0_), 
        .B(KeyArray_S01reg_gff_1_SFF_0_QD), .S(n189), .Z(
        KeyArray_S01reg_gff_1_SFF_0_n6) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_0_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2020), 
        .B(new_AGEMA_signal_2888), .S(n189), .Z(new_AGEMA_signal_3275) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS01ser[0]), .B(KeyArray_outS11ser[0]), .S(n163), .Z(
        KeyArray_S01reg_gff_1_SFF_0_QD) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2444), .B(new_AGEMA_signal_2515), .S(n163), .Z(
        new_AGEMA_signal_2888) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_1_U1_Ins_0_U1 ( .A(KeyArray_outS01ser_1_), 
        .B(KeyArray_S01reg_gff_1_SFF_1_QD), .S(n189), .Z(
        KeyArray_S01reg_gff_1_SFF_1_n6) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2018), 
        .B(new_AGEMA_signal_2889), .S(n189), .Z(new_AGEMA_signal_3276) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS01ser[1]), .B(KeyArray_outS11ser[1]), .S(n161), .Z(
        KeyArray_S01reg_gff_1_SFF_1_QD) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2447), .B(new_AGEMA_signal_2518), .S(n161), .Z(
        new_AGEMA_signal_2889) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_2_U1_Ins_0_U1 ( .A(KeyArray_outS01ser_2_), 
        .B(KeyArray_S01reg_gff_1_SFF_2_QD), .S(n188), .Z(
        KeyArray_S01reg_gff_1_SFF_2_n6) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2016), 
        .B(new_AGEMA_signal_2890), .S(n188), .Z(new_AGEMA_signal_3277) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS01ser[2]), .B(KeyArray_outS11ser[2]), .S(n164), .Z(
        KeyArray_S01reg_gff_1_SFF_2_QD) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2450), .B(new_AGEMA_signal_2521), .S(n164), .Z(
        new_AGEMA_signal_2890) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_3_U1_Ins_0_U1 ( .A(KeyArray_outS01ser_3_), 
        .B(KeyArray_S01reg_gff_1_SFF_3_QD), .S(n188), .Z(
        KeyArray_S01reg_gff_1_SFF_3_n6) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_3_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2014), 
        .B(new_AGEMA_signal_2891), .S(n188), .Z(new_AGEMA_signal_3278) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS01ser[3]), .B(KeyArray_outS11ser[3]), .S(n167), .Z(
        KeyArray_S01reg_gff_1_SFF_3_QD) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2453), .B(new_AGEMA_signal_2524), .S(n167), .Z(
        new_AGEMA_signal_2891) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_4_U1_Ins_0_U1 ( .A(KeyArray_outS01ser_4_), 
        .B(KeyArray_S01reg_gff_1_SFF_4_QD), .S(n188), .Z(
        KeyArray_S01reg_gff_1_SFF_4_n6) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2012), 
        .B(new_AGEMA_signal_2892), .S(n188), .Z(new_AGEMA_signal_3279) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS01ser[4]), .B(KeyArray_outS11ser[4]), .S(n171), .Z(
        KeyArray_S01reg_gff_1_SFF_4_QD) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2456), .B(new_AGEMA_signal_2527), .S(n171), .Z(
        new_AGEMA_signal_2892) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_5_U1_Ins_0_U1 ( .A(KeyArray_outS01ser_5_), 
        .B(KeyArray_S01reg_gff_1_SFF_5_QD), .S(n188), .Z(
        KeyArray_S01reg_gff_1_SFF_5_n6) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2010), 
        .B(new_AGEMA_signal_2893), .S(n188), .Z(new_AGEMA_signal_3280) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS01ser[5]), .B(KeyArray_outS11ser[5]), .S(n170), .Z(
        KeyArray_S01reg_gff_1_SFF_5_QD) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2459), .B(new_AGEMA_signal_2530), .S(n170), .Z(
        new_AGEMA_signal_2893) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_6_U1_Ins_0_U1 ( .A(KeyArray_outS01ser_6_), 
        .B(KeyArray_S01reg_gff_1_SFF_6_QD), .S(n188), .Z(
        KeyArray_S01reg_gff_1_SFF_6_n6) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2008), 
        .B(new_AGEMA_signal_2894), .S(n188), .Z(new_AGEMA_signal_3281) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS01ser[6]), .B(KeyArray_outS11ser[6]), .S(n169), .Z(
        KeyArray_S01reg_gff_1_SFF_6_QD) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2462), .B(new_AGEMA_signal_2533), .S(n169), .Z(
        new_AGEMA_signal_2894) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_7_U1_Ins_0_U1 ( .A(KeyArray_outS01ser_7_), 
        .B(KeyArray_S01reg_gff_1_SFF_7_QD), .S(n188), .Z(
        KeyArray_S01reg_gff_1_SFF_7_n6) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2006), 
        .B(new_AGEMA_signal_2895), .S(n188), .Z(new_AGEMA_signal_3282) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS01ser[7]), .B(KeyArray_outS11ser[7]), .S(n168), .Z(
        KeyArray_S01reg_gff_1_SFF_7_QD) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2465), .B(new_AGEMA_signal_2536), .S(n168), .Z(
        new_AGEMA_signal_2895) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_0_U1_Ins_0_U1 ( .A(KeyArray_outS02ser[0]), 
        .B(KeyArray_S02reg_gff_1_SFF_0_QD), .S(n187), .Z(
        KeyArray_S02reg_gff_1_SFF_0_n6) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_0_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2443), 
        .B(new_AGEMA_signal_2896), .S(n187), .Z(new_AGEMA_signal_3283) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS02ser[0]), .B(KeyArray_outS12ser[0]), .S(n172), .Z(
        KeyArray_S02reg_gff_1_SFF_0_QD) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2468), .B(new_AGEMA_signal_2539), .S(n172), .Z(
        new_AGEMA_signal_2896) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_1_U1_Ins_0_U1 ( .A(KeyArray_outS02ser[1]), 
        .B(KeyArray_S02reg_gff_1_SFF_1_QD), .S(n188), .Z(
        KeyArray_S02reg_gff_1_SFF_1_n6) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2446), 
        .B(new_AGEMA_signal_2897), .S(n188), .Z(new_AGEMA_signal_3284) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS02ser[1]), .B(KeyArray_outS12ser[1]), .S(n165), .Z(
        KeyArray_S02reg_gff_1_SFF_1_QD) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2471), .B(new_AGEMA_signal_2542), .S(n165), .Z(
        new_AGEMA_signal_2897) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_2_U1_Ins_0_U1 ( .A(KeyArray_outS02ser[2]), 
        .B(KeyArray_S02reg_gff_1_SFF_2_QD), .S(n187), .Z(
        KeyArray_S02reg_gff_1_SFF_2_n6) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2449), 
        .B(new_AGEMA_signal_2898), .S(n187), .Z(new_AGEMA_signal_3285) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS02ser[2]), .B(KeyArray_outS12ser[2]), .S(n164), .Z(
        KeyArray_S02reg_gff_1_SFF_2_QD) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2474), .B(new_AGEMA_signal_2545), .S(n164), .Z(
        new_AGEMA_signal_2898) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_3_U1_Ins_0_U1 ( .A(KeyArray_outS02ser[3]), 
        .B(KeyArray_S02reg_gff_1_SFF_3_QD), .S(n187), .Z(
        KeyArray_S02reg_gff_1_SFF_3_n6) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_3_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2452), 
        .B(new_AGEMA_signal_2899), .S(n187), .Z(new_AGEMA_signal_3286) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS02ser[3]), .B(KeyArray_outS12ser[3]), .S(n165), .Z(
        KeyArray_S02reg_gff_1_SFF_3_QD) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2477), .B(new_AGEMA_signal_2548), .S(n165), .Z(
        new_AGEMA_signal_2899) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_4_U1_Ins_0_U1 ( .A(KeyArray_outS02ser[4]), 
        .B(KeyArray_S02reg_gff_1_SFF_4_QD), .S(n187), .Z(
        KeyArray_S02reg_gff_1_SFF_4_n6) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2455), 
        .B(new_AGEMA_signal_2900), .S(n187), .Z(new_AGEMA_signal_3287) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS02ser[4]), .B(KeyArray_outS12ser[4]), .S(n166), .Z(
        KeyArray_S02reg_gff_1_SFF_4_QD) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2480), .B(new_AGEMA_signal_2551), .S(n166), .Z(
        new_AGEMA_signal_2900) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_5_U1_Ins_0_U1 ( .A(KeyArray_outS02ser[5]), 
        .B(KeyArray_S02reg_gff_1_SFF_5_QD), .S(n187), .Z(
        KeyArray_S02reg_gff_1_SFF_5_n6) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2458), 
        .B(new_AGEMA_signal_2901), .S(n187), .Z(new_AGEMA_signal_3288) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS02ser[5]), .B(KeyArray_outS12ser[5]), .S(n167), .Z(
        KeyArray_S02reg_gff_1_SFF_5_QD) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2483), .B(new_AGEMA_signal_2554), .S(n167), .Z(
        new_AGEMA_signal_2901) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_6_U1_Ins_0_U1 ( .A(KeyArray_outS02ser[6]), 
        .B(KeyArray_S02reg_gff_1_SFF_6_QD), .S(n187), .Z(
        KeyArray_S02reg_gff_1_SFF_6_n6) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2461), 
        .B(new_AGEMA_signal_2902), .S(n187), .Z(new_AGEMA_signal_3289) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS02ser[6]), .B(KeyArray_outS12ser[6]), .S(n171), .Z(
        KeyArray_S02reg_gff_1_SFF_6_QD) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2486), .B(new_AGEMA_signal_2557), .S(n171), .Z(
        new_AGEMA_signal_2902) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_7_U1_Ins_0_U1 ( .A(KeyArray_outS02ser[7]), 
        .B(KeyArray_S02reg_gff_1_SFF_7_QD), .S(n187), .Z(
        KeyArray_S02reg_gff_1_SFF_7_n6) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2464), 
        .B(new_AGEMA_signal_2903), .S(n187), .Z(new_AGEMA_signal_3290) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS02ser[7]), .B(KeyArray_outS12ser[7]), .S(n170), .Z(
        KeyArray_S02reg_gff_1_SFF_7_QD) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2489), .B(new_AGEMA_signal_2560), .S(n170), .Z(
        new_AGEMA_signal_2903) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_0_U1_Ins_0_U1 ( .A(KeyArray_outS03ser[0]), 
        .B(KeyArray_S03reg_gff_1_SFF_0_QD), .S(n185), .Z(
        KeyArray_S03reg_gff_1_SFF_0_n6) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_0_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2467), 
        .B(new_AGEMA_signal_2904), .S(n185), .Z(new_AGEMA_signal_3291) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS03ser[0]), .B(keySBIn[0]), .S(n169), .Z(
        KeyArray_S03reg_gff_1_SFF_0_QD) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2492), .B(new_AGEMA_signal_2563), .S(n169), .Z(
        new_AGEMA_signal_2904) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_1_U1_Ins_0_U1 ( .A(KeyArray_outS03ser[1]), 
        .B(KeyArray_S03reg_gff_1_SFF_1_QD), .S(n178), .Z(
        KeyArray_S03reg_gff_1_SFF_1_n6) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2470), 
        .B(new_AGEMA_signal_2905), .S(n178), .Z(new_AGEMA_signal_3292) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS03ser[1]), .B(keySBIn[1]), .S(n172), .Z(
        KeyArray_S03reg_gff_1_SFF_1_QD) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2495), .B(new_AGEMA_signal_2566), .S(n172), .Z(
        new_AGEMA_signal_2905) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_2_U1_Ins_0_U1 ( .A(KeyArray_outS03ser[2]), 
        .B(KeyArray_S03reg_gff_1_SFF_2_QD), .S(n187), .Z(
        KeyArray_S03reg_gff_1_SFF_2_n6) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2473), 
        .B(new_AGEMA_signal_2906), .S(n187), .Z(new_AGEMA_signal_3293) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS03ser[2]), .B(keySBIn[2]), .S(n168), .Z(
        KeyArray_S03reg_gff_1_SFF_2_QD) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2498), .B(new_AGEMA_signal_2569), .S(n168), .Z(
        new_AGEMA_signal_2906) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_3_U1_Ins_0_U1 ( .A(KeyArray_outS03ser[3]), 
        .B(KeyArray_S03reg_gff_1_SFF_3_QD), .S(n182), .Z(
        KeyArray_S03reg_gff_1_SFF_3_n6) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_3_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2476), 
        .B(new_AGEMA_signal_2907), .S(n182), .Z(new_AGEMA_signal_3294) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS03ser[3]), .B(keySBIn[3]), .S(n163), .Z(
        KeyArray_S03reg_gff_1_SFF_3_QD) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2501), .B(new_AGEMA_signal_2572), .S(n163), .Z(
        new_AGEMA_signal_2907) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_4_U1_Ins_0_U1 ( .A(KeyArray_outS03ser[4]), 
        .B(KeyArray_S03reg_gff_1_SFF_4_QD), .S(n186), .Z(
        KeyArray_S03reg_gff_1_SFF_4_n6) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2479), 
        .B(new_AGEMA_signal_2908), .S(n186), .Z(new_AGEMA_signal_3295) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS03ser[4]), .B(keySBIn[4]), .S(n166), .Z(
        KeyArray_S03reg_gff_1_SFF_4_QD) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2504), .B(new_AGEMA_signal_2575), .S(n166), .Z(
        new_AGEMA_signal_2908) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_5_U1_Ins_0_U1 ( .A(KeyArray_outS03ser[5]), 
        .B(KeyArray_S03reg_gff_1_SFF_5_QD), .S(n183), .Z(
        KeyArray_S03reg_gff_1_SFF_5_n5) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2482), 
        .B(new_AGEMA_signal_2909), .S(n183), .Z(new_AGEMA_signal_3296) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS03ser[5]), .B(keySBIn[5]), .S(n160), .Z(
        KeyArray_S03reg_gff_1_SFF_5_QD) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2507), .B(new_AGEMA_signal_2578), .S(n160), .Z(
        new_AGEMA_signal_2909) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_6_U1_Ins_0_U1 ( .A(KeyArray_outS03ser[6]), 
        .B(KeyArray_S03reg_gff_1_SFF_6_QD), .S(n179), .Z(
        KeyArray_S03reg_gff_1_SFF_6_n5) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2485), 
        .B(new_AGEMA_signal_2910), .S(n179), .Z(new_AGEMA_signal_3297) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS03ser[6]), .B(keySBIn[6]), .S(n164), .Z(
        KeyArray_S03reg_gff_1_SFF_6_QD) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2510), .B(new_AGEMA_signal_2581), .S(n164), .Z(
        new_AGEMA_signal_2910) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_7_U1_Ins_0_U1 ( .A(KeyArray_outS03ser[7]), 
        .B(KeyArray_S03reg_gff_1_SFF_7_QD), .S(n186), .Z(
        KeyArray_S03reg_gff_1_SFF_7_n5) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2488), 
        .B(new_AGEMA_signal_2911), .S(n186), .Z(new_AGEMA_signal_3298) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS03ser[7]), .B(keySBIn[7]), .S(n165), .Z(
        KeyArray_S03reg_gff_1_SFF_7_QD) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2513), .B(new_AGEMA_signal_2584), .S(n165), .Z(
        new_AGEMA_signal_2911) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_0_U1_Ins_0_U1 ( .A(KeyArray_outS10ser[0]), 
        .B(KeyArray_S10reg_gff_1_SFF_0_QD), .S(n186), .Z(
        KeyArray_S10reg_gff_1_SFF_0_n5) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_0_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2491), 
        .B(new_AGEMA_signal_2912), .S(n186), .Z(new_AGEMA_signal_3299) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS10ser[0]), .B(KeyArray_outS20ser[0]), .S(n166), .Z(
        KeyArray_S10reg_gff_1_SFF_0_QD) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2516), .B(new_AGEMA_signal_2587), .S(n166), .Z(
        new_AGEMA_signal_2912) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_1_U1_Ins_0_U1 ( .A(KeyArray_outS10ser[1]), 
        .B(KeyArray_S10reg_gff_1_SFF_1_QD), .S(n186), .Z(
        KeyArray_S10reg_gff_1_SFF_1_n5) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2494), 
        .B(new_AGEMA_signal_2913), .S(n186), .Z(new_AGEMA_signal_3300) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS10ser[1]), .B(KeyArray_outS20ser[1]), .S(n167), .Z(
        KeyArray_S10reg_gff_1_SFF_1_QD) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2519), .B(new_AGEMA_signal_2590), .S(n167), .Z(
        new_AGEMA_signal_2913) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_2_U1_Ins_0_U1 ( .A(KeyArray_outS10ser[2]), 
        .B(KeyArray_S10reg_gff_1_SFF_2_QD), .S(n186), .Z(
        KeyArray_S10reg_gff_1_SFF_2_n5) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2497), 
        .B(new_AGEMA_signal_2914), .S(n186), .Z(new_AGEMA_signal_3301) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS10ser[2]), .B(KeyArray_outS20ser[2]), .S(n171), .Z(
        KeyArray_S10reg_gff_1_SFF_2_QD) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2522), .B(new_AGEMA_signal_2593), .S(n171), .Z(
        new_AGEMA_signal_2914) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_3_U1_Ins_0_U1 ( .A(KeyArray_outS10ser[3]), 
        .B(KeyArray_S10reg_gff_1_SFF_3_QD), .S(n186), .Z(
        KeyArray_S10reg_gff_1_SFF_3_n5) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_3_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2500), 
        .B(new_AGEMA_signal_2915), .S(n186), .Z(new_AGEMA_signal_3302) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS10ser[3]), .B(KeyArray_outS20ser[3]), .S(n170), .Z(
        KeyArray_S10reg_gff_1_SFF_3_QD) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2525), .B(new_AGEMA_signal_2596), .S(n170), .Z(
        new_AGEMA_signal_2915) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_4_U1_Ins_0_U1 ( .A(KeyArray_outS10ser[4]), 
        .B(KeyArray_S10reg_gff_1_SFF_4_QD), .S(n186), .Z(
        KeyArray_S10reg_gff_1_SFF_4_n5) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2503), 
        .B(new_AGEMA_signal_2916), .S(n186), .Z(new_AGEMA_signal_3303) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS10ser[4]), .B(KeyArray_outS20ser[4]), .S(n169), .Z(
        KeyArray_S10reg_gff_1_SFF_4_QD) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2528), .B(new_AGEMA_signal_2599), .S(n169), .Z(
        new_AGEMA_signal_2916) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_5_U1_Ins_0_U1 ( .A(KeyArray_outS10ser[5]), 
        .B(KeyArray_S10reg_gff_1_SFF_5_QD), .S(n186), .Z(
        KeyArray_S10reg_gff_1_SFF_5_n5) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2506), 
        .B(new_AGEMA_signal_2917), .S(n186), .Z(new_AGEMA_signal_3304) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS10ser[5]), .B(KeyArray_outS20ser[5]), .S(n168), .Z(
        KeyArray_S10reg_gff_1_SFF_5_QD) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2531), .B(new_AGEMA_signal_2602), .S(n168), .Z(
        new_AGEMA_signal_2917) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_6_U1_Ins_0_U1 ( .A(KeyArray_outS10ser[6]), 
        .B(KeyArray_S10reg_gff_1_SFF_6_QD), .S(n185), .Z(
        KeyArray_S10reg_gff_1_SFF_6_n5) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2509), 
        .B(new_AGEMA_signal_2918), .S(n185), .Z(new_AGEMA_signal_3305) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS10ser[6]), .B(KeyArray_outS20ser[6]), .S(n172), .Z(
        KeyArray_S10reg_gff_1_SFF_6_QD) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2534), .B(new_AGEMA_signal_2605), .S(n172), .Z(
        new_AGEMA_signal_2918) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_7_U1_Ins_0_U1 ( .A(KeyArray_outS10ser[7]), 
        .B(KeyArray_S10reg_gff_1_SFF_7_QD), .S(n185), .Z(
        KeyArray_S10reg_gff_1_SFF_7_n5) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2512), 
        .B(new_AGEMA_signal_2919), .S(n185), .Z(new_AGEMA_signal_3306) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS10ser[7]), .B(KeyArray_outS20ser[7]), .S(n174), .Z(
        KeyArray_S10reg_gff_1_SFF_7_QD) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2537), .B(new_AGEMA_signal_2608), .S(n174), .Z(
        new_AGEMA_signal_2919) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_0_U1_Ins_0_U1 ( .A(KeyArray_outS11ser[0]), 
        .B(KeyArray_S11reg_gff_1_SFF_0_QD), .S(n185), .Z(
        KeyArray_S11reg_gff_1_SFF_0_n6) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_0_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2515), 
        .B(new_AGEMA_signal_2920), .S(n185), .Z(new_AGEMA_signal_3307) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS11ser[0]), .B(KeyArray_outS21ser[0]), .S(n173), .Z(
        KeyArray_S11reg_gff_1_SFF_0_QD) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2540), .B(new_AGEMA_signal_2611), .S(n173), .Z(
        new_AGEMA_signal_2920) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_1_U1_Ins_0_U1 ( .A(KeyArray_outS11ser[1]), 
        .B(KeyArray_S11reg_gff_1_SFF_1_QD), .S(n185), .Z(
        KeyArray_S11reg_gff_1_SFF_1_n6) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2518), 
        .B(new_AGEMA_signal_2921), .S(n185), .Z(new_AGEMA_signal_3308) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS11ser[1]), .B(KeyArray_outS21ser[1]), .S(n173), .Z(
        KeyArray_S11reg_gff_1_SFF_1_QD) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2543), .B(new_AGEMA_signal_2614), .S(n173), .Z(
        new_AGEMA_signal_2921) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_2_U1_Ins_0_U1 ( .A(KeyArray_outS11ser[2]), 
        .B(KeyArray_S11reg_gff_1_SFF_2_QD), .S(n185), .Z(
        KeyArray_S11reg_gff_1_SFF_2_n6) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2521), 
        .B(new_AGEMA_signal_2922), .S(n185), .Z(new_AGEMA_signal_3309) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS11ser[2]), .B(KeyArray_outS21ser[2]), .S(n173), .Z(
        KeyArray_S11reg_gff_1_SFF_2_QD) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2546), .B(new_AGEMA_signal_2617), .S(n173), .Z(
        new_AGEMA_signal_2922) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_3_U1_Ins_0_U1 ( .A(KeyArray_outS11ser[3]), 
        .B(KeyArray_S11reg_gff_1_SFF_3_QD), .S(n185), .Z(
        KeyArray_S11reg_gff_1_SFF_3_n6) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_3_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2524), 
        .B(new_AGEMA_signal_2923), .S(n185), .Z(new_AGEMA_signal_3310) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS11ser[3]), .B(KeyArray_outS21ser[3]), .S(n175), .Z(
        KeyArray_S11reg_gff_1_SFF_3_QD) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2549), .B(new_AGEMA_signal_2620), .S(n175), .Z(
        new_AGEMA_signal_2923) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_4_U1_Ins_0_U1 ( .A(KeyArray_outS11ser[4]), 
        .B(KeyArray_S11reg_gff_1_SFF_4_QD), .S(n185), .Z(
        KeyArray_S11reg_gff_1_SFF_4_n6) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2527), 
        .B(new_AGEMA_signal_2924), .S(n185), .Z(new_AGEMA_signal_3311) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS11ser[4]), .B(KeyArray_outS21ser[4]), .S(n162), .Z(
        KeyArray_S11reg_gff_1_SFF_4_QD) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2552), .B(new_AGEMA_signal_2623), .S(n162), .Z(
        new_AGEMA_signal_2924) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_5_U1_Ins_0_U1 ( .A(KeyArray_outS11ser[5]), 
        .B(KeyArray_S11reg_gff_1_SFF_5_QD), .S(n184), .Z(
        KeyArray_S11reg_gff_1_SFF_5_n6) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2530), 
        .B(new_AGEMA_signal_2925), .S(n184), .Z(new_AGEMA_signal_3312) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS11ser[5]), .B(KeyArray_outS21ser[5]), .S(n160), .Z(
        KeyArray_S11reg_gff_1_SFF_5_QD) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2555), .B(new_AGEMA_signal_2626), .S(n160), .Z(
        new_AGEMA_signal_2925) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_6_U1_Ins_0_U1 ( .A(KeyArray_outS11ser[6]), 
        .B(KeyArray_S11reg_gff_1_SFF_6_QD), .S(n184), .Z(
        KeyArray_S11reg_gff_1_SFF_6_n6) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2533), 
        .B(new_AGEMA_signal_2926), .S(n184), .Z(new_AGEMA_signal_3313) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS11ser[6]), .B(KeyArray_outS21ser[6]), .S(n164), .Z(
        KeyArray_S11reg_gff_1_SFF_6_QD) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2558), .B(new_AGEMA_signal_2629), .S(n164), .Z(
        new_AGEMA_signal_2926) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_7_U1_Ins_0_U1 ( .A(KeyArray_outS11ser[7]), 
        .B(KeyArray_S11reg_gff_1_SFF_7_QD), .S(n184), .Z(
        KeyArray_S11reg_gff_1_SFF_7_n6) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2536), 
        .B(new_AGEMA_signal_2927), .S(n184), .Z(new_AGEMA_signal_3314) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS11ser[7]), .B(KeyArray_outS21ser[7]), .S(n164), .Z(
        KeyArray_S11reg_gff_1_SFF_7_QD) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2561), .B(new_AGEMA_signal_2632), .S(n164), .Z(
        new_AGEMA_signal_2927) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_0_U1_Ins_0_U1 ( .A(KeyArray_outS12ser[0]), 
        .B(KeyArray_S12reg_gff_1_SFF_0_QD), .S(n184), .Z(
        KeyArray_S12reg_gff_1_SFF_0_n6) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_0_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2539), 
        .B(new_AGEMA_signal_2928), .S(n184), .Z(new_AGEMA_signal_3093) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS12ser[0]), .B(KeyArray_outS22ser[0]), .S(n164), .Z(
        KeyArray_S12reg_gff_1_SFF_0_QD) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2564), .B(new_AGEMA_signal_2635), .S(n164), .Z(
        new_AGEMA_signal_2928) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_1_U1_Ins_0_U1 ( .A(KeyArray_outS12ser[1]), 
        .B(KeyArray_S12reg_gff_1_SFF_1_QD), .S(n184), .Z(
        KeyArray_S12reg_gff_1_SFF_1_n6) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2542), 
        .B(new_AGEMA_signal_2929), .S(n184), .Z(new_AGEMA_signal_3094) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS12ser[1]), .B(KeyArray_outS22ser[1]), .S(n164), .Z(
        KeyArray_S12reg_gff_1_SFF_1_QD) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2567), .B(new_AGEMA_signal_2638), .S(n164), .Z(
        new_AGEMA_signal_2929) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_2_U1_Ins_0_U1 ( .A(KeyArray_outS12ser[2]), 
        .B(KeyArray_S12reg_gff_1_SFF_2_QD), .S(n184), .Z(
        KeyArray_S12reg_gff_1_SFF_2_n6) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2545), 
        .B(new_AGEMA_signal_2930), .S(n184), .Z(new_AGEMA_signal_3095) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS12ser[2]), .B(KeyArray_outS22ser[2]), .S(n164), .Z(
        KeyArray_S12reg_gff_1_SFF_2_QD) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2570), .B(new_AGEMA_signal_2641), .S(n164), .Z(
        new_AGEMA_signal_2930) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_3_U1_Ins_0_U1 ( .A(KeyArray_outS12ser[3]), 
        .B(KeyArray_S12reg_gff_1_SFF_3_QD), .S(n184), .Z(
        KeyArray_S12reg_gff_1_SFF_3_n6) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_3_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2548), 
        .B(new_AGEMA_signal_2931), .S(n184), .Z(new_AGEMA_signal_3096) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS12ser[3]), .B(KeyArray_outS22ser[3]), .S(n164), .Z(
        KeyArray_S12reg_gff_1_SFF_3_QD) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2573), .B(new_AGEMA_signal_2644), .S(n164), .Z(
        new_AGEMA_signal_2931) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_4_U1_Ins_0_U1 ( .A(KeyArray_outS12ser[4]), 
        .B(KeyArray_S12reg_gff_1_SFF_4_QD), .S(n188), .Z(
        KeyArray_S12reg_gff_1_SFF_4_n6) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2551), 
        .B(new_AGEMA_signal_2932), .S(n188), .Z(new_AGEMA_signal_3097) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS12ser[4]), .B(KeyArray_outS22ser[4]), .S(n164), .Z(
        KeyArray_S12reg_gff_1_SFF_4_QD) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2576), .B(new_AGEMA_signal_2647), .S(n164), .Z(
        new_AGEMA_signal_2932) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_5_U1_Ins_0_U1 ( .A(KeyArray_outS12ser[5]), 
        .B(KeyArray_S12reg_gff_1_SFF_5_QD), .S(n181), .Z(
        KeyArray_S12reg_gff_1_SFF_5_n6) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2554), 
        .B(new_AGEMA_signal_2933), .S(n181), .Z(new_AGEMA_signal_3098) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS12ser[5]), .B(KeyArray_outS22ser[5]), .S(n165), .Z(
        KeyArray_S12reg_gff_1_SFF_5_QD) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2579), .B(new_AGEMA_signal_2650), .S(n165), .Z(
        new_AGEMA_signal_2933) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_6_U1_Ins_0_U1 ( .A(KeyArray_outS12ser[6]), 
        .B(KeyArray_S12reg_gff_1_SFF_6_QD), .S(n189), .Z(
        KeyArray_S12reg_gff_1_SFF_6_n6) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2557), 
        .B(new_AGEMA_signal_2934), .S(n189), .Z(new_AGEMA_signal_3099) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS12ser[6]), .B(KeyArray_outS22ser[6]), .S(n165), .Z(
        KeyArray_S12reg_gff_1_SFF_6_QD) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2582), .B(new_AGEMA_signal_2653), .S(n165), .Z(
        new_AGEMA_signal_2934) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_7_U1_Ins_0_U1 ( .A(KeyArray_outS12ser[7]), 
        .B(KeyArray_S12reg_gff_1_SFF_7_QD), .S(n184), .Z(
        KeyArray_S12reg_gff_1_SFF_7_n6) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2560), 
        .B(new_AGEMA_signal_2935), .S(n184), .Z(new_AGEMA_signal_3100) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS12ser[7]), .B(KeyArray_outS22ser[7]), .S(n165), .Z(
        KeyArray_S12reg_gff_1_SFF_7_QD) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2585), .B(new_AGEMA_signal_2656), .S(n165), .Z(
        new_AGEMA_signal_2935) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_0_U1_Ins_0_U1 ( .A(keySBIn[0]), .B(
        KeyArray_S13reg_gff_1_SFF_0_QD), .S(n180), .Z(
        KeyArray_S13reg_gff_1_SFF_0_n6) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_0_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2563), 
        .B(new_AGEMA_signal_2936), .S(n180), .Z(new_AGEMA_signal_3101) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS13ser[0]), .B(KeyArray_outS23ser[0]), .S(n165), .Z(
        KeyArray_S13reg_gff_1_SFF_0_QD) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2588), .B(new_AGEMA_signal_2659), .S(n165), .Z(
        new_AGEMA_signal_2936) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_1_U1_Ins_0_U1 ( .A(keySBIn[1]), .B(
        KeyArray_S13reg_gff_1_SFF_1_QD), .S(n182), .Z(
        KeyArray_S13reg_gff_1_SFF_1_n6) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2566), 
        .B(new_AGEMA_signal_2937), .S(n182), .Z(new_AGEMA_signal_3102) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS13ser[1]), .B(KeyArray_outS23ser[1]), .S(n165), .Z(
        KeyArray_S13reg_gff_1_SFF_1_QD) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2591), .B(new_AGEMA_signal_2662), .S(n165), .Z(
        new_AGEMA_signal_2937) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_2_U1_Ins_0_U1 ( .A(keySBIn[2]), .B(
        KeyArray_S13reg_gff_1_SFF_2_QD), .S(n188), .Z(
        KeyArray_S13reg_gff_1_SFF_2_n6) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2569), 
        .B(new_AGEMA_signal_2938), .S(n188), .Z(new_AGEMA_signal_3103) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS13ser[2]), .B(KeyArray_outS23ser[2]), .S(n165), .Z(
        KeyArray_S13reg_gff_1_SFF_2_QD) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2594), .B(new_AGEMA_signal_2665), .S(n165), .Z(
        new_AGEMA_signal_2938) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_3_U1_Ins_0_U1 ( .A(keySBIn[3]), .B(
        KeyArray_S13reg_gff_1_SFF_3_QD), .S(n183), .Z(
        KeyArray_S13reg_gff_1_SFF_3_n6) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_3_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2572), 
        .B(new_AGEMA_signal_2939), .S(n183), .Z(new_AGEMA_signal_3104) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS13ser[3]), .B(KeyArray_outS23ser[3]), .S(n165), .Z(
        KeyArray_S13reg_gff_1_SFF_3_QD) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2597), .B(new_AGEMA_signal_2668), .S(n165), .Z(
        new_AGEMA_signal_2939) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_4_U1_Ins_0_U1 ( .A(keySBIn[4]), .B(
        KeyArray_S13reg_gff_1_SFF_4_QD), .S(n183), .Z(
        KeyArray_S13reg_gff_1_SFF_4_n6) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2575), 
        .B(new_AGEMA_signal_2940), .S(n183), .Z(new_AGEMA_signal_3105) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS13ser[4]), .B(KeyArray_outS23ser[4]), .S(n166), .Z(
        KeyArray_S13reg_gff_1_SFF_4_QD) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2600), .B(new_AGEMA_signal_2671), .S(n166), .Z(
        new_AGEMA_signal_2940) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_5_U1_Ins_0_U1 ( .A(keySBIn[5]), .B(
        KeyArray_S13reg_gff_1_SFF_5_QD), .S(n183), .Z(
        KeyArray_S13reg_gff_1_SFF_5_n5) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2578), 
        .B(new_AGEMA_signal_2941), .S(n183), .Z(new_AGEMA_signal_3106) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS13ser[5]), .B(KeyArray_outS23ser[5]), .S(n166), .Z(
        KeyArray_S13reg_gff_1_SFF_5_QD) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2603), .B(new_AGEMA_signal_2674), .S(n166), .Z(
        new_AGEMA_signal_2941) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_6_U1_Ins_0_U1 ( .A(keySBIn[6]), .B(
        KeyArray_S13reg_gff_1_SFF_6_QD), .S(n183), .Z(
        KeyArray_S13reg_gff_1_SFF_6_n5) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2581), 
        .B(new_AGEMA_signal_2942), .S(n183), .Z(new_AGEMA_signal_3107) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS13ser[6]), .B(KeyArray_outS23ser[6]), .S(n166), .Z(
        KeyArray_S13reg_gff_1_SFF_6_QD) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2606), .B(new_AGEMA_signal_2677), .S(n166), .Z(
        new_AGEMA_signal_2942) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_7_U1_Ins_0_U1 ( .A(keySBIn[7]), .B(
        KeyArray_S13reg_gff_1_SFF_7_QD), .S(n183), .Z(
        KeyArray_S13reg_gff_1_SFF_7_n5) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2584), 
        .B(new_AGEMA_signal_2943), .S(n183), .Z(new_AGEMA_signal_3108) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS13ser[7]), .B(KeyArray_outS23ser[7]), .S(n166), .Z(
        KeyArray_S13reg_gff_1_SFF_7_QD) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2609), .B(new_AGEMA_signal_2680), .S(n166), .Z(
        new_AGEMA_signal_2943) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_0_U1_Ins_0_U1 ( .A(KeyArray_outS20ser[0]), 
        .B(KeyArray_S20reg_gff_1_SFF_0_QD), .S(n183), .Z(
        KeyArray_S20reg_gff_1_SFF_0_n5) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_0_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2587), 
        .B(new_AGEMA_signal_2944), .S(n183), .Z(new_AGEMA_signal_3315) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS20ser[0]), .B(KeyArray_outS30ser[0]), .S(n166), .Z(
        KeyArray_S20reg_gff_1_SFF_0_QD) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2612), .B(new_AGEMA_signal_2683), .S(n166), .Z(
        new_AGEMA_signal_2944) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_1_U1_Ins_0_U1 ( .A(KeyArray_outS20ser[1]), 
        .B(KeyArray_S20reg_gff_1_SFF_1_QD), .S(n182), .Z(
        KeyArray_S20reg_gff_1_SFF_1_n5) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2590), 
        .B(new_AGEMA_signal_2945), .S(n182), .Z(new_AGEMA_signal_3316) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS20ser[1]), .B(KeyArray_outS30ser[1]), .S(n166), .Z(
        KeyArray_S20reg_gff_1_SFF_1_QD) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2615), .B(new_AGEMA_signal_2686), .S(n166), .Z(
        new_AGEMA_signal_2945) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_2_U1_Ins_0_U1 ( .A(KeyArray_outS20ser[2]), 
        .B(KeyArray_S20reg_gff_1_SFF_2_QD), .S(n182), .Z(
        KeyArray_S20reg_gff_1_SFF_2_n5) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2593), 
        .B(new_AGEMA_signal_2946), .S(n182), .Z(new_AGEMA_signal_3317) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS20ser[2]), .B(KeyArray_outS30ser[2]), .S(n166), .Z(
        KeyArray_S20reg_gff_1_SFF_2_QD) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2618), .B(new_AGEMA_signal_2689), .S(n166), .Z(
        new_AGEMA_signal_2946) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_3_U1_Ins_0_U1 ( .A(KeyArray_outS20ser[3]), 
        .B(KeyArray_S20reg_gff_1_SFF_3_QD), .S(n182), .Z(
        KeyArray_S20reg_gff_1_SFF_3_n5) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_3_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2596), 
        .B(new_AGEMA_signal_2947), .S(n182), .Z(new_AGEMA_signal_3318) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS20ser[3]), .B(KeyArray_outS30ser[3]), .S(n167), .Z(
        KeyArray_S20reg_gff_1_SFF_3_QD) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2621), .B(new_AGEMA_signal_2692), .S(n167), .Z(
        new_AGEMA_signal_2947) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_4_U1_Ins_0_U1 ( .A(KeyArray_outS20ser[4]), 
        .B(KeyArray_S20reg_gff_1_SFF_4_QD), .S(n182), .Z(
        KeyArray_S20reg_gff_1_SFF_4_n5) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2599), 
        .B(new_AGEMA_signal_2948), .S(n182), .Z(new_AGEMA_signal_3319) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS20ser[4]), .B(KeyArray_outS30ser[4]), .S(n167), .Z(
        KeyArray_S20reg_gff_1_SFF_4_QD) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2624), .B(new_AGEMA_signal_2695), .S(n167), .Z(
        new_AGEMA_signal_2948) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_5_U1_Ins_0_U1 ( .A(KeyArray_outS20ser[5]), 
        .B(KeyArray_S20reg_gff_1_SFF_5_QD), .S(n182), .Z(
        KeyArray_S20reg_gff_1_SFF_5_n5) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2602), 
        .B(new_AGEMA_signal_2949), .S(n182), .Z(new_AGEMA_signal_3320) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS20ser[5]), .B(KeyArray_outS30ser[5]), .S(n167), .Z(
        KeyArray_S20reg_gff_1_SFF_5_QD) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2627), .B(new_AGEMA_signal_2698), .S(n167), .Z(
        new_AGEMA_signal_2949) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_6_U1_Ins_0_U1 ( .A(KeyArray_outS20ser[6]), 
        .B(KeyArray_S20reg_gff_1_SFF_6_QD), .S(n182), .Z(
        KeyArray_S20reg_gff_1_SFF_6_n5) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2605), 
        .B(new_AGEMA_signal_2950), .S(n182), .Z(new_AGEMA_signal_3321) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS20ser[6]), .B(KeyArray_outS30ser[6]), .S(n167), .Z(
        KeyArray_S20reg_gff_1_SFF_6_QD) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2630), .B(new_AGEMA_signal_2701), .S(n167), .Z(
        new_AGEMA_signal_2950) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_7_U1_Ins_0_U1 ( .A(KeyArray_outS20ser[7]), 
        .B(KeyArray_S20reg_gff_1_SFF_7_QD), .S(n182), .Z(
        KeyArray_S20reg_gff_1_SFF_7_n5) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2608), 
        .B(new_AGEMA_signal_2951), .S(n182), .Z(new_AGEMA_signal_3322) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS20ser[7]), .B(KeyArray_outS30ser[7]), .S(n167), .Z(
        KeyArray_S20reg_gff_1_SFF_7_QD) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2633), .B(new_AGEMA_signal_2704), .S(n167), .Z(
        new_AGEMA_signal_2951) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_0_U1_Ins_0_U1 ( .A(KeyArray_outS21ser[0]), 
        .B(KeyArray_S21reg_gff_1_SFF_0_QD), .S(n181), .Z(
        KeyArray_S21reg_gff_1_SFF_0_n6) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_0_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2611), 
        .B(new_AGEMA_signal_2952), .S(n181), .Z(new_AGEMA_signal_3323) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS21ser[0]), .B(KeyArray_outS31ser[0]), .S(n167), .Z(
        KeyArray_S21reg_gff_1_SFF_0_QD) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2636), .B(new_AGEMA_signal_2707), .S(n167), .Z(
        new_AGEMA_signal_2952) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_1_U1_Ins_0_U1 ( .A(KeyArray_outS21ser[1]), 
        .B(KeyArray_S21reg_gff_1_SFF_1_QD), .S(n181), .Z(
        KeyArray_S21reg_gff_1_SFF_1_n6) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2614), 
        .B(new_AGEMA_signal_2953), .S(n181), .Z(new_AGEMA_signal_3324) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS21ser[1]), .B(KeyArray_outS31ser[1]), .S(n167), .Z(
        KeyArray_S21reg_gff_1_SFF_1_QD) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2639), .B(new_AGEMA_signal_2710), .S(n167), .Z(
        new_AGEMA_signal_2953) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_2_U1_Ins_0_U1 ( .A(KeyArray_outS21ser[2]), 
        .B(KeyArray_S21reg_gff_1_SFF_2_QD), .S(n181), .Z(
        KeyArray_S21reg_gff_1_SFF_2_n6) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2617), 
        .B(new_AGEMA_signal_2954), .S(n181), .Z(new_AGEMA_signal_3325) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS21ser[2]), .B(KeyArray_outS31ser[2]), .S(n168), .Z(
        KeyArray_S21reg_gff_1_SFF_2_QD) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2642), .B(new_AGEMA_signal_2713), .S(n168), .Z(
        new_AGEMA_signal_2954) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_3_U1_Ins_0_U1 ( .A(KeyArray_outS21ser[3]), 
        .B(KeyArray_S21reg_gff_1_SFF_3_QD), .S(n181), .Z(
        KeyArray_S21reg_gff_1_SFF_3_n6) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_3_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2620), 
        .B(new_AGEMA_signal_2955), .S(n181), .Z(new_AGEMA_signal_3326) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS21ser[3]), .B(KeyArray_outS31ser[3]), .S(n168), .Z(
        KeyArray_S21reg_gff_1_SFF_3_QD) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2645), .B(new_AGEMA_signal_2716), .S(n168), .Z(
        new_AGEMA_signal_2955) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_4_U1_Ins_0_U1 ( .A(KeyArray_outS21ser[4]), 
        .B(KeyArray_S21reg_gff_1_SFF_4_QD), .S(n181), .Z(
        KeyArray_S21reg_gff_1_SFF_4_n6) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2623), 
        .B(new_AGEMA_signal_2956), .S(n181), .Z(new_AGEMA_signal_3327) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS21ser[4]), .B(KeyArray_outS31ser[4]), .S(n168), .Z(
        KeyArray_S21reg_gff_1_SFF_4_QD) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2648), .B(new_AGEMA_signal_2719), .S(n168), .Z(
        new_AGEMA_signal_2956) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_5_U1_Ins_0_U1 ( .A(KeyArray_outS21ser[5]), 
        .B(KeyArray_S21reg_gff_1_SFF_5_QD), .S(n181), .Z(
        KeyArray_S21reg_gff_1_SFF_5_n6) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2626), 
        .B(new_AGEMA_signal_2957), .S(n181), .Z(new_AGEMA_signal_3328) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS21ser[5]), .B(KeyArray_outS31ser[5]), .S(n168), .Z(
        KeyArray_S21reg_gff_1_SFF_5_QD) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2651), .B(new_AGEMA_signal_2722), .S(n168), .Z(
        new_AGEMA_signal_2957) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_6_U1_Ins_0_U1 ( .A(KeyArray_outS21ser[6]), 
        .B(KeyArray_S21reg_gff_1_SFF_6_QD), .S(n181), .Z(
        KeyArray_S21reg_gff_1_SFF_6_n6) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2629), 
        .B(new_AGEMA_signal_2958), .S(n181), .Z(new_AGEMA_signal_3329) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS21ser[6]), .B(KeyArray_outS31ser[6]), .S(n168), .Z(
        KeyArray_S21reg_gff_1_SFF_6_QD) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2654), .B(new_AGEMA_signal_2725), .S(n168), .Z(
        new_AGEMA_signal_2958) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_7_U1_Ins_0_U1 ( .A(KeyArray_outS21ser[7]), 
        .B(KeyArray_S21reg_gff_1_SFF_7_QD), .S(n180), .Z(
        KeyArray_S21reg_gff_1_SFF_7_n6) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2632), 
        .B(new_AGEMA_signal_2959), .S(n180), .Z(new_AGEMA_signal_3330) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS21ser[7]), .B(KeyArray_outS31ser[7]), .S(n168), .Z(
        KeyArray_S21reg_gff_1_SFF_7_QD) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2657), .B(new_AGEMA_signal_2728), .S(n168), .Z(
        new_AGEMA_signal_2959) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_0_U1_Ins_0_U1 ( .A(KeyArray_outS22ser[0]), 
        .B(KeyArray_S22reg_gff_1_SFF_0_QD), .S(n180), .Z(
        KeyArray_S22reg_gff_1_SFF_0_n6) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_0_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2635), 
        .B(new_AGEMA_signal_2960), .S(n180), .Z(new_AGEMA_signal_3331) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS22ser[0]), .B(KeyArray_outS32ser[0]), .S(n168), .Z(
        KeyArray_S22reg_gff_1_SFF_0_QD) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2660), .B(new_AGEMA_signal_2731), .S(n168), .Z(
        new_AGEMA_signal_2960) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_1_U1_Ins_0_U1 ( .A(KeyArray_outS22ser[1]), 
        .B(KeyArray_S22reg_gff_1_SFF_1_QD), .S(n180), .Z(
        KeyArray_S22reg_gff_1_SFF_1_n6) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2638), 
        .B(new_AGEMA_signal_2961), .S(n180), .Z(new_AGEMA_signal_3332) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS22ser[1]), .B(KeyArray_outS32ser[1]), .S(n169), .Z(
        KeyArray_S22reg_gff_1_SFF_1_QD) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2663), .B(new_AGEMA_signal_2734), .S(n169), .Z(
        new_AGEMA_signal_2961) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_2_U1_Ins_0_U1 ( .A(KeyArray_outS22ser[2]), 
        .B(KeyArray_S22reg_gff_1_SFF_2_QD), .S(n180), .Z(
        KeyArray_S22reg_gff_1_SFF_2_n6) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2641), 
        .B(new_AGEMA_signal_2962), .S(n180), .Z(new_AGEMA_signal_3333) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS22ser[2]), .B(KeyArray_outS32ser[2]), .S(n169), .Z(
        KeyArray_S22reg_gff_1_SFF_2_QD) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2666), .B(new_AGEMA_signal_2737), .S(n169), .Z(
        new_AGEMA_signal_2962) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_3_U1_Ins_0_U1 ( .A(KeyArray_outS22ser[3]), 
        .B(KeyArray_S22reg_gff_1_SFF_3_QD), .S(n180), .Z(
        KeyArray_S22reg_gff_1_SFF_3_n6) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_3_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2644), 
        .B(new_AGEMA_signal_2963), .S(n180), .Z(new_AGEMA_signal_3334) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS22ser[3]), .B(KeyArray_outS32ser[3]), .S(n169), .Z(
        KeyArray_S22reg_gff_1_SFF_3_QD) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2669), .B(new_AGEMA_signal_2740), .S(n169), .Z(
        new_AGEMA_signal_2963) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_4_U1_Ins_0_U1 ( .A(KeyArray_outS22ser[4]), 
        .B(KeyArray_S22reg_gff_1_SFF_4_QD), .S(n180), .Z(
        KeyArray_S22reg_gff_1_SFF_4_n6) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2647), 
        .B(new_AGEMA_signal_2964), .S(n180), .Z(new_AGEMA_signal_3335) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS22ser[4]), .B(KeyArray_outS32ser[4]), .S(n169), .Z(
        KeyArray_S22reg_gff_1_SFF_4_QD) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2672), .B(new_AGEMA_signal_2743), .S(n169), .Z(
        new_AGEMA_signal_2964) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_5_U1_Ins_0_U1 ( .A(KeyArray_outS22ser[5]), 
        .B(KeyArray_S22reg_gff_1_SFF_5_QD), .S(n180), .Z(
        KeyArray_S22reg_gff_1_SFF_5_n6) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2650), 
        .B(new_AGEMA_signal_2965), .S(n180), .Z(new_AGEMA_signal_3336) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS22ser[5]), .B(KeyArray_outS32ser[5]), .S(n169), .Z(
        KeyArray_S22reg_gff_1_SFF_5_QD) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2675), .B(new_AGEMA_signal_2746), .S(n169), .Z(
        new_AGEMA_signal_2965) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_6_U1_Ins_0_U1 ( .A(KeyArray_outS22ser[6]), 
        .B(KeyArray_S22reg_gff_1_SFF_6_QD), .S(n177), .Z(
        KeyArray_S22reg_gff_1_SFF_6_n6) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2653), 
        .B(new_AGEMA_signal_2966), .S(n177), .Z(new_AGEMA_signal_3337) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS22ser[6]), .B(KeyArray_outS32ser[6]), .S(n169), .Z(
        KeyArray_S22reg_gff_1_SFF_6_QD) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2678), .B(new_AGEMA_signal_2749), .S(n169), .Z(
        new_AGEMA_signal_2966) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_7_U1_Ins_0_U1 ( .A(KeyArray_outS22ser[7]), 
        .B(KeyArray_S22reg_gff_1_SFF_7_QD), .S(n181), .Z(
        KeyArray_S22reg_gff_1_SFF_7_n6) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2656), 
        .B(new_AGEMA_signal_2967), .S(n181), .Z(new_AGEMA_signal_3338) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS22ser[7]), .B(KeyArray_outS32ser[7]), .S(n169), .Z(
        KeyArray_S22reg_gff_1_SFF_7_QD) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2681), .B(new_AGEMA_signal_2752), .S(n169), .Z(
        new_AGEMA_signal_2967) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_0_U1_Ins_0_U1 ( .A(KeyArray_outS23ser[0]), 
        .B(KeyArray_S23reg_gff_1_SFF_0_QD), .S(n189), .Z(
        KeyArray_S23reg_gff_1_SFF_0_n6) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_0_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2659), 
        .B(new_AGEMA_signal_2968), .S(n189), .Z(new_AGEMA_signal_3339) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS23ser[0]), .B(KeyArray_outS33ser[0]), .S(n170), .Z(
        KeyArray_S23reg_gff_1_SFF_0_QD) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2684), .B(new_AGEMA_signal_2755), .S(n170), .Z(
        new_AGEMA_signal_2968) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_1_U1_Ins_0_U1 ( .A(KeyArray_outS23ser[1]), 
        .B(KeyArray_S23reg_gff_1_SFF_1_QD), .S(n184), .Z(
        KeyArray_S23reg_gff_1_SFF_1_n6) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2662), 
        .B(new_AGEMA_signal_2969), .S(n184), .Z(new_AGEMA_signal_3340) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS23ser[1]), .B(KeyArray_outS33ser[1]), .S(n170), .Z(
        KeyArray_S23reg_gff_1_SFF_1_QD) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2687), .B(new_AGEMA_signal_2758), .S(n170), .Z(
        new_AGEMA_signal_2969) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_2_U1_Ins_0_U1 ( .A(KeyArray_outS23ser[2]), 
        .B(KeyArray_S23reg_gff_1_SFF_2_QD), .S(n180), .Z(
        KeyArray_S23reg_gff_1_SFF_2_n6) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2665), 
        .B(new_AGEMA_signal_2970), .S(n180), .Z(new_AGEMA_signal_3341) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS23ser[2]), .B(KeyArray_outS33ser[2]), .S(n170), .Z(
        KeyArray_S23reg_gff_1_SFF_2_QD) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2690), .B(new_AGEMA_signal_2761), .S(n170), .Z(
        new_AGEMA_signal_2970) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_3_U1_Ins_0_U1 ( .A(KeyArray_outS23ser[3]), 
        .B(KeyArray_S23reg_gff_1_SFF_3_QD), .S(n178), .Z(
        KeyArray_S23reg_gff_1_SFF_3_n6) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_3_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2668), 
        .B(new_AGEMA_signal_2971), .S(n178), .Z(new_AGEMA_signal_3342) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS23ser[3]), .B(KeyArray_outS33ser[3]), .S(n170), .Z(
        KeyArray_S23reg_gff_1_SFF_3_QD) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2693), .B(new_AGEMA_signal_2764), .S(n170), .Z(
        new_AGEMA_signal_2971) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_4_U1_Ins_0_U1 ( .A(KeyArray_outS23ser[4]), 
        .B(KeyArray_S23reg_gff_1_SFF_4_QD), .S(n185), .Z(
        KeyArray_S23reg_gff_1_SFF_4_n6) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2671), 
        .B(new_AGEMA_signal_2972), .S(n185), .Z(new_AGEMA_signal_3343) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS23ser[4]), .B(KeyArray_outS33ser[4]), .S(n170), .Z(
        KeyArray_S23reg_gff_1_SFF_4_QD) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2696), .B(new_AGEMA_signal_2767), .S(n170), .Z(
        new_AGEMA_signal_2972) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_5_U1_Ins_0_U1 ( .A(KeyArray_outS23ser[5]), 
        .B(KeyArray_S23reg_gff_1_SFF_5_QD), .S(n179), .Z(
        KeyArray_S23reg_gff_1_SFF_5_n5) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2674), 
        .B(new_AGEMA_signal_2973), .S(n179), .Z(new_AGEMA_signal_3344) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS23ser[5]), .B(KeyArray_outS33ser[5]), .S(n170), .Z(
        KeyArray_S23reg_gff_1_SFF_5_QD) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2699), .B(new_AGEMA_signal_2770), .S(n170), .Z(
        new_AGEMA_signal_2973) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_6_U1_Ins_0_U1 ( .A(KeyArray_outS23ser[6]), 
        .B(KeyArray_S23reg_gff_1_SFF_6_QD), .S(n179), .Z(
        KeyArray_S23reg_gff_1_SFF_6_n5) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2677), 
        .B(new_AGEMA_signal_2974), .S(n179), .Z(new_AGEMA_signal_3345) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS23ser[6]), .B(KeyArray_outS33ser[6]), .S(n170), .Z(
        KeyArray_S23reg_gff_1_SFF_6_QD) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2702), .B(new_AGEMA_signal_2773), .S(n170), .Z(
        new_AGEMA_signal_2974) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_7_U1_Ins_0_U1 ( .A(KeyArray_outS23ser[7]), 
        .B(KeyArray_S23reg_gff_1_SFF_7_QD), .S(n179), .Z(
        KeyArray_S23reg_gff_1_SFF_7_n5) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2680), 
        .B(new_AGEMA_signal_2975), .S(n179), .Z(new_AGEMA_signal_3346) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS23ser[7]), .B(KeyArray_outS33ser[7]), .S(n171), .Z(
        KeyArray_S23reg_gff_1_SFF_7_QD) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2705), .B(new_AGEMA_signal_2776), .S(n171), .Z(
        new_AGEMA_signal_2975) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_0_U1_Ins_0_U1 ( .A(KeyArray_outS31ser[0]), 
        .B(KeyArray_S31reg_gff_1_SFF_0_QD), .S(n179), .Z(
        KeyArray_S31reg_gff_1_SFF_0_n6) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_0_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2707), 
        .B(new_AGEMA_signal_2976), .S(n179), .Z(new_AGEMA_signal_3347) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS31ser[0]), .B(KeyArray_outS01ser_0_), .S(n171), .Z(
        KeyArray_S31reg_gff_1_SFF_0_QD) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2732), .B(new_AGEMA_signal_2020), .S(n171), .Z(
        new_AGEMA_signal_2976) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_1_U1_Ins_0_U1 ( .A(KeyArray_outS31ser[1]), 
        .B(KeyArray_S31reg_gff_1_SFF_1_QD), .S(n179), .Z(
        KeyArray_S31reg_gff_1_SFF_1_n6) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2710), 
        .B(new_AGEMA_signal_2977), .S(n179), .Z(new_AGEMA_signal_3348) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS31ser[1]), .B(KeyArray_outS01ser_1_), .S(n171), .Z(
        KeyArray_S31reg_gff_1_SFF_1_QD) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2735), .B(new_AGEMA_signal_2018), .S(n171), .Z(
        new_AGEMA_signal_2977) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_2_U1_Ins_0_U1 ( .A(KeyArray_outS31ser[2]), 
        .B(KeyArray_S31reg_gff_1_SFF_2_QD), .S(n179), .Z(
        KeyArray_S31reg_gff_1_SFF_2_n6) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2713), 
        .B(new_AGEMA_signal_2978), .S(n179), .Z(new_AGEMA_signal_3349) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS31ser[2]), .B(KeyArray_outS01ser_2_), .S(n171), .Z(
        KeyArray_S31reg_gff_1_SFF_2_QD) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2738), .B(new_AGEMA_signal_2016), .S(n171), .Z(
        new_AGEMA_signal_2978) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_3_U1_Ins_0_U1 ( .A(KeyArray_outS31ser[3]), 
        .B(KeyArray_S31reg_gff_1_SFF_3_QD), .S(n179), .Z(
        KeyArray_S31reg_gff_1_SFF_3_n6) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_3_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2716), 
        .B(new_AGEMA_signal_2979), .S(n179), .Z(new_AGEMA_signal_3350) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS31ser[3]), .B(KeyArray_outS01ser_3_), .S(n171), .Z(
        KeyArray_S31reg_gff_1_SFF_3_QD) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2741), .B(new_AGEMA_signal_2014), .S(n171), .Z(
        new_AGEMA_signal_2979) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_4_U1_Ins_0_U1 ( .A(KeyArray_outS31ser[4]), 
        .B(KeyArray_S31reg_gff_1_SFF_4_QD), .S(n178), .Z(
        KeyArray_S31reg_gff_1_SFF_4_n6) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2719), 
        .B(new_AGEMA_signal_2980), .S(n178), .Z(new_AGEMA_signal_3351) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS31ser[4]), .B(KeyArray_outS01ser_4_), .S(n171), .Z(
        KeyArray_S31reg_gff_1_SFF_4_QD) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2744), .B(new_AGEMA_signal_2012), .S(n171), .Z(
        new_AGEMA_signal_2980) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_5_U1_Ins_0_U1 ( .A(KeyArray_outS31ser[5]), 
        .B(KeyArray_S31reg_gff_1_SFF_5_QD), .S(n183), .Z(
        KeyArray_S31reg_gff_1_SFF_5_n6) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2722), 
        .B(new_AGEMA_signal_2981), .S(n183), .Z(new_AGEMA_signal_3352) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS31ser[5]), .B(KeyArray_outS01ser_5_), .S(n171), .Z(
        KeyArray_S31reg_gff_1_SFF_5_QD) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2747), .B(new_AGEMA_signal_2010), .S(n171), .Z(
        new_AGEMA_signal_2981) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_6_U1_Ins_0_U1 ( .A(KeyArray_outS31ser[6]), 
        .B(KeyArray_S31reg_gff_1_SFF_6_QD), .S(n178), .Z(
        KeyArray_S31reg_gff_1_SFF_6_n6) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2725), 
        .B(new_AGEMA_signal_2982), .S(n178), .Z(new_AGEMA_signal_3353) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS31ser[6]), .B(KeyArray_outS01ser_6_), .S(n172), .Z(
        KeyArray_S31reg_gff_1_SFF_6_QD) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2750), .B(new_AGEMA_signal_2008), .S(n172), .Z(
        new_AGEMA_signal_2982) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_7_U1_Ins_0_U1 ( .A(KeyArray_outS31ser[7]), 
        .B(KeyArray_S31reg_gff_1_SFF_7_QD), .S(n178), .Z(
        KeyArray_S31reg_gff_1_SFF_7_n6) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2728), 
        .B(new_AGEMA_signal_2983), .S(n178), .Z(new_AGEMA_signal_3354) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS31ser[7]), .B(KeyArray_outS01ser_7_), .S(n172), .Z(
        KeyArray_S31reg_gff_1_SFF_7_QD) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2753), .B(new_AGEMA_signal_2006), .S(n172), .Z(
        new_AGEMA_signal_2983) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_0_U1_Ins_0_U1 ( .A(KeyArray_outS32ser[0]), 
        .B(KeyArray_S32reg_gff_1_SFF_0_QD), .S(n178), .Z(
        KeyArray_S32reg_gff_1_SFF_0_n6) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_0_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2731), 
        .B(new_AGEMA_signal_2984), .S(n178), .Z(new_AGEMA_signal_3355) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS32ser[0]), .B(KeyArray_outS02ser[0]), .S(n172), .Z(
        KeyArray_S32reg_gff_1_SFF_0_QD) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2756), .B(new_AGEMA_signal_2443), .S(n172), .Z(
        new_AGEMA_signal_2984) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_1_U1_Ins_0_U1 ( .A(KeyArray_outS32ser[1]), 
        .B(KeyArray_S32reg_gff_1_SFF_1_QD), .S(n178), .Z(
        KeyArray_S32reg_gff_1_SFF_1_n6) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2734), 
        .B(new_AGEMA_signal_2985), .S(n178), .Z(new_AGEMA_signal_3356) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS32ser[1]), .B(KeyArray_outS02ser[1]), .S(n172), .Z(
        KeyArray_S32reg_gff_1_SFF_1_QD) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2759), .B(new_AGEMA_signal_2446), .S(n172), .Z(
        new_AGEMA_signal_2985) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_2_U1_Ins_0_U1 ( .A(KeyArray_outS32ser[2]), 
        .B(KeyArray_S32reg_gff_1_SFF_2_QD), .S(n178), .Z(
        KeyArray_S32reg_gff_1_SFF_2_n6) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2737), 
        .B(new_AGEMA_signal_2986), .S(n178), .Z(new_AGEMA_signal_3357) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS32ser[2]), .B(KeyArray_outS02ser[2]), .S(n172), .Z(
        KeyArray_S32reg_gff_1_SFF_2_QD) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2762), .B(new_AGEMA_signal_2449), .S(n172), .Z(
        new_AGEMA_signal_2986) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_3_U1_Ins_0_U1 ( .A(KeyArray_outS32ser[3]), 
        .B(KeyArray_S32reg_gff_1_SFF_3_QD), .S(n178), .Z(
        KeyArray_S32reg_gff_1_SFF_3_n6) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_3_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2740), 
        .B(new_AGEMA_signal_2987), .S(n178), .Z(new_AGEMA_signal_3358) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS32ser[3]), .B(KeyArray_outS02ser[3]), .S(n172), .Z(
        KeyArray_S32reg_gff_1_SFF_3_QD) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2765), .B(new_AGEMA_signal_2452), .S(n172), .Z(
        new_AGEMA_signal_2987) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_4_U1_Ins_0_U1 ( .A(KeyArray_outS32ser[4]), 
        .B(KeyArray_S32reg_gff_1_SFF_4_QD), .S(n177), .Z(
        KeyArray_S32reg_gff_1_SFF_4_n6) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2743), 
        .B(new_AGEMA_signal_2988), .S(n177), .Z(new_AGEMA_signal_3359) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS32ser[4]), .B(KeyArray_outS02ser[4]), .S(n172), .Z(
        KeyArray_S32reg_gff_1_SFF_4_QD) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2768), .B(new_AGEMA_signal_2455), .S(n172), .Z(
        new_AGEMA_signal_2988) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_5_U1_Ins_0_U1 ( .A(KeyArray_outS32ser[5]), 
        .B(KeyArray_S32reg_gff_1_SFF_5_QD), .S(n177), .Z(
        KeyArray_S32reg_gff_1_SFF_5_n6) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2746), 
        .B(new_AGEMA_signal_2989), .S(n177), .Z(new_AGEMA_signal_3360) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS32ser[5]), .B(KeyArray_outS02ser[5]), .S(n175), .Z(
        KeyArray_S32reg_gff_1_SFF_5_QD) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2771), .B(new_AGEMA_signal_2458), .S(n175), .Z(
        new_AGEMA_signal_2989) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_6_U1_Ins_0_U1 ( .A(KeyArray_outS32ser[6]), 
        .B(KeyArray_S32reg_gff_1_SFF_6_QD), .S(n177), .Z(
        KeyArray_S32reg_gff_1_SFF_6_n5) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2749), 
        .B(new_AGEMA_signal_2990), .S(n177), .Z(new_AGEMA_signal_3361) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS32ser[6]), .B(KeyArray_outS02ser[6]), .S(n162), .Z(
        KeyArray_S32reg_gff_1_SFF_6_QD) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2774), .B(new_AGEMA_signal_2461), .S(n162), .Z(
        new_AGEMA_signal_2990) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_7_U1_Ins_0_U1 ( .A(KeyArray_outS32ser[7]), 
        .B(KeyArray_S32reg_gff_1_SFF_7_QD), .S(n177), .Z(
        KeyArray_S32reg_gff_1_SFF_7_n5) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2752), 
        .B(new_AGEMA_signal_2991), .S(n177), .Z(new_AGEMA_signal_3362) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS32ser[7]), .B(KeyArray_outS02ser[7]), .S(n175), .Z(
        KeyArray_S32reg_gff_1_SFF_7_QD) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2777), .B(new_AGEMA_signal_2464), .S(n175), .Z(
        new_AGEMA_signal_2991) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_0_U1_Ins_0_U1 ( .A(KeyArray_outS33ser[0]), 
        .B(KeyArray_S33reg_gff_1_SFF_0_QD), .S(n177), .Z(
        KeyArray_S33reg_gff_1_SFF_0_n5) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_0_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2755), 
        .B(new_AGEMA_signal_2992), .S(n177), .Z(new_AGEMA_signal_3363) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS33ser[0]), .B(KeyArray_outS03ser[0]), .S(n162), .Z(
        KeyArray_S33reg_gff_1_SFF_0_QD) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2779), .B(new_AGEMA_signal_2467), .S(n162), .Z(
        new_AGEMA_signal_2992) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_1_U1_Ins_0_U1 ( .A(KeyArray_outS33ser[1]), 
        .B(KeyArray_S33reg_gff_1_SFF_1_QD), .S(n177), .Z(
        KeyArray_S33reg_gff_1_SFF_1_n5) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2758), 
        .B(new_AGEMA_signal_2993), .S(n177), .Z(new_AGEMA_signal_3364) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS33ser[1]), .B(KeyArray_outS03ser[1]), .S(n176), .Z(
        KeyArray_S33reg_gff_1_SFF_1_QD) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2781), .B(new_AGEMA_signal_2470), .S(n176), .Z(
        new_AGEMA_signal_2993) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_2_U1_Ins_0_U1 ( .A(KeyArray_outS33ser[2]), 
        .B(KeyArray_S33reg_gff_1_SFF_2_QD), .S(n177), .Z(
        KeyArray_S33reg_gff_1_SFF_2_n5) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2761), 
        .B(new_AGEMA_signal_2994), .S(n177), .Z(new_AGEMA_signal_3365) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS33ser[2]), .B(KeyArray_outS03ser[2]), .S(n176), .Z(
        KeyArray_S33reg_gff_1_SFF_2_QD) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2783), .B(new_AGEMA_signal_2473), .S(n176), .Z(
        new_AGEMA_signal_2994) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_3_U1_Ins_0_U1 ( .A(KeyArray_outS33ser[3]), 
        .B(KeyArray_S33reg_gff_1_SFF_3_QD), .S(n178), .Z(
        KeyArray_S33reg_gff_1_SFF_3_n5) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_3_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2764), 
        .B(new_AGEMA_signal_2995), .S(n178), .Z(new_AGEMA_signal_3366) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS33ser[3]), .B(KeyArray_outS03ser[3]), .S(n176), .Z(
        KeyArray_S33reg_gff_1_SFF_3_QD) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2785), .B(new_AGEMA_signal_2476), .S(n176), .Z(
        new_AGEMA_signal_2995) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_4_U1_Ins_0_U1 ( .A(KeyArray_outS33ser[4]), 
        .B(KeyArray_S33reg_gff_1_SFF_4_QD), .S(n185), .Z(
        KeyArray_S33reg_gff_1_SFF_4_n5) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2767), 
        .B(new_AGEMA_signal_2996), .S(n185), .Z(new_AGEMA_signal_3367) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS33ser[4]), .B(KeyArray_outS03ser[4]), .S(n173), .Z(
        KeyArray_S33reg_gff_1_SFF_4_QD) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2787), .B(new_AGEMA_signal_2479), .S(n173), .Z(
        new_AGEMA_signal_2996) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_5_U1_Ins_0_U1 ( .A(KeyArray_outS33ser[5]), 
        .B(KeyArray_S33reg_gff_1_SFF_5_QD), .S(n190), .Z(
        KeyArray_S33reg_gff_1_SFF_5_n5) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2770), 
        .B(new_AGEMA_signal_2997), .S(n190), .Z(new_AGEMA_signal_3368) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS33ser[5]), .B(KeyArray_outS03ser[5]), .S(n173), .Z(
        KeyArray_S33reg_gff_1_SFF_5_QD) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2789), .B(new_AGEMA_signal_2482), .S(n173), .Z(
        new_AGEMA_signal_2997) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_6_U1_Ins_0_U1 ( .A(KeyArray_outS33ser[6]), 
        .B(KeyArray_S33reg_gff_1_SFF_6_QD), .S(n182), .Z(
        KeyArray_S33reg_gff_1_SFF_6_n5) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2773), 
        .B(new_AGEMA_signal_2998), .S(n182), .Z(new_AGEMA_signal_3369) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS33ser[6]), .B(KeyArray_outS03ser[6]), .S(n173), .Z(
        KeyArray_S33reg_gff_1_SFF_6_QD) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2791), .B(new_AGEMA_signal_2485), .S(n173), .Z(
        new_AGEMA_signal_2998) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_7_U1_Ins_0_U1 ( .A(KeyArray_outS33ser[7]), 
        .B(KeyArray_S33reg_gff_1_SFF_7_QD), .S(n187), .Z(
        KeyArray_S33reg_gff_1_SFF_7_n5) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2776), 
        .B(new_AGEMA_signal_2999), .S(n187), .Z(new_AGEMA_signal_3370) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS33ser[7]), .B(KeyArray_outS03ser[7]), .S(n173), .Z(
        KeyArray_S33reg_gff_1_SFF_7_QD) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2793), .B(new_AGEMA_signal_2488), .S(n173), .Z(
        new_AGEMA_signal_2999) );
  MUX2_X1 KeyArray_MUX_selXOR_mux_inst_0_U1_Ins_0_U1 ( .A(
        KeyArray_outS01ser_0_), .B(KeyArray_outS01ser_XOR_00[0]), .S(intselXOR), .Z(KeyArray_outS01ser_p[0]) );
  MUX2_X1 KeyArray_MUX_selXOR_mux_inst_0_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2020), .B(new_AGEMA_signal_2021), .S(intselXOR), .Z(
        new_AGEMA_signal_3109) );
  MUX2_X1 KeyArray_MUX_selXOR_mux_inst_1_U1_Ins_0_U1 ( .A(
        KeyArray_outS01ser_1_), .B(KeyArray_outS01ser_XOR_00[1]), .S(intselXOR), .Z(KeyArray_outS01ser_p[1]) );
  MUX2_X1 KeyArray_MUX_selXOR_mux_inst_1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2018), .B(new_AGEMA_signal_2019), .S(intselXOR), .Z(
        new_AGEMA_signal_3110) );
  MUX2_X1 KeyArray_MUX_selXOR_mux_inst_2_U1_Ins_0_U1 ( .A(
        KeyArray_outS01ser_2_), .B(KeyArray_outS01ser_XOR_00[2]), .S(intselXOR), .Z(KeyArray_outS01ser_p[2]) );
  MUX2_X1 KeyArray_MUX_selXOR_mux_inst_2_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2016), .B(new_AGEMA_signal_2017), .S(intselXOR), .Z(
        new_AGEMA_signal_3111) );
  MUX2_X1 KeyArray_MUX_selXOR_mux_inst_3_U1_Ins_0_U1 ( .A(
        KeyArray_outS01ser_3_), .B(KeyArray_outS01ser_XOR_00[3]), .S(intselXOR), .Z(KeyArray_outS01ser_p[3]) );
  MUX2_X1 KeyArray_MUX_selXOR_mux_inst_3_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2014), .B(new_AGEMA_signal_2015), .S(intselXOR), .Z(
        new_AGEMA_signal_3112) );
  MUX2_X1 KeyArray_MUX_selXOR_mux_inst_4_U1_Ins_0_U1 ( .A(
        KeyArray_outS01ser_4_), .B(KeyArray_outS01ser_XOR_00[4]), .S(intselXOR), .Z(KeyArray_outS01ser_p[4]) );
  MUX2_X1 KeyArray_MUX_selXOR_mux_inst_4_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2012), .B(new_AGEMA_signal_2013), .S(intselXOR), .Z(
        new_AGEMA_signal_3113) );
  MUX2_X1 KeyArray_MUX_selXOR_mux_inst_5_U1_Ins_0_U1 ( .A(
        KeyArray_outS01ser_5_), .B(KeyArray_outS01ser_XOR_00[5]), .S(intselXOR), .Z(KeyArray_outS01ser_p[5]) );
  MUX2_X1 KeyArray_MUX_selXOR_mux_inst_5_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2010), .B(new_AGEMA_signal_2011), .S(intselXOR), .Z(
        new_AGEMA_signal_3114) );
  MUX2_X1 KeyArray_MUX_selXOR_mux_inst_6_U1_Ins_0_U1 ( .A(
        KeyArray_outS01ser_6_), .B(KeyArray_outS01ser_XOR_00[6]), .S(intselXOR), .Z(KeyArray_outS01ser_p[6]) );
  MUX2_X1 KeyArray_MUX_selXOR_mux_inst_6_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2008), .B(new_AGEMA_signal_2009), .S(intselXOR), .Z(
        new_AGEMA_signal_3115) );
  MUX2_X1 KeyArray_MUX_selXOR_mux_inst_7_U1_Ins_0_U1 ( .A(
        KeyArray_outS01ser_7_), .B(KeyArray_outS01ser_XOR_00[7]), .S(intselXOR), .Z(KeyArray_outS01ser_p[7]) );
  MUX2_X1 KeyArray_MUX_selXOR_mux_inst_7_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2006), .B(new_AGEMA_signal_2007), .S(intselXOR), .Z(
        new_AGEMA_signal_3116) );
  MUX2_X1 KeyArray_MUX_inS00ser_mux_inst_0_U1_Ins_0_U1 ( .A(key_s0[120]), .B(
        KeyArray_outS01ser_p[0]), .S(n206), .Z(KeyArray_inS00ser[0]) );
  MUX2_X1 KeyArray_MUX_inS00ser_mux_inst_0_U1_Ins_1_U1 ( .A(key_s1[120]), .B(
        new_AGEMA_signal_3109), .S(n206), .Z(new_AGEMA_signal_3247) );
  MUX2_X1 KeyArray_MUX_inS00ser_mux_inst_1_U1_Ins_0_U1 ( .A(key_s0[121]), .B(
        KeyArray_outS01ser_p[1]), .S(n211), .Z(KeyArray_inS00ser[1]) );
  MUX2_X1 KeyArray_MUX_inS00ser_mux_inst_1_U1_Ins_1_U1 ( .A(key_s1[121]), .B(
        new_AGEMA_signal_3110), .S(n211), .Z(new_AGEMA_signal_3249) );
  MUX2_X1 KeyArray_MUX_inS00ser_mux_inst_2_U1_Ins_0_U1 ( .A(key_s0[122]), .B(
        KeyArray_outS01ser_p[2]), .S(n207), .Z(KeyArray_inS00ser[2]) );
  MUX2_X1 KeyArray_MUX_inS00ser_mux_inst_2_U1_Ins_1_U1 ( .A(key_s1[122]), .B(
        new_AGEMA_signal_3111), .S(n207), .Z(new_AGEMA_signal_3251) );
  MUX2_X1 KeyArray_MUX_inS00ser_mux_inst_3_U1_Ins_0_U1 ( .A(key_s0[123]), .B(
        KeyArray_outS01ser_p[3]), .S(n212), .Z(KeyArray_inS00ser[3]) );
  MUX2_X1 KeyArray_MUX_inS00ser_mux_inst_3_U1_Ins_1_U1 ( .A(key_s1[123]), .B(
        new_AGEMA_signal_3112), .S(n212), .Z(new_AGEMA_signal_3253) );
  MUX2_X1 KeyArray_MUX_inS00ser_mux_inst_4_U1_Ins_0_U1 ( .A(key_s0[124]), .B(
        KeyArray_outS01ser_p[4]), .S(n220), .Z(KeyArray_inS00ser[4]) );
  MUX2_X1 KeyArray_MUX_inS00ser_mux_inst_4_U1_Ins_1_U1 ( .A(key_s1[124]), .B(
        new_AGEMA_signal_3113), .S(n220), .Z(new_AGEMA_signal_3255) );
  MUX2_X1 KeyArray_MUX_inS00ser_mux_inst_5_U1_Ins_0_U1 ( .A(key_s0[125]), .B(
        KeyArray_outS01ser_p[5]), .S(n219), .Z(KeyArray_inS00ser[5]) );
  MUX2_X1 KeyArray_MUX_inS00ser_mux_inst_5_U1_Ins_1_U1 ( .A(key_s1[125]), .B(
        new_AGEMA_signal_3114), .S(n219), .Z(new_AGEMA_signal_3257) );
  MUX2_X1 KeyArray_MUX_inS00ser_mux_inst_6_U1_Ins_0_U1 ( .A(key_s0[126]), .B(
        KeyArray_outS01ser_p[6]), .S(n222), .Z(KeyArray_inS00ser[6]) );
  MUX2_X1 KeyArray_MUX_inS00ser_mux_inst_6_U1_Ins_1_U1 ( .A(key_s1[126]), .B(
        new_AGEMA_signal_3115), .S(n222), .Z(new_AGEMA_signal_3259) );
  MUX2_X1 KeyArray_MUX_inS00ser_mux_inst_7_U1_Ins_0_U1 ( .A(key_s0[127]), .B(
        KeyArray_outS01ser_p[7]), .S(n221), .Z(KeyArray_inS00ser[7]) );
  MUX2_X1 KeyArray_MUX_inS00ser_mux_inst_7_U1_Ins_1_U1 ( .A(key_s1[127]), .B(
        new_AGEMA_signal_3116), .S(n221), .Z(new_AGEMA_signal_3261) );
  MUX2_X1 KeyArray_MUX_inS01ser_mux_inst_0_U1_Ins_0_U1 ( .A(key_s0[112]), .B(
        KeyArray_outS02ser[0]), .S(n213), .Z(KeyArray_inS01ser[0]) );
  MUX2_X1 KeyArray_MUX_inS01ser_mux_inst_0_U1_Ins_1_U1 ( .A(key_s1[112]), .B(
        new_AGEMA_signal_2443), .S(n213), .Z(new_AGEMA_signal_2444) );
  MUX2_X1 KeyArray_MUX_inS01ser_mux_inst_1_U1_Ins_0_U1 ( .A(key_s0[113]), .B(
        KeyArray_outS02ser[1]), .S(n218), .Z(KeyArray_inS01ser[1]) );
  MUX2_X1 KeyArray_MUX_inS01ser_mux_inst_1_U1_Ins_1_U1 ( .A(key_s1[113]), .B(
        new_AGEMA_signal_2446), .S(n218), .Z(new_AGEMA_signal_2447) );
  MUX2_X1 KeyArray_MUX_inS01ser_mux_inst_2_U1_Ins_0_U1 ( .A(key_s0[114]), .B(
        KeyArray_outS02ser[2]), .S(n217), .Z(KeyArray_inS01ser[2]) );
  MUX2_X1 KeyArray_MUX_inS01ser_mux_inst_2_U1_Ins_1_U1 ( .A(key_s1[114]), .B(
        new_AGEMA_signal_2449), .S(n217), .Z(new_AGEMA_signal_2450) );
  MUX2_X1 KeyArray_MUX_inS01ser_mux_inst_3_U1_Ins_0_U1 ( .A(key_s0[115]), .B(
        KeyArray_outS02ser[3]), .S(n216), .Z(KeyArray_inS01ser[3]) );
  MUX2_X1 KeyArray_MUX_inS01ser_mux_inst_3_U1_Ins_1_U1 ( .A(key_s1[115]), .B(
        new_AGEMA_signal_2452), .S(n216), .Z(new_AGEMA_signal_2453) );
  MUX2_X1 KeyArray_MUX_inS01ser_mux_inst_4_U1_Ins_0_U1 ( .A(key_s0[116]), .B(
        KeyArray_outS02ser[4]), .S(n215), .Z(KeyArray_inS01ser[4]) );
  MUX2_X1 KeyArray_MUX_inS01ser_mux_inst_4_U1_Ins_1_U1 ( .A(key_s1[116]), .B(
        new_AGEMA_signal_2455), .S(n215), .Z(new_AGEMA_signal_2456) );
  MUX2_X1 KeyArray_MUX_inS01ser_mux_inst_5_U1_Ins_0_U1 ( .A(key_s0[117]), .B(
        KeyArray_outS02ser[5]), .S(n208), .Z(KeyArray_inS01ser[5]) );
  MUX2_X1 KeyArray_MUX_inS01ser_mux_inst_5_U1_Ins_1_U1 ( .A(key_s1[117]), .B(
        new_AGEMA_signal_2458), .S(n208), .Z(new_AGEMA_signal_2459) );
  MUX2_X1 KeyArray_MUX_inS01ser_mux_inst_6_U1_Ins_0_U1 ( .A(key_s0[118]), .B(
        KeyArray_outS02ser[6]), .S(n213), .Z(KeyArray_inS01ser[6]) );
  MUX2_X1 KeyArray_MUX_inS01ser_mux_inst_6_U1_Ins_1_U1 ( .A(key_s1[118]), .B(
        new_AGEMA_signal_2461), .S(n213), .Z(new_AGEMA_signal_2462) );
  MUX2_X1 KeyArray_MUX_inS01ser_mux_inst_7_U1_Ins_0_U1 ( .A(key_s0[119]), .B(
        KeyArray_outS02ser[7]), .S(n205), .Z(KeyArray_inS01ser[7]) );
  MUX2_X1 KeyArray_MUX_inS01ser_mux_inst_7_U1_Ins_1_U1 ( .A(key_s1[119]), .B(
        new_AGEMA_signal_2464), .S(n205), .Z(new_AGEMA_signal_2465) );
  MUX2_X1 KeyArray_MUX_inS02ser_mux_inst_0_U1_Ins_0_U1 ( .A(key_s0[104]), .B(
        KeyArray_outS03ser[0]), .S(n205), .Z(KeyArray_inS02ser[0]) );
  MUX2_X1 KeyArray_MUX_inS02ser_mux_inst_0_U1_Ins_1_U1 ( .A(key_s1[104]), .B(
        new_AGEMA_signal_2467), .S(n205), .Z(new_AGEMA_signal_2468) );
  MUX2_X1 KeyArray_MUX_inS02ser_mux_inst_1_U1_Ins_0_U1 ( .A(key_s0[105]), .B(
        KeyArray_outS03ser[1]), .S(n205), .Z(KeyArray_inS02ser[1]) );
  MUX2_X1 KeyArray_MUX_inS02ser_mux_inst_1_U1_Ins_1_U1 ( .A(key_s1[105]), .B(
        new_AGEMA_signal_2470), .S(n205), .Z(new_AGEMA_signal_2471) );
  MUX2_X1 KeyArray_MUX_inS02ser_mux_inst_2_U1_Ins_0_U1 ( .A(key_s0[106]), .B(
        KeyArray_outS03ser[2]), .S(n205), .Z(KeyArray_inS02ser[2]) );
  MUX2_X1 KeyArray_MUX_inS02ser_mux_inst_2_U1_Ins_1_U1 ( .A(key_s1[106]), .B(
        new_AGEMA_signal_2473), .S(n205), .Z(new_AGEMA_signal_2474) );
  MUX2_X1 KeyArray_MUX_inS02ser_mux_inst_3_U1_Ins_0_U1 ( .A(key_s0[107]), .B(
        KeyArray_outS03ser[3]), .S(n205), .Z(KeyArray_inS02ser[3]) );
  MUX2_X1 KeyArray_MUX_inS02ser_mux_inst_3_U1_Ins_1_U1 ( .A(key_s1[107]), .B(
        new_AGEMA_signal_2476), .S(n205), .Z(new_AGEMA_signal_2477) );
  MUX2_X1 KeyArray_MUX_inS02ser_mux_inst_4_U1_Ins_0_U1 ( .A(key_s0[108]), .B(
        KeyArray_outS03ser[4]), .S(n205), .Z(KeyArray_inS02ser[4]) );
  MUX2_X1 KeyArray_MUX_inS02ser_mux_inst_4_U1_Ins_1_U1 ( .A(key_s1[108]), .B(
        new_AGEMA_signal_2479), .S(n205), .Z(new_AGEMA_signal_2480) );
  MUX2_X1 KeyArray_MUX_inS02ser_mux_inst_5_U1_Ins_0_U1 ( .A(key_s0[109]), .B(
        KeyArray_outS03ser[5]), .S(n205), .Z(KeyArray_inS02ser[5]) );
  MUX2_X1 KeyArray_MUX_inS02ser_mux_inst_5_U1_Ins_1_U1 ( .A(key_s1[109]), .B(
        new_AGEMA_signal_2482), .S(n205), .Z(new_AGEMA_signal_2483) );
  MUX2_X1 KeyArray_MUX_inS02ser_mux_inst_6_U1_Ins_0_U1 ( .A(key_s0[110]), .B(
        KeyArray_outS03ser[6]), .S(n206), .Z(KeyArray_inS02ser[6]) );
  MUX2_X1 KeyArray_MUX_inS02ser_mux_inst_6_U1_Ins_1_U1 ( .A(key_s1[110]), .B(
        new_AGEMA_signal_2485), .S(n206), .Z(new_AGEMA_signal_2486) );
  MUX2_X1 KeyArray_MUX_inS02ser_mux_inst_7_U1_Ins_0_U1 ( .A(key_s0[111]), .B(
        KeyArray_outS03ser[7]), .S(n206), .Z(KeyArray_inS02ser[7]) );
  MUX2_X1 KeyArray_MUX_inS02ser_mux_inst_7_U1_Ins_1_U1 ( .A(key_s1[111]), .B(
        new_AGEMA_signal_2488), .S(n206), .Z(new_AGEMA_signal_2489) );
  MUX2_X1 KeyArray_MUX_inS03ser_mux_inst_0_U1_Ins_0_U1 ( .A(key_s0[96]), .B(
        KeyArray_outS10ser[0]), .S(n206), .Z(KeyArray_inS03ser[0]) );
  MUX2_X1 KeyArray_MUX_inS03ser_mux_inst_0_U1_Ins_1_U1 ( .A(key_s1[96]), .B(
        new_AGEMA_signal_2491), .S(n206), .Z(new_AGEMA_signal_2492) );
  MUX2_X1 KeyArray_MUX_inS03ser_mux_inst_1_U1_Ins_0_U1 ( .A(key_s0[97]), .B(
        KeyArray_outS10ser[1]), .S(n206), .Z(KeyArray_inS03ser[1]) );
  MUX2_X1 KeyArray_MUX_inS03ser_mux_inst_1_U1_Ins_1_U1 ( .A(key_s1[97]), .B(
        new_AGEMA_signal_2494), .S(n206), .Z(new_AGEMA_signal_2495) );
  MUX2_X1 KeyArray_MUX_inS03ser_mux_inst_2_U1_Ins_0_U1 ( .A(key_s0[98]), .B(
        KeyArray_outS10ser[2]), .S(n206), .Z(KeyArray_inS03ser[2]) );
  MUX2_X1 KeyArray_MUX_inS03ser_mux_inst_2_U1_Ins_1_U1 ( .A(key_s1[98]), .B(
        new_AGEMA_signal_2497), .S(n206), .Z(new_AGEMA_signal_2498) );
  MUX2_X1 KeyArray_MUX_inS03ser_mux_inst_3_U1_Ins_0_U1 ( .A(key_s0[99]), .B(
        KeyArray_outS10ser[3]), .S(n206), .Z(KeyArray_inS03ser[3]) );
  MUX2_X1 KeyArray_MUX_inS03ser_mux_inst_3_U1_Ins_1_U1 ( .A(key_s1[99]), .B(
        new_AGEMA_signal_2500), .S(n206), .Z(new_AGEMA_signal_2501) );
  MUX2_X1 KeyArray_MUX_inS03ser_mux_inst_4_U1_Ins_0_U1 ( .A(key_s0[100]), .B(
        KeyArray_outS10ser[4]), .S(n206), .Z(KeyArray_inS03ser[4]) );
  MUX2_X1 KeyArray_MUX_inS03ser_mux_inst_4_U1_Ins_1_U1 ( .A(key_s1[100]), .B(
        new_AGEMA_signal_2503), .S(n206), .Z(new_AGEMA_signal_2504) );
  MUX2_X1 KeyArray_MUX_inS03ser_mux_inst_5_U1_Ins_0_U1 ( .A(key_s0[101]), .B(
        KeyArray_outS10ser[5]), .S(n207), .Z(KeyArray_inS03ser[5]) );
  MUX2_X1 KeyArray_MUX_inS03ser_mux_inst_5_U1_Ins_1_U1 ( .A(key_s1[101]), .B(
        new_AGEMA_signal_2506), .S(n207), .Z(new_AGEMA_signal_2507) );
  MUX2_X1 KeyArray_MUX_inS03ser_mux_inst_6_U1_Ins_0_U1 ( .A(key_s0[102]), .B(
        KeyArray_outS10ser[6]), .S(n207), .Z(KeyArray_inS03ser[6]) );
  MUX2_X1 KeyArray_MUX_inS03ser_mux_inst_6_U1_Ins_1_U1 ( .A(key_s1[102]), .B(
        new_AGEMA_signal_2509), .S(n207), .Z(new_AGEMA_signal_2510) );
  MUX2_X1 KeyArray_MUX_inS03ser_mux_inst_7_U1_Ins_0_U1 ( .A(key_s0[103]), .B(
        KeyArray_outS10ser[7]), .S(n207), .Z(KeyArray_inS03ser[7]) );
  MUX2_X1 KeyArray_MUX_inS03ser_mux_inst_7_U1_Ins_1_U1 ( .A(key_s1[103]), .B(
        new_AGEMA_signal_2512), .S(n207), .Z(new_AGEMA_signal_2513) );
  MUX2_X1 KeyArray_MUX_inS10ser_mux_inst_0_U1_Ins_0_U1 ( .A(key_s0[88]), .B(
        KeyArray_outS11ser[0]), .S(n207), .Z(KeyArray_inS10ser[0]) );
  MUX2_X1 KeyArray_MUX_inS10ser_mux_inst_0_U1_Ins_1_U1 ( .A(key_s1[88]), .B(
        new_AGEMA_signal_2515), .S(n207), .Z(new_AGEMA_signal_2516) );
  MUX2_X1 KeyArray_MUX_inS10ser_mux_inst_1_U1_Ins_0_U1 ( .A(key_s0[89]), .B(
        KeyArray_outS11ser[1]), .S(n207), .Z(KeyArray_inS10ser[1]) );
  MUX2_X1 KeyArray_MUX_inS10ser_mux_inst_1_U1_Ins_1_U1 ( .A(key_s1[89]), .B(
        new_AGEMA_signal_2518), .S(n207), .Z(new_AGEMA_signal_2519) );
  MUX2_X1 KeyArray_MUX_inS10ser_mux_inst_2_U1_Ins_0_U1 ( .A(key_s0[90]), .B(
        KeyArray_outS11ser[2]), .S(n207), .Z(KeyArray_inS10ser[2]) );
  MUX2_X1 KeyArray_MUX_inS10ser_mux_inst_2_U1_Ins_1_U1 ( .A(key_s1[90]), .B(
        new_AGEMA_signal_2521), .S(n207), .Z(new_AGEMA_signal_2522) );
  MUX2_X1 KeyArray_MUX_inS10ser_mux_inst_3_U1_Ins_0_U1 ( .A(key_s0[91]), .B(
        KeyArray_outS11ser[3]), .S(n207), .Z(KeyArray_inS10ser[3]) );
  MUX2_X1 KeyArray_MUX_inS10ser_mux_inst_3_U1_Ins_1_U1 ( .A(key_s1[91]), .B(
        new_AGEMA_signal_2524), .S(n207), .Z(new_AGEMA_signal_2525) );
  MUX2_X1 KeyArray_MUX_inS10ser_mux_inst_4_U1_Ins_0_U1 ( .A(key_s0[92]), .B(
        KeyArray_outS11ser[4]), .S(n208), .Z(KeyArray_inS10ser[4]) );
  MUX2_X1 KeyArray_MUX_inS10ser_mux_inst_4_U1_Ins_1_U1 ( .A(key_s1[92]), .B(
        new_AGEMA_signal_2527), .S(n208), .Z(new_AGEMA_signal_2528) );
  MUX2_X1 KeyArray_MUX_inS10ser_mux_inst_5_U1_Ins_0_U1 ( .A(key_s0[93]), .B(
        KeyArray_outS11ser[5]), .S(n208), .Z(KeyArray_inS10ser[5]) );
  MUX2_X1 KeyArray_MUX_inS10ser_mux_inst_5_U1_Ins_1_U1 ( .A(key_s1[93]), .B(
        new_AGEMA_signal_2530), .S(n208), .Z(new_AGEMA_signal_2531) );
  MUX2_X1 KeyArray_MUX_inS10ser_mux_inst_6_U1_Ins_0_U1 ( .A(key_s0[94]), .B(
        KeyArray_outS11ser[6]), .S(n208), .Z(KeyArray_inS10ser[6]) );
  MUX2_X1 KeyArray_MUX_inS10ser_mux_inst_6_U1_Ins_1_U1 ( .A(key_s1[94]), .B(
        new_AGEMA_signal_2533), .S(n208), .Z(new_AGEMA_signal_2534) );
  MUX2_X1 KeyArray_MUX_inS10ser_mux_inst_7_U1_Ins_0_U1 ( .A(key_s0[95]), .B(
        KeyArray_outS11ser[7]), .S(n208), .Z(KeyArray_inS10ser[7]) );
  MUX2_X1 KeyArray_MUX_inS10ser_mux_inst_7_U1_Ins_1_U1 ( .A(key_s1[95]), .B(
        new_AGEMA_signal_2536), .S(n208), .Z(new_AGEMA_signal_2537) );
  MUX2_X1 KeyArray_MUX_inS11ser_mux_inst_0_U1_Ins_0_U1 ( .A(key_s0[80]), .B(
        KeyArray_outS12ser[0]), .S(n208), .Z(KeyArray_inS11ser[0]) );
  MUX2_X1 KeyArray_MUX_inS11ser_mux_inst_0_U1_Ins_1_U1 ( .A(key_s1[80]), .B(
        new_AGEMA_signal_2539), .S(n208), .Z(new_AGEMA_signal_2540) );
  MUX2_X1 KeyArray_MUX_inS11ser_mux_inst_1_U1_Ins_0_U1 ( .A(key_s0[81]), .B(
        KeyArray_outS12ser[1]), .S(n208), .Z(KeyArray_inS11ser[1]) );
  MUX2_X1 KeyArray_MUX_inS11ser_mux_inst_1_U1_Ins_1_U1 ( .A(key_s1[81]), .B(
        new_AGEMA_signal_2542), .S(n208), .Z(new_AGEMA_signal_2543) );
  MUX2_X1 KeyArray_MUX_inS11ser_mux_inst_2_U1_Ins_0_U1 ( .A(key_s0[82]), .B(
        KeyArray_outS12ser[2]), .S(n208), .Z(KeyArray_inS11ser[2]) );
  MUX2_X1 KeyArray_MUX_inS11ser_mux_inst_2_U1_Ins_1_U1 ( .A(key_s1[82]), .B(
        new_AGEMA_signal_2545), .S(n208), .Z(new_AGEMA_signal_2546) );
  MUX2_X1 KeyArray_MUX_inS11ser_mux_inst_3_U1_Ins_0_U1 ( .A(key_s0[83]), .B(
        KeyArray_outS12ser[3]), .S(n209), .Z(KeyArray_inS11ser[3]) );
  MUX2_X1 KeyArray_MUX_inS11ser_mux_inst_3_U1_Ins_1_U1 ( .A(key_s1[83]), .B(
        new_AGEMA_signal_2548), .S(n209), .Z(new_AGEMA_signal_2549) );
  MUX2_X1 KeyArray_MUX_inS11ser_mux_inst_4_U1_Ins_0_U1 ( .A(key_s0[84]), .B(
        KeyArray_outS12ser[4]), .S(n209), .Z(KeyArray_inS11ser[4]) );
  MUX2_X1 KeyArray_MUX_inS11ser_mux_inst_4_U1_Ins_1_U1 ( .A(key_s1[84]), .B(
        new_AGEMA_signal_2551), .S(n209), .Z(new_AGEMA_signal_2552) );
  MUX2_X1 KeyArray_MUX_inS11ser_mux_inst_5_U1_Ins_0_U1 ( .A(key_s0[85]), .B(
        KeyArray_outS12ser[5]), .S(n209), .Z(KeyArray_inS11ser[5]) );
  MUX2_X1 KeyArray_MUX_inS11ser_mux_inst_5_U1_Ins_1_U1 ( .A(key_s1[85]), .B(
        new_AGEMA_signal_2554), .S(n209), .Z(new_AGEMA_signal_2555) );
  MUX2_X1 KeyArray_MUX_inS11ser_mux_inst_6_U1_Ins_0_U1 ( .A(key_s0[86]), .B(
        KeyArray_outS12ser[6]), .S(n209), .Z(KeyArray_inS11ser[6]) );
  MUX2_X1 KeyArray_MUX_inS11ser_mux_inst_6_U1_Ins_1_U1 ( .A(key_s1[86]), .B(
        new_AGEMA_signal_2557), .S(n209), .Z(new_AGEMA_signal_2558) );
  MUX2_X1 KeyArray_MUX_inS11ser_mux_inst_7_U1_Ins_0_U1 ( .A(key_s0[87]), .B(
        KeyArray_outS12ser[7]), .S(n209), .Z(KeyArray_inS11ser[7]) );
  MUX2_X1 KeyArray_MUX_inS11ser_mux_inst_7_U1_Ins_1_U1 ( .A(key_s1[87]), .B(
        new_AGEMA_signal_2560), .S(n209), .Z(new_AGEMA_signal_2561) );
  MUX2_X1 KeyArray_MUX_inS12ser_mux_inst_0_U1_Ins_0_U1 ( .A(key_s0[72]), .B(
        keySBIn[0]), .S(n209), .Z(KeyArray_inS12ser[0]) );
  MUX2_X1 KeyArray_MUX_inS12ser_mux_inst_0_U1_Ins_1_U1 ( .A(key_s1[72]), .B(
        new_AGEMA_signal_2563), .S(n209), .Z(new_AGEMA_signal_2564) );
  MUX2_X1 KeyArray_MUX_inS12ser_mux_inst_1_U1_Ins_0_U1 ( .A(key_s0[73]), .B(
        keySBIn[1]), .S(n209), .Z(KeyArray_inS12ser[1]) );
  MUX2_X1 KeyArray_MUX_inS12ser_mux_inst_1_U1_Ins_1_U1 ( .A(key_s1[73]), .B(
        new_AGEMA_signal_2566), .S(n209), .Z(new_AGEMA_signal_2567) );
  MUX2_X1 KeyArray_MUX_inS12ser_mux_inst_2_U1_Ins_0_U1 ( .A(key_s0[74]), .B(
        keySBIn[2]), .S(n210), .Z(KeyArray_inS12ser[2]) );
  MUX2_X1 KeyArray_MUX_inS12ser_mux_inst_2_U1_Ins_1_U1 ( .A(key_s1[74]), .B(
        new_AGEMA_signal_2569), .S(n210), .Z(new_AGEMA_signal_2570) );
  MUX2_X1 KeyArray_MUX_inS12ser_mux_inst_3_U1_Ins_0_U1 ( .A(key_s0[75]), .B(
        keySBIn[3]), .S(n210), .Z(KeyArray_inS12ser[3]) );
  MUX2_X1 KeyArray_MUX_inS12ser_mux_inst_3_U1_Ins_1_U1 ( .A(key_s1[75]), .B(
        new_AGEMA_signal_2572), .S(n210), .Z(new_AGEMA_signal_2573) );
  MUX2_X1 KeyArray_MUX_inS12ser_mux_inst_4_U1_Ins_0_U1 ( .A(key_s0[76]), .B(
        keySBIn[4]), .S(n210), .Z(KeyArray_inS12ser[4]) );
  MUX2_X1 KeyArray_MUX_inS12ser_mux_inst_4_U1_Ins_1_U1 ( .A(key_s1[76]), .B(
        new_AGEMA_signal_2575), .S(n210), .Z(new_AGEMA_signal_2576) );
  MUX2_X1 KeyArray_MUX_inS12ser_mux_inst_5_U1_Ins_0_U1 ( .A(key_s0[77]), .B(
        keySBIn[5]), .S(n210), .Z(KeyArray_inS12ser[5]) );
  MUX2_X1 KeyArray_MUX_inS12ser_mux_inst_5_U1_Ins_1_U1 ( .A(key_s1[77]), .B(
        new_AGEMA_signal_2578), .S(n210), .Z(new_AGEMA_signal_2579) );
  MUX2_X1 KeyArray_MUX_inS12ser_mux_inst_6_U1_Ins_0_U1 ( .A(key_s0[78]), .B(
        keySBIn[6]), .S(n210), .Z(KeyArray_inS12ser[6]) );
  MUX2_X1 KeyArray_MUX_inS12ser_mux_inst_6_U1_Ins_1_U1 ( .A(key_s1[78]), .B(
        new_AGEMA_signal_2581), .S(n210), .Z(new_AGEMA_signal_2582) );
  MUX2_X1 KeyArray_MUX_inS12ser_mux_inst_7_U1_Ins_0_U1 ( .A(key_s0[79]), .B(
        keySBIn[7]), .S(n210), .Z(KeyArray_inS12ser[7]) );
  MUX2_X1 KeyArray_MUX_inS12ser_mux_inst_7_U1_Ins_1_U1 ( .A(key_s1[79]), .B(
        new_AGEMA_signal_2584), .S(n210), .Z(new_AGEMA_signal_2585) );
  MUX2_X1 KeyArray_MUX_inS13ser_mux_inst_0_U1_Ins_0_U1 ( .A(key_s0[64]), .B(
        KeyArray_outS20ser[0]), .S(n210), .Z(KeyArray_inS13ser[0]) );
  MUX2_X1 KeyArray_MUX_inS13ser_mux_inst_0_U1_Ins_1_U1 ( .A(key_s1[64]), .B(
        new_AGEMA_signal_2587), .S(n210), .Z(new_AGEMA_signal_2588) );
  MUX2_X1 KeyArray_MUX_inS13ser_mux_inst_1_U1_Ins_0_U1 ( .A(key_s0[65]), .B(
        KeyArray_outS20ser[1]), .S(n211), .Z(KeyArray_inS13ser[1]) );
  MUX2_X1 KeyArray_MUX_inS13ser_mux_inst_1_U1_Ins_1_U1 ( .A(key_s1[65]), .B(
        new_AGEMA_signal_2590), .S(n211), .Z(new_AGEMA_signal_2591) );
  MUX2_X1 KeyArray_MUX_inS13ser_mux_inst_2_U1_Ins_0_U1 ( .A(key_s0[66]), .B(
        KeyArray_outS20ser[2]), .S(n211), .Z(KeyArray_inS13ser[2]) );
  MUX2_X1 KeyArray_MUX_inS13ser_mux_inst_2_U1_Ins_1_U1 ( .A(key_s1[66]), .B(
        new_AGEMA_signal_2593), .S(n211), .Z(new_AGEMA_signal_2594) );
  MUX2_X1 KeyArray_MUX_inS13ser_mux_inst_3_U1_Ins_0_U1 ( .A(key_s0[67]), .B(
        KeyArray_outS20ser[3]), .S(n211), .Z(KeyArray_inS13ser[3]) );
  MUX2_X1 KeyArray_MUX_inS13ser_mux_inst_3_U1_Ins_1_U1 ( .A(key_s1[67]), .B(
        new_AGEMA_signal_2596), .S(n211), .Z(new_AGEMA_signal_2597) );
  MUX2_X1 KeyArray_MUX_inS13ser_mux_inst_4_U1_Ins_0_U1 ( .A(key_s0[68]), .B(
        KeyArray_outS20ser[4]), .S(n211), .Z(KeyArray_inS13ser[4]) );
  MUX2_X1 KeyArray_MUX_inS13ser_mux_inst_4_U1_Ins_1_U1 ( .A(key_s1[68]), .B(
        new_AGEMA_signal_2599), .S(n211), .Z(new_AGEMA_signal_2600) );
  MUX2_X1 KeyArray_MUX_inS13ser_mux_inst_5_U1_Ins_0_U1 ( .A(key_s0[69]), .B(
        KeyArray_outS20ser[5]), .S(n211), .Z(KeyArray_inS13ser[5]) );
  MUX2_X1 KeyArray_MUX_inS13ser_mux_inst_5_U1_Ins_1_U1 ( .A(key_s1[69]), .B(
        new_AGEMA_signal_2602), .S(n211), .Z(new_AGEMA_signal_2603) );
  MUX2_X1 KeyArray_MUX_inS13ser_mux_inst_6_U1_Ins_0_U1 ( .A(key_s0[70]), .B(
        KeyArray_outS20ser[6]), .S(n211), .Z(KeyArray_inS13ser[6]) );
  MUX2_X1 KeyArray_MUX_inS13ser_mux_inst_6_U1_Ins_1_U1 ( .A(key_s1[70]), .B(
        new_AGEMA_signal_2605), .S(n211), .Z(new_AGEMA_signal_2606) );
  MUX2_X1 KeyArray_MUX_inS13ser_mux_inst_7_U1_Ins_0_U1 ( .A(key_s0[71]), .B(
        KeyArray_outS20ser[7]), .S(n211), .Z(KeyArray_inS13ser[7]) );
  MUX2_X1 KeyArray_MUX_inS13ser_mux_inst_7_U1_Ins_1_U1 ( .A(key_s1[71]), .B(
        new_AGEMA_signal_2608), .S(n211), .Z(new_AGEMA_signal_2609) );
  MUX2_X1 KeyArray_MUX_inS20ser_mux_inst_0_U1_Ins_0_U1 ( .A(key_s0[56]), .B(
        KeyArray_outS21ser[0]), .S(n212), .Z(KeyArray_inS20ser[0]) );
  MUX2_X1 KeyArray_MUX_inS20ser_mux_inst_0_U1_Ins_1_U1 ( .A(key_s1[56]), .B(
        new_AGEMA_signal_2611), .S(n212), .Z(new_AGEMA_signal_2612) );
  MUX2_X1 KeyArray_MUX_inS20ser_mux_inst_1_U1_Ins_0_U1 ( .A(key_s0[57]), .B(
        KeyArray_outS21ser[1]), .S(n212), .Z(KeyArray_inS20ser[1]) );
  MUX2_X1 KeyArray_MUX_inS20ser_mux_inst_1_U1_Ins_1_U1 ( .A(key_s1[57]), .B(
        new_AGEMA_signal_2614), .S(n212), .Z(new_AGEMA_signal_2615) );
  MUX2_X1 KeyArray_MUX_inS20ser_mux_inst_2_U1_Ins_0_U1 ( .A(key_s0[58]), .B(
        KeyArray_outS21ser[2]), .S(n212), .Z(KeyArray_inS20ser[2]) );
  MUX2_X1 KeyArray_MUX_inS20ser_mux_inst_2_U1_Ins_1_U1 ( .A(key_s1[58]), .B(
        new_AGEMA_signal_2617), .S(n212), .Z(new_AGEMA_signal_2618) );
  MUX2_X1 KeyArray_MUX_inS20ser_mux_inst_3_U1_Ins_0_U1 ( .A(key_s0[59]), .B(
        KeyArray_outS21ser[3]), .S(n212), .Z(KeyArray_inS20ser[3]) );
  MUX2_X1 KeyArray_MUX_inS20ser_mux_inst_3_U1_Ins_1_U1 ( .A(key_s1[59]), .B(
        new_AGEMA_signal_2620), .S(n212), .Z(new_AGEMA_signal_2621) );
  MUX2_X1 KeyArray_MUX_inS20ser_mux_inst_4_U1_Ins_0_U1 ( .A(key_s0[60]), .B(
        KeyArray_outS21ser[4]), .S(n212), .Z(KeyArray_inS20ser[4]) );
  MUX2_X1 KeyArray_MUX_inS20ser_mux_inst_4_U1_Ins_1_U1 ( .A(key_s1[60]), .B(
        new_AGEMA_signal_2623), .S(n212), .Z(new_AGEMA_signal_2624) );
  MUX2_X1 KeyArray_MUX_inS20ser_mux_inst_5_U1_Ins_0_U1 ( .A(key_s0[61]), .B(
        KeyArray_outS21ser[5]), .S(n212), .Z(KeyArray_inS20ser[5]) );
  MUX2_X1 KeyArray_MUX_inS20ser_mux_inst_5_U1_Ins_1_U1 ( .A(key_s1[61]), .B(
        new_AGEMA_signal_2626), .S(n212), .Z(new_AGEMA_signal_2627) );
  MUX2_X1 KeyArray_MUX_inS20ser_mux_inst_6_U1_Ins_0_U1 ( .A(key_s0[62]), .B(
        KeyArray_outS21ser[6]), .S(n212), .Z(KeyArray_inS20ser[6]) );
  MUX2_X1 KeyArray_MUX_inS20ser_mux_inst_6_U1_Ins_1_U1 ( .A(key_s1[62]), .B(
        new_AGEMA_signal_2629), .S(n212), .Z(new_AGEMA_signal_2630) );
  MUX2_X1 KeyArray_MUX_inS20ser_mux_inst_7_U1_Ins_0_U1 ( .A(key_s0[63]), .B(
        KeyArray_outS21ser[7]), .S(n213), .Z(KeyArray_inS20ser[7]) );
  MUX2_X1 KeyArray_MUX_inS20ser_mux_inst_7_U1_Ins_1_U1 ( .A(key_s1[63]), .B(
        new_AGEMA_signal_2632), .S(n213), .Z(new_AGEMA_signal_2633) );
  MUX2_X1 KeyArray_MUX_inS21ser_mux_inst_0_U1_Ins_0_U1 ( .A(key_s0[48]), .B(
        KeyArray_outS22ser[0]), .S(n213), .Z(KeyArray_inS21ser[0]) );
  MUX2_X1 KeyArray_MUX_inS21ser_mux_inst_0_U1_Ins_1_U1 ( .A(key_s1[48]), .B(
        new_AGEMA_signal_2635), .S(n213), .Z(new_AGEMA_signal_2636) );
  MUX2_X1 KeyArray_MUX_inS21ser_mux_inst_1_U1_Ins_0_U1 ( .A(key_s0[49]), .B(
        KeyArray_outS22ser[1]), .S(n213), .Z(KeyArray_inS21ser[1]) );
  MUX2_X1 KeyArray_MUX_inS21ser_mux_inst_1_U1_Ins_1_U1 ( .A(key_s1[49]), .B(
        new_AGEMA_signal_2638), .S(n213), .Z(new_AGEMA_signal_2639) );
  MUX2_X1 KeyArray_MUX_inS21ser_mux_inst_2_U1_Ins_0_U1 ( .A(key_s0[50]), .B(
        KeyArray_outS22ser[2]), .S(n213), .Z(KeyArray_inS21ser[2]) );
  MUX2_X1 KeyArray_MUX_inS21ser_mux_inst_2_U1_Ins_1_U1 ( .A(key_s1[50]), .B(
        new_AGEMA_signal_2641), .S(n213), .Z(new_AGEMA_signal_2642) );
  MUX2_X1 KeyArray_MUX_inS21ser_mux_inst_3_U1_Ins_0_U1 ( .A(key_s0[51]), .B(
        KeyArray_outS22ser[3]), .S(n213), .Z(KeyArray_inS21ser[3]) );
  MUX2_X1 KeyArray_MUX_inS21ser_mux_inst_3_U1_Ins_1_U1 ( .A(key_s1[51]), .B(
        new_AGEMA_signal_2644), .S(n213), .Z(new_AGEMA_signal_2645) );
  MUX2_X1 KeyArray_MUX_inS21ser_mux_inst_4_U1_Ins_0_U1 ( .A(key_s0[52]), .B(
        KeyArray_outS22ser[4]), .S(n213), .Z(KeyArray_inS21ser[4]) );
  MUX2_X1 KeyArray_MUX_inS21ser_mux_inst_4_U1_Ins_1_U1 ( .A(key_s1[52]), .B(
        new_AGEMA_signal_2647), .S(n213), .Z(new_AGEMA_signal_2648) );
  MUX2_X1 KeyArray_MUX_inS21ser_mux_inst_5_U1_Ins_0_U1 ( .A(key_s0[53]), .B(
        KeyArray_outS22ser[5]), .S(n214), .Z(KeyArray_inS21ser[5]) );
  MUX2_X1 KeyArray_MUX_inS21ser_mux_inst_5_U1_Ins_1_U1 ( .A(key_s1[53]), .B(
        new_AGEMA_signal_2650), .S(n214), .Z(new_AGEMA_signal_2651) );
  MUX2_X1 KeyArray_MUX_inS21ser_mux_inst_6_U1_Ins_0_U1 ( .A(key_s0[54]), .B(
        KeyArray_outS22ser[6]), .S(n216), .Z(KeyArray_inS21ser[6]) );
  MUX2_X1 KeyArray_MUX_inS21ser_mux_inst_6_U1_Ins_1_U1 ( .A(key_s1[54]), .B(
        new_AGEMA_signal_2653), .S(n216), .Z(new_AGEMA_signal_2654) );
  MUX2_X1 KeyArray_MUX_inS21ser_mux_inst_7_U1_Ins_0_U1 ( .A(key_s0[55]), .B(
        KeyArray_outS22ser[7]), .S(n214), .Z(KeyArray_inS21ser[7]) );
  MUX2_X1 KeyArray_MUX_inS21ser_mux_inst_7_U1_Ins_1_U1 ( .A(key_s1[55]), .B(
        new_AGEMA_signal_2656), .S(n214), .Z(new_AGEMA_signal_2657) );
  MUX2_X1 KeyArray_MUX_inS22ser_mux_inst_0_U1_Ins_0_U1 ( .A(key_s0[40]), .B(
        KeyArray_outS23ser[0]), .S(n214), .Z(KeyArray_inS22ser[0]) );
  MUX2_X1 KeyArray_MUX_inS22ser_mux_inst_0_U1_Ins_1_U1 ( .A(key_s1[40]), .B(
        new_AGEMA_signal_2659), .S(n214), .Z(new_AGEMA_signal_2660) );
  MUX2_X1 KeyArray_MUX_inS22ser_mux_inst_1_U1_Ins_0_U1 ( .A(key_s0[41]), .B(
        KeyArray_outS23ser[1]), .S(n214), .Z(KeyArray_inS22ser[1]) );
  MUX2_X1 KeyArray_MUX_inS22ser_mux_inst_1_U1_Ins_1_U1 ( .A(key_s1[41]), .B(
        new_AGEMA_signal_2662), .S(n214), .Z(new_AGEMA_signal_2663) );
  MUX2_X1 KeyArray_MUX_inS22ser_mux_inst_2_U1_Ins_0_U1 ( .A(key_s0[42]), .B(
        KeyArray_outS23ser[2]), .S(n214), .Z(KeyArray_inS22ser[2]) );
  MUX2_X1 KeyArray_MUX_inS22ser_mux_inst_2_U1_Ins_1_U1 ( .A(key_s1[42]), .B(
        new_AGEMA_signal_2665), .S(n214), .Z(new_AGEMA_signal_2666) );
  MUX2_X1 KeyArray_MUX_inS22ser_mux_inst_3_U1_Ins_0_U1 ( .A(key_s0[43]), .B(
        KeyArray_outS23ser[3]), .S(n214), .Z(KeyArray_inS22ser[3]) );
  MUX2_X1 KeyArray_MUX_inS22ser_mux_inst_3_U1_Ins_1_U1 ( .A(key_s1[43]), .B(
        new_AGEMA_signal_2668), .S(n214), .Z(new_AGEMA_signal_2669) );
  MUX2_X1 KeyArray_MUX_inS22ser_mux_inst_4_U1_Ins_0_U1 ( .A(key_s0[44]), .B(
        KeyArray_outS23ser[4]), .S(n214), .Z(KeyArray_inS22ser[4]) );
  MUX2_X1 KeyArray_MUX_inS22ser_mux_inst_4_U1_Ins_1_U1 ( .A(key_s1[44]), .B(
        new_AGEMA_signal_2671), .S(n214), .Z(new_AGEMA_signal_2672) );
  MUX2_X1 KeyArray_MUX_inS22ser_mux_inst_5_U1_Ins_0_U1 ( .A(key_s0[45]), .B(
        KeyArray_outS23ser[5]), .S(nReset), .Z(KeyArray_inS22ser[5]) );
  MUX2_X1 KeyArray_MUX_inS22ser_mux_inst_5_U1_Ins_1_U1 ( .A(key_s1[45]), .B(
        new_AGEMA_signal_2674), .S(nReset), .Z(new_AGEMA_signal_2675) );
  MUX2_X1 KeyArray_MUX_inS22ser_mux_inst_6_U1_Ins_0_U1 ( .A(key_s0[46]), .B(
        KeyArray_outS23ser[6]), .S(nReset), .Z(KeyArray_inS22ser[6]) );
  MUX2_X1 KeyArray_MUX_inS22ser_mux_inst_6_U1_Ins_1_U1 ( .A(key_s1[46]), .B(
        new_AGEMA_signal_2677), .S(nReset), .Z(new_AGEMA_signal_2678) );
  MUX2_X1 KeyArray_MUX_inS22ser_mux_inst_7_U1_Ins_0_U1 ( .A(key_s0[47]), .B(
        KeyArray_outS23ser[7]), .S(nReset), .Z(KeyArray_inS22ser[7]) );
  MUX2_X1 KeyArray_MUX_inS22ser_mux_inst_7_U1_Ins_1_U1 ( .A(key_s1[47]), .B(
        new_AGEMA_signal_2680), .S(nReset), .Z(new_AGEMA_signal_2681) );
  MUX2_X1 KeyArray_MUX_inS23ser_mux_inst_0_U1_Ins_0_U1 ( .A(key_s0[32]), .B(
        KeyArray_outS30ser[0]), .S(nReset), .Z(KeyArray_inS23ser[0]) );
  MUX2_X1 KeyArray_MUX_inS23ser_mux_inst_0_U1_Ins_1_U1 ( .A(key_s1[32]), .B(
        new_AGEMA_signal_2683), .S(nReset), .Z(new_AGEMA_signal_2684) );
  MUX2_X1 KeyArray_MUX_inS23ser_mux_inst_1_U1_Ins_0_U1 ( .A(key_s0[33]), .B(
        KeyArray_outS30ser[1]), .S(nReset), .Z(KeyArray_inS23ser[1]) );
  MUX2_X1 KeyArray_MUX_inS23ser_mux_inst_1_U1_Ins_1_U1 ( .A(key_s1[33]), .B(
        new_AGEMA_signal_2686), .S(nReset), .Z(new_AGEMA_signal_2687) );
  MUX2_X1 KeyArray_MUX_inS23ser_mux_inst_2_U1_Ins_0_U1 ( .A(key_s0[34]), .B(
        KeyArray_outS30ser[2]), .S(nReset), .Z(KeyArray_inS23ser[2]) );
  MUX2_X1 KeyArray_MUX_inS23ser_mux_inst_2_U1_Ins_1_U1 ( .A(key_s1[34]), .B(
        new_AGEMA_signal_2689), .S(nReset), .Z(new_AGEMA_signal_2690) );
  MUX2_X1 KeyArray_MUX_inS23ser_mux_inst_3_U1_Ins_0_U1 ( .A(key_s0[35]), .B(
        KeyArray_outS30ser[3]), .S(nReset), .Z(KeyArray_inS23ser[3]) );
  MUX2_X1 KeyArray_MUX_inS23ser_mux_inst_3_U1_Ins_1_U1 ( .A(key_s1[35]), .B(
        new_AGEMA_signal_2692), .S(nReset), .Z(new_AGEMA_signal_2693) );
  MUX2_X1 KeyArray_MUX_inS23ser_mux_inst_4_U1_Ins_0_U1 ( .A(key_s0[36]), .B(
        KeyArray_outS30ser[4]), .S(n215), .Z(KeyArray_inS23ser[4]) );
  MUX2_X1 KeyArray_MUX_inS23ser_mux_inst_4_U1_Ins_1_U1 ( .A(key_s1[36]), .B(
        new_AGEMA_signal_2695), .S(n215), .Z(new_AGEMA_signal_2696) );
  MUX2_X1 KeyArray_MUX_inS23ser_mux_inst_5_U1_Ins_0_U1 ( .A(key_s0[37]), .B(
        KeyArray_outS30ser[5]), .S(n215), .Z(KeyArray_inS23ser[5]) );
  MUX2_X1 KeyArray_MUX_inS23ser_mux_inst_5_U1_Ins_1_U1 ( .A(key_s1[37]), .B(
        new_AGEMA_signal_2698), .S(n215), .Z(new_AGEMA_signal_2699) );
  MUX2_X1 KeyArray_MUX_inS23ser_mux_inst_6_U1_Ins_0_U1 ( .A(key_s0[38]), .B(
        KeyArray_outS30ser[6]), .S(n215), .Z(KeyArray_inS23ser[6]) );
  MUX2_X1 KeyArray_MUX_inS23ser_mux_inst_6_U1_Ins_1_U1 ( .A(key_s1[38]), .B(
        new_AGEMA_signal_2701), .S(n215), .Z(new_AGEMA_signal_2702) );
  MUX2_X1 KeyArray_MUX_inS23ser_mux_inst_7_U1_Ins_0_U1 ( .A(key_s0[39]), .B(
        KeyArray_outS30ser[7]), .S(n215), .Z(KeyArray_inS23ser[7]) );
  MUX2_X1 KeyArray_MUX_inS23ser_mux_inst_7_U1_Ins_1_U1 ( .A(key_s1[39]), .B(
        new_AGEMA_signal_2704), .S(n215), .Z(new_AGEMA_signal_2705) );
  MUX2_X1 KeyArray_MUX_inS30ser_mux_inst_0_U1_Ins_0_U1 ( .A(key_s0[24]), .B(
        KeyArray_outS31ser[0]), .S(n215), .Z(KeyArray_inS30ser[0]) );
  MUX2_X1 KeyArray_MUX_inS30ser_mux_inst_0_U1_Ins_1_U1 ( .A(key_s1[24]), .B(
        new_AGEMA_signal_2707), .S(n215), .Z(new_AGEMA_signal_2708) );
  MUX2_X1 KeyArray_MUX_inS30ser_mux_inst_1_U1_Ins_0_U1 ( .A(key_s0[25]), .B(
        KeyArray_outS31ser[1]), .S(n215), .Z(KeyArray_inS30ser[1]) );
  MUX2_X1 KeyArray_MUX_inS30ser_mux_inst_1_U1_Ins_1_U1 ( .A(key_s1[25]), .B(
        new_AGEMA_signal_2710), .S(n215), .Z(new_AGEMA_signal_2711) );
  MUX2_X1 KeyArray_MUX_inS30ser_mux_inst_2_U1_Ins_0_U1 ( .A(key_s0[26]), .B(
        KeyArray_outS31ser[2]), .S(n215), .Z(KeyArray_inS30ser[2]) );
  MUX2_X1 KeyArray_MUX_inS30ser_mux_inst_2_U1_Ins_1_U1 ( .A(key_s1[26]), .B(
        new_AGEMA_signal_2713), .S(n215), .Z(new_AGEMA_signal_2714) );
  MUX2_X1 KeyArray_MUX_inS30ser_mux_inst_3_U1_Ins_0_U1 ( .A(key_s0[27]), .B(
        KeyArray_outS31ser[3]), .S(n216), .Z(KeyArray_inS30ser[3]) );
  MUX2_X1 KeyArray_MUX_inS30ser_mux_inst_3_U1_Ins_1_U1 ( .A(key_s1[27]), .B(
        new_AGEMA_signal_2716), .S(n216), .Z(new_AGEMA_signal_2717) );
  MUX2_X1 KeyArray_MUX_inS30ser_mux_inst_4_U1_Ins_0_U1 ( .A(key_s0[28]), .B(
        KeyArray_outS31ser[4]), .S(n216), .Z(KeyArray_inS30ser[4]) );
  MUX2_X1 KeyArray_MUX_inS30ser_mux_inst_4_U1_Ins_1_U1 ( .A(key_s1[28]), .B(
        new_AGEMA_signal_2719), .S(n216), .Z(new_AGEMA_signal_2720) );
  MUX2_X1 KeyArray_MUX_inS30ser_mux_inst_5_U1_Ins_0_U1 ( .A(key_s0[29]), .B(
        KeyArray_outS31ser[5]), .S(n216), .Z(KeyArray_inS30ser[5]) );
  MUX2_X1 KeyArray_MUX_inS30ser_mux_inst_5_U1_Ins_1_U1 ( .A(key_s1[29]), .B(
        new_AGEMA_signal_2722), .S(n216), .Z(new_AGEMA_signal_2723) );
  MUX2_X1 KeyArray_MUX_inS30ser_mux_inst_6_U1_Ins_0_U1 ( .A(key_s0[30]), .B(
        KeyArray_outS31ser[6]), .S(n216), .Z(KeyArray_inS30ser[6]) );
  MUX2_X1 KeyArray_MUX_inS30ser_mux_inst_6_U1_Ins_1_U1 ( .A(key_s1[30]), .B(
        new_AGEMA_signal_2725), .S(n216), .Z(new_AGEMA_signal_2726) );
  MUX2_X1 KeyArray_MUX_inS30ser_mux_inst_7_U1_Ins_0_U1 ( .A(key_s0[31]), .B(
        KeyArray_outS31ser[7]), .S(n216), .Z(KeyArray_inS30ser[7]) );
  MUX2_X1 KeyArray_MUX_inS30ser_mux_inst_7_U1_Ins_1_U1 ( .A(key_s1[31]), .B(
        new_AGEMA_signal_2728), .S(n216), .Z(new_AGEMA_signal_2729) );
  MUX2_X1 KeyArray_MUX_inS31ser_mux_inst_0_U1_Ins_0_U1 ( .A(key_s0[16]), .B(
        KeyArray_outS32ser[0]), .S(n216), .Z(KeyArray_inS31ser[0]) );
  MUX2_X1 KeyArray_MUX_inS31ser_mux_inst_0_U1_Ins_1_U1 ( .A(key_s1[16]), .B(
        new_AGEMA_signal_2731), .S(n216), .Z(new_AGEMA_signal_2732) );
  MUX2_X1 KeyArray_MUX_inS31ser_mux_inst_1_U1_Ins_0_U1 ( .A(key_s0[17]), .B(
        KeyArray_outS32ser[1]), .S(n216), .Z(KeyArray_inS31ser[1]) );
  MUX2_X1 KeyArray_MUX_inS31ser_mux_inst_1_U1_Ins_1_U1 ( .A(key_s1[17]), .B(
        new_AGEMA_signal_2734), .S(n216), .Z(new_AGEMA_signal_2735) );
  MUX2_X1 KeyArray_MUX_inS31ser_mux_inst_2_U1_Ins_0_U1 ( .A(key_s0[18]), .B(
        KeyArray_outS32ser[2]), .S(n217), .Z(KeyArray_inS31ser[2]) );
  MUX2_X1 KeyArray_MUX_inS31ser_mux_inst_2_U1_Ins_1_U1 ( .A(key_s1[18]), .B(
        new_AGEMA_signal_2737), .S(n217), .Z(new_AGEMA_signal_2738) );
  MUX2_X1 KeyArray_MUX_inS31ser_mux_inst_3_U1_Ins_0_U1 ( .A(key_s0[19]), .B(
        KeyArray_outS32ser[3]), .S(n217), .Z(KeyArray_inS31ser[3]) );
  MUX2_X1 KeyArray_MUX_inS31ser_mux_inst_3_U1_Ins_1_U1 ( .A(key_s1[19]), .B(
        new_AGEMA_signal_2740), .S(n217), .Z(new_AGEMA_signal_2741) );
  MUX2_X1 KeyArray_MUX_inS31ser_mux_inst_4_U1_Ins_0_U1 ( .A(key_s0[20]), .B(
        KeyArray_outS32ser[4]), .S(n217), .Z(KeyArray_inS31ser[4]) );
  MUX2_X1 KeyArray_MUX_inS31ser_mux_inst_4_U1_Ins_1_U1 ( .A(key_s1[20]), .B(
        new_AGEMA_signal_2743), .S(n217), .Z(new_AGEMA_signal_2744) );
  MUX2_X1 KeyArray_MUX_inS31ser_mux_inst_5_U1_Ins_0_U1 ( .A(key_s0[21]), .B(
        KeyArray_outS32ser[5]), .S(n217), .Z(KeyArray_inS31ser[5]) );
  MUX2_X1 KeyArray_MUX_inS31ser_mux_inst_5_U1_Ins_1_U1 ( .A(key_s1[21]), .B(
        new_AGEMA_signal_2746), .S(n217), .Z(new_AGEMA_signal_2747) );
  MUX2_X1 KeyArray_MUX_inS31ser_mux_inst_6_U1_Ins_0_U1 ( .A(key_s0[22]), .B(
        KeyArray_outS32ser[6]), .S(n217), .Z(KeyArray_inS31ser[6]) );
  MUX2_X1 KeyArray_MUX_inS31ser_mux_inst_6_U1_Ins_1_U1 ( .A(key_s1[22]), .B(
        new_AGEMA_signal_2749), .S(n217), .Z(new_AGEMA_signal_2750) );
  MUX2_X1 KeyArray_MUX_inS31ser_mux_inst_7_U1_Ins_0_U1 ( .A(key_s0[23]), .B(
        KeyArray_outS32ser[7]), .S(n217), .Z(KeyArray_inS31ser[7]) );
  MUX2_X1 KeyArray_MUX_inS31ser_mux_inst_7_U1_Ins_1_U1 ( .A(key_s1[23]), .B(
        new_AGEMA_signal_2752), .S(n217), .Z(new_AGEMA_signal_2753) );
  MUX2_X1 KeyArray_MUX_inS32ser_mux_inst_0_U1_Ins_0_U1 ( .A(key_s0[8]), .B(
        KeyArray_outS33ser[0]), .S(n217), .Z(KeyArray_inS32ser[0]) );
  MUX2_X1 KeyArray_MUX_inS32ser_mux_inst_0_U1_Ins_1_U1 ( .A(key_s1[8]), .B(
        new_AGEMA_signal_2755), .S(n217), .Z(new_AGEMA_signal_2756) );
  MUX2_X1 KeyArray_MUX_inS32ser_mux_inst_1_U1_Ins_0_U1 ( .A(key_s0[9]), .B(
        KeyArray_outS33ser[1]), .S(n218), .Z(KeyArray_inS32ser[1]) );
  MUX2_X1 KeyArray_MUX_inS32ser_mux_inst_1_U1_Ins_1_U1 ( .A(key_s1[9]), .B(
        new_AGEMA_signal_2758), .S(n218), .Z(new_AGEMA_signal_2759) );
  MUX2_X1 KeyArray_MUX_inS32ser_mux_inst_2_U1_Ins_0_U1 ( .A(key_s0[10]), .B(
        KeyArray_outS33ser[2]), .S(n218), .Z(KeyArray_inS32ser[2]) );
  MUX2_X1 KeyArray_MUX_inS32ser_mux_inst_2_U1_Ins_1_U1 ( .A(key_s1[10]), .B(
        new_AGEMA_signal_2761), .S(n218), .Z(new_AGEMA_signal_2762) );
  MUX2_X1 KeyArray_MUX_inS32ser_mux_inst_3_U1_Ins_0_U1 ( .A(key_s0[11]), .B(
        KeyArray_outS33ser[3]), .S(n218), .Z(KeyArray_inS32ser[3]) );
  MUX2_X1 KeyArray_MUX_inS32ser_mux_inst_3_U1_Ins_1_U1 ( .A(key_s1[11]), .B(
        new_AGEMA_signal_2764), .S(n218), .Z(new_AGEMA_signal_2765) );
  MUX2_X1 KeyArray_MUX_inS32ser_mux_inst_4_U1_Ins_0_U1 ( .A(key_s0[12]), .B(
        KeyArray_outS33ser[4]), .S(n218), .Z(KeyArray_inS32ser[4]) );
  MUX2_X1 KeyArray_MUX_inS32ser_mux_inst_4_U1_Ins_1_U1 ( .A(key_s1[12]), .B(
        new_AGEMA_signal_2767), .S(n218), .Z(new_AGEMA_signal_2768) );
  MUX2_X1 KeyArray_MUX_inS32ser_mux_inst_5_U1_Ins_0_U1 ( .A(key_s0[13]), .B(
        KeyArray_outS33ser[5]), .S(n218), .Z(KeyArray_inS32ser[5]) );
  MUX2_X1 KeyArray_MUX_inS32ser_mux_inst_5_U1_Ins_1_U1 ( .A(key_s1[13]), .B(
        new_AGEMA_signal_2770), .S(n218), .Z(new_AGEMA_signal_2771) );
  MUX2_X1 KeyArray_MUX_inS32ser_mux_inst_6_U1_Ins_0_U1 ( .A(key_s0[14]), .B(
        KeyArray_outS33ser[6]), .S(n218), .Z(KeyArray_inS32ser[6]) );
  MUX2_X1 KeyArray_MUX_inS32ser_mux_inst_6_U1_Ins_1_U1 ( .A(key_s1[14]), .B(
        new_AGEMA_signal_2773), .S(n218), .Z(new_AGEMA_signal_2774) );
  MUX2_X1 KeyArray_MUX_inS32ser_mux_inst_7_U1_Ins_0_U1 ( .A(key_s0[15]), .B(
        KeyArray_outS33ser[7]), .S(n218), .Z(KeyArray_inS32ser[7]) );
  MUX2_X1 KeyArray_MUX_inS32ser_mux_inst_7_U1_Ins_1_U1 ( .A(key_s1[15]), .B(
        new_AGEMA_signal_2776), .S(n218), .Z(new_AGEMA_signal_2777) );
  MUX2_X1 KeyArray_MUX_inS33ser_mux_inst_0_U1_Ins_0_U1 ( .A(key_s0[0]), .B(
        keyStateIn[0]), .S(n216), .Z(KeyArray_inS33ser[0]) );
  MUX2_X1 KeyArray_MUX_inS33ser_mux_inst_0_U1_Ins_1_U1 ( .A(key_s1[0]), .B(
        new_AGEMA_signal_1983), .S(n216), .Z(new_AGEMA_signal_2779) );
  MUX2_X1 KeyArray_MUX_inS33ser_mux_inst_1_U1_Ins_0_U1 ( .A(key_s0[1]), .B(
        keyStateIn[1]), .S(n215), .Z(KeyArray_inS33ser[1]) );
  MUX2_X1 KeyArray_MUX_inS33ser_mux_inst_1_U1_Ins_1_U1 ( .A(key_s1[1]), .B(
        new_AGEMA_signal_1986), .S(n215), .Z(new_AGEMA_signal_2781) );
  MUX2_X1 KeyArray_MUX_inS33ser_mux_inst_2_U1_Ins_0_U1 ( .A(key_s0[2]), .B(
        keyStateIn[2]), .S(n215), .Z(KeyArray_inS33ser[2]) );
  MUX2_X1 KeyArray_MUX_inS33ser_mux_inst_2_U1_Ins_1_U1 ( .A(key_s1[2]), .B(
        new_AGEMA_signal_1989), .S(n215), .Z(new_AGEMA_signal_2783) );
  MUX2_X1 KeyArray_MUX_inS33ser_mux_inst_3_U1_Ins_0_U1 ( .A(key_s0[3]), .B(
        keyStateIn[3]), .S(n217), .Z(KeyArray_inS33ser[3]) );
  MUX2_X1 KeyArray_MUX_inS33ser_mux_inst_3_U1_Ins_1_U1 ( .A(key_s1[3]), .B(
        new_AGEMA_signal_1992), .S(n217), .Z(new_AGEMA_signal_2785) );
  MUX2_X1 KeyArray_MUX_inS33ser_mux_inst_4_U1_Ins_0_U1 ( .A(key_s0[4]), .B(
        keyStateIn[4]), .S(n205), .Z(KeyArray_inS33ser[4]) );
  MUX2_X1 KeyArray_MUX_inS33ser_mux_inst_4_U1_Ins_1_U1 ( .A(key_s1[4]), .B(
        new_AGEMA_signal_1995), .S(n205), .Z(new_AGEMA_signal_2787) );
  MUX2_X1 KeyArray_MUX_inS33ser_mux_inst_5_U1_Ins_0_U1 ( .A(key_s0[5]), .B(
        keyStateIn[5]), .S(n218), .Z(KeyArray_inS33ser[5]) );
  MUX2_X1 KeyArray_MUX_inS33ser_mux_inst_5_U1_Ins_1_U1 ( .A(key_s1[5]), .B(
        new_AGEMA_signal_1998), .S(n218), .Z(new_AGEMA_signal_2789) );
  MUX2_X1 KeyArray_MUX_inS33ser_mux_inst_6_U1_Ins_0_U1 ( .A(key_s0[6]), .B(
        keyStateIn[6]), .S(n217), .Z(KeyArray_inS33ser[6]) );
  MUX2_X1 KeyArray_MUX_inS33ser_mux_inst_6_U1_Ins_1_U1 ( .A(key_s1[6]), .B(
        new_AGEMA_signal_2001), .S(n217), .Z(new_AGEMA_signal_2791) );
  MUX2_X1 KeyArray_MUX_inS33ser_mux_inst_7_U1_Ins_0_U1 ( .A(key_s0[7]), .B(
        keyStateIn[7]), .S(n214), .Z(KeyArray_inS33ser[7]) );
  MUX2_X1 KeyArray_MUX_inS33ser_mux_inst_7_U1_Ins_1_U1 ( .A(key_s1[7]), .B(
        new_AGEMA_signal_2004), .S(n214), .Z(new_AGEMA_signal_2793) );
  XNOR2_X1 MixColumns_line0_U24_Ins0_U1 ( .A(MixColumns_line0_n16), .B(
        MixColumns_line0_n15), .ZN(MCout[31]) );
  XOR2_X1 MixColumns_line0_U24_Ins_1_U1 ( .A(new_AGEMA_signal_2122), .B(
        new_AGEMA_signal_2024), .Z(new_AGEMA_signal_2794) );
  XNOR2_X1 MixColumns_line0_U23_Ins0_U1 ( .A(ciphertext_s0[63]), .B(
        ciphertext_s0[31]), .ZN(MixColumns_line0_n15) );
  XOR2_X1 MixColumns_line0_U23_Ins_1_U1 ( .A(ciphertext_s1[63]), .B(
        ciphertext_s1[31]), .Z(new_AGEMA_signal_2024) );
  XOR2_X1 MixColumns_line0_U22_Ins_0_U1 ( .A(ciphertext_s0[126]), .B(
        MixColumns_line0_S13[7]), .Z(MixColumns_line0_n16) );
  XOR2_X1 MixColumns_line0_U22_Ins_1_U1 ( .A(ciphertext_s1[126]), .B(
        new_AGEMA_signal_2051), .Z(new_AGEMA_signal_2122) );
  XNOR2_X1 MixColumns_line0_U21_Ins0_U1 ( .A(MixColumns_line0_n14), .B(
        MixColumns_line0_n13), .ZN(MCout[30]) );
  XOR2_X1 MixColumns_line0_U21_Ins_1_U1 ( .A(new_AGEMA_signal_2123), .B(
        new_AGEMA_signal_2027), .Z(new_AGEMA_signal_2795) );
  XNOR2_X1 MixColumns_line0_U20_Ins0_U1 ( .A(ciphertext_s0[62]), .B(
        ciphertext_s0[30]), .ZN(MixColumns_line0_n13) );
  XOR2_X1 MixColumns_line0_U20_Ins_1_U1 ( .A(ciphertext_s1[62]), .B(
        ciphertext_s1[30]), .Z(new_AGEMA_signal_2027) );
  XOR2_X1 MixColumns_line0_U19_Ins_0_U1 ( .A(ciphertext_s0[125]), .B(
        MixColumns_line0_S13[6]), .Z(MixColumns_line0_n14) );
  XOR2_X1 MixColumns_line0_U19_Ins_1_U1 ( .A(ciphertext_s1[125]), .B(
        new_AGEMA_signal_2053), .Z(new_AGEMA_signal_2123) );
  XNOR2_X1 MixColumns_line0_U18_Ins0_U1 ( .A(MixColumns_line0_n12), .B(
        MixColumns_line0_n11), .ZN(MCout[29]) );
  XOR2_X1 MixColumns_line0_U18_Ins_1_U1 ( .A(new_AGEMA_signal_2124), .B(
        new_AGEMA_signal_2030), .Z(new_AGEMA_signal_2796) );
  XNOR2_X1 MixColumns_line0_U17_Ins0_U1 ( .A(ciphertext_s0[61]), .B(
        ciphertext_s0[29]), .ZN(MixColumns_line0_n11) );
  XOR2_X1 MixColumns_line0_U17_Ins_1_U1 ( .A(ciphertext_s1[61]), .B(
        ciphertext_s1[29]), .Z(new_AGEMA_signal_2030) );
  XOR2_X1 MixColumns_line0_U16_Ins_0_U1 ( .A(ciphertext_s0[124]), .B(
        MixColumns_line0_S13[5]), .Z(MixColumns_line0_n12) );
  XOR2_X1 MixColumns_line0_U16_Ins_1_U1 ( .A(ciphertext_s1[124]), .B(
        new_AGEMA_signal_2055), .Z(new_AGEMA_signal_2124) );
  XNOR2_X1 MixColumns_line0_U15_Ins0_U1 ( .A(MixColumns_line0_n10), .B(
        MixColumns_line0_n9), .ZN(MCout[28]) );
  XOR2_X1 MixColumns_line0_U15_Ins_1_U1 ( .A(new_AGEMA_signal_2797), .B(
        new_AGEMA_signal_2033), .Z(new_AGEMA_signal_2838) );
  XNOR2_X1 MixColumns_line0_U14_Ins0_U1 ( .A(ciphertext_s0[60]), .B(
        ciphertext_s0[28]), .ZN(MixColumns_line0_n9) );
  XOR2_X1 MixColumns_line0_U14_Ins_1_U1 ( .A(ciphertext_s1[60]), .B(
        ciphertext_s1[28]), .Z(new_AGEMA_signal_2033) );
  XOR2_X1 MixColumns_line0_U13_Ins_0_U1 ( .A(MixColumns_line0_S02[4]), .B(
        MixColumns_line0_S13[4]), .Z(MixColumns_line0_n10) );
  XOR2_X1 MixColumns_line0_U13_Ins_1_U1 ( .A(new_AGEMA_signal_2046), .B(
        new_AGEMA_signal_2127), .Z(new_AGEMA_signal_2797) );
  XNOR2_X1 MixColumns_line0_U12_Ins0_U1 ( .A(MixColumns_line0_n8), .B(
        MixColumns_line0_n7), .ZN(MCout[27]) );
  XOR2_X1 MixColumns_line0_U12_Ins_1_U1 ( .A(new_AGEMA_signal_2798), .B(
        new_AGEMA_signal_2036), .Z(new_AGEMA_signal_2839) );
  XNOR2_X1 MixColumns_line0_U11_Ins0_U1 ( .A(ciphertext_s0[59]), .B(
        ciphertext_s0[27]), .ZN(MixColumns_line0_n7) );
  XOR2_X1 MixColumns_line0_U11_Ins_1_U1 ( .A(ciphertext_s1[59]), .B(
        ciphertext_s1[27]), .Z(new_AGEMA_signal_2036) );
  XOR2_X1 MixColumns_line0_U10_Ins_0_U1 ( .A(MixColumns_line0_S02[3]), .B(
        MixColumns_line0_S13[3]), .Z(MixColumns_line0_n8) );
  XOR2_X1 MixColumns_line0_U10_Ins_1_U1 ( .A(new_AGEMA_signal_2047), .B(
        new_AGEMA_signal_2128), .Z(new_AGEMA_signal_2798) );
  XNOR2_X1 MixColumns_line0_U9_Ins0_U1 ( .A(MixColumns_line0_n6), .B(
        MixColumns_line0_n5), .ZN(MCout[26]) );
  XOR2_X1 MixColumns_line0_U9_Ins_1_U1 ( .A(new_AGEMA_signal_2125), .B(
        new_AGEMA_signal_2039), .Z(new_AGEMA_signal_2799) );
  XNOR2_X1 MixColumns_line0_U8_Ins0_U1 ( .A(ciphertext_s0[58]), .B(
        ciphertext_s0[26]), .ZN(MixColumns_line0_n5) );
  XOR2_X1 MixColumns_line0_U8_Ins_1_U1 ( .A(ciphertext_s1[58]), .B(
        ciphertext_s1[26]), .Z(new_AGEMA_signal_2039) );
  XOR2_X1 MixColumns_line0_U7_Ins_0_U1 ( .A(ciphertext_s0[121]), .B(
        MixColumns_line0_S13[2]), .Z(MixColumns_line0_n6) );
  XOR2_X1 MixColumns_line0_U7_Ins_1_U1 ( .A(ciphertext_s1[121]), .B(
        new_AGEMA_signal_2058), .Z(new_AGEMA_signal_2125) );
  XNOR2_X1 MixColumns_line0_U6_Ins0_U1 ( .A(MixColumns_line0_n4), .B(
        MixColumns_line0_n3), .ZN(MCout[25]) );
  XOR2_X1 MixColumns_line0_U6_Ins_1_U1 ( .A(new_AGEMA_signal_2800), .B(
        new_AGEMA_signal_2042), .Z(new_AGEMA_signal_2840) );
  XNOR2_X1 MixColumns_line0_U5_Ins0_U1 ( .A(ciphertext_s0[25]), .B(
        ciphertext_s0[57]), .ZN(MixColumns_line0_n3) );
  XOR2_X1 MixColumns_line0_U5_Ins_1_U1 ( .A(ciphertext_s1[25]), .B(
        ciphertext_s1[57]), .Z(new_AGEMA_signal_2042) );
  XOR2_X1 MixColumns_line0_U4_Ins_0_U1 ( .A(MixColumns_line0_S02_1), .B(
        MixColumns_line0_S13[1]), .Z(MixColumns_line0_n4) );
  XOR2_X1 MixColumns_line0_U4_Ins_1_U1 ( .A(new_AGEMA_signal_2048), .B(
        new_AGEMA_signal_2129), .Z(new_AGEMA_signal_2800) );
  XNOR2_X1 MixColumns_line0_U3_Ins0_U1 ( .A(MixColumns_line0_n2), .B(
        MixColumns_line0_n1), .ZN(MCout[24]) );
  XOR2_X1 MixColumns_line0_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2126), .B(
        new_AGEMA_signal_2045), .Z(new_AGEMA_signal_2801) );
  XNOR2_X1 MixColumns_line0_U2_Ins0_U1 ( .A(ciphertext_s0[24]), .B(
        ciphertext_s0[56]), .ZN(MixColumns_line0_n1) );
  XOR2_X1 MixColumns_line0_U2_Ins_1_U1 ( .A(ciphertext_s1[24]), .B(
        ciphertext_s1[56]), .Z(new_AGEMA_signal_2045) );
  XOR2_X1 MixColumns_line0_U1_Ins_0_U1 ( .A(ciphertext_s0[127]), .B(
        MixColumns_line0_S13[0]), .Z(MixColumns_line0_n2) );
  XOR2_X1 MixColumns_line0_U1_Ins_1_U1 ( .A(ciphertext_s1[127]), .B(
        new_AGEMA_signal_2060), .Z(new_AGEMA_signal_2126) );
  XOR2_X1 MixColumns_line0_timesTWO_U3_Ins_0_U1 ( .A(ciphertext_s0[127]), .B(
        ciphertext_s0[123]), .Z(MixColumns_line0_S02[4]) );
  XOR2_X1 MixColumns_line0_timesTWO_U3_Ins_1_U1 ( .A(ciphertext_s1[127]), .B(
        ciphertext_s1[123]), .Z(new_AGEMA_signal_2046) );
  XOR2_X1 MixColumns_line0_timesTWO_U2_Ins_0_U1 ( .A(ciphertext_s0[127]), .B(
        ciphertext_s0[122]), .Z(MixColumns_line0_S02[3]) );
  XOR2_X1 MixColumns_line0_timesTWO_U2_Ins_1_U1 ( .A(ciphertext_s1[127]), .B(
        ciphertext_s1[122]), .Z(new_AGEMA_signal_2047) );
  XOR2_X1 MixColumns_line0_timesTWO_U1_Ins_0_U1 ( .A(ciphertext_s0[127]), .B(
        ciphertext_s0[120]), .Z(MixColumns_line0_S02_1) );
  XOR2_X1 MixColumns_line0_timesTWO_U1_Ins_1_U1 ( .A(ciphertext_s1[127]), .B(
        ciphertext_s1[120]), .Z(new_AGEMA_signal_2048) );
  XOR2_X1 MixColumns_line0_timesTHREE_U8_Ins_0_U1 ( .A(ciphertext_s0[95]), .B(
        ciphertext_s0[94]), .Z(MixColumns_line0_S13[7]) );
  XOR2_X1 MixColumns_line0_timesTHREE_U8_Ins_1_U1 ( .A(ciphertext_s1[95]), .B(
        ciphertext_s1[94]), .Z(new_AGEMA_signal_2051) );
  XOR2_X1 MixColumns_line0_timesTHREE_U7_Ins_0_U1 ( .A(ciphertext_s0[94]), .B(
        ciphertext_s0[93]), .Z(MixColumns_line0_S13[6]) );
  XOR2_X1 MixColumns_line0_timesTHREE_U7_Ins_1_U1 ( .A(ciphertext_s1[94]), .B(
        ciphertext_s1[93]), .Z(new_AGEMA_signal_2053) );
  XOR2_X1 MixColumns_line0_timesTHREE_U6_Ins_0_U1 ( .A(ciphertext_s0[93]), .B(
        ciphertext_s0[92]), .Z(MixColumns_line0_S13[5]) );
  XOR2_X1 MixColumns_line0_timesTHREE_U6_Ins_1_U1 ( .A(ciphertext_s1[93]), .B(
        ciphertext_s1[92]), .Z(new_AGEMA_signal_2055) );
  XOR2_X1 MixColumns_line0_timesTHREE_U5_Ins_0_U1 ( .A(ciphertext_s0[92]), .B(
        MixColumns_line0_timesTHREE_input2[4]), .Z(MixColumns_line0_S13[4]) );
  XOR2_X1 MixColumns_line0_timesTHREE_U5_Ins_1_U1 ( .A(ciphertext_s1[92]), .B(
        new_AGEMA_signal_2062), .Z(new_AGEMA_signal_2127) );
  XOR2_X1 MixColumns_line0_timesTHREE_U4_Ins_0_U1 ( .A(ciphertext_s0[91]), .B(
        MixColumns_line0_timesTHREE_input2[3]), .Z(MixColumns_line0_S13[3]) );
  XOR2_X1 MixColumns_line0_timesTHREE_U4_Ins_1_U1 ( .A(ciphertext_s1[91]), .B(
        new_AGEMA_signal_2063), .Z(new_AGEMA_signal_2128) );
  XOR2_X1 MixColumns_line0_timesTHREE_U3_Ins_0_U1 ( .A(ciphertext_s0[90]), .B(
        ciphertext_s0[89]), .Z(MixColumns_line0_S13[2]) );
  XOR2_X1 MixColumns_line0_timesTHREE_U3_Ins_1_U1 ( .A(ciphertext_s1[90]), .B(
        ciphertext_s1[89]), .Z(new_AGEMA_signal_2058) );
  XOR2_X1 MixColumns_line0_timesTHREE_U2_Ins_0_U1 ( .A(ciphertext_s0[89]), .B(
        MixColumns_line0_timesTHREE_input2_1), .Z(MixColumns_line0_S13[1]) );
  XOR2_X1 MixColumns_line0_timesTHREE_U2_Ins_1_U1 ( .A(ciphertext_s1[89]), .B(
        new_AGEMA_signal_2064), .Z(new_AGEMA_signal_2129) );
  XOR2_X1 MixColumns_line0_timesTHREE_U1_Ins_0_U1 ( .A(ciphertext_s0[88]), .B(
        ciphertext_s0[95]), .Z(MixColumns_line0_S13[0]) );
  XOR2_X1 MixColumns_line0_timesTHREE_U1_Ins_1_U1 ( .A(ciphertext_s1[88]), .B(
        ciphertext_s1[95]), .Z(new_AGEMA_signal_2060) );
  XOR2_X1 MixColumns_line0_timesTHREE_timesTWO_U3_Ins_0_U1 ( .A(
        ciphertext_s0[95]), .B(ciphertext_s0[91]), .Z(
        MixColumns_line0_timesTHREE_input2[4]) );
  XOR2_X1 MixColumns_line0_timesTHREE_timesTWO_U3_Ins_1_U1 ( .A(
        ciphertext_s1[95]), .B(ciphertext_s1[91]), .Z(new_AGEMA_signal_2062)
         );
  XOR2_X1 MixColumns_line0_timesTHREE_timesTWO_U2_Ins_0_U1 ( .A(
        ciphertext_s0[95]), .B(ciphertext_s0[90]), .Z(
        MixColumns_line0_timesTHREE_input2[3]) );
  XOR2_X1 MixColumns_line0_timesTHREE_timesTWO_U2_Ins_1_U1 ( .A(
        ciphertext_s1[95]), .B(ciphertext_s1[90]), .Z(new_AGEMA_signal_2063)
         );
  XOR2_X1 MixColumns_line0_timesTHREE_timesTWO_U1_Ins_0_U1 ( .A(
        ciphertext_s0[95]), .B(ciphertext_s0[88]), .Z(
        MixColumns_line0_timesTHREE_input2_1) );
  XOR2_X1 MixColumns_line0_timesTHREE_timesTWO_U1_Ins_1_U1 ( .A(
        ciphertext_s1[95]), .B(ciphertext_s1[88]), .Z(new_AGEMA_signal_2064)
         );
  XNOR2_X1 MixColumns_line1_U24_Ins0_U1 ( .A(MixColumns_line1_n16), .B(
        MixColumns_line1_n15), .ZN(MCout[23]) );
  XOR2_X1 MixColumns_line1_U24_Ins_1_U1 ( .A(new_AGEMA_signal_2130), .B(
        new_AGEMA_signal_2065), .Z(new_AGEMA_signal_2802) );
  XNOR2_X1 MixColumns_line1_U23_Ins0_U1 ( .A(ciphertext_s0[31]), .B(
        ciphertext_s0[127]), .ZN(MixColumns_line1_n15) );
  XOR2_X1 MixColumns_line1_U23_Ins_1_U1 ( .A(ciphertext_s1[31]), .B(
        ciphertext_s1[127]), .Z(new_AGEMA_signal_2065) );
  XOR2_X1 MixColumns_line1_U22_Ins_0_U1 ( .A(ciphertext_s0[94]), .B(
        MixColumns_line1_S13[7]), .Z(MixColumns_line1_n16) );
  XOR2_X1 MixColumns_line1_U22_Ins_1_U1 ( .A(ciphertext_s1[94]), .B(
        new_AGEMA_signal_2076), .Z(new_AGEMA_signal_2130) );
  XNOR2_X1 MixColumns_line1_U21_Ins0_U1 ( .A(MixColumns_line1_n14), .B(
        MixColumns_line1_n13), .ZN(MCout[22]) );
  XOR2_X1 MixColumns_line1_U21_Ins_1_U1 ( .A(new_AGEMA_signal_2131), .B(
        new_AGEMA_signal_2066), .Z(new_AGEMA_signal_2803) );
  XNOR2_X1 MixColumns_line1_U20_Ins0_U1 ( .A(ciphertext_s0[30]), .B(
        ciphertext_s0[126]), .ZN(MixColumns_line1_n13) );
  XOR2_X1 MixColumns_line1_U20_Ins_1_U1 ( .A(ciphertext_s1[30]), .B(
        ciphertext_s1[126]), .Z(new_AGEMA_signal_2066) );
  XOR2_X1 MixColumns_line1_U19_Ins_0_U1 ( .A(ciphertext_s0[93]), .B(
        MixColumns_line1_S13[6]), .Z(MixColumns_line1_n14) );
  XOR2_X1 MixColumns_line1_U19_Ins_1_U1 ( .A(ciphertext_s1[93]), .B(
        new_AGEMA_signal_2077), .Z(new_AGEMA_signal_2131) );
  XNOR2_X1 MixColumns_line1_U18_Ins0_U1 ( .A(MixColumns_line1_n12), .B(
        MixColumns_line1_n11), .ZN(MCout[21]) );
  XOR2_X1 MixColumns_line1_U18_Ins_1_U1 ( .A(new_AGEMA_signal_2132), .B(
        new_AGEMA_signal_2067), .Z(new_AGEMA_signal_2804) );
  XNOR2_X1 MixColumns_line1_U17_Ins0_U1 ( .A(ciphertext_s0[29]), .B(
        ciphertext_s0[125]), .ZN(MixColumns_line1_n11) );
  XOR2_X1 MixColumns_line1_U17_Ins_1_U1 ( .A(ciphertext_s1[29]), .B(
        ciphertext_s1[125]), .Z(new_AGEMA_signal_2067) );
  XOR2_X1 MixColumns_line1_U16_Ins_0_U1 ( .A(ciphertext_s0[92]), .B(
        MixColumns_line1_S13[5]), .Z(MixColumns_line1_n12) );
  XOR2_X1 MixColumns_line1_U16_Ins_1_U1 ( .A(ciphertext_s1[92]), .B(
        new_AGEMA_signal_2078), .Z(new_AGEMA_signal_2132) );
  XNOR2_X1 MixColumns_line1_U15_Ins0_U1 ( .A(MixColumns_line1_n10), .B(
        MixColumns_line1_n9), .ZN(MCout[20]) );
  XOR2_X1 MixColumns_line1_U15_Ins_1_U1 ( .A(new_AGEMA_signal_2805), .B(
        new_AGEMA_signal_2068), .Z(new_AGEMA_signal_2841) );
  XNOR2_X1 MixColumns_line1_U14_Ins0_U1 ( .A(ciphertext_s0[28]), .B(
        ciphertext_s0[124]), .ZN(MixColumns_line1_n9) );
  XOR2_X1 MixColumns_line1_U14_Ins_1_U1 ( .A(ciphertext_s1[28]), .B(
        ciphertext_s1[124]), .Z(new_AGEMA_signal_2068) );
  XOR2_X1 MixColumns_line1_U13_Ins_0_U1 ( .A(MixColumns_line1_S02_4_), .B(
        MixColumns_line1_S13[4]), .Z(MixColumns_line1_n10) );
  XOR2_X1 MixColumns_line1_U13_Ins_1_U1 ( .A(new_AGEMA_signal_2073), .B(
        new_AGEMA_signal_2135), .Z(new_AGEMA_signal_2805) );
  XNOR2_X1 MixColumns_line1_U12_Ins0_U1 ( .A(MixColumns_line1_n8), .B(
        MixColumns_line1_n7), .ZN(MCout[19]) );
  XOR2_X1 MixColumns_line1_U12_Ins_1_U1 ( .A(new_AGEMA_signal_2806), .B(
        new_AGEMA_signal_2069), .Z(new_AGEMA_signal_2842) );
  XNOR2_X1 MixColumns_line1_U11_Ins0_U1 ( .A(ciphertext_s0[27]), .B(
        ciphertext_s0[123]), .ZN(MixColumns_line1_n7) );
  XOR2_X1 MixColumns_line1_U11_Ins_1_U1 ( .A(ciphertext_s1[27]), .B(
        ciphertext_s1[123]), .Z(new_AGEMA_signal_2069) );
  XOR2_X1 MixColumns_line1_U10_Ins_0_U1 ( .A(MixColumns_line1_S02_3_), .B(
        MixColumns_line1_S13[3]), .Z(MixColumns_line1_n8) );
  XOR2_X1 MixColumns_line1_U10_Ins_1_U1 ( .A(new_AGEMA_signal_2074), .B(
        new_AGEMA_signal_2136), .Z(new_AGEMA_signal_2806) );
  XNOR2_X1 MixColumns_line1_U9_Ins0_U1 ( .A(MixColumns_line1_n6), .B(
        MixColumns_line1_n5), .ZN(MCout[18]) );
  XOR2_X1 MixColumns_line1_U9_Ins_1_U1 ( .A(new_AGEMA_signal_2133), .B(
        new_AGEMA_signal_2070), .Z(new_AGEMA_signal_2807) );
  XNOR2_X1 MixColumns_line1_U8_Ins0_U1 ( .A(ciphertext_s0[26]), .B(
        ciphertext_s0[122]), .ZN(MixColumns_line1_n5) );
  XOR2_X1 MixColumns_line1_U8_Ins_1_U1 ( .A(ciphertext_s1[26]), .B(
        ciphertext_s1[122]), .Z(new_AGEMA_signal_2070) );
  XOR2_X1 MixColumns_line1_U7_Ins_0_U1 ( .A(ciphertext_s0[89]), .B(
        MixColumns_line1_S13[2]), .Z(MixColumns_line1_n6) );
  XOR2_X1 MixColumns_line1_U7_Ins_1_U1 ( .A(ciphertext_s1[89]), .B(
        new_AGEMA_signal_2079), .Z(new_AGEMA_signal_2133) );
  XNOR2_X1 MixColumns_line1_U6_Ins0_U1 ( .A(MixColumns_line1_n4), .B(
        MixColumns_line1_n3), .ZN(MCout[17]) );
  XOR2_X1 MixColumns_line1_U6_Ins_1_U1 ( .A(new_AGEMA_signal_2808), .B(
        new_AGEMA_signal_2071), .Z(new_AGEMA_signal_2843) );
  XNOR2_X1 MixColumns_line1_U5_Ins0_U1 ( .A(ciphertext_s0[121]), .B(
        ciphertext_s0[25]), .ZN(MixColumns_line1_n3) );
  XOR2_X1 MixColumns_line1_U5_Ins_1_U1 ( .A(ciphertext_s1[121]), .B(
        ciphertext_s1[25]), .Z(new_AGEMA_signal_2071) );
  XOR2_X1 MixColumns_line1_U4_Ins_0_U1 ( .A(MixColumns_line1_S02_1_), .B(
        MixColumns_line1_S13[1]), .Z(MixColumns_line1_n4) );
  XOR2_X1 MixColumns_line1_U4_Ins_1_U1 ( .A(new_AGEMA_signal_2075), .B(
        new_AGEMA_signal_2137), .Z(new_AGEMA_signal_2808) );
  XNOR2_X1 MixColumns_line1_U3_Ins0_U1 ( .A(MixColumns_line1_n2), .B(
        MixColumns_line1_n1), .ZN(MCout[16]) );
  XOR2_X1 MixColumns_line1_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2134), .B(
        new_AGEMA_signal_2072), .Z(new_AGEMA_signal_2809) );
  XNOR2_X1 MixColumns_line1_U2_Ins0_U1 ( .A(ciphertext_s0[120]), .B(
        ciphertext_s0[24]), .ZN(MixColumns_line1_n1) );
  XOR2_X1 MixColumns_line1_U2_Ins_1_U1 ( .A(ciphertext_s1[120]), .B(
        ciphertext_s1[24]), .Z(new_AGEMA_signal_2072) );
  XOR2_X1 MixColumns_line1_U1_Ins_0_U1 ( .A(ciphertext_s0[95]), .B(
        MixColumns_line1_S13[0]), .Z(MixColumns_line1_n2) );
  XOR2_X1 MixColumns_line1_U1_Ins_1_U1 ( .A(ciphertext_s1[95]), .B(
        new_AGEMA_signal_2080), .Z(new_AGEMA_signal_2134) );
  XOR2_X1 MixColumns_line1_timesTWO_U3_Ins_0_U1 ( .A(ciphertext_s0[95]), .B(
        ciphertext_s0[91]), .Z(MixColumns_line1_S02_4_) );
  XOR2_X1 MixColumns_line1_timesTWO_U3_Ins_1_U1 ( .A(ciphertext_s1[95]), .B(
        ciphertext_s1[91]), .Z(new_AGEMA_signal_2073) );
  XOR2_X1 MixColumns_line1_timesTWO_U2_Ins_0_U1 ( .A(ciphertext_s0[95]), .B(
        ciphertext_s0[90]), .Z(MixColumns_line1_S02_3_) );
  XOR2_X1 MixColumns_line1_timesTWO_U2_Ins_1_U1 ( .A(ciphertext_s1[95]), .B(
        ciphertext_s1[90]), .Z(new_AGEMA_signal_2074) );
  XOR2_X1 MixColumns_line1_timesTWO_U1_Ins_0_U1 ( .A(ciphertext_s0[95]), .B(
        ciphertext_s0[88]), .Z(MixColumns_line1_S02_1_) );
  XOR2_X1 MixColumns_line1_timesTWO_U1_Ins_1_U1 ( .A(ciphertext_s1[95]), .B(
        ciphertext_s1[88]), .Z(new_AGEMA_signal_2075) );
  XOR2_X1 MixColumns_line1_timesTHREE_U8_Ins_0_U1 ( .A(ciphertext_s0[63]), .B(
        ciphertext_s0[62]), .Z(MixColumns_line1_S13[7]) );
  XOR2_X1 MixColumns_line1_timesTHREE_U8_Ins_1_U1 ( .A(ciphertext_s1[63]), .B(
        ciphertext_s1[62]), .Z(new_AGEMA_signal_2076) );
  XOR2_X1 MixColumns_line1_timesTHREE_U7_Ins_0_U1 ( .A(ciphertext_s0[62]), .B(
        ciphertext_s0[61]), .Z(MixColumns_line1_S13[6]) );
  XOR2_X1 MixColumns_line1_timesTHREE_U7_Ins_1_U1 ( .A(ciphertext_s1[62]), .B(
        ciphertext_s1[61]), .Z(new_AGEMA_signal_2077) );
  XOR2_X1 MixColumns_line1_timesTHREE_U6_Ins_0_U1 ( .A(ciphertext_s0[61]), .B(
        ciphertext_s0[60]), .Z(MixColumns_line1_S13[5]) );
  XOR2_X1 MixColumns_line1_timesTHREE_U6_Ins_1_U1 ( .A(ciphertext_s1[61]), .B(
        ciphertext_s1[60]), .Z(new_AGEMA_signal_2078) );
  XOR2_X1 MixColumns_line1_timesTHREE_U5_Ins_0_U1 ( .A(ciphertext_s0[60]), .B(
        MixColumns_line1_timesTHREE_input2[4]), .Z(MixColumns_line1_S13[4]) );
  XOR2_X1 MixColumns_line1_timesTHREE_U5_Ins_1_U1 ( .A(ciphertext_s1[60]), .B(
        new_AGEMA_signal_2081), .Z(new_AGEMA_signal_2135) );
  XOR2_X1 MixColumns_line1_timesTHREE_U4_Ins_0_U1 ( .A(ciphertext_s0[59]), .B(
        MixColumns_line1_timesTHREE_input2[3]), .Z(MixColumns_line1_S13[3]) );
  XOR2_X1 MixColumns_line1_timesTHREE_U4_Ins_1_U1 ( .A(ciphertext_s1[59]), .B(
        new_AGEMA_signal_2082), .Z(new_AGEMA_signal_2136) );
  XOR2_X1 MixColumns_line1_timesTHREE_U3_Ins_0_U1 ( .A(ciphertext_s0[58]), .B(
        ciphertext_s0[57]), .Z(MixColumns_line1_S13[2]) );
  XOR2_X1 MixColumns_line1_timesTHREE_U3_Ins_1_U1 ( .A(ciphertext_s1[58]), .B(
        ciphertext_s1[57]), .Z(new_AGEMA_signal_2079) );
  XOR2_X1 MixColumns_line1_timesTHREE_U2_Ins_0_U1 ( .A(ciphertext_s0[57]), .B(
        MixColumns_line1_timesTHREE_input2_1), .Z(MixColumns_line1_S13[1]) );
  XOR2_X1 MixColumns_line1_timesTHREE_U2_Ins_1_U1 ( .A(ciphertext_s1[57]), .B(
        new_AGEMA_signal_2083), .Z(new_AGEMA_signal_2137) );
  XOR2_X1 MixColumns_line1_timesTHREE_U1_Ins_0_U1 ( .A(ciphertext_s0[56]), .B(
        ciphertext_s0[63]), .Z(MixColumns_line1_S13[0]) );
  XOR2_X1 MixColumns_line1_timesTHREE_U1_Ins_1_U1 ( .A(ciphertext_s1[56]), .B(
        ciphertext_s1[63]), .Z(new_AGEMA_signal_2080) );
  XOR2_X1 MixColumns_line1_timesTHREE_timesTWO_U3_Ins_0_U1 ( .A(
        ciphertext_s0[63]), .B(ciphertext_s0[59]), .Z(
        MixColumns_line1_timesTHREE_input2[4]) );
  XOR2_X1 MixColumns_line1_timesTHREE_timesTWO_U3_Ins_1_U1 ( .A(
        ciphertext_s1[63]), .B(ciphertext_s1[59]), .Z(new_AGEMA_signal_2081)
         );
  XOR2_X1 MixColumns_line1_timesTHREE_timesTWO_U2_Ins_0_U1 ( .A(
        ciphertext_s0[63]), .B(ciphertext_s0[58]), .Z(
        MixColumns_line1_timesTHREE_input2[3]) );
  XOR2_X1 MixColumns_line1_timesTHREE_timesTWO_U2_Ins_1_U1 ( .A(
        ciphertext_s1[63]), .B(ciphertext_s1[58]), .Z(new_AGEMA_signal_2082)
         );
  XOR2_X1 MixColumns_line1_timesTHREE_timesTWO_U1_Ins_0_U1 ( .A(
        ciphertext_s0[63]), .B(ciphertext_s0[56]), .Z(
        MixColumns_line1_timesTHREE_input2_1) );
  XOR2_X1 MixColumns_line1_timesTHREE_timesTWO_U1_Ins_1_U1 ( .A(
        ciphertext_s1[63]), .B(ciphertext_s1[56]), .Z(new_AGEMA_signal_2083)
         );
  XNOR2_X1 MixColumns_line2_U24_Ins0_U1 ( .A(MixColumns_line2_n16), .B(
        MixColumns_line2_n15), .ZN(MCout[15]) );
  XOR2_X1 MixColumns_line2_U24_Ins_1_U1 ( .A(new_AGEMA_signal_2138), .B(
        new_AGEMA_signal_2084), .Z(new_AGEMA_signal_2810) );
  XNOR2_X1 MixColumns_line2_U23_Ins0_U1 ( .A(ciphertext_s0[127]), .B(
        ciphertext_s0[95]), .ZN(MixColumns_line2_n15) );
  XOR2_X1 MixColumns_line2_U23_Ins_1_U1 ( .A(ciphertext_s1[127]), .B(
        ciphertext_s1[95]), .Z(new_AGEMA_signal_2084) );
  XOR2_X1 MixColumns_line2_U22_Ins_0_U1 ( .A(ciphertext_s0[62]), .B(
        MixColumns_line2_S13[7]), .Z(MixColumns_line2_n16) );
  XOR2_X1 MixColumns_line2_U22_Ins_1_U1 ( .A(ciphertext_s1[62]), .B(
        new_AGEMA_signal_2095), .Z(new_AGEMA_signal_2138) );
  XNOR2_X1 MixColumns_line2_U21_Ins0_U1 ( .A(MixColumns_line2_n14), .B(
        MixColumns_line2_n13), .ZN(MCout[14]) );
  XOR2_X1 MixColumns_line2_U21_Ins_1_U1 ( .A(new_AGEMA_signal_2139), .B(
        new_AGEMA_signal_2085), .Z(new_AGEMA_signal_2811) );
  XNOR2_X1 MixColumns_line2_U20_Ins0_U1 ( .A(ciphertext_s0[126]), .B(
        ciphertext_s0[94]), .ZN(MixColumns_line2_n13) );
  XOR2_X1 MixColumns_line2_U20_Ins_1_U1 ( .A(ciphertext_s1[126]), .B(
        ciphertext_s1[94]), .Z(new_AGEMA_signal_2085) );
  XOR2_X1 MixColumns_line2_U19_Ins_0_U1 ( .A(ciphertext_s0[61]), .B(
        MixColumns_line2_S13[6]), .Z(MixColumns_line2_n14) );
  XOR2_X1 MixColumns_line2_U19_Ins_1_U1 ( .A(ciphertext_s1[61]), .B(
        new_AGEMA_signal_2096), .Z(new_AGEMA_signal_2139) );
  XNOR2_X1 MixColumns_line2_U18_Ins0_U1 ( .A(MixColumns_line2_n12), .B(
        MixColumns_line2_n11), .ZN(MCout[13]) );
  XOR2_X1 MixColumns_line2_U18_Ins_1_U1 ( .A(new_AGEMA_signal_2140), .B(
        new_AGEMA_signal_2086), .Z(new_AGEMA_signal_2812) );
  XNOR2_X1 MixColumns_line2_U17_Ins0_U1 ( .A(ciphertext_s0[125]), .B(
        ciphertext_s0[93]), .ZN(MixColumns_line2_n11) );
  XOR2_X1 MixColumns_line2_U17_Ins_1_U1 ( .A(ciphertext_s1[125]), .B(
        ciphertext_s1[93]), .Z(new_AGEMA_signal_2086) );
  XOR2_X1 MixColumns_line2_U16_Ins_0_U1 ( .A(ciphertext_s0[60]), .B(
        MixColumns_line2_S13[5]), .Z(MixColumns_line2_n12) );
  XOR2_X1 MixColumns_line2_U16_Ins_1_U1 ( .A(ciphertext_s1[60]), .B(
        new_AGEMA_signal_2097), .Z(new_AGEMA_signal_2140) );
  XNOR2_X1 MixColumns_line2_U15_Ins0_U1 ( .A(MixColumns_line2_n10), .B(
        MixColumns_line2_n9), .ZN(MCout[12]) );
  XOR2_X1 MixColumns_line2_U15_Ins_1_U1 ( .A(new_AGEMA_signal_2813), .B(
        new_AGEMA_signal_2087), .Z(new_AGEMA_signal_2844) );
  XNOR2_X1 MixColumns_line2_U14_Ins0_U1 ( .A(ciphertext_s0[124]), .B(
        ciphertext_s0[92]), .ZN(MixColumns_line2_n9) );
  XOR2_X1 MixColumns_line2_U14_Ins_1_U1 ( .A(ciphertext_s1[124]), .B(
        ciphertext_s1[92]), .Z(new_AGEMA_signal_2087) );
  XOR2_X1 MixColumns_line2_U13_Ins_0_U1 ( .A(MixColumns_line2_S02_4_), .B(
        MixColumns_line2_S13[4]), .Z(MixColumns_line2_n10) );
  XOR2_X1 MixColumns_line2_U13_Ins_1_U1 ( .A(new_AGEMA_signal_2092), .B(
        new_AGEMA_signal_2143), .Z(new_AGEMA_signal_2813) );
  XNOR2_X1 MixColumns_line2_U12_Ins0_U1 ( .A(MixColumns_line2_n8), .B(
        MixColumns_line2_n7), .ZN(MCout[11]) );
  XOR2_X1 MixColumns_line2_U12_Ins_1_U1 ( .A(new_AGEMA_signal_2814), .B(
        new_AGEMA_signal_2088), .Z(new_AGEMA_signal_2845) );
  XNOR2_X1 MixColumns_line2_U11_Ins0_U1 ( .A(ciphertext_s0[123]), .B(
        ciphertext_s0[91]), .ZN(MixColumns_line2_n7) );
  XOR2_X1 MixColumns_line2_U11_Ins_1_U1 ( .A(ciphertext_s1[123]), .B(
        ciphertext_s1[91]), .Z(new_AGEMA_signal_2088) );
  XOR2_X1 MixColumns_line2_U10_Ins_0_U1 ( .A(MixColumns_line2_S02_3_), .B(
        MixColumns_line2_S13[3]), .Z(MixColumns_line2_n8) );
  XOR2_X1 MixColumns_line2_U10_Ins_1_U1 ( .A(new_AGEMA_signal_2093), .B(
        new_AGEMA_signal_2144), .Z(new_AGEMA_signal_2814) );
  XNOR2_X1 MixColumns_line2_U9_Ins0_U1 ( .A(MixColumns_line2_n6), .B(
        MixColumns_line2_n5), .ZN(MCout[10]) );
  XOR2_X1 MixColumns_line2_U9_Ins_1_U1 ( .A(new_AGEMA_signal_2141), .B(
        new_AGEMA_signal_2089), .Z(new_AGEMA_signal_2815) );
  XNOR2_X1 MixColumns_line2_U8_Ins0_U1 ( .A(ciphertext_s0[122]), .B(
        ciphertext_s0[90]), .ZN(MixColumns_line2_n5) );
  XOR2_X1 MixColumns_line2_U8_Ins_1_U1 ( .A(ciphertext_s1[122]), .B(
        ciphertext_s1[90]), .Z(new_AGEMA_signal_2089) );
  XOR2_X1 MixColumns_line2_U7_Ins_0_U1 ( .A(ciphertext_s0[57]), .B(
        MixColumns_line2_S13[2]), .Z(MixColumns_line2_n6) );
  XOR2_X1 MixColumns_line2_U7_Ins_1_U1 ( .A(ciphertext_s1[57]), .B(
        new_AGEMA_signal_2098), .Z(new_AGEMA_signal_2141) );
  XNOR2_X1 MixColumns_line2_U6_Ins0_U1 ( .A(MixColumns_line2_n4), .B(
        MixColumns_line2_n3), .ZN(MCout[9]) );
  XOR2_X1 MixColumns_line2_U6_Ins_1_U1 ( .A(new_AGEMA_signal_2816), .B(
        new_AGEMA_signal_2090), .Z(new_AGEMA_signal_2846) );
  XNOR2_X1 MixColumns_line2_U5_Ins0_U1 ( .A(ciphertext_s0[89]), .B(
        ciphertext_s0[121]), .ZN(MixColumns_line2_n3) );
  XOR2_X1 MixColumns_line2_U5_Ins_1_U1 ( .A(ciphertext_s1[89]), .B(
        ciphertext_s1[121]), .Z(new_AGEMA_signal_2090) );
  XOR2_X1 MixColumns_line2_U4_Ins_0_U1 ( .A(MixColumns_line2_S02_1_), .B(
        MixColumns_line2_S13[1]), .Z(MixColumns_line2_n4) );
  XOR2_X1 MixColumns_line2_U4_Ins_1_U1 ( .A(new_AGEMA_signal_2094), .B(
        new_AGEMA_signal_2145), .Z(new_AGEMA_signal_2816) );
  XNOR2_X1 MixColumns_line2_U3_Ins0_U1 ( .A(MixColumns_line2_n2), .B(
        MixColumns_line2_n1), .ZN(MCout[8]) );
  XOR2_X1 MixColumns_line2_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2142), .B(
        new_AGEMA_signal_2091), .Z(new_AGEMA_signal_2817) );
  XNOR2_X1 MixColumns_line2_U2_Ins0_U1 ( .A(ciphertext_s0[88]), .B(
        ciphertext_s0[120]), .ZN(MixColumns_line2_n1) );
  XOR2_X1 MixColumns_line2_U2_Ins_1_U1 ( .A(ciphertext_s1[88]), .B(
        ciphertext_s1[120]), .Z(new_AGEMA_signal_2091) );
  XOR2_X1 MixColumns_line2_U1_Ins_0_U1 ( .A(ciphertext_s0[63]), .B(
        MixColumns_line2_S13[0]), .Z(MixColumns_line2_n2) );
  XOR2_X1 MixColumns_line2_U1_Ins_1_U1 ( .A(ciphertext_s1[63]), .B(
        new_AGEMA_signal_2099), .Z(new_AGEMA_signal_2142) );
  XOR2_X1 MixColumns_line2_timesTWO_U3_Ins_0_U1 ( .A(ciphertext_s0[63]), .B(
        ciphertext_s0[59]), .Z(MixColumns_line2_S02_4_) );
  XOR2_X1 MixColumns_line2_timesTWO_U3_Ins_1_U1 ( .A(ciphertext_s1[63]), .B(
        ciphertext_s1[59]), .Z(new_AGEMA_signal_2092) );
  XOR2_X1 MixColumns_line2_timesTWO_U2_Ins_0_U1 ( .A(ciphertext_s0[63]), .B(
        ciphertext_s0[58]), .Z(MixColumns_line2_S02_3_) );
  XOR2_X1 MixColumns_line2_timesTWO_U2_Ins_1_U1 ( .A(ciphertext_s1[63]), .B(
        ciphertext_s1[58]), .Z(new_AGEMA_signal_2093) );
  XOR2_X1 MixColumns_line2_timesTWO_U1_Ins_0_U1 ( .A(ciphertext_s0[63]), .B(
        ciphertext_s0[56]), .Z(MixColumns_line2_S02_1_) );
  XOR2_X1 MixColumns_line2_timesTWO_U1_Ins_1_U1 ( .A(ciphertext_s1[63]), .B(
        ciphertext_s1[56]), .Z(new_AGEMA_signal_2094) );
  XOR2_X1 MixColumns_line2_timesTHREE_U8_Ins_0_U1 ( .A(ciphertext_s0[31]), .B(
        ciphertext_s0[30]), .Z(MixColumns_line2_S13[7]) );
  XOR2_X1 MixColumns_line2_timesTHREE_U8_Ins_1_U1 ( .A(ciphertext_s1[31]), .B(
        ciphertext_s1[30]), .Z(new_AGEMA_signal_2095) );
  XOR2_X1 MixColumns_line2_timesTHREE_U7_Ins_0_U1 ( .A(ciphertext_s0[30]), .B(
        ciphertext_s0[29]), .Z(MixColumns_line2_S13[6]) );
  XOR2_X1 MixColumns_line2_timesTHREE_U7_Ins_1_U1 ( .A(ciphertext_s1[30]), .B(
        ciphertext_s1[29]), .Z(new_AGEMA_signal_2096) );
  XOR2_X1 MixColumns_line2_timesTHREE_U6_Ins_0_U1 ( .A(ciphertext_s0[29]), .B(
        ciphertext_s0[28]), .Z(MixColumns_line2_S13[5]) );
  XOR2_X1 MixColumns_line2_timesTHREE_U6_Ins_1_U1 ( .A(ciphertext_s1[29]), .B(
        ciphertext_s1[28]), .Z(new_AGEMA_signal_2097) );
  XOR2_X1 MixColumns_line2_timesTHREE_U5_Ins_0_U1 ( .A(ciphertext_s0[28]), .B(
        MixColumns_line2_timesTHREE_input2[4]), .Z(MixColumns_line2_S13[4]) );
  XOR2_X1 MixColumns_line2_timesTHREE_U5_Ins_1_U1 ( .A(ciphertext_s1[28]), .B(
        new_AGEMA_signal_2100), .Z(new_AGEMA_signal_2143) );
  XOR2_X1 MixColumns_line2_timesTHREE_U4_Ins_0_U1 ( .A(ciphertext_s0[27]), .B(
        MixColumns_line2_timesTHREE_input2[3]), .Z(MixColumns_line2_S13[3]) );
  XOR2_X1 MixColumns_line2_timesTHREE_U4_Ins_1_U1 ( .A(ciphertext_s1[27]), .B(
        new_AGEMA_signal_2101), .Z(new_AGEMA_signal_2144) );
  XOR2_X1 MixColumns_line2_timesTHREE_U3_Ins_0_U1 ( .A(ciphertext_s0[26]), .B(
        ciphertext_s0[25]), .Z(MixColumns_line2_S13[2]) );
  XOR2_X1 MixColumns_line2_timesTHREE_U3_Ins_1_U1 ( .A(ciphertext_s1[26]), .B(
        ciphertext_s1[25]), .Z(new_AGEMA_signal_2098) );
  XOR2_X1 MixColumns_line2_timesTHREE_U2_Ins_0_U1 ( .A(ciphertext_s0[25]), .B(
        MixColumns_line2_timesTHREE_input2_1), .Z(MixColumns_line2_S13[1]) );
  XOR2_X1 MixColumns_line2_timesTHREE_U2_Ins_1_U1 ( .A(ciphertext_s1[25]), .B(
        new_AGEMA_signal_2102), .Z(new_AGEMA_signal_2145) );
  XOR2_X1 MixColumns_line2_timesTHREE_U1_Ins_0_U1 ( .A(ciphertext_s0[24]), .B(
        ciphertext_s0[31]), .Z(MixColumns_line2_S13[0]) );
  XOR2_X1 MixColumns_line2_timesTHREE_U1_Ins_1_U1 ( .A(ciphertext_s1[24]), .B(
        ciphertext_s1[31]), .Z(new_AGEMA_signal_2099) );
  XOR2_X1 MixColumns_line2_timesTHREE_timesTWO_U3_Ins_0_U1 ( .A(
        ciphertext_s0[31]), .B(ciphertext_s0[27]), .Z(
        MixColumns_line2_timesTHREE_input2[4]) );
  XOR2_X1 MixColumns_line2_timesTHREE_timesTWO_U3_Ins_1_U1 ( .A(
        ciphertext_s1[31]), .B(ciphertext_s1[27]), .Z(new_AGEMA_signal_2100)
         );
  XOR2_X1 MixColumns_line2_timesTHREE_timesTWO_U2_Ins_0_U1 ( .A(
        ciphertext_s0[31]), .B(ciphertext_s0[26]), .Z(
        MixColumns_line2_timesTHREE_input2[3]) );
  XOR2_X1 MixColumns_line2_timesTHREE_timesTWO_U2_Ins_1_U1 ( .A(
        ciphertext_s1[31]), .B(ciphertext_s1[26]), .Z(new_AGEMA_signal_2101)
         );
  XOR2_X1 MixColumns_line2_timesTHREE_timesTWO_U1_Ins_0_U1 ( .A(
        ciphertext_s0[31]), .B(ciphertext_s0[24]), .Z(
        MixColumns_line2_timesTHREE_input2_1) );
  XOR2_X1 MixColumns_line2_timesTHREE_timesTWO_U1_Ins_1_U1 ( .A(
        ciphertext_s1[31]), .B(ciphertext_s1[24]), .Z(new_AGEMA_signal_2102)
         );
  XNOR2_X1 MixColumns_line3_U24_Ins0_U1 ( .A(MixColumns_line3_n16), .B(
        MixColumns_line3_n15), .ZN(MCout[7]) );
  XOR2_X1 MixColumns_line3_U24_Ins_1_U1 ( .A(new_AGEMA_signal_2146), .B(
        new_AGEMA_signal_2103), .Z(new_AGEMA_signal_2818) );
  XNOR2_X1 MixColumns_line3_U23_Ins0_U1 ( .A(ciphertext_s0[95]), .B(
        ciphertext_s0[63]), .ZN(MixColumns_line3_n15) );
  XOR2_X1 MixColumns_line3_U23_Ins_1_U1 ( .A(ciphertext_s1[95]), .B(
        ciphertext_s1[63]), .Z(new_AGEMA_signal_2103) );
  XOR2_X1 MixColumns_line3_U22_Ins_0_U1 ( .A(ciphertext_s0[30]), .B(
        MixColumns_line3_S13[7]), .Z(MixColumns_line3_n16) );
  XOR2_X1 MixColumns_line3_U22_Ins_1_U1 ( .A(ciphertext_s1[30]), .B(
        new_AGEMA_signal_2114), .Z(new_AGEMA_signal_2146) );
  XNOR2_X1 MixColumns_line3_U21_Ins0_U1 ( .A(MixColumns_line3_n14), .B(
        MixColumns_line3_n13), .ZN(MCout[6]) );
  XOR2_X1 MixColumns_line3_U21_Ins_1_U1 ( .A(new_AGEMA_signal_2147), .B(
        new_AGEMA_signal_2104), .Z(new_AGEMA_signal_2819) );
  XNOR2_X1 MixColumns_line3_U20_Ins0_U1 ( .A(ciphertext_s0[94]), .B(
        ciphertext_s0[62]), .ZN(MixColumns_line3_n13) );
  XOR2_X1 MixColumns_line3_U20_Ins_1_U1 ( .A(ciphertext_s1[94]), .B(
        ciphertext_s1[62]), .Z(new_AGEMA_signal_2104) );
  XOR2_X1 MixColumns_line3_U19_Ins_0_U1 ( .A(ciphertext_s0[29]), .B(
        MixColumns_line3_S13[6]), .Z(MixColumns_line3_n14) );
  XOR2_X1 MixColumns_line3_U19_Ins_1_U1 ( .A(ciphertext_s1[29]), .B(
        new_AGEMA_signal_2115), .Z(new_AGEMA_signal_2147) );
  XNOR2_X1 MixColumns_line3_U18_Ins0_U1 ( .A(MixColumns_line3_n12), .B(
        MixColumns_line3_n11), .ZN(MCout[5]) );
  XOR2_X1 MixColumns_line3_U18_Ins_1_U1 ( .A(new_AGEMA_signal_2148), .B(
        new_AGEMA_signal_2105), .Z(new_AGEMA_signal_2820) );
  XNOR2_X1 MixColumns_line3_U17_Ins0_U1 ( .A(ciphertext_s0[93]), .B(
        ciphertext_s0[61]), .ZN(MixColumns_line3_n11) );
  XOR2_X1 MixColumns_line3_U17_Ins_1_U1 ( .A(ciphertext_s1[93]), .B(
        ciphertext_s1[61]), .Z(new_AGEMA_signal_2105) );
  XOR2_X1 MixColumns_line3_U16_Ins_0_U1 ( .A(ciphertext_s0[28]), .B(
        MixColumns_line3_S13[5]), .Z(MixColumns_line3_n12) );
  XOR2_X1 MixColumns_line3_U16_Ins_1_U1 ( .A(ciphertext_s1[28]), .B(
        new_AGEMA_signal_2116), .Z(new_AGEMA_signal_2148) );
  XNOR2_X1 MixColumns_line3_U15_Ins0_U1 ( .A(MixColumns_line3_n10), .B(
        MixColumns_line3_n9), .ZN(MCout[4]) );
  XOR2_X1 MixColumns_line3_U15_Ins_1_U1 ( .A(new_AGEMA_signal_2821), .B(
        new_AGEMA_signal_2106), .Z(new_AGEMA_signal_2847) );
  XNOR2_X1 MixColumns_line3_U14_Ins0_U1 ( .A(ciphertext_s0[92]), .B(
        ciphertext_s0[60]), .ZN(MixColumns_line3_n9) );
  XOR2_X1 MixColumns_line3_U14_Ins_1_U1 ( .A(ciphertext_s1[92]), .B(
        ciphertext_s1[60]), .Z(new_AGEMA_signal_2106) );
  XOR2_X1 MixColumns_line3_U13_Ins_0_U1 ( .A(MixColumns_line3_S02_4_), .B(
        MixColumns_line3_S13[4]), .Z(MixColumns_line3_n10) );
  XOR2_X1 MixColumns_line3_U13_Ins_1_U1 ( .A(new_AGEMA_signal_2111), .B(
        new_AGEMA_signal_2151), .Z(new_AGEMA_signal_2821) );
  XNOR2_X1 MixColumns_line3_U12_Ins0_U1 ( .A(MixColumns_line3_n8), .B(
        MixColumns_line3_n7), .ZN(MCout[3]) );
  XOR2_X1 MixColumns_line3_U12_Ins_1_U1 ( .A(new_AGEMA_signal_2822), .B(
        new_AGEMA_signal_2107), .Z(new_AGEMA_signal_2848) );
  XNOR2_X1 MixColumns_line3_U11_Ins0_U1 ( .A(ciphertext_s0[91]), .B(
        ciphertext_s0[59]), .ZN(MixColumns_line3_n7) );
  XOR2_X1 MixColumns_line3_U11_Ins_1_U1 ( .A(ciphertext_s1[91]), .B(
        ciphertext_s1[59]), .Z(new_AGEMA_signal_2107) );
  XOR2_X1 MixColumns_line3_U10_Ins_0_U1 ( .A(MixColumns_line3_S02_3_), .B(
        MixColumns_line3_S13[3]), .Z(MixColumns_line3_n8) );
  XOR2_X1 MixColumns_line3_U10_Ins_1_U1 ( .A(new_AGEMA_signal_2112), .B(
        new_AGEMA_signal_2152), .Z(new_AGEMA_signal_2822) );
  XNOR2_X1 MixColumns_line3_U9_Ins0_U1 ( .A(MixColumns_line3_n6), .B(
        MixColumns_line3_n5), .ZN(MCout[2]) );
  XOR2_X1 MixColumns_line3_U9_Ins_1_U1 ( .A(new_AGEMA_signal_2149), .B(
        new_AGEMA_signal_2108), .Z(new_AGEMA_signal_2823) );
  XNOR2_X1 MixColumns_line3_U8_Ins0_U1 ( .A(ciphertext_s0[90]), .B(
        ciphertext_s0[58]), .ZN(MixColumns_line3_n5) );
  XOR2_X1 MixColumns_line3_U8_Ins_1_U1 ( .A(ciphertext_s1[90]), .B(
        ciphertext_s1[58]), .Z(new_AGEMA_signal_2108) );
  XOR2_X1 MixColumns_line3_U7_Ins_0_U1 ( .A(ciphertext_s0[25]), .B(
        MixColumns_line3_S13[2]), .Z(MixColumns_line3_n6) );
  XOR2_X1 MixColumns_line3_U7_Ins_1_U1 ( .A(ciphertext_s1[25]), .B(
        new_AGEMA_signal_2117), .Z(new_AGEMA_signal_2149) );
  XNOR2_X1 MixColumns_line3_U6_Ins0_U1 ( .A(MixColumns_line3_n4), .B(
        MixColumns_line3_n3), .ZN(MCout[1]) );
  XOR2_X1 MixColumns_line3_U6_Ins_1_U1 ( .A(new_AGEMA_signal_2824), .B(
        new_AGEMA_signal_2109), .Z(new_AGEMA_signal_2849) );
  XNOR2_X1 MixColumns_line3_U5_Ins0_U1 ( .A(ciphertext_s0[57]), .B(
        ciphertext_s0[89]), .ZN(MixColumns_line3_n3) );
  XOR2_X1 MixColumns_line3_U5_Ins_1_U1 ( .A(ciphertext_s1[57]), .B(
        ciphertext_s1[89]), .Z(new_AGEMA_signal_2109) );
  XOR2_X1 MixColumns_line3_U4_Ins_0_U1 ( .A(MixColumns_line3_S02_1_), .B(
        MixColumns_line3_S13[1]), .Z(MixColumns_line3_n4) );
  XOR2_X1 MixColumns_line3_U4_Ins_1_U1 ( .A(new_AGEMA_signal_2113), .B(
        new_AGEMA_signal_2153), .Z(new_AGEMA_signal_2824) );
  XNOR2_X1 MixColumns_line3_U3_Ins0_U1 ( .A(MixColumns_line3_n2), .B(
        MixColumns_line3_n1), .ZN(MCout[0]) );
  XOR2_X1 MixColumns_line3_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2150), .B(
        new_AGEMA_signal_2110), .Z(new_AGEMA_signal_2825) );
  XNOR2_X1 MixColumns_line3_U2_Ins0_U1 ( .A(ciphertext_s0[56]), .B(
        ciphertext_s0[88]), .ZN(MixColumns_line3_n1) );
  XOR2_X1 MixColumns_line3_U2_Ins_1_U1 ( .A(ciphertext_s1[56]), .B(
        ciphertext_s1[88]), .Z(new_AGEMA_signal_2110) );
  XOR2_X1 MixColumns_line3_U1_Ins_0_U1 ( .A(ciphertext_s0[31]), .B(
        MixColumns_line3_S13[0]), .Z(MixColumns_line3_n2) );
  XOR2_X1 MixColumns_line3_U1_Ins_1_U1 ( .A(ciphertext_s1[31]), .B(
        new_AGEMA_signal_2118), .Z(new_AGEMA_signal_2150) );
  XOR2_X1 MixColumns_line3_timesTWO_U3_Ins_0_U1 ( .A(ciphertext_s0[31]), .B(
        ciphertext_s0[27]), .Z(MixColumns_line3_S02_4_) );
  XOR2_X1 MixColumns_line3_timesTWO_U3_Ins_1_U1 ( .A(ciphertext_s1[31]), .B(
        ciphertext_s1[27]), .Z(new_AGEMA_signal_2111) );
  XOR2_X1 MixColumns_line3_timesTWO_U2_Ins_0_U1 ( .A(ciphertext_s0[31]), .B(
        ciphertext_s0[26]), .Z(MixColumns_line3_S02_3_) );
  XOR2_X1 MixColumns_line3_timesTWO_U2_Ins_1_U1 ( .A(ciphertext_s1[31]), .B(
        ciphertext_s1[26]), .Z(new_AGEMA_signal_2112) );
  XOR2_X1 MixColumns_line3_timesTWO_U1_Ins_0_U1 ( .A(ciphertext_s0[31]), .B(
        ciphertext_s0[24]), .Z(MixColumns_line3_S02_1_) );
  XOR2_X1 MixColumns_line3_timesTWO_U1_Ins_1_U1 ( .A(ciphertext_s1[31]), .B(
        ciphertext_s1[24]), .Z(new_AGEMA_signal_2113) );
  XOR2_X1 MixColumns_line3_timesTHREE_U8_Ins_0_U1 ( .A(ciphertext_s0[127]), 
        .B(ciphertext_s0[126]), .Z(MixColumns_line3_S13[7]) );
  XOR2_X1 MixColumns_line3_timesTHREE_U8_Ins_1_U1 ( .A(ciphertext_s1[127]), 
        .B(ciphertext_s1[126]), .Z(new_AGEMA_signal_2114) );
  XOR2_X1 MixColumns_line3_timesTHREE_U7_Ins_0_U1 ( .A(ciphertext_s0[126]), 
        .B(ciphertext_s0[125]), .Z(MixColumns_line3_S13[6]) );
  XOR2_X1 MixColumns_line3_timesTHREE_U7_Ins_1_U1 ( .A(ciphertext_s1[126]), 
        .B(ciphertext_s1[125]), .Z(new_AGEMA_signal_2115) );
  XOR2_X1 MixColumns_line3_timesTHREE_U6_Ins_0_U1 ( .A(ciphertext_s0[125]), 
        .B(ciphertext_s0[124]), .Z(MixColumns_line3_S13[5]) );
  XOR2_X1 MixColumns_line3_timesTHREE_U6_Ins_1_U1 ( .A(ciphertext_s1[125]), 
        .B(ciphertext_s1[124]), .Z(new_AGEMA_signal_2116) );
  XOR2_X1 MixColumns_line3_timesTHREE_U5_Ins_0_U1 ( .A(ciphertext_s0[124]), 
        .B(MixColumns_line3_timesTHREE_input2_4_), .Z(MixColumns_line3_S13[4])
         );
  XOR2_X1 MixColumns_line3_timesTHREE_U5_Ins_1_U1 ( .A(ciphertext_s1[124]), 
        .B(new_AGEMA_signal_2119), .Z(new_AGEMA_signal_2151) );
  XOR2_X1 MixColumns_line3_timesTHREE_U4_Ins_0_U1 ( .A(ciphertext_s0[123]), 
        .B(MixColumns_line3_timesTHREE_input2_3_), .Z(MixColumns_line3_S13[3])
         );
  XOR2_X1 MixColumns_line3_timesTHREE_U4_Ins_1_U1 ( .A(ciphertext_s1[123]), 
        .B(new_AGEMA_signal_2120), .Z(new_AGEMA_signal_2152) );
  XOR2_X1 MixColumns_line3_timesTHREE_U3_Ins_0_U1 ( .A(ciphertext_s0[122]), 
        .B(ciphertext_s0[121]), .Z(MixColumns_line3_S13[2]) );
  XOR2_X1 MixColumns_line3_timesTHREE_U3_Ins_1_U1 ( .A(ciphertext_s1[122]), 
        .B(ciphertext_s1[121]), .Z(new_AGEMA_signal_2117) );
  XOR2_X1 MixColumns_line3_timesTHREE_U2_Ins_0_U1 ( .A(ciphertext_s0[121]), 
        .B(MixColumns_line3_timesTHREE_input2_1_), .Z(MixColumns_line3_S13[1])
         );
  XOR2_X1 MixColumns_line3_timesTHREE_U2_Ins_1_U1 ( .A(ciphertext_s1[121]), 
        .B(new_AGEMA_signal_2121), .Z(new_AGEMA_signal_2153) );
  XOR2_X1 MixColumns_line3_timesTHREE_U1_Ins_0_U1 ( .A(ciphertext_s0[120]), 
        .B(ciphertext_s0[127]), .Z(MixColumns_line3_S13[0]) );
  XOR2_X1 MixColumns_line3_timesTHREE_U1_Ins_1_U1 ( .A(ciphertext_s1[120]), 
        .B(ciphertext_s1[127]), .Z(new_AGEMA_signal_2118) );
  XOR2_X1 MixColumns_line3_timesTHREE_timesTWO_U3_Ins_0_U1 ( .A(
        ciphertext_s0[127]), .B(ciphertext_s0[123]), .Z(
        MixColumns_line3_timesTHREE_input2_4_) );
  XOR2_X1 MixColumns_line3_timesTHREE_timesTWO_U3_Ins_1_U1 ( .A(
        ciphertext_s1[127]), .B(ciphertext_s1[123]), .Z(new_AGEMA_signal_2119)
         );
  XOR2_X1 MixColumns_line3_timesTHREE_timesTWO_U2_Ins_0_U1 ( .A(
        ciphertext_s0[127]), .B(ciphertext_s0[122]), .Z(
        MixColumns_line3_timesTHREE_input2_3_) );
  XOR2_X1 MixColumns_line3_timesTHREE_timesTWO_U2_Ins_1_U1 ( .A(
        ciphertext_s1[127]), .B(ciphertext_s1[122]), .Z(new_AGEMA_signal_2120)
         );
  XOR2_X1 MixColumns_line3_timesTHREE_timesTWO_U1_Ins_0_U1 ( .A(
        ciphertext_s0[127]), .B(ciphertext_s0[120]), .Z(
        MixColumns_line3_timesTHREE_input2_1_) );
  XOR2_X1 MixColumns_line3_timesTHREE_timesTWO_U1_Ins_1_U1 ( .A(
        ciphertext_s1[127]), .B(ciphertext_s1[120]), .Z(new_AGEMA_signal_2121)
         );
  MUX2_X1 MUX_SboxIn_mux_inst_0_U1_Ins_0_U1 ( .A(StateOutXORroundKey[0]), .B(
        keySBIn[0]), .S(n173), .Z(SboxIn[0]) );
  MUX2_X1 MUX_SboxIn_mux_inst_0_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1984), .B(
        new_AGEMA_signal_2563), .S(n173), .Z(new_AGEMA_signal_2826) );
  MUX2_X1 MUX_SboxIn_mux_inst_1_U1_Ins_0_U1 ( .A(StateOutXORroundKey[1]), .B(
        keySBIn[1]), .S(n173), .Z(SboxIn[1]) );
  MUX2_X1 MUX_SboxIn_mux_inst_1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1987), .B(
        new_AGEMA_signal_2566), .S(n173), .Z(new_AGEMA_signal_2827) );
  MUX2_X1 MUX_SboxIn_mux_inst_2_U1_Ins_0_U1 ( .A(StateOutXORroundKey[2]), .B(
        keySBIn[2]), .S(n173), .Z(SboxIn[2]) );
  MUX2_X1 MUX_SboxIn_mux_inst_2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1990), .B(
        new_AGEMA_signal_2569), .S(n173), .Z(new_AGEMA_signal_2828) );
  MUX2_X1 MUX_SboxIn_mux_inst_3_U1_Ins_0_U1 ( .A(StateOutXORroundKey[3]), .B(
        keySBIn[3]), .S(n174), .Z(SboxIn[3]) );
  MUX2_X1 MUX_SboxIn_mux_inst_3_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1993), .B(
        new_AGEMA_signal_2572), .S(n174), .Z(new_AGEMA_signal_2829) );
  MUX2_X1 MUX_SboxIn_mux_inst_4_U1_Ins_0_U1 ( .A(StateOutXORroundKey[4]), .B(
        keySBIn[4]), .S(n174), .Z(SboxIn[4]) );
  MUX2_X1 MUX_SboxIn_mux_inst_4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1996), .B(
        new_AGEMA_signal_2575), .S(n174), .Z(new_AGEMA_signal_2830) );
  MUX2_X1 MUX_SboxIn_mux_inst_5_U1_Ins_0_U1 ( .A(StateOutXORroundKey[5]), .B(
        keySBIn[5]), .S(n174), .Z(SboxIn[5]) );
  MUX2_X1 MUX_SboxIn_mux_inst_5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1999), .B(
        new_AGEMA_signal_2578), .S(n174), .Z(new_AGEMA_signal_2831) );
  MUX2_X1 MUX_SboxIn_mux_inst_6_U1_Ins_0_U1 ( .A(StateOutXORroundKey[6]), .B(
        keySBIn[6]), .S(n174), .Z(SboxIn[6]) );
  MUX2_X1 MUX_SboxIn_mux_inst_6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2002), .B(
        new_AGEMA_signal_2581), .S(n174), .Z(new_AGEMA_signal_2832) );
  MUX2_X1 MUX_SboxIn_mux_inst_7_U1_Ins_0_U1 ( .A(StateOutXORroundKey[7]), .B(
        keySBIn[7]), .S(n174), .Z(SboxIn[7]) );
  MUX2_X1 MUX_SboxIn_mux_inst_7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2005), .B(
        new_AGEMA_signal_2584), .S(n174), .Z(new_AGEMA_signal_2833) );
  XOR2_X2 Inst_bSbox_XOR_T1_U1_Ins_0_U1 ( .A(SboxIn[7]), .B(SboxIn[4]), .Z(
        Inst_bSbox_T1) );
  XOR2_X1 Inst_bSbox_XOR_T1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2833), .B(
        new_AGEMA_signal_2830), .Z(new_AGEMA_signal_2850) );
  XOR2_X1 Inst_bSbox_XOR_T2_U1_Ins_0_U1 ( .A(SboxIn[7]), .B(SboxIn[2]), .Z(
        Inst_bSbox_T2) );
  XOR2_X1 Inst_bSbox_XOR_T2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2833), .B(
        new_AGEMA_signal_2828), .Z(new_AGEMA_signal_2851) );
  XOR2_X1 Inst_bSbox_XOR_T3_U1_Ins_0_U1 ( .A(SboxIn[7]), .B(SboxIn[1]), .Z(
        Inst_bSbox_T3) );
  XOR2_X1 Inst_bSbox_XOR_T3_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2833), .B(
        new_AGEMA_signal_2827), .Z(new_AGEMA_signal_2852) );
  XOR2_X1 Inst_bSbox_XOR_T4_U1_Ins_0_U1 ( .A(SboxIn[4]), .B(SboxIn[2]), .Z(
        Inst_bSbox_T4) );
  XOR2_X1 Inst_bSbox_XOR_T4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2830), .B(
        new_AGEMA_signal_2828), .Z(new_AGEMA_signal_2853) );
  XOR2_X1 Inst_bSbox_XOR_T5_U1_Ins_0_U1 ( .A(SboxIn[3]), .B(SboxIn[1]), .Z(
        Inst_bSbox_T5) );
  XOR2_X1 Inst_bSbox_XOR_T5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2829), .B(
        new_AGEMA_signal_2827), .Z(new_AGEMA_signal_2854) );
  XOR2_X2 Inst_bSbox_XOR_T6_U1_Ins_0_U1 ( .A(Inst_bSbox_T1), .B(Inst_bSbox_T5), 
        .Z(Inst_bSbox_T6) );
  INV_X1 Inst_bSbox_XOR_T6_U1_Ins_1_U2 ( .A(Inst_bSbox_XOR_T6_U1_Ins_1_n2), 
        .ZN(new_AGEMA_signal_3000) );
  XNOR2_X1 Inst_bSbox_XOR_T6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2850), .B(
        new_AGEMA_signal_2854), .ZN(Inst_bSbox_XOR_T6_U1_Ins_1_n2) );
  XOR2_X1 Inst_bSbox_XOR_T7_U1_Ins_0_U1 ( .A(SboxIn[6]), .B(SboxIn[5]), .Z(
        Inst_bSbox_T7) );
  XOR2_X1 Inst_bSbox_XOR_T7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2832), .B(
        new_AGEMA_signal_2831), .Z(new_AGEMA_signal_2855) );
  XOR2_X1 Inst_bSbox_XOR_T8_U1_Ins_0_U1 ( .A(SboxIn[0]), .B(Inst_bSbox_T6), 
        .Z(Inst_bSbox_T8) );
  XOR2_X1 Inst_bSbox_XOR_T8_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2826), .B(
        new_AGEMA_signal_3000), .Z(new_AGEMA_signal_3032) );
  XOR2_X1 Inst_bSbox_XOR_T9_U1_Ins_0_U1 ( .A(SboxIn[0]), .B(Inst_bSbox_T7), 
        .Z(Inst_bSbox_T9) );
  XOR2_X1 Inst_bSbox_XOR_T9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2826), .B(
        new_AGEMA_signal_2855), .Z(new_AGEMA_signal_3001) );
  XOR2_X1 Inst_bSbox_XOR_T10_U1_Ins_0_U1 ( .A(Inst_bSbox_T6), .B(Inst_bSbox_T7), .Z(Inst_bSbox_T10) );
  XOR2_X1 Inst_bSbox_XOR_T10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3000), .B(
        new_AGEMA_signal_2855), .Z(new_AGEMA_signal_3033) );
  XOR2_X1 Inst_bSbox_XOR_T11_U1_Ins_0_U1 ( .A(SboxIn[6]), .B(SboxIn[2]), .Z(
        Inst_bSbox_T11) );
  XOR2_X1 Inst_bSbox_XOR_T11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2832), .B(
        new_AGEMA_signal_2828), .Z(new_AGEMA_signal_2856) );
  XOR2_X1 Inst_bSbox_XOR_T12_U1_Ins_0_U1 ( .A(SboxIn[5]), .B(SboxIn[2]), .Z(
        Inst_bSbox_T12) );
  XOR2_X1 Inst_bSbox_XOR_T12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2831), .B(
        new_AGEMA_signal_2828), .Z(new_AGEMA_signal_2857) );
  XOR2_X1 Inst_bSbox_XOR_T13_U1_Ins_0_U1 ( .A(Inst_bSbox_T3), .B(Inst_bSbox_T4), .Z(Inst_bSbox_T13) );
  XOR2_X1 Inst_bSbox_XOR_T13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2852), .B(
        new_AGEMA_signal_2853), .Z(new_AGEMA_signal_3002) );
  XOR2_X1 Inst_bSbox_XOR_T14_U1_Ins_0_U1 ( .A(Inst_bSbox_T6), .B(
        Inst_bSbox_T11), .Z(Inst_bSbox_T14) );
  XOR2_X1 Inst_bSbox_XOR_T14_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3000), .B(
        new_AGEMA_signal_2856), .Z(new_AGEMA_signal_3034) );
  XOR2_X1 Inst_bSbox_XOR_T15_U1_Ins_0_U1 ( .A(Inst_bSbox_T5), .B(
        Inst_bSbox_T11), .Z(Inst_bSbox_T15) );
  XOR2_X1 Inst_bSbox_XOR_T15_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2854), .B(
        new_AGEMA_signal_2856), .Z(new_AGEMA_signal_3003) );
  XOR2_X2 Inst_bSbox_XOR_T16_U1_Ins_0_U1 ( .A(Inst_bSbox_T5), .B(
        Inst_bSbox_T12), .Z(Inst_bSbox_T16) );
  XOR2_X1 Inst_bSbox_XOR_T16_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2854), .B(
        new_AGEMA_signal_2857), .Z(new_AGEMA_signal_3004) );
  XOR2_X1 Inst_bSbox_XOR_T17_U1_Ins_0_U1 ( .A(Inst_bSbox_T9), .B(
        Inst_bSbox_T16), .Z(Inst_bSbox_T17) );
  XOR2_X1 Inst_bSbox_XOR_T17_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3001), .B(
        new_AGEMA_signal_3004), .Z(new_AGEMA_signal_3035) );
  XOR2_X1 Inst_bSbox_XOR_T18_U1_Ins_0_U1 ( .A(SboxIn[4]), .B(SboxIn[0]), .Z(
        Inst_bSbox_T18) );
  XOR2_X1 Inst_bSbox_XOR_T18_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2830), .B(
        new_AGEMA_signal_2826), .Z(new_AGEMA_signal_2858) );
  XOR2_X1 Inst_bSbox_XOR_T19_U1_Ins_0_U1 ( .A(Inst_bSbox_T7), .B(
        Inst_bSbox_T18), .Z(Inst_bSbox_T19) );
  XOR2_X1 Inst_bSbox_XOR_T19_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2855), .B(
        new_AGEMA_signal_2858), .Z(new_AGEMA_signal_3005) );
  XOR2_X1 Inst_bSbox_XOR_T20_U1_Ins_0_U1 ( .A(Inst_bSbox_T1), .B(
        Inst_bSbox_T19), .Z(Inst_bSbox_T20) );
  XOR2_X1 Inst_bSbox_XOR_T20_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2850), .B(
        new_AGEMA_signal_3005), .Z(new_AGEMA_signal_3036) );
  XOR2_X1 Inst_bSbox_XOR_T21_U1_Ins_0_U1 ( .A(SboxIn[1]), .B(SboxIn[0]), .Z(
        Inst_bSbox_T21) );
  XOR2_X1 Inst_bSbox_XOR_T21_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2827), .B(
        new_AGEMA_signal_2826), .Z(new_AGEMA_signal_2859) );
  XOR2_X1 Inst_bSbox_XOR_T22_U1_Ins_0_U1 ( .A(Inst_bSbox_T7), .B(
        Inst_bSbox_T21), .Z(Inst_bSbox_T22) );
  XOR2_X1 Inst_bSbox_XOR_T22_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2855), .B(
        new_AGEMA_signal_2859), .Z(new_AGEMA_signal_3006) );
  XOR2_X1 Inst_bSbox_XOR_T23_U1_Ins_0_U1 ( .A(Inst_bSbox_T2), .B(
        Inst_bSbox_T22), .Z(Inst_bSbox_T23) );
  XOR2_X1 Inst_bSbox_XOR_T23_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2851), .B(
        new_AGEMA_signal_3006), .Z(new_AGEMA_signal_3037) );
  XOR2_X1 Inst_bSbox_XOR_T24_U1_Ins_0_U1 ( .A(Inst_bSbox_T2), .B(
        Inst_bSbox_T10), .Z(Inst_bSbox_T24) );
  XOR2_X1 Inst_bSbox_XOR_T24_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2851), .B(
        new_AGEMA_signal_3033), .Z(new_AGEMA_signal_3117) );
  XOR2_X1 Inst_bSbox_XOR_T25_U1_Ins_0_U1 ( .A(Inst_bSbox_T20), .B(
        Inst_bSbox_T17), .Z(Inst_bSbox_T25) );
  XOR2_X1 Inst_bSbox_XOR_T25_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3036), .B(
        new_AGEMA_signal_3035), .Z(new_AGEMA_signal_3118) );
  XOR2_X1 Inst_bSbox_XOR_T26_U1_Ins_0_U1 ( .A(Inst_bSbox_T3), .B(
        Inst_bSbox_T16), .Z(Inst_bSbox_T26) );
  XOR2_X1 Inst_bSbox_XOR_T26_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2852), .B(
        new_AGEMA_signal_3004), .Z(new_AGEMA_signal_3038) );
  XOR2_X1 Inst_bSbox_XOR_T27_U1_Ins_0_U1 ( .A(Inst_bSbox_T1), .B(
        Inst_bSbox_T12), .Z(Inst_bSbox_T27) );
  XOR2_X1 Inst_bSbox_XOR_T27_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2850), .B(
        new_AGEMA_signal_2857), .Z(new_AGEMA_signal_3007) );
  NOR2_X1 ClockGatingInst_U9 ( .A1(start), .A2(ClockGatingInst_n9), .ZN(
        ClockGatingInst_n4) );
  NOR2_X1 ClockGatingInst_U8 ( .A1(start), .A2(ClockGatingInst_n8), .ZN(
        ClockGatingInst_n3) );
  NOR2_X1 ClockGatingInst_U7 ( .A1(start), .A2(ClockGatingInst_n7), .ZN(
        ClockGatingInst_n2) );
  NOR2_X1 ClockGatingInst_U6 ( .A1(start), .A2(ClockGatingInst_n6), .ZN(
        ClockGatingInst_n1) );
  NAND2_X1 ClockGatingInst_U5 ( .A1(ClockGatingInst_n10), .A2(
        ClockGatingInst_n5), .ZN(ClockGatingInst_N7) );
  INV_X1 ClockGatingInst_U4 ( .A(start), .ZN(ClockGatingInst_n5) );
  AND2_X1 ClockGatingInst_U3 ( .A1(ClockGatingInst_LatchedEnable), .A2(clk), 
        .ZN(clk_gated) );
  DFF_X1 ClockGatingInst_ShiftRegister_reg_2_ ( .D(ClockGatingInst_n1), .CK(
        clk), .Q(), .QN(ClockGatingInst_n7) );
  DFF_X1 ClockGatingInst_ShiftRegister_reg_3_ ( .D(ClockGatingInst_n2), .CK(
        clk), .Q(), .QN(ClockGatingInst_n8) );
  DFF_X1 ClockGatingInst_ShiftRegister_reg_4_ ( .D(ClockGatingInst_n3), .CK(
        clk), .Q(), .QN(ClockGatingInst_n9) );
  DFF_X1 ClockGatingInst_ShiftRegister_reg_5_ ( .D(ClockGatingInst_n4), .CK(
        clk), .Q(ClockGatingInst_ShiftRegister_5_), .QN(ClockGatingInst_n10)
         );
  DLL_X1 ClockGatingInst_LatchedEnable_reg ( .D(ClockGatingInst_N7), .GN(clk), 
        .Q(ClockGatingInst_LatchedEnable) );
  DLL_X1 ClockGatingInst_Synch_reg ( .D(ClockGatingInst_ShiftRegister_5_), 
        .GN(clk), .Q(Synch) );
  DFF_X1 ClockGatingInst_ShiftRegister_reg_1_ ( .D(ClockGatingInst_N7), .CK(
        clk), .Q(), .QN(ClockGatingInst_n6) );
  OAI21_X1 Inst_bSbox_AND_M1_U1_U4 ( .B1(new_AGEMA_signal_3002), .B2(
        Inst_bSbox_AND_M1_U1_n3), .A(Inst_bSbox_AND_M1_U1_n2), .ZN(
        Inst_bSbox_AND_M1_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M1_U1_U3 ( .B1(new_AGEMA_signal_3000), .B2(Fresh[1]), .C1(Inst_bSbox_AND_M1_U1_n1), .C2(Fresh[3]), .A(new_AGEMA_signal_3002), .ZN(
        Inst_bSbox_AND_M1_U1_n2) );
  AOI22_X1 Inst_bSbox_AND_M1_U1_U2 ( .A1(new_AGEMA_signal_3000), .A2(Fresh[2]), 
        .B1(Fresh[0]), .B2(Inst_bSbox_AND_M1_U1_n1), .ZN(
        Inst_bSbox_AND_M1_U1_n3) );
  INV_X1 Inst_bSbox_AND_M1_U1_U1 ( .A(new_AGEMA_signal_3000), .ZN(
        Inst_bSbox_AND_M1_U1_n1) );
  DFF_X1 Inst_bSbox_AND_M1_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3002), .CK(clk), .Q(Inst_bSbox_AND_M1_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M1_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3000), .CK(clk), .Q(Inst_bSbox_AND_M1_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M1_U1_Step1_ins_U9 ( .A(Fresh[3]), .B(
        Inst_bSbox_AND_M1_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M1_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M1_U1_Step1_ins_U8 ( .A1(Inst_bSbox_T13), .A2(
        Inst_bSbox_T6), .ZN(Inst_bSbox_AND_M1_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M1_U1_Step1_ins_U7 ( .A(Fresh[2]), .B(
        Inst_bSbox_AND_M1_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M1_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M1_U1_Step1_ins_U6 ( .A1(Inst_bSbox_T6), .A2(
        Inst_bSbox_AND_M1_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M1_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M1_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M1_U1_Step1_ins_n14), .B(Fresh[1]), .ZN(
        Inst_bSbox_AND_M1_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M1_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M1_U1_Step1_ins_n15), .A2(Inst_bSbox_T6), .ZN(
        Inst_bSbox_AND_M1_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M1_U1_Step1_ins_U3 ( .A(Inst_bSbox_T13), .ZN(
        Inst_bSbox_AND_M1_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M1_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M1_U1_Step1_ins_n13), .B(Fresh[0]), .ZN(
        Inst_bSbox_AND_M1_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M1_U1_Step1_ins_U1 ( .A1(Inst_bSbox_T6), .A2(
        Inst_bSbox_T13), .ZN(Inst_bSbox_AND_M1_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M1_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M1_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M1_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M1_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M1_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M1_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M1_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M1_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M1_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M1_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M1_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M1_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M1_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M1_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M1_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M1_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3039) );
  OAI221_X1 Inst_bSbox_AND_M1_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M1_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M1_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M1_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M1_U1_Step1_reg[3]), .A(Inst_bSbox_AND_M1_U1_in1_reg[1]), .ZN(Inst_bSbox_AND_M1_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M1_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M1_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M1_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M1_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M1_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M1_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M1_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M1_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M1_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M1_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M1_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M1), .QN()
         );
  OAI21_X1 Inst_bSbox_AND_M2_U1_U4 ( .B1(new_AGEMA_signal_3037), .B2(
        Inst_bSbox_AND_M2_U1_n11), .A(Inst_bSbox_AND_M2_U1_n10), .ZN(
        Inst_bSbox_AND_M2_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M2_U1_U3 ( .B1(new_AGEMA_signal_3032), .B2(Fresh[5]), .C1(Inst_bSbox_AND_M2_U1_n9), .C2(Fresh[7]), .A(new_AGEMA_signal_3037), .ZN(
        Inst_bSbox_AND_M2_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M2_U1_U2 ( .A1(new_AGEMA_signal_3032), .A2(Fresh[6]), 
        .B1(Fresh[4]), .B2(Inst_bSbox_AND_M2_U1_n9), .ZN(
        Inst_bSbox_AND_M2_U1_n11) );
  INV_X1 Inst_bSbox_AND_M2_U1_U1 ( .A(new_AGEMA_signal_3032), .ZN(
        Inst_bSbox_AND_M2_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M2_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3037), .CK(clk), .Q(Inst_bSbox_AND_M2_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M2_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3032), .CK(clk), .Q(Inst_bSbox_AND_M2_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M2_U1_Step1_ins_U9 ( .A(Fresh[7]), .B(
        Inst_bSbox_AND_M2_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M2_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M2_U1_Step1_ins_U8 ( .A1(Inst_bSbox_T23), .A2(
        Inst_bSbox_T8), .ZN(Inst_bSbox_AND_M2_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M2_U1_Step1_ins_U7 ( .A(Fresh[6]), .B(
        Inst_bSbox_AND_M2_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M2_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M2_U1_Step1_ins_U6 ( .A1(Inst_bSbox_T8), .A2(
        Inst_bSbox_AND_M2_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M2_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M2_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M2_U1_Step1_ins_n14), .B(Fresh[5]), .ZN(
        Inst_bSbox_AND_M2_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M2_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M2_U1_Step1_ins_n15), .A2(Inst_bSbox_T8), .ZN(
        Inst_bSbox_AND_M2_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M2_U1_Step1_ins_U3 ( .A(Inst_bSbox_T23), .ZN(
        Inst_bSbox_AND_M2_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M2_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M2_U1_Step1_ins_n13), .B(Fresh[4]), .ZN(
        Inst_bSbox_AND_M2_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M2_U1_Step1_ins_U1 ( .A1(Inst_bSbox_T8), .A2(
        Inst_bSbox_T23), .ZN(Inst_bSbox_AND_M2_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M2_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M2_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M2_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M2_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M2_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M2_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M2_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M2_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M2_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M2_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M2_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M2_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M2_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M2_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M2_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M2_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3119) );
  OAI221_X1 Inst_bSbox_AND_M2_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M2_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M2_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M2_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M2_U1_Step1_reg[3]), .A(Inst_bSbox_AND_M2_U1_in1_reg[1]), .ZN(Inst_bSbox_AND_M2_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M2_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M2_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M2_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M2_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M2_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M2_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M2_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M2_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M2_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M2_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M2_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M2), .QN()
         );
  XOR2_X1 Inst_bSbox_XOR_M3_U1_Ins_0_U1 ( .A(Inst_bSbox_T14), .B(Inst_bSbox_M1), .Z(Inst_bSbox_M3) );
  XOR2_X1 Inst_bSbox_XOR_M3_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3034), .B(
        new_AGEMA_signal_3039), .Z(new_AGEMA_signal_3120) );
  OAI21_X1 Inst_bSbox_AND_M4_U1_U4 ( .B1(new_AGEMA_signal_3005), .B2(
        Inst_bSbox_AND_M4_U1_n11), .A(Inst_bSbox_AND_M4_U1_n10), .ZN(
        Inst_bSbox_AND_M4_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M4_U1_U3 ( .B1(new_AGEMA_signal_2826), .B2(Fresh[9]), .C1(Inst_bSbox_AND_M4_U1_n9), .C2(Fresh[11]), .A(new_AGEMA_signal_3005), 
        .ZN(Inst_bSbox_AND_M4_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M4_U1_U2 ( .A1(new_AGEMA_signal_2826), .A2(Fresh[10]), .B1(Fresh[8]), .B2(Inst_bSbox_AND_M4_U1_n9), .ZN(Inst_bSbox_AND_M4_U1_n11)
         );
  INV_X1 Inst_bSbox_AND_M4_U1_U1 ( .A(new_AGEMA_signal_2826), .ZN(
        Inst_bSbox_AND_M4_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M4_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3005), .CK(clk), .Q(Inst_bSbox_AND_M4_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M4_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_2826), .CK(clk), .Q(Inst_bSbox_AND_M4_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M4_U1_Step1_ins_U9 ( .A(Fresh[11]), .B(
        Inst_bSbox_AND_M4_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M4_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M4_U1_Step1_ins_U8 ( .A1(Inst_bSbox_T19), .A2(
        SboxIn[0]), .ZN(Inst_bSbox_AND_M4_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M4_U1_Step1_ins_U7 ( .A(Fresh[10]), .B(
        Inst_bSbox_AND_M4_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M4_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M4_U1_Step1_ins_U6 ( .A1(SboxIn[0]), .A2(
        Inst_bSbox_AND_M4_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M4_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M4_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M4_U1_Step1_ins_n14), .B(Fresh[9]), .ZN(
        Inst_bSbox_AND_M4_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M4_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M4_U1_Step1_ins_n15), .A2(SboxIn[0]), .ZN(
        Inst_bSbox_AND_M4_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M4_U1_Step1_ins_U3 ( .A(Inst_bSbox_T19), .ZN(
        Inst_bSbox_AND_M4_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M4_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M4_U1_Step1_ins_n13), .B(Fresh[8]), .ZN(
        Inst_bSbox_AND_M4_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M4_U1_Step1_ins_U1 ( .A1(SboxIn[0]), .A2(
        Inst_bSbox_T19), .ZN(Inst_bSbox_AND_M4_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M4_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M4_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M4_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M4_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M4_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M4_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M4_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M4_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M4_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M4_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M4_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M4_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M4_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M4_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M4_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M4_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3040) );
  OAI221_X1 Inst_bSbox_AND_M4_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M4_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M4_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M4_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M4_U1_Step1_reg[3]), .A(Inst_bSbox_AND_M4_U1_in1_reg[1]), .ZN(Inst_bSbox_AND_M4_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M4_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M4_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M4_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M4_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M4_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M4_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M4_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M4_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M4_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M4_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M4_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M4), .QN()
         );
  XOR2_X1 Inst_bSbox_XOR_M5_U1_Ins_0_U1 ( .A(Inst_bSbox_M4), .B(Inst_bSbox_M1), 
        .Z(Inst_bSbox_M5) );
  XOR2_X1 Inst_bSbox_XOR_M5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3040), .B(
        new_AGEMA_signal_3039), .Z(new_AGEMA_signal_3121) );
  OAI21_X1 Inst_bSbox_AND_M6_U1_U4 ( .B1(new_AGEMA_signal_2852), .B2(
        Inst_bSbox_AND_M6_U1_n11), .A(Inst_bSbox_AND_M6_U1_n10), .ZN(
        Inst_bSbox_AND_M6_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M6_U1_U3 ( .B1(new_AGEMA_signal_3004), .B2(
        Fresh[13]), .C1(Inst_bSbox_AND_M6_U1_n9), .C2(Fresh[15]), .A(
        new_AGEMA_signal_2852), .ZN(Inst_bSbox_AND_M6_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M6_U1_U2 ( .A1(new_AGEMA_signal_3004), .A2(Fresh[14]), .B1(Fresh[12]), .B2(Inst_bSbox_AND_M6_U1_n9), .ZN(Inst_bSbox_AND_M6_U1_n11)
         );
  INV_X1 Inst_bSbox_AND_M6_U1_U1 ( .A(new_AGEMA_signal_3004), .ZN(
        Inst_bSbox_AND_M6_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M6_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_2852), .CK(clk), .Q(Inst_bSbox_AND_M6_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M6_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3004), .CK(clk), .Q(Inst_bSbox_AND_M6_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M6_U1_Step1_ins_U9 ( .A(Fresh[15]), .B(
        Inst_bSbox_AND_M6_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M6_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M6_U1_Step1_ins_U8 ( .A1(Inst_bSbox_T3), .A2(
        Inst_bSbox_T16), .ZN(Inst_bSbox_AND_M6_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M6_U1_Step1_ins_U7 ( .A(Fresh[14]), .B(
        Inst_bSbox_AND_M6_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M6_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M6_U1_Step1_ins_U6 ( .A1(Inst_bSbox_T16), .A2(
        Inst_bSbox_AND_M6_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M6_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M6_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M6_U1_Step1_ins_n14), .B(Fresh[13]), .ZN(
        Inst_bSbox_AND_M6_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M6_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M6_U1_Step1_ins_n15), .A2(Inst_bSbox_T16), .ZN(
        Inst_bSbox_AND_M6_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M6_U1_Step1_ins_U3 ( .A(Inst_bSbox_T3), .ZN(
        Inst_bSbox_AND_M6_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M6_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M6_U1_Step1_ins_n13), .B(Fresh[12]), .ZN(
        Inst_bSbox_AND_M6_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M6_U1_Step1_ins_U1 ( .A1(Inst_bSbox_T16), .A2(
        Inst_bSbox_T3), .ZN(Inst_bSbox_AND_M6_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M6_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M6_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M6_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M6_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M6_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M6_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M6_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M6_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M6_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M6_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M6_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M6_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M6_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M6_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M6_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M6_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3041) );
  OAI221_X1 Inst_bSbox_AND_M6_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M6_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M6_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M6_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M6_U1_Step1_reg[3]), .A(Inst_bSbox_AND_M6_U1_in1_reg[1]), .ZN(Inst_bSbox_AND_M6_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M6_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M6_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M6_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M6_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M6_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M6_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M6_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M6_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M6_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M6_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M6_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M6), .QN()
         );
  OAI21_X1 Inst_bSbox_AND_M7_U1_U4 ( .B1(new_AGEMA_signal_3006), .B2(
        Inst_bSbox_AND_M7_U1_n11), .A(Inst_bSbox_AND_M7_U1_n10), .ZN(
        Inst_bSbox_AND_M7_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M7_U1_U3 ( .B1(new_AGEMA_signal_3001), .B2(
        Fresh[17]), .C1(Inst_bSbox_AND_M7_U1_n9), .C2(Fresh[19]), .A(
        new_AGEMA_signal_3006), .ZN(Inst_bSbox_AND_M7_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M7_U1_U2 ( .A1(new_AGEMA_signal_3001), .A2(Fresh[18]), .B1(Fresh[16]), .B2(Inst_bSbox_AND_M7_U1_n9), .ZN(Inst_bSbox_AND_M7_U1_n11)
         );
  INV_X1 Inst_bSbox_AND_M7_U1_U1 ( .A(new_AGEMA_signal_3001), .ZN(
        Inst_bSbox_AND_M7_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M7_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3006), .CK(clk), .Q(Inst_bSbox_AND_M7_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M7_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3001), .CK(clk), .Q(Inst_bSbox_AND_M7_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M7_U1_Step1_ins_U9 ( .A(Fresh[19]), .B(
        Inst_bSbox_AND_M7_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M7_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M7_U1_Step1_ins_U8 ( .A1(Inst_bSbox_T22), .A2(
        Inst_bSbox_T9), .ZN(Inst_bSbox_AND_M7_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M7_U1_Step1_ins_U7 ( .A(Fresh[18]), .B(
        Inst_bSbox_AND_M7_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M7_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M7_U1_Step1_ins_U6 ( .A1(Inst_bSbox_T9), .A2(
        Inst_bSbox_AND_M7_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M7_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M7_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M7_U1_Step1_ins_n14), .B(Fresh[17]), .ZN(
        Inst_bSbox_AND_M7_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M7_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M7_U1_Step1_ins_n15), .A2(Inst_bSbox_T9), .ZN(
        Inst_bSbox_AND_M7_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M7_U1_Step1_ins_U3 ( .A(Inst_bSbox_T22), .ZN(
        Inst_bSbox_AND_M7_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M7_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M7_U1_Step1_ins_n13), .B(Fresh[16]), .ZN(
        Inst_bSbox_AND_M7_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M7_U1_Step1_ins_U1 ( .A1(Inst_bSbox_T9), .A2(
        Inst_bSbox_T22), .ZN(Inst_bSbox_AND_M7_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M7_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M7_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M7_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M7_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M7_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M7_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M7_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M7_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M7_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M7_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M7_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M7_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M7_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M7_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M7_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M7_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3042) );
  OAI221_X1 Inst_bSbox_AND_M7_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M7_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M7_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M7_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M7_U1_Step1_reg[3]), .A(Inst_bSbox_AND_M7_U1_in1_reg[1]), .ZN(Inst_bSbox_AND_M7_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M7_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M7_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M7_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M7_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M7_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M7_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M7_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M7_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M7_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M7_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M7_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M7), .QN()
         );
  XOR2_X1 Inst_bSbox_XOR_M8_U1_Ins_0_U1 ( .A(Inst_bSbox_T26), .B(Inst_bSbox_M6), .Z(Inst_bSbox_M8) );
  XOR2_X1 Inst_bSbox_XOR_M8_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3038), .B(
        new_AGEMA_signal_3041), .Z(new_AGEMA_signal_3122) );
  OAI21_X1 Inst_bSbox_AND_M9_U1_U4 ( .B1(new_AGEMA_signal_3036), .B2(
        Inst_bSbox_AND_M9_U1_n11), .A(Inst_bSbox_AND_M9_U1_n10), .ZN(
        Inst_bSbox_AND_M9_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M9_U1_U3 ( .B1(new_AGEMA_signal_3035), .B2(
        Fresh[21]), .C1(Inst_bSbox_AND_M9_U1_n9), .C2(Fresh[23]), .A(
        new_AGEMA_signal_3036), .ZN(Inst_bSbox_AND_M9_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M9_U1_U2 ( .A1(new_AGEMA_signal_3035), .A2(Fresh[22]), .B1(Fresh[20]), .B2(Inst_bSbox_AND_M9_U1_n9), .ZN(Inst_bSbox_AND_M9_U1_n11)
         );
  INV_X1 Inst_bSbox_AND_M9_U1_U1 ( .A(new_AGEMA_signal_3035), .ZN(
        Inst_bSbox_AND_M9_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M9_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3036), .CK(clk), .Q(Inst_bSbox_AND_M9_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M9_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3035), .CK(clk), .Q(Inst_bSbox_AND_M9_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M9_U1_Step1_ins_U9 ( .A(Fresh[23]), .B(
        Inst_bSbox_AND_M9_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M9_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M9_U1_Step1_ins_U8 ( .A1(Inst_bSbox_T20), .A2(
        Inst_bSbox_T17), .ZN(Inst_bSbox_AND_M9_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M9_U1_Step1_ins_U7 ( .A(Fresh[22]), .B(
        Inst_bSbox_AND_M9_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M9_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M9_U1_Step1_ins_U6 ( .A1(Inst_bSbox_T17), .A2(
        Inst_bSbox_AND_M9_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M9_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M9_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M9_U1_Step1_ins_n14), .B(Fresh[21]), .ZN(
        Inst_bSbox_AND_M9_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M9_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M9_U1_Step1_ins_n15), .A2(Inst_bSbox_T17), .ZN(
        Inst_bSbox_AND_M9_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M9_U1_Step1_ins_U3 ( .A(Inst_bSbox_T20), .ZN(
        Inst_bSbox_AND_M9_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M9_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M9_U1_Step1_ins_n13), .B(Fresh[20]), .ZN(
        Inst_bSbox_AND_M9_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M9_U1_Step1_ins_U1 ( .A1(Inst_bSbox_T17), .A2(
        Inst_bSbox_T20), .ZN(Inst_bSbox_AND_M9_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M9_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M9_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M9_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M9_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M9_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M9_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M9_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M9_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M9_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M9_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M9_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M9_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M9_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M9_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M9_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M9_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3123) );
  OAI221_X1 Inst_bSbox_AND_M9_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M9_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M9_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M9_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M9_U1_Step1_reg[3]), .A(Inst_bSbox_AND_M9_U1_in1_reg[1]), .ZN(Inst_bSbox_AND_M9_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M9_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M9_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M9_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M9_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M9_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M9_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M9_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M9_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M9_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M9_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M9_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M9), .QN()
         );
  XOR2_X1 Inst_bSbox_XOR_M10_U1_Ins_0_U1 ( .A(Inst_bSbox_M9), .B(Inst_bSbox_M6), .Z(Inst_bSbox_M10) );
  XOR2_X1 Inst_bSbox_XOR_M10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3123), .B(
        new_AGEMA_signal_3041), .Z(new_AGEMA_signal_3262) );
  OAI21_X1 Inst_bSbox_AND_M11_U1_U4 ( .B1(new_AGEMA_signal_2850), .B2(
        Inst_bSbox_AND_M11_U1_n11), .A(Inst_bSbox_AND_M11_U1_n10), .ZN(
        Inst_bSbox_AND_M11_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M11_U1_U3 ( .B1(new_AGEMA_signal_3003), .B2(
        Fresh[25]), .C1(Inst_bSbox_AND_M11_U1_n9), .C2(Fresh[27]), .A(
        new_AGEMA_signal_2850), .ZN(Inst_bSbox_AND_M11_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M11_U1_U2 ( .A1(new_AGEMA_signal_3003), .A2(
        Fresh[26]), .B1(Fresh[24]), .B2(Inst_bSbox_AND_M11_U1_n9), .ZN(
        Inst_bSbox_AND_M11_U1_n11) );
  INV_X1 Inst_bSbox_AND_M11_U1_U1 ( .A(new_AGEMA_signal_3003), .ZN(
        Inst_bSbox_AND_M11_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M11_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_2850), .CK(clk), .Q(Inst_bSbox_AND_M11_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M11_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3003), .CK(clk), .Q(Inst_bSbox_AND_M11_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M11_U1_Step1_ins_U9 ( .A(Fresh[27]), .B(
        Inst_bSbox_AND_M11_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M11_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M11_U1_Step1_ins_U8 ( .A1(Inst_bSbox_T1), .A2(
        Inst_bSbox_T15), .ZN(Inst_bSbox_AND_M11_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M11_U1_Step1_ins_U7 ( .A(Fresh[26]), .B(
        Inst_bSbox_AND_M11_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M11_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M11_U1_Step1_ins_U6 ( .A1(Inst_bSbox_T15), .A2(
        Inst_bSbox_AND_M11_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M11_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M11_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M11_U1_Step1_ins_n14), .B(Fresh[25]), .ZN(
        Inst_bSbox_AND_M11_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M11_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M11_U1_Step1_ins_n15), .A2(Inst_bSbox_T15), .ZN(
        Inst_bSbox_AND_M11_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M11_U1_Step1_ins_U3 ( .A(Inst_bSbox_T1), .ZN(
        Inst_bSbox_AND_M11_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M11_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M11_U1_Step1_ins_n13), .B(Fresh[24]), .ZN(
        Inst_bSbox_AND_M11_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M11_U1_Step1_ins_U1 ( .A1(Inst_bSbox_T15), .A2(
        Inst_bSbox_T1), .ZN(Inst_bSbox_AND_M11_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M11_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M11_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M11_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M11_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M11_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M11_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M11_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M11_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M11_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M11_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M11_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M11_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M11_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M11_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M11_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M11_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3043) );
  OAI221_X1 Inst_bSbox_AND_M11_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M11_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M11_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M11_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M11_U1_Step1_reg[3]), .A(
        Inst_bSbox_AND_M11_U1_in1_reg[1]), .ZN(
        Inst_bSbox_AND_M11_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M11_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M11_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M11_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M11_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M11_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M11_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M11_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M11_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M11_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M11_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M11_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M11), 
        .QN() );
  OAI21_X1 Inst_bSbox_AND_M12_U1_U4 ( .B1(new_AGEMA_signal_2853), .B2(
        Inst_bSbox_AND_M12_U1_n11), .A(Inst_bSbox_AND_M12_U1_n10), .ZN(
        Inst_bSbox_AND_M12_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M12_U1_U3 ( .B1(new_AGEMA_signal_3007), .B2(
        Fresh[29]), .C1(Inst_bSbox_AND_M12_U1_n9), .C2(Fresh[31]), .A(
        new_AGEMA_signal_2853), .ZN(Inst_bSbox_AND_M12_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M12_U1_U2 ( .A1(new_AGEMA_signal_3007), .A2(
        Fresh[30]), .B1(Fresh[28]), .B2(Inst_bSbox_AND_M12_U1_n9), .ZN(
        Inst_bSbox_AND_M12_U1_n11) );
  INV_X1 Inst_bSbox_AND_M12_U1_U1 ( .A(new_AGEMA_signal_3007), .ZN(
        Inst_bSbox_AND_M12_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M12_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_2853), .CK(clk), .Q(Inst_bSbox_AND_M12_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M12_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3007), .CK(clk), .Q(Inst_bSbox_AND_M12_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M12_U1_Step1_ins_U9 ( .A(Fresh[31]), .B(
        Inst_bSbox_AND_M12_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M12_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M12_U1_Step1_ins_U8 ( .A1(Inst_bSbox_T4), .A2(
        Inst_bSbox_T27), .ZN(Inst_bSbox_AND_M12_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M12_U1_Step1_ins_U7 ( .A(Fresh[30]), .B(
        Inst_bSbox_AND_M12_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M12_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M12_U1_Step1_ins_U6 ( .A1(Inst_bSbox_T27), .A2(
        Inst_bSbox_AND_M12_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M12_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M12_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M12_U1_Step1_ins_n14), .B(Fresh[29]), .ZN(
        Inst_bSbox_AND_M12_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M12_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M12_U1_Step1_ins_n15), .A2(Inst_bSbox_T27), .ZN(
        Inst_bSbox_AND_M12_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M12_U1_Step1_ins_U3 ( .A(Inst_bSbox_T4), .ZN(
        Inst_bSbox_AND_M12_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M12_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M12_U1_Step1_ins_n13), .B(Fresh[28]), .ZN(
        Inst_bSbox_AND_M12_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M12_U1_Step1_ins_U1 ( .A1(Inst_bSbox_T27), .A2(
        Inst_bSbox_T4), .ZN(Inst_bSbox_AND_M12_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M12_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M12_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M12_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M12_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M12_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M12_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M12_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M12_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M12_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M12_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M12_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M12_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M12_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M12_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M12_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M12_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3044) );
  OAI221_X1 Inst_bSbox_AND_M12_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M12_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M12_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M12_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M12_U1_Step1_reg[3]), .A(
        Inst_bSbox_AND_M12_U1_in1_reg[1]), .ZN(
        Inst_bSbox_AND_M12_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M12_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M12_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M12_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M12_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M12_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M12_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M12_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M12_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M12_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M12_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M12_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M12), 
        .QN() );
  XOR2_X1 Inst_bSbox_XOR_M13_U1_Ins_0_U1 ( .A(Inst_bSbox_M12), .B(
        Inst_bSbox_M11), .Z(Inst_bSbox_M13) );
  XOR2_X1 Inst_bSbox_XOR_M13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3044), .B(
        new_AGEMA_signal_3043), .Z(new_AGEMA_signal_3124) );
  OAI21_X1 Inst_bSbox_AND_M14_U1_U4 ( .B1(new_AGEMA_signal_2851), .B2(
        Inst_bSbox_AND_M14_U1_n11), .A(Inst_bSbox_AND_M14_U1_n10), .ZN(
        Inst_bSbox_AND_M14_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M14_U1_U3 ( .B1(new_AGEMA_signal_3033), .B2(
        Fresh[33]), .C1(Inst_bSbox_AND_M14_U1_n9), .C2(Fresh[35]), .A(
        new_AGEMA_signal_2851), .ZN(Inst_bSbox_AND_M14_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M14_U1_U2 ( .A1(new_AGEMA_signal_3033), .A2(
        Fresh[34]), .B1(Fresh[32]), .B2(Inst_bSbox_AND_M14_U1_n9), .ZN(
        Inst_bSbox_AND_M14_U1_n11) );
  INV_X1 Inst_bSbox_AND_M14_U1_U1 ( .A(new_AGEMA_signal_3033), .ZN(
        Inst_bSbox_AND_M14_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M14_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_2851), .CK(clk), .Q(Inst_bSbox_AND_M14_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M14_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3033), .CK(clk), .Q(Inst_bSbox_AND_M14_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M14_U1_Step1_ins_U9 ( .A(Fresh[35]), .B(
        Inst_bSbox_AND_M14_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M14_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M14_U1_Step1_ins_U8 ( .A1(Inst_bSbox_T2), .A2(
        Inst_bSbox_T10), .ZN(Inst_bSbox_AND_M14_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M14_U1_Step1_ins_U7 ( .A(Fresh[34]), .B(
        Inst_bSbox_AND_M14_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M14_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M14_U1_Step1_ins_U6 ( .A1(Inst_bSbox_T10), .A2(
        Inst_bSbox_AND_M14_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M14_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M14_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M14_U1_Step1_ins_n14), .B(Fresh[33]), .ZN(
        Inst_bSbox_AND_M14_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M14_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M14_U1_Step1_ins_n15), .A2(Inst_bSbox_T10), .ZN(
        Inst_bSbox_AND_M14_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M14_U1_Step1_ins_U3 ( .A(Inst_bSbox_T2), .ZN(
        Inst_bSbox_AND_M14_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M14_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M14_U1_Step1_ins_n13), .B(Fresh[32]), .ZN(
        Inst_bSbox_AND_M14_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M14_U1_Step1_ins_U1 ( .A1(Inst_bSbox_T10), .A2(
        Inst_bSbox_T2), .ZN(Inst_bSbox_AND_M14_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M14_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M14_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M14_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M14_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M14_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M14_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M14_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M14_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M14_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M14_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M14_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M14_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M14_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M14_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M14_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M14_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3125) );
  OAI221_X1 Inst_bSbox_AND_M14_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M14_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M14_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M14_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M14_U1_Step1_reg[3]), .A(
        Inst_bSbox_AND_M14_U1_in1_reg[1]), .ZN(
        Inst_bSbox_AND_M14_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M14_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M14_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M14_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M14_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M14_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M14_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M14_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M14_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M14_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M14_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M14_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M14), 
        .QN() );
  XOR2_X1 Inst_bSbox_XOR_M15_U1_Ins_0_U1 ( .A(Inst_bSbox_M14), .B(
        Inst_bSbox_M11), .Z(Inst_bSbox_M15) );
  XOR2_X1 Inst_bSbox_XOR_M15_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3125), .B(
        new_AGEMA_signal_3043), .Z(new_AGEMA_signal_3263) );
  XOR2_X1 Inst_bSbox_XOR_M16_U1_Ins_0_U1 ( .A(Inst_bSbox_M3), .B(Inst_bSbox_M2), .Z(Inst_bSbox_M16) );
  XOR2_X1 Inst_bSbox_XOR_M16_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3120), .B(
        new_AGEMA_signal_3119), .Z(new_AGEMA_signal_3264) );
  XOR2_X1 Inst_bSbox_XOR_M17_U1_Ins_0_U1 ( .A(Inst_bSbox_M5), .B(
        Inst_bSbox_T24), .Z(Inst_bSbox_M17) );
  XOR2_X1 Inst_bSbox_XOR_M17_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3121), .B(
        new_AGEMA_signal_3117), .Z(new_AGEMA_signal_3265) );
  XOR2_X1 Inst_bSbox_XOR_M18_U1_Ins_0_U1 ( .A(Inst_bSbox_M8), .B(Inst_bSbox_M7), .Z(Inst_bSbox_M18) );
  XOR2_X1 Inst_bSbox_XOR_M18_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3122), .B(
        new_AGEMA_signal_3042), .Z(new_AGEMA_signal_3266) );
  XOR2_X1 Inst_bSbox_XOR_M19_U1_Ins_0_U1 ( .A(Inst_bSbox_M10), .B(
        Inst_bSbox_M15), .Z(Inst_bSbox_M19) );
  XOR2_X1 Inst_bSbox_XOR_M19_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3262), .B(
        new_AGEMA_signal_3263), .Z(new_AGEMA_signal_3371) );
  XOR2_X1 Inst_bSbox_XOR_M20_U1_Ins_0_U1 ( .A(Inst_bSbox_M16), .B(
        Inst_bSbox_M13), .Z(Inst_bSbox_M20) );
  XOR2_X1 Inst_bSbox_XOR_M20_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3264), .B(
        new_AGEMA_signal_3124), .Z(new_AGEMA_signal_3372) );
  XOR2_X1 Inst_bSbox_XOR_M21_U1_Ins_0_U1 ( .A(Inst_bSbox_M17), .B(
        Inst_bSbox_M15), .Z(Inst_bSbox_M21) );
  XOR2_X1 Inst_bSbox_XOR_M21_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3265), .B(
        new_AGEMA_signal_3263), .Z(new_AGEMA_signal_3373) );
  XOR2_X1 Inst_bSbox_XOR_M22_U1_Ins_0_U1 ( .A(Inst_bSbox_M18), .B(
        Inst_bSbox_M13), .Z(Inst_bSbox_M22) );
  XOR2_X1 Inst_bSbox_XOR_M22_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3266), .B(
        new_AGEMA_signal_3124), .Z(new_AGEMA_signal_3374) );
  XOR2_X1 Inst_bSbox_XOR_M23_U1_Ins_0_U1 ( .A(Inst_bSbox_M19), .B(
        Inst_bSbox_T25), .Z(Inst_bSbox_M23) );
  XOR2_X1 Inst_bSbox_XOR_M23_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3371), .B(
        new_AGEMA_signal_3118), .Z(new_AGEMA_signal_3383) );
  XOR2_X1 Inst_bSbox_XOR_M24_U1_Ins_0_U1 ( .A(Inst_bSbox_M22), .B(
        Inst_bSbox_M23), .Z(Inst_bSbox_M24) );
  XOR2_X1 Inst_bSbox_XOR_M24_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3374), .B(
        new_AGEMA_signal_3383), .Z(new_AGEMA_signal_3387) );
  XOR2_X1 Inst_bSbox_XOR_M27_U1_Ins_0_U1 ( .A(Inst_bSbox_M20), .B(
        Inst_bSbox_M21), .Z(Inst_bSbox_M27) );
  XOR2_X1 Inst_bSbox_XOR_M27_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3372), .B(
        new_AGEMA_signal_3373), .Z(new_AGEMA_signal_3385) );
  OAI21_X1 Inst_bSbox_AND_M25_U1_U4 ( .B1(new_AGEMA_signal_3374), .B2(
        Inst_bSbox_AND_M25_U1_n11), .A(Inst_bSbox_AND_M25_U1_n10), .ZN(
        Inst_bSbox_AND_M25_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M25_U1_U3 ( .B1(new_AGEMA_signal_3372), .B2(
        Fresh[37]), .C1(Inst_bSbox_AND_M25_U1_n9), .C2(Fresh[39]), .A(
        new_AGEMA_signal_3374), .ZN(Inst_bSbox_AND_M25_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M25_U1_U2 ( .A1(new_AGEMA_signal_3372), .A2(
        Fresh[38]), .B1(Fresh[36]), .B2(Inst_bSbox_AND_M25_U1_n9), .ZN(
        Inst_bSbox_AND_M25_U1_n11) );
  INV_X1 Inst_bSbox_AND_M25_U1_U1 ( .A(new_AGEMA_signal_3372), .ZN(
        Inst_bSbox_AND_M25_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M25_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3374), .CK(clk), .Q(Inst_bSbox_AND_M25_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M25_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3372), .CK(clk), .Q(Inst_bSbox_AND_M25_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M25_U1_Step1_ins_U9 ( .A(Fresh[39]), .B(
        Inst_bSbox_AND_M25_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M25_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M25_U1_Step1_ins_U8 ( .A1(Inst_bSbox_M22), .A2(
        Inst_bSbox_M20), .ZN(Inst_bSbox_AND_M25_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M25_U1_Step1_ins_U7 ( .A(Fresh[38]), .B(
        Inst_bSbox_AND_M25_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M25_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M25_U1_Step1_ins_U6 ( .A1(Inst_bSbox_M20), .A2(
        Inst_bSbox_AND_M25_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M25_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M25_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M25_U1_Step1_ins_n14), .B(Fresh[37]), .ZN(
        Inst_bSbox_AND_M25_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M25_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M25_U1_Step1_ins_n15), .A2(Inst_bSbox_M20), .ZN(
        Inst_bSbox_AND_M25_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M25_U1_Step1_ins_U3 ( .A(Inst_bSbox_M22), .ZN(
        Inst_bSbox_AND_M25_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M25_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M25_U1_Step1_ins_n13), .B(Fresh[36]), .ZN(
        Inst_bSbox_AND_M25_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M25_U1_Step1_ins_U1 ( .A1(Inst_bSbox_M20), .A2(
        Inst_bSbox_M22), .ZN(Inst_bSbox_AND_M25_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M25_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M25_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M25_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M25_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M25_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M25_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M25_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M25_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M25_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M25_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M25_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M25_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M25_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M25_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M25_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M25_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3384) );
  OAI221_X1 Inst_bSbox_AND_M25_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M25_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M25_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M25_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M25_U1_Step1_reg[3]), .A(
        Inst_bSbox_AND_M25_U1_in1_reg[1]), .ZN(
        Inst_bSbox_AND_M25_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M25_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M25_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M25_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M25_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M25_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M25_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M25_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M25_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M25_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M25_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M25_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M25), 
        .QN() );
  XOR2_X1 Inst_bSbox_XOR_M26_U1_Ins_0_U1 ( .A(Inst_bSbox_M21), .B(
        Inst_bSbox_M25), .Z(Inst_bSbox_M26) );
  XOR2_X1 Inst_bSbox_XOR_M26_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3373), .B(
        new_AGEMA_signal_3384), .Z(new_AGEMA_signal_3388) );
  XOR2_X1 Inst_bSbox_XOR_M28_U1_Ins_0_U1 ( .A(Inst_bSbox_M23), .B(
        Inst_bSbox_M25), .Z(Inst_bSbox_M28) );
  XOR2_X1 Inst_bSbox_XOR_M28_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3383), .B(
        new_AGEMA_signal_3384), .Z(new_AGEMA_signal_3389) );
  OAI21_X1 Inst_bSbox_AND_M31_U1_U4 ( .B1(new_AGEMA_signal_3372), .B2(
        Inst_bSbox_AND_M31_U1_n11), .A(Inst_bSbox_AND_M31_U1_n10), .ZN(
        Inst_bSbox_AND_M31_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M31_U1_U3 ( .B1(new_AGEMA_signal_3383), .B2(
        Fresh[41]), .C1(Inst_bSbox_AND_M31_U1_n9), .C2(Fresh[43]), .A(
        new_AGEMA_signal_3372), .ZN(Inst_bSbox_AND_M31_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M31_U1_U2 ( .A1(new_AGEMA_signal_3383), .A2(
        Fresh[42]), .B1(Fresh[40]), .B2(Inst_bSbox_AND_M31_U1_n9), .ZN(
        Inst_bSbox_AND_M31_U1_n11) );
  INV_X1 Inst_bSbox_AND_M31_U1_U1 ( .A(new_AGEMA_signal_3383), .ZN(
        Inst_bSbox_AND_M31_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M31_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3372), .CK(clk), .Q(Inst_bSbox_AND_M31_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M31_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3383), .CK(clk), .Q(Inst_bSbox_AND_M31_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M31_U1_Step1_ins_U9 ( .A(Fresh[43]), .B(
        Inst_bSbox_AND_M31_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M31_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M31_U1_Step1_ins_U8 ( .A1(Inst_bSbox_M20), .A2(
        Inst_bSbox_M23), .ZN(Inst_bSbox_AND_M31_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M31_U1_Step1_ins_U7 ( .A(Fresh[42]), .B(
        Inst_bSbox_AND_M31_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M31_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M31_U1_Step1_ins_U6 ( .A1(Inst_bSbox_M23), .A2(
        Inst_bSbox_AND_M31_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M31_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M31_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M31_U1_Step1_ins_n14), .B(Fresh[41]), .ZN(
        Inst_bSbox_AND_M31_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M31_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M31_U1_Step1_ins_n15), .A2(Inst_bSbox_M23), .ZN(
        Inst_bSbox_AND_M31_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M31_U1_Step1_ins_U3 ( .A(Inst_bSbox_M20), .ZN(
        Inst_bSbox_AND_M31_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M31_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M31_U1_Step1_ins_n13), .B(Fresh[40]), .ZN(
        Inst_bSbox_AND_M31_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M31_U1_Step1_ins_U1 ( .A1(Inst_bSbox_M23), .A2(
        Inst_bSbox_M20), .ZN(Inst_bSbox_AND_M31_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M31_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M31_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M31_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M31_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M31_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M31_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M31_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M31_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M31_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M31_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M31_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M31_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M31_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M31_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M31_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M31_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3390) );
  OAI221_X1 Inst_bSbox_AND_M31_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M31_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M31_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M31_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M31_U1_Step1_reg[3]), .A(
        Inst_bSbox_AND_M31_U1_in1_reg[1]), .ZN(
        Inst_bSbox_AND_M31_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M31_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M31_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M31_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M31_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M31_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M31_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M31_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M31_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M31_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M31_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M31_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M31), 
        .QN() );
  XOR2_X1 Inst_bSbox_XOR_M33_U1_Ins_0_U1 ( .A(Inst_bSbox_M27), .B(
        Inst_bSbox_M25), .Z(Inst_bSbox_M33) );
  XOR2_X1 Inst_bSbox_XOR_M33_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3385), .B(
        new_AGEMA_signal_3384), .Z(new_AGEMA_signal_3391) );
  OAI21_X1 Inst_bSbox_AND_M34_U1_U4 ( .B1(new_AGEMA_signal_3373), .B2(
        Inst_bSbox_AND_M34_U1_n11), .A(Inst_bSbox_AND_M34_U1_n10), .ZN(
        Inst_bSbox_AND_M34_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M34_U1_U3 ( .B1(new_AGEMA_signal_3374), .B2(
        Fresh[45]), .C1(Inst_bSbox_AND_M34_U1_n9), .C2(Fresh[47]), .A(
        new_AGEMA_signal_3373), .ZN(Inst_bSbox_AND_M34_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M34_U1_U2 ( .A1(new_AGEMA_signal_3374), .A2(
        Fresh[46]), .B1(Fresh[44]), .B2(Inst_bSbox_AND_M34_U1_n9), .ZN(
        Inst_bSbox_AND_M34_U1_n11) );
  INV_X1 Inst_bSbox_AND_M34_U1_U1 ( .A(new_AGEMA_signal_3374), .ZN(
        Inst_bSbox_AND_M34_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M34_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3373), .CK(clk), .Q(Inst_bSbox_AND_M34_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M34_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3374), .CK(clk), .Q(Inst_bSbox_AND_M34_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M34_U1_Step1_ins_U9 ( .A(Fresh[47]), .B(
        Inst_bSbox_AND_M34_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M34_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M34_U1_Step1_ins_U8 ( .A1(Inst_bSbox_M21), .A2(
        Inst_bSbox_M22), .ZN(Inst_bSbox_AND_M34_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M34_U1_Step1_ins_U7 ( .A(Fresh[46]), .B(
        Inst_bSbox_AND_M34_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M34_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M34_U1_Step1_ins_U6 ( .A1(Inst_bSbox_M22), .A2(
        Inst_bSbox_AND_M34_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M34_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M34_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M34_U1_Step1_ins_n14), .B(Fresh[45]), .ZN(
        Inst_bSbox_AND_M34_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M34_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M34_U1_Step1_ins_n15), .A2(Inst_bSbox_M22), .ZN(
        Inst_bSbox_AND_M34_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M34_U1_Step1_ins_U3 ( .A(Inst_bSbox_M21), .ZN(
        Inst_bSbox_AND_M34_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M34_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M34_U1_Step1_ins_n13), .B(Fresh[44]), .ZN(
        Inst_bSbox_AND_M34_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M34_U1_Step1_ins_U1 ( .A1(Inst_bSbox_M22), .A2(
        Inst_bSbox_M21), .ZN(Inst_bSbox_AND_M34_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M34_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M34_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M34_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M34_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M34_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M34_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M34_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M34_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M34_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M34_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M34_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M34_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M34_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M34_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M34_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M34_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3386) );
  OAI221_X1 Inst_bSbox_AND_M34_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M34_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M34_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M34_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M34_U1_Step1_reg[3]), .A(
        Inst_bSbox_AND_M34_U1_in1_reg[1]), .ZN(
        Inst_bSbox_AND_M34_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M34_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M34_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M34_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M34_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M34_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M34_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M34_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M34_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M34_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M34_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M34_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M34), 
        .QN() );
  XOR2_X1 Inst_bSbox_XOR_M36_U1_Ins_0_U1 ( .A(Inst_bSbox_M24), .B(
        Inst_bSbox_M25), .Z(Inst_bSbox_M36) );
  XOR2_X1 Inst_bSbox_XOR_M36_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3387), .B(
        new_AGEMA_signal_3384), .Z(new_AGEMA_signal_3396) );
  OAI21_X1 Inst_bSbox_AND_M29_U1_U4 ( .B1(new_AGEMA_signal_3389), .B2(
        Inst_bSbox_AND_M29_U1_n11), .A(Inst_bSbox_AND_M29_U1_n10), .ZN(
        Inst_bSbox_AND_M29_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M29_U1_U3 ( .B1(new_AGEMA_signal_3385), .B2(
        Fresh[49]), .C1(Inst_bSbox_AND_M29_U1_n9), .C2(Fresh[51]), .A(
        new_AGEMA_signal_3389), .ZN(Inst_bSbox_AND_M29_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M29_U1_U2 ( .A1(new_AGEMA_signal_3385), .A2(
        Fresh[50]), .B1(Fresh[48]), .B2(Inst_bSbox_AND_M29_U1_n9), .ZN(
        Inst_bSbox_AND_M29_U1_n11) );
  INV_X1 Inst_bSbox_AND_M29_U1_U1 ( .A(new_AGEMA_signal_3385), .ZN(
        Inst_bSbox_AND_M29_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M29_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3389), .CK(clk), .Q(Inst_bSbox_AND_M29_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M29_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3385), .CK(clk), .Q(Inst_bSbox_AND_M29_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M29_U1_Step1_ins_U9 ( .A(Fresh[51]), .B(
        Inst_bSbox_AND_M29_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M29_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M29_U1_Step1_ins_U8 ( .A1(Inst_bSbox_M28), .A2(
        Inst_bSbox_M27), .ZN(Inst_bSbox_AND_M29_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M29_U1_Step1_ins_U7 ( .A(Fresh[50]), .B(
        Inst_bSbox_AND_M29_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M29_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M29_U1_Step1_ins_U6 ( .A1(Inst_bSbox_M27), .A2(
        Inst_bSbox_AND_M29_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M29_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M29_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M29_U1_Step1_ins_n14), .B(Fresh[49]), .ZN(
        Inst_bSbox_AND_M29_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M29_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M29_U1_Step1_ins_n15), .A2(Inst_bSbox_M27), .ZN(
        Inst_bSbox_AND_M29_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M29_U1_Step1_ins_U3 ( .A(Inst_bSbox_M28), .ZN(
        Inst_bSbox_AND_M29_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M29_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M29_U1_Step1_ins_n13), .B(Fresh[48]), .ZN(
        Inst_bSbox_AND_M29_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M29_U1_Step1_ins_U1 ( .A1(Inst_bSbox_M27), .A2(
        Inst_bSbox_M28), .ZN(Inst_bSbox_AND_M29_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M29_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M29_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M29_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M29_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M29_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M29_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M29_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M29_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M29_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M29_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M29_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M29_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M29_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M29_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M29_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M29_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3392) );
  OAI221_X1 Inst_bSbox_AND_M29_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M29_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M29_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M29_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M29_U1_Step1_reg[3]), .A(
        Inst_bSbox_AND_M29_U1_in1_reg[1]), .ZN(
        Inst_bSbox_AND_M29_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M29_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M29_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M29_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M29_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M29_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M29_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M29_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M29_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M29_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M29_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M29_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M29), 
        .QN() );
  OAI21_X1 Inst_bSbox_AND_M30_U1_U4 ( .B1(new_AGEMA_signal_3388), .B2(
        Inst_bSbox_AND_M30_U1_n11), .A(Inst_bSbox_AND_M30_U1_n10), .ZN(
        Inst_bSbox_AND_M30_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M30_U1_U3 ( .B1(new_AGEMA_signal_3387), .B2(
        Fresh[53]), .C1(Inst_bSbox_AND_M30_U1_n9), .C2(Fresh[55]), .A(
        new_AGEMA_signal_3388), .ZN(Inst_bSbox_AND_M30_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M30_U1_U2 ( .A1(new_AGEMA_signal_3387), .A2(
        Fresh[54]), .B1(Fresh[52]), .B2(Inst_bSbox_AND_M30_U1_n9), .ZN(
        Inst_bSbox_AND_M30_U1_n11) );
  INV_X1 Inst_bSbox_AND_M30_U1_U1 ( .A(new_AGEMA_signal_3387), .ZN(
        Inst_bSbox_AND_M30_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M30_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3388), .CK(clk), .Q(Inst_bSbox_AND_M30_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M30_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3387), .CK(clk), .Q(Inst_bSbox_AND_M30_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M30_U1_Step1_ins_U9 ( .A(Fresh[55]), .B(
        Inst_bSbox_AND_M30_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M30_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M30_U1_Step1_ins_U8 ( .A1(Inst_bSbox_M26), .A2(
        Inst_bSbox_M24), .ZN(Inst_bSbox_AND_M30_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M30_U1_Step1_ins_U7 ( .A(Fresh[54]), .B(
        Inst_bSbox_AND_M30_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M30_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M30_U1_Step1_ins_U6 ( .A1(Inst_bSbox_M24), .A2(
        Inst_bSbox_AND_M30_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M30_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M30_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M30_U1_Step1_ins_n14), .B(Fresh[53]), .ZN(
        Inst_bSbox_AND_M30_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M30_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M30_U1_Step1_ins_n15), .A2(Inst_bSbox_M24), .ZN(
        Inst_bSbox_AND_M30_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M30_U1_Step1_ins_U3 ( .A(Inst_bSbox_M26), .ZN(
        Inst_bSbox_AND_M30_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M30_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M30_U1_Step1_ins_n13), .B(Fresh[52]), .ZN(
        Inst_bSbox_AND_M30_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M30_U1_Step1_ins_U1 ( .A1(Inst_bSbox_M24), .A2(
        Inst_bSbox_M26), .ZN(Inst_bSbox_AND_M30_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M30_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M30_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M30_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M30_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M30_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M30_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M30_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M30_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M30_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M30_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M30_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M30_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M30_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M30_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M30_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M30_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3393) );
  OAI221_X1 Inst_bSbox_AND_M30_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M30_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M30_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M30_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M30_U1_Step1_reg[3]), .A(
        Inst_bSbox_AND_M30_U1_in1_reg[1]), .ZN(
        Inst_bSbox_AND_M30_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M30_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M30_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M30_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M30_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M30_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M30_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M30_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M30_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M30_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M30_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M30_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M30), 
        .QN() );
  OAI21_X1 Inst_bSbox_AND_M32_U1_U4 ( .B1(new_AGEMA_signal_3385), .B2(
        Inst_bSbox_AND_M32_U1_n11), .A(Inst_bSbox_AND_M32_U1_n10), .ZN(
        Inst_bSbox_AND_M32_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M32_U1_U3 ( .B1(new_AGEMA_signal_3390), .B2(
        Fresh[57]), .C1(Inst_bSbox_AND_M32_U1_n9), .C2(Fresh[59]), .A(
        new_AGEMA_signal_3385), .ZN(Inst_bSbox_AND_M32_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M32_U1_U2 ( .A1(new_AGEMA_signal_3390), .A2(
        Fresh[58]), .B1(Fresh[56]), .B2(Inst_bSbox_AND_M32_U1_n9), .ZN(
        Inst_bSbox_AND_M32_U1_n11) );
  INV_X1 Inst_bSbox_AND_M32_U1_U1 ( .A(new_AGEMA_signal_3390), .ZN(
        Inst_bSbox_AND_M32_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M32_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3385), .CK(clk), .Q(Inst_bSbox_AND_M32_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M32_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3390), .CK(clk), .Q(Inst_bSbox_AND_M32_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M32_U1_Step1_ins_U9 ( .A(Fresh[59]), .B(
        Inst_bSbox_AND_M32_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M32_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M32_U1_Step1_ins_U8 ( .A1(Inst_bSbox_M27), .A2(
        Inst_bSbox_M31), .ZN(Inst_bSbox_AND_M32_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M32_U1_Step1_ins_U7 ( .A(Fresh[58]), .B(
        Inst_bSbox_AND_M32_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M32_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M32_U1_Step1_ins_U6 ( .A1(Inst_bSbox_M31), .A2(
        Inst_bSbox_AND_M32_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M32_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M32_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M32_U1_Step1_ins_n14), .B(Fresh[57]), .ZN(
        Inst_bSbox_AND_M32_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M32_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M32_U1_Step1_ins_n15), .A2(Inst_bSbox_M31), .ZN(
        Inst_bSbox_AND_M32_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M32_U1_Step1_ins_U3 ( .A(Inst_bSbox_M27), .ZN(
        Inst_bSbox_AND_M32_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M32_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M32_U1_Step1_ins_n13), .B(Fresh[56]), .ZN(
        Inst_bSbox_AND_M32_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M32_U1_Step1_ins_U1 ( .A1(Inst_bSbox_M31), .A2(
        Inst_bSbox_M27), .ZN(Inst_bSbox_AND_M32_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M32_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M32_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M32_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M32_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M32_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M32_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M32_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M32_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M32_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M32_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M32_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M32_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M32_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M32_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M32_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M32_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3394) );
  OAI221_X1 Inst_bSbox_AND_M32_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M32_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M32_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M32_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M32_U1_Step1_reg[3]), .A(
        Inst_bSbox_AND_M32_U1_in1_reg[1]), .ZN(
        Inst_bSbox_AND_M32_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M32_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M32_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M32_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M32_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M32_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M32_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M32_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M32_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M32_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M32_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M32_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M32), 
        .QN() );
  OAI21_X1 Inst_bSbox_AND_M35_U1_U4 ( .B1(new_AGEMA_signal_3387), .B2(
        Inst_bSbox_AND_M35_U1_n11), .A(Inst_bSbox_AND_M35_U1_n10), .ZN(
        Inst_bSbox_AND_M35_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M35_U1_U3 ( .B1(new_AGEMA_signal_3386), .B2(
        Fresh[61]), .C1(Inst_bSbox_AND_M35_U1_n9), .C2(Fresh[63]), .A(
        new_AGEMA_signal_3387), .ZN(Inst_bSbox_AND_M35_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M35_U1_U2 ( .A1(new_AGEMA_signal_3386), .A2(
        Fresh[62]), .B1(Fresh[60]), .B2(Inst_bSbox_AND_M35_U1_n9), .ZN(
        Inst_bSbox_AND_M35_U1_n11) );
  INV_X1 Inst_bSbox_AND_M35_U1_U1 ( .A(new_AGEMA_signal_3386), .ZN(
        Inst_bSbox_AND_M35_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M35_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3387), .CK(clk), .Q(Inst_bSbox_AND_M35_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M35_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3386), .CK(clk), .Q(Inst_bSbox_AND_M35_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M35_U1_Step1_ins_U9 ( .A(Fresh[63]), .B(
        Inst_bSbox_AND_M35_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M35_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M35_U1_Step1_ins_U8 ( .A1(Inst_bSbox_M24), .A2(
        Inst_bSbox_M34), .ZN(Inst_bSbox_AND_M35_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M35_U1_Step1_ins_U7 ( .A(Fresh[62]), .B(
        Inst_bSbox_AND_M35_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M35_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M35_U1_Step1_ins_U6 ( .A1(Inst_bSbox_M34), .A2(
        Inst_bSbox_AND_M35_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M35_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M35_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M35_U1_Step1_ins_n14), .B(Fresh[61]), .ZN(
        Inst_bSbox_AND_M35_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M35_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M35_U1_Step1_ins_n15), .A2(Inst_bSbox_M34), .ZN(
        Inst_bSbox_AND_M35_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M35_U1_Step1_ins_U3 ( .A(Inst_bSbox_M24), .ZN(
        Inst_bSbox_AND_M35_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M35_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M35_U1_Step1_ins_n13), .B(Fresh[60]), .ZN(
        Inst_bSbox_AND_M35_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M35_U1_Step1_ins_U1 ( .A1(Inst_bSbox_M34), .A2(
        Inst_bSbox_M24), .ZN(Inst_bSbox_AND_M35_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M35_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M35_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M35_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M35_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M35_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M35_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M35_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M35_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M35_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M35_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M35_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M35_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M35_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M35_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M35_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M35_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3395) );
  OAI221_X1 Inst_bSbox_AND_M35_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M35_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M35_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M35_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M35_U1_Step1_reg[3]), .A(
        Inst_bSbox_AND_M35_U1_in1_reg[1]), .ZN(
        Inst_bSbox_AND_M35_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M35_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M35_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M35_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M35_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M35_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M35_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M35_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M35_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M35_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M35_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M35_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M35), 
        .QN() );
  XOR2_X1 Inst_bSbox_XOR_M37_U1_Ins_0_U1 ( .A(Inst_bSbox_M21), .B(
        Inst_bSbox_M29), .Z(Inst_bSbox_M37) );
  XOR2_X1 Inst_bSbox_XOR_M37_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3373), .B(
        new_AGEMA_signal_3392), .Z(new_AGEMA_signal_3397) );
  XOR2_X1 Inst_bSbox_XOR_M38_U1_Ins_0_U1 ( .A(Inst_bSbox_M32), .B(
        Inst_bSbox_M33), .Z(Inst_bSbox_M38) );
  XOR2_X1 Inst_bSbox_XOR_M38_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3394), .B(
        new_AGEMA_signal_3391), .Z(new_AGEMA_signal_3398) );
  XOR2_X1 Inst_bSbox_XOR_M39_U1_Ins_0_U1 ( .A(Inst_bSbox_M23), .B(
        Inst_bSbox_M30), .Z(Inst_bSbox_M39) );
  XOR2_X1 Inst_bSbox_XOR_M39_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3383), .B(
        new_AGEMA_signal_3393), .Z(new_AGEMA_signal_3399) );
  XOR2_X1 Inst_bSbox_XOR_M40_U1_Ins_0_U1 ( .A(Inst_bSbox_M35), .B(
        Inst_bSbox_M36), .Z(Inst_bSbox_M40) );
  XOR2_X1 Inst_bSbox_XOR_M40_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3395), .B(
        new_AGEMA_signal_3396), .Z(new_AGEMA_signal_3400) );
  XOR2_X1 Inst_bSbox_XOR_M41_U1_Ins_0_U1 ( .A(Inst_bSbox_M38), .B(
        Inst_bSbox_M40), .Z(Inst_bSbox_M41) );
  XOR2_X1 Inst_bSbox_XOR_M41_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3398), .B(
        new_AGEMA_signal_3400), .Z(new_AGEMA_signal_3401) );
  XOR2_X1 Inst_bSbox_XOR_M42_U1_Ins_0_U1 ( .A(Inst_bSbox_M37), .B(
        Inst_bSbox_M39), .Z(Inst_bSbox_M42) );
  XOR2_X1 Inst_bSbox_XOR_M42_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3397), .B(
        new_AGEMA_signal_3399), .Z(new_AGEMA_signal_3402) );
  XOR2_X1 Inst_bSbox_XOR_M43_U1_Ins_0_U1 ( .A(Inst_bSbox_M37), .B(
        Inst_bSbox_M38), .Z(Inst_bSbox_M43) );
  XOR2_X1 Inst_bSbox_XOR_M43_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3397), .B(
        new_AGEMA_signal_3398), .Z(new_AGEMA_signal_3403) );
  XOR2_X1 Inst_bSbox_XOR_M44_U1_Ins_0_U1 ( .A(Inst_bSbox_M39), .B(
        Inst_bSbox_M40), .Z(Inst_bSbox_M44) );
  XOR2_X1 Inst_bSbox_XOR_M44_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3399), .B(
        new_AGEMA_signal_3400), .Z(new_AGEMA_signal_3404) );
  XOR2_X1 Inst_bSbox_XOR_M45_U1_Ins_0_U1 ( .A(Inst_bSbox_M42), .B(
        Inst_bSbox_M41), .Z(Inst_bSbox_M45) );
  XOR2_X1 Inst_bSbox_XOR_M45_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3402), .B(
        new_AGEMA_signal_3401), .Z(new_AGEMA_signal_3413) );
  MUX2_X1 MUX_StateIn_mux_inst_0_U1_Ins_0_U1 ( .A(SboxOut[0]), .B(
        StateOutXORroundKey[0]), .S(n159), .Z(StateIn[0]) );
  MUX2_X1 MUX_StateIn_mux_inst_0_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3454), .B(
        new_AGEMA_signal_1984), .S(n159), .Z(new_AGEMA_signal_3455) );
  MUX2_X1 MUX_StateIn_mux_inst_1_U1_Ins_0_U1 ( .A(SboxOut[1]), .B(
        StateOutXORroundKey[1]), .S(n159), .Z(StateIn[1]) );
  MUX2_X1 MUX_StateIn_mux_inst_1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3463), .B(
        new_AGEMA_signal_1987), .S(n159), .Z(new_AGEMA_signal_3464) );
  MUX2_X1 MUX_StateIn_mux_inst_2_U1_Ins_0_U1 ( .A(SboxOut[2]), .B(
        StateOutXORroundKey[2]), .S(n159), .Z(StateIn[2]) );
  MUX2_X1 MUX_StateIn_mux_inst_2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3462), .B(
        new_AGEMA_signal_1990), .S(n159), .Z(new_AGEMA_signal_3465) );
  MUX2_X1 MUX_StateIn_mux_inst_3_U1_Ins_0_U1 ( .A(SboxOut[3]), .B(
        StateOutXORroundKey[3]), .S(n141), .Z(StateIn[3]) );
  MUX2_X1 MUX_StateIn_mux_inst_3_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3461), .B(
        new_AGEMA_signal_1993), .S(n141), .Z(new_AGEMA_signal_3466) );
  MUX2_X1 MUX_StateIn_mux_inst_4_U1_Ins_0_U1 ( .A(SboxOut[4]), .B(
        StateOutXORroundKey[4]), .S(n141), .Z(StateIn[4]) );
  MUX2_X1 MUX_StateIn_mux_inst_4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3460), .B(
        new_AGEMA_signal_1996), .S(n141), .Z(new_AGEMA_signal_3467) );
  MUX2_X1 MUX_StateIn_mux_inst_5_U1_Ins_0_U1 ( .A(SboxOut[5]), .B(
        StateOutXORroundKey[5]), .S(n141), .Z(StateIn[5]) );
  MUX2_X1 MUX_StateIn_mux_inst_5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3459), .B(
        new_AGEMA_signal_1999), .S(n141), .Z(new_AGEMA_signal_3468) );
  MUX2_X1 MUX_StateIn_mux_inst_6_U1_Ins_0_U1 ( .A(SboxOut[6]), .B(
        StateOutXORroundKey[6]), .S(n141), .Z(StateIn[6]) );
  MUX2_X1 MUX_StateIn_mux_inst_6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3458), .B(
        new_AGEMA_signal_2002), .S(n141), .Z(new_AGEMA_signal_3469) );
  MUX2_X1 MUX_StateIn_mux_inst_7_U1_Ins_0_U1 ( .A(SboxOut[7]), .B(
        StateOutXORroundKey[7]), .S(n141), .Z(StateIn[7]) );
  MUX2_X1 MUX_StateIn_mux_inst_7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3457), .B(
        new_AGEMA_signal_2005), .S(n141), .Z(new_AGEMA_signal_3470) );
  MUX2_X1 stateArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS33ser[0]), .B(ciphertext_s0[8]), .S(n197), .Z(
        stateArray_S33reg_gff_1_SFF_0_QD) );
  MUX2_X1 stateArray_S33reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3488), .B(ciphertext_s1[8]), .S(n197), .Z(
        new_AGEMA_signal_3497) );
  MUX2_X1 stateArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS33ser[1]), .B(ciphertext_s0[9]), .S(n191), .Z(
        stateArray_S33reg_gff_1_SFF_1_QD) );
  MUX2_X1 stateArray_S33reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3499), .B(ciphertext_s1[9]), .S(n191), .Z(
        new_AGEMA_signal_3520) );
  MUX2_X1 stateArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS33ser[2]), .B(ciphertext_s0[10]), .S(n197), .Z(
        stateArray_S33reg_gff_1_SFF_2_QD) );
  MUX2_X1 stateArray_S33reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3501), .B(ciphertext_s1[10]), .S(n197), .Z(
        new_AGEMA_signal_3521) );
  MUX2_X1 stateArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS33ser[3]), .B(ciphertext_s0[11]), .S(n192), .Z(
        stateArray_S33reg_gff_1_SFF_3_QD) );
  MUX2_X1 stateArray_S33reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3503), .B(ciphertext_s1[11]), .S(n192), .Z(
        new_AGEMA_signal_3522) );
  MUX2_X1 stateArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS33ser[4]), .B(ciphertext_s0[12]), .S(n192), .Z(
        stateArray_S33reg_gff_1_SFF_4_QD) );
  MUX2_X1 stateArray_S33reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3505), .B(ciphertext_s1[12]), .S(n192), .Z(
        new_AGEMA_signal_3523) );
  MUX2_X1 stateArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS33ser[5]), .B(ciphertext_s0[13]), .S(n192), .Z(
        stateArray_S33reg_gff_1_SFF_5_QD) );
  MUX2_X1 stateArray_S33reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3507), .B(ciphertext_s1[13]), .S(n192), .Z(
        new_AGEMA_signal_3524) );
  MUX2_X1 stateArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS33ser[6]), .B(ciphertext_s0[14]), .S(n191), .Z(
        stateArray_S33reg_gff_1_SFF_6_QD) );
  MUX2_X1 stateArray_S33reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3509), .B(ciphertext_s1[14]), .S(n191), .Z(
        new_AGEMA_signal_3525) );
  MUX2_X1 stateArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A(
        stateArray_inS33ser[7]), .B(ciphertext_s0[15]), .S(n191), .Z(
        stateArray_S33reg_gff_1_SFF_7_QD) );
  MUX2_X1 stateArray_S33reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3511), .B(ciphertext_s1[15]), .S(n191), .Z(
        new_AGEMA_signal_3526) );
  MUX2_X1 stateArray_MUX_input_MC_mux_inst_0_U1_Ins_0_U1 ( .A(StateIn[0]), .B(
        StateInMC[0]), .S(n174), .Z(stateArray_input_MC[0]) );
  MUX2_X1 stateArray_MUX_input_MC_mux_inst_0_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3455), .B(new_AGEMA_signal_2860), .S(n174), .Z(
        new_AGEMA_signal_3471) );
  MUX2_X1 stateArray_MUX_input_MC_mux_inst_1_U1_Ins_0_U1 ( .A(StateIn[1]), .B(
        StateInMC[1]), .S(n174), .Z(stateArray_input_MC[1]) );
  MUX2_X1 stateArray_MUX_input_MC_mux_inst_1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3464), .B(new_AGEMA_signal_2861), .S(n174), .Z(
        new_AGEMA_signal_3480) );
  MUX2_X1 stateArray_MUX_input_MC_mux_inst_2_U1_Ins_0_U1 ( .A(StateIn[2]), .B(
        StateInMC[2]), .S(n175), .Z(stateArray_input_MC[2]) );
  MUX2_X1 stateArray_MUX_input_MC_mux_inst_2_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3465), .B(new_AGEMA_signal_2834), .S(n175), .Z(
        new_AGEMA_signal_3481) );
  MUX2_X1 stateArray_MUX_input_MC_mux_inst_3_U1_Ins_0_U1 ( .A(StateIn[3]), .B(
        StateInMC[3]), .S(n175), .Z(stateArray_input_MC[3]) );
  MUX2_X1 stateArray_MUX_input_MC_mux_inst_3_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3466), .B(new_AGEMA_signal_2862), .S(n175), .Z(
        new_AGEMA_signal_3482) );
  MUX2_X1 stateArray_MUX_input_MC_mux_inst_4_U1_Ins_0_U1 ( .A(StateIn[4]), .B(
        StateInMC[4]), .S(n175), .Z(stateArray_input_MC[4]) );
  MUX2_X1 stateArray_MUX_input_MC_mux_inst_4_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3467), .B(new_AGEMA_signal_2863), .S(n175), .Z(
        new_AGEMA_signal_3483) );
  MUX2_X1 stateArray_MUX_input_MC_mux_inst_5_U1_Ins_0_U1 ( .A(StateIn[5]), .B(
        StateInMC[5]), .S(n175), .Z(stateArray_input_MC[5]) );
  MUX2_X1 stateArray_MUX_input_MC_mux_inst_5_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3468), .B(new_AGEMA_signal_2835), .S(n175), .Z(
        new_AGEMA_signal_3484) );
  MUX2_X1 stateArray_MUX_input_MC_mux_inst_6_U1_Ins_0_U1 ( .A(StateIn[6]), .B(
        StateInMC[6]), .S(n175), .Z(stateArray_input_MC[6]) );
  MUX2_X1 stateArray_MUX_input_MC_mux_inst_6_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3469), .B(new_AGEMA_signal_2836), .S(n175), .Z(
        new_AGEMA_signal_3485) );
  MUX2_X1 stateArray_MUX_input_MC_mux_inst_7_U1_Ins_0_U1 ( .A(StateIn[7]), .B(
        StateInMC[7]), .S(n175), .Z(stateArray_input_MC[7]) );
  MUX2_X1 stateArray_MUX_input_MC_mux_inst_7_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_3470), .B(new_AGEMA_signal_2837), .S(n175), .Z(
        new_AGEMA_signal_3486) );
  MUX2_X1 stateArray_MUX_inS33ser_mux_inst_0_U1_Ins_0_U1 ( .A(plaintext_s0[0]), 
        .B(stateArray_input_MC[0]), .S(n211), .Z(stateArray_inS33ser[0]) );
  MUX2_X1 stateArray_MUX_inS33ser_mux_inst_0_U1_Ins_1_U1 ( .A(plaintext_s1[0]), 
        .B(new_AGEMA_signal_3471), .S(n211), .Z(new_AGEMA_signal_3488) );
  MUX2_X1 stateArray_MUX_inS33ser_mux_inst_1_U1_Ins_0_U1 ( .A(plaintext_s0[1]), 
        .B(stateArray_input_MC[1]), .S(n212), .Z(stateArray_inS33ser[1]) );
  MUX2_X1 stateArray_MUX_inS33ser_mux_inst_1_U1_Ins_1_U1 ( .A(plaintext_s1[1]), 
        .B(new_AGEMA_signal_3480), .S(n212), .Z(new_AGEMA_signal_3499) );
  MUX2_X1 stateArray_MUX_inS33ser_mux_inst_2_U1_Ins_0_U1 ( .A(plaintext_s0[2]), 
        .B(stateArray_input_MC[2]), .S(n206), .Z(stateArray_inS33ser[2]) );
  MUX2_X1 stateArray_MUX_inS33ser_mux_inst_2_U1_Ins_1_U1 ( .A(plaintext_s1[2]), 
        .B(new_AGEMA_signal_3481), .S(n206), .Z(new_AGEMA_signal_3501) );
  MUX2_X1 stateArray_MUX_inS33ser_mux_inst_3_U1_Ins_0_U1 ( .A(plaintext_s0[3]), 
        .B(stateArray_input_MC[3]), .S(n207), .Z(stateArray_inS33ser[3]) );
  MUX2_X1 stateArray_MUX_inS33ser_mux_inst_3_U1_Ins_1_U1 ( .A(plaintext_s1[3]), 
        .B(new_AGEMA_signal_3482), .S(n207), .Z(new_AGEMA_signal_3503) );
  MUX2_X1 stateArray_MUX_inS33ser_mux_inst_4_U1_Ins_0_U1 ( .A(plaintext_s0[4]), 
        .B(stateArray_input_MC[4]), .S(n209), .Z(stateArray_inS33ser[4]) );
  MUX2_X1 stateArray_MUX_inS33ser_mux_inst_4_U1_Ins_1_U1 ( .A(plaintext_s1[4]), 
        .B(new_AGEMA_signal_3483), .S(n209), .Z(new_AGEMA_signal_3505) );
  MUX2_X1 stateArray_MUX_inS33ser_mux_inst_5_U1_Ins_0_U1 ( .A(plaintext_s0[5]), 
        .B(stateArray_input_MC[5]), .S(n210), .Z(stateArray_inS33ser[5]) );
  MUX2_X1 stateArray_MUX_inS33ser_mux_inst_5_U1_Ins_1_U1 ( .A(plaintext_s1[5]), 
        .B(new_AGEMA_signal_3484), .S(n210), .Z(new_AGEMA_signal_3507) );
  MUX2_X1 stateArray_MUX_inS33ser_mux_inst_6_U1_Ins_0_U1 ( .A(plaintext_s0[6]), 
        .B(stateArray_input_MC[6]), .S(n219), .Z(stateArray_inS33ser[6]) );
  MUX2_X1 stateArray_MUX_inS33ser_mux_inst_6_U1_Ins_1_U1 ( .A(plaintext_s1[6]), 
        .B(new_AGEMA_signal_3485), .S(n219), .Z(new_AGEMA_signal_3509) );
  MUX2_X1 stateArray_MUX_inS33ser_mux_inst_7_U1_Ins_0_U1 ( .A(plaintext_s0[7]), 
        .B(stateArray_input_MC[7]), .S(n220), .Z(stateArray_inS33ser[7]) );
  MUX2_X1 stateArray_MUX_inS33ser_mux_inst_7_U1_Ins_1_U1 ( .A(plaintext_s1[7]), 
        .B(new_AGEMA_signal_3486), .S(n220), .Z(new_AGEMA_signal_3511) );
  XNOR2_X1 KeyArray_U42_Ins0_U1 ( .A(KeyArray_n55), .B(keyStateIn[7]), .ZN(
        KeyArray_inS30par[7]) );
  XOR2_X1 KeyArray_U42_Ins_1_U1 ( .A(new_AGEMA_signal_3472), .B(
        new_AGEMA_signal_2004), .Z(new_AGEMA_signal_3489) );
  XNOR2_X1 KeyArray_U41_Ins0_U1 ( .A(roundConstant[7]), .B(SboxOut[7]), .ZN(
        KeyArray_n55) );
  XOR2_X1 KeyArray_U41_Ins_1_U1 ( .A(1'b0), .B(new_AGEMA_signal_3457), .Z(
        new_AGEMA_signal_3472) );
  XNOR2_X1 KeyArray_U40_Ins0_U1 ( .A(KeyArray_n54), .B(keyStateIn[6]), .ZN(
        KeyArray_inS30par[6]) );
  XOR2_X1 KeyArray_U40_Ins_1_U1 ( .A(new_AGEMA_signal_3473), .B(
        new_AGEMA_signal_2001), .Z(new_AGEMA_signal_3490) );
  XNOR2_X1 KeyArray_U39_Ins0_U1 ( .A(roundConstant[6]), .B(SboxOut[6]), .ZN(
        KeyArray_n54) );
  XOR2_X1 KeyArray_U39_Ins_1_U1 ( .A(1'b0), .B(new_AGEMA_signal_3458), .Z(
        new_AGEMA_signal_3473) );
  XNOR2_X1 KeyArray_U38_Ins0_U1 ( .A(KeyArray_n53), .B(keyStateIn[5]), .ZN(
        KeyArray_inS30par[5]) );
  XOR2_X1 KeyArray_U38_Ins_1_U1 ( .A(new_AGEMA_signal_3474), .B(
        new_AGEMA_signal_1998), .Z(new_AGEMA_signal_3491) );
  XNOR2_X1 KeyArray_U37_Ins0_U1 ( .A(roundConstant[5]), .B(SboxOut[5]), .ZN(
        KeyArray_n53) );
  XOR2_X1 KeyArray_U37_Ins_1_U1 ( .A(1'b0), .B(new_AGEMA_signal_3459), .Z(
        new_AGEMA_signal_3474) );
  XNOR2_X1 KeyArray_U36_Ins0_U1 ( .A(KeyArray_n52), .B(keyStateIn[4]), .ZN(
        KeyArray_inS30par[4]) );
  XOR2_X1 KeyArray_U36_Ins_1_U1 ( .A(new_AGEMA_signal_3475), .B(
        new_AGEMA_signal_1995), .Z(new_AGEMA_signal_3492) );
  XNOR2_X1 KeyArray_U35_Ins0_U1 ( .A(roundConstant[4]), .B(SboxOut[4]), .ZN(
        KeyArray_n52) );
  XOR2_X1 KeyArray_U35_Ins_1_U1 ( .A(1'b0), .B(new_AGEMA_signal_3460), .Z(
        new_AGEMA_signal_3475) );
  XNOR2_X1 KeyArray_U34_Ins0_U1 ( .A(KeyArray_n51), .B(keyStateIn[3]), .ZN(
        KeyArray_inS30par[3]) );
  XOR2_X1 KeyArray_U34_Ins_1_U1 ( .A(new_AGEMA_signal_3476), .B(
        new_AGEMA_signal_1992), .Z(new_AGEMA_signal_3493) );
  XNOR2_X1 KeyArray_U33_Ins0_U1 ( .A(roundConstant[3]), .B(SboxOut[3]), .ZN(
        KeyArray_n51) );
  XOR2_X1 KeyArray_U33_Ins_1_U1 ( .A(1'b0), .B(new_AGEMA_signal_3461), .Z(
        new_AGEMA_signal_3476) );
  XNOR2_X1 KeyArray_U32_Ins0_U1 ( .A(KeyArray_n50), .B(keyStateIn[2]), .ZN(
        KeyArray_inS30par[2]) );
  XOR2_X1 KeyArray_U32_Ins_1_U1 ( .A(new_AGEMA_signal_3477), .B(
        new_AGEMA_signal_1989), .Z(new_AGEMA_signal_3494) );
  XNOR2_X1 KeyArray_U31_Ins0_U1 ( .A(roundConstant[2]), .B(SboxOut[2]), .ZN(
        KeyArray_n50) );
  XOR2_X1 KeyArray_U31_Ins_1_U1 ( .A(1'b0), .B(new_AGEMA_signal_3462), .Z(
        new_AGEMA_signal_3477) );
  XNOR2_X1 KeyArray_U30_Ins0_U1 ( .A(KeyArray_n49), .B(keyStateIn[1]), .ZN(
        KeyArray_inS30par[1]) );
  XOR2_X1 KeyArray_U30_Ins_1_U1 ( .A(new_AGEMA_signal_3478), .B(
        new_AGEMA_signal_1986), .Z(new_AGEMA_signal_3495) );
  XNOR2_X1 KeyArray_U29_Ins0_U1 ( .A(roundConstant[1]), .B(SboxOut[1]), .ZN(
        KeyArray_n49) );
  XOR2_X1 KeyArray_U29_Ins_1_U1 ( .A(1'b0), .B(new_AGEMA_signal_3463), .Z(
        new_AGEMA_signal_3478) );
  XNOR2_X1 KeyArray_U28_Ins0_U1 ( .A(KeyArray_n48), .B(keyStateIn[0]), .ZN(
        KeyArray_inS30par[0]) );
  XOR2_X1 KeyArray_U28_Ins_1_U1 ( .A(new_AGEMA_signal_3456), .B(
        new_AGEMA_signal_1983), .Z(new_AGEMA_signal_3479) );
  XNOR2_X1 KeyArray_U27_Ins0_U1 ( .A(roundConstant[0]), .B(SboxOut[0]), .ZN(
        KeyArray_n48) );
  XOR2_X1 KeyArray_U27_Ins_1_U1 ( .A(1'b0), .B(new_AGEMA_signal_3454), .Z(
        new_AGEMA_signal_3456) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_0_U1_Ins_0_U1 ( .A(KeyArray_outS30ser[0]), 
        .B(KeyArray_S30reg_gff_1_SFF_0_QD), .S(n186), .Z(
        KeyArray_S30reg_gff_1_SFF_0_n5) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_0_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2683), 
        .B(new_AGEMA_signal_3496), .S(n186), .Z(new_AGEMA_signal_3512) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS30ser[0]), .B(KeyArray_inS30par[0]), .S(n175), .Z(
        KeyArray_S30reg_gff_1_SFF_0_QD) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2708), .B(new_AGEMA_signal_3479), .S(n175), .Z(
        new_AGEMA_signal_3496) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_1_U1_Ins_0_U1 ( .A(KeyArray_outS30ser[1]), 
        .B(KeyArray_S30reg_gff_1_SFF_1_QD), .S(n179), .Z(
        KeyArray_S30reg_gff_1_SFF_1_n5) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2686), 
        .B(new_AGEMA_signal_3513), .S(n179), .Z(new_AGEMA_signal_3527) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS30ser[1]), .B(KeyArray_inS30par[1]), .S(n176), .Z(
        KeyArray_S30reg_gff_1_SFF_1_QD) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2711), .B(new_AGEMA_signal_3495), .S(n176), .Z(
        new_AGEMA_signal_3513) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_2_U1_Ins_0_U1 ( .A(KeyArray_outS30ser[2]), 
        .B(KeyArray_S30reg_gff_1_SFF_2_QD), .S(n183), .Z(
        KeyArray_S30reg_gff_1_SFF_2_n5) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2689), 
        .B(new_AGEMA_signal_3514), .S(n183), .Z(new_AGEMA_signal_3528) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS30ser[2]), .B(KeyArray_inS30par[2]), .S(n176), .Z(
        KeyArray_S30reg_gff_1_SFF_2_QD) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2714), .B(new_AGEMA_signal_3494), .S(n176), .Z(
        new_AGEMA_signal_3514) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_3_U1_Ins_0_U1 ( .A(KeyArray_outS30ser[3]), 
        .B(KeyArray_S30reg_gff_1_SFF_3_QD), .S(n190), .Z(
        KeyArray_S30reg_gff_1_SFF_3_n5) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_3_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2692), 
        .B(new_AGEMA_signal_3515), .S(n190), .Z(new_AGEMA_signal_3529) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS30ser[3]), .B(KeyArray_inS30par[3]), .S(n176), .Z(
        KeyArray_S30reg_gff_1_SFF_3_QD) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2717), .B(new_AGEMA_signal_3493), .S(n176), .Z(
        new_AGEMA_signal_3515) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_4_U1_Ins_0_U1 ( .A(KeyArray_outS30ser[4]), 
        .B(KeyArray_S30reg_gff_1_SFF_4_QD), .S(n190), .Z(
        KeyArray_S30reg_gff_1_SFF_4_n5) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2695), 
        .B(new_AGEMA_signal_3516), .S(n190), .Z(new_AGEMA_signal_3530) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS30ser[4]), .B(KeyArray_inS30par[4]), .S(n176), .Z(
        KeyArray_S30reg_gff_1_SFF_4_QD) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2720), .B(new_AGEMA_signal_3492), .S(n176), .Z(
        new_AGEMA_signal_3516) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_5_U1_Ins_0_U1 ( .A(KeyArray_outS30ser[5]), 
        .B(KeyArray_S30reg_gff_1_SFF_5_QD), .S(n188), .Z(
        KeyArray_S30reg_gff_1_SFF_5_n5) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2698), 
        .B(new_AGEMA_signal_3517), .S(n188), .Z(new_AGEMA_signal_3531) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS30ser[5]), .B(KeyArray_inS30par[5]), .S(n176), .Z(
        KeyArray_S30reg_gff_1_SFF_5_QD) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2723), .B(new_AGEMA_signal_3491), .S(n176), .Z(
        new_AGEMA_signal_3517) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_6_U1_Ins_0_U1 ( .A(KeyArray_outS30ser[6]), 
        .B(KeyArray_S30reg_gff_1_SFF_6_QD), .S(n181), .Z(
        KeyArray_S30reg_gff_1_SFF_6_n5) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2701), 
        .B(new_AGEMA_signal_3518), .S(n181), .Z(new_AGEMA_signal_3532) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS30ser[6]), .B(KeyArray_inS30par[6]), .S(n176), .Z(
        KeyArray_S30reg_gff_1_SFF_6_QD) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2726), .B(new_AGEMA_signal_3490), .S(n176), .Z(
        new_AGEMA_signal_3518) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_7_U1_Ins_0_U1 ( .A(KeyArray_outS30ser[7]), 
        .B(KeyArray_S30reg_gff_1_SFF_7_QD), .S(n189), .Z(
        KeyArray_S30reg_gff_1_SFF_7_n5) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2704), 
        .B(new_AGEMA_signal_3519), .S(n189), .Z(new_AGEMA_signal_3533) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_0_U1 ( .A(
        KeyArray_inS30ser[7]), .B(KeyArray_inS30par[7]), .S(n176), .Z(
        KeyArray_S30reg_gff_1_SFF_7_QD) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2729), .B(new_AGEMA_signal_3489), .S(n176), .Z(
        new_AGEMA_signal_3519) );
  OAI21_X1 Inst_bSbox_AND_M46_U1_U4 ( .B1(new_AGEMA_signal_3404), .B2(
        Inst_bSbox_AND_M46_U1_n11), .A(Inst_bSbox_AND_M46_U1_n10), .ZN(
        Inst_bSbox_AND_M46_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M46_U1_U3 ( .B1(new_AGEMA_signal_3000), .B2(
        Fresh[65]), .C1(Inst_bSbox_AND_M46_U1_n9), .C2(Fresh[67]), .A(
        new_AGEMA_signal_3404), .ZN(Inst_bSbox_AND_M46_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M46_U1_U2 ( .A1(new_AGEMA_signal_3000), .A2(
        Fresh[66]), .B1(Fresh[64]), .B2(Inst_bSbox_AND_M46_U1_n9), .ZN(
        Inst_bSbox_AND_M46_U1_n11) );
  INV_X1 Inst_bSbox_AND_M46_U1_U1 ( .A(new_AGEMA_signal_3000), .ZN(
        Inst_bSbox_AND_M46_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M46_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3404), .CK(clk), .Q(Inst_bSbox_AND_M46_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M46_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3000), .CK(clk), .Q(Inst_bSbox_AND_M46_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M46_U1_Step1_ins_U9 ( .A(Fresh[67]), .B(
        Inst_bSbox_AND_M46_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M46_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M46_U1_Step1_ins_U8 ( .A1(Inst_bSbox_M44), .A2(
        Inst_bSbox_T6), .ZN(Inst_bSbox_AND_M46_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M46_U1_Step1_ins_U7 ( .A(Fresh[66]), .B(
        Inst_bSbox_AND_M46_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M46_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M46_U1_Step1_ins_U6 ( .A1(Inst_bSbox_T6), .A2(
        Inst_bSbox_AND_M46_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M46_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M46_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M46_U1_Step1_ins_n14), .B(Fresh[65]), .ZN(
        Inst_bSbox_AND_M46_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M46_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M46_U1_Step1_ins_n15), .A2(Inst_bSbox_T6), .ZN(
        Inst_bSbox_AND_M46_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M46_U1_Step1_ins_U3 ( .A(Inst_bSbox_M44), .ZN(
        Inst_bSbox_AND_M46_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M46_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M46_U1_Step1_ins_n13), .B(Fresh[64]), .ZN(
        Inst_bSbox_AND_M46_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M46_U1_Step1_ins_U1 ( .A1(Inst_bSbox_T6), .A2(
        Inst_bSbox_M44), .ZN(Inst_bSbox_AND_M46_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M46_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M46_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M46_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M46_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M46_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M46_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M46_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M46_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M46_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M46_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M46_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M46_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M46_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M46_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M46_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M46_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3414) );
  OAI221_X1 Inst_bSbox_AND_M46_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M46_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M46_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M46_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M46_U1_Step1_reg[3]), .A(
        Inst_bSbox_AND_M46_U1_in1_reg[1]), .ZN(
        Inst_bSbox_AND_M46_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M46_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M46_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M46_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M46_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M46_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M46_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M46_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M46_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M46_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M46_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M46_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M46), 
        .QN() );
  OAI21_X1 Inst_bSbox_AND_M47_U1_U4 ( .B1(new_AGEMA_signal_3400), .B2(
        Inst_bSbox_AND_M47_U1_n11), .A(Inst_bSbox_AND_M47_U1_n10), .ZN(
        Inst_bSbox_AND_M47_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M47_U1_U3 ( .B1(new_AGEMA_signal_3032), .B2(
        Fresh[69]), .C1(Inst_bSbox_AND_M47_U1_n9), .C2(Fresh[71]), .A(
        new_AGEMA_signal_3400), .ZN(Inst_bSbox_AND_M47_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M47_U1_U2 ( .A1(new_AGEMA_signal_3032), .A2(
        Fresh[70]), .B1(Fresh[68]), .B2(Inst_bSbox_AND_M47_U1_n9), .ZN(
        Inst_bSbox_AND_M47_U1_n11) );
  INV_X1 Inst_bSbox_AND_M47_U1_U1 ( .A(new_AGEMA_signal_3032), .ZN(
        Inst_bSbox_AND_M47_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M47_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3400), .CK(clk), .Q(Inst_bSbox_AND_M47_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M47_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3032), .CK(clk), .Q(Inst_bSbox_AND_M47_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M47_U1_Step1_ins_U9 ( .A(Fresh[71]), .B(
        Inst_bSbox_AND_M47_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M47_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M47_U1_Step1_ins_U8 ( .A1(Inst_bSbox_M40), .A2(
        Inst_bSbox_T8), .ZN(Inst_bSbox_AND_M47_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M47_U1_Step1_ins_U7 ( .A(Fresh[70]), .B(
        Inst_bSbox_AND_M47_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M47_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M47_U1_Step1_ins_U6 ( .A1(Inst_bSbox_T8), .A2(
        Inst_bSbox_AND_M47_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M47_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M47_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M47_U1_Step1_ins_n14), .B(Fresh[69]), .ZN(
        Inst_bSbox_AND_M47_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M47_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M47_U1_Step1_ins_n15), .A2(Inst_bSbox_T8), .ZN(
        Inst_bSbox_AND_M47_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M47_U1_Step1_ins_U3 ( .A(Inst_bSbox_M40), .ZN(
        Inst_bSbox_AND_M47_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M47_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M47_U1_Step1_ins_n13), .B(Fresh[68]), .ZN(
        Inst_bSbox_AND_M47_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M47_U1_Step1_ins_U1 ( .A1(Inst_bSbox_T8), .A2(
        Inst_bSbox_M40), .ZN(Inst_bSbox_AND_M47_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M47_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M47_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M47_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M47_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M47_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M47_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M47_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M47_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M47_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M47_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M47_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M47_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M47_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M47_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M47_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M47_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3405) );
  OAI221_X1 Inst_bSbox_AND_M47_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M47_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M47_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M47_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M47_U1_Step1_reg[3]), .A(
        Inst_bSbox_AND_M47_U1_in1_reg[1]), .ZN(
        Inst_bSbox_AND_M47_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M47_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M47_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M47_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M47_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M47_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M47_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M47_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M47_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M47_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M47_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M47_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M47), 
        .QN() );
  OAI21_X1 Inst_bSbox_AND_M48_U1_U4 ( .B1(new_AGEMA_signal_3399), .B2(
        Inst_bSbox_AND_M48_U1_n11), .A(Inst_bSbox_AND_M48_U1_n10), .ZN(
        Inst_bSbox_AND_M48_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M48_U1_U3 ( .B1(new_AGEMA_signal_2826), .B2(
        Fresh[73]), .C1(Inst_bSbox_AND_M48_U1_n9), .C2(Fresh[75]), .A(
        new_AGEMA_signal_3399), .ZN(Inst_bSbox_AND_M48_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M48_U1_U2 ( .A1(new_AGEMA_signal_2826), .A2(
        Fresh[74]), .B1(Fresh[72]), .B2(Inst_bSbox_AND_M48_U1_n9), .ZN(
        Inst_bSbox_AND_M48_U1_n11) );
  INV_X1 Inst_bSbox_AND_M48_U1_U1 ( .A(new_AGEMA_signal_2826), .ZN(
        Inst_bSbox_AND_M48_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M48_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3399), .CK(clk), .Q(Inst_bSbox_AND_M48_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M48_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_2826), .CK(clk), .Q(Inst_bSbox_AND_M48_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M48_U1_Step1_ins_U9 ( .A(Fresh[75]), .B(
        Inst_bSbox_AND_M48_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M48_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M48_U1_Step1_ins_U8 ( .A1(Inst_bSbox_M39), .A2(
        SboxIn[0]), .ZN(Inst_bSbox_AND_M48_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M48_U1_Step1_ins_U7 ( .A(Fresh[74]), .B(
        Inst_bSbox_AND_M48_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M48_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M48_U1_Step1_ins_U6 ( .A1(SboxIn[0]), .A2(
        Inst_bSbox_AND_M48_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M48_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M48_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M48_U1_Step1_ins_n14), .B(Fresh[73]), .ZN(
        Inst_bSbox_AND_M48_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M48_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M48_U1_Step1_ins_n15), .A2(SboxIn[0]), .ZN(
        Inst_bSbox_AND_M48_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M48_U1_Step1_ins_U3 ( .A(Inst_bSbox_M39), .ZN(
        Inst_bSbox_AND_M48_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M48_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M48_U1_Step1_ins_n13), .B(Fresh[72]), .ZN(
        Inst_bSbox_AND_M48_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M48_U1_Step1_ins_U1 ( .A1(SboxIn[0]), .A2(
        Inst_bSbox_M39), .ZN(Inst_bSbox_AND_M48_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M48_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M48_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M48_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M48_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M48_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M48_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M48_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M48_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M48_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M48_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M48_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M48_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M48_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M48_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M48_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M48_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3406) );
  OAI221_X1 Inst_bSbox_AND_M48_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M48_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M48_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M48_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M48_U1_Step1_reg[3]), .A(
        Inst_bSbox_AND_M48_U1_in1_reg[1]), .ZN(
        Inst_bSbox_AND_M48_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M48_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M48_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M48_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M48_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M48_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M48_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M48_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M48_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M48_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M48_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M48_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M48), 
        .QN() );
  OAI21_X1 Inst_bSbox_AND_M49_U1_U4 ( .B1(new_AGEMA_signal_3403), .B2(
        Inst_bSbox_AND_M49_U1_n11), .A(Inst_bSbox_AND_M49_U1_n10), .ZN(
        Inst_bSbox_AND_M49_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M49_U1_U3 ( .B1(new_AGEMA_signal_3004), .B2(
        Fresh[77]), .C1(Inst_bSbox_AND_M49_U1_n9), .C2(Fresh[79]), .A(
        new_AGEMA_signal_3403), .ZN(Inst_bSbox_AND_M49_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M49_U1_U2 ( .A1(new_AGEMA_signal_3004), .A2(
        Fresh[78]), .B1(Fresh[76]), .B2(Inst_bSbox_AND_M49_U1_n9), .ZN(
        Inst_bSbox_AND_M49_U1_n11) );
  INV_X1 Inst_bSbox_AND_M49_U1_U1 ( .A(new_AGEMA_signal_3004), .ZN(
        Inst_bSbox_AND_M49_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M49_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3403), .CK(clk), .Q(Inst_bSbox_AND_M49_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M49_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3004), .CK(clk), .Q(Inst_bSbox_AND_M49_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M49_U1_Step1_ins_U9 ( .A(Fresh[79]), .B(
        Inst_bSbox_AND_M49_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M49_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M49_U1_Step1_ins_U8 ( .A1(Inst_bSbox_M43), .A2(
        Inst_bSbox_T16), .ZN(Inst_bSbox_AND_M49_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M49_U1_Step1_ins_U7 ( .A(Fresh[78]), .B(
        Inst_bSbox_AND_M49_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M49_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M49_U1_Step1_ins_U6 ( .A1(Inst_bSbox_T16), .A2(
        Inst_bSbox_AND_M49_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M49_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M49_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M49_U1_Step1_ins_n14), .B(Fresh[77]), .ZN(
        Inst_bSbox_AND_M49_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M49_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M49_U1_Step1_ins_n15), .A2(Inst_bSbox_T16), .ZN(
        Inst_bSbox_AND_M49_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M49_U1_Step1_ins_U3 ( .A(Inst_bSbox_M43), .ZN(
        Inst_bSbox_AND_M49_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M49_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M49_U1_Step1_ins_n13), .B(Fresh[76]), .ZN(
        Inst_bSbox_AND_M49_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M49_U1_Step1_ins_U1 ( .A1(Inst_bSbox_T16), .A2(
        Inst_bSbox_M43), .ZN(Inst_bSbox_AND_M49_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M49_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M49_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M49_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M49_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M49_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M49_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M49_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M49_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M49_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M49_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M49_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M49_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M49_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M49_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M49_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M49_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3415) );
  OAI221_X1 Inst_bSbox_AND_M49_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M49_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M49_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M49_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M49_U1_Step1_reg[3]), .A(
        Inst_bSbox_AND_M49_U1_in1_reg[1]), .ZN(
        Inst_bSbox_AND_M49_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M49_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M49_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M49_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M49_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M49_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M49_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M49_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M49_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M49_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M49_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M49_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M49), 
        .QN() );
  OAI21_X1 Inst_bSbox_AND_M50_U1_U4 ( .B1(new_AGEMA_signal_3398), .B2(
        Inst_bSbox_AND_M50_U1_n11), .A(Inst_bSbox_AND_M50_U1_n10), .ZN(
        Inst_bSbox_AND_M50_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M50_U1_U3 ( .B1(new_AGEMA_signal_3001), .B2(
        Fresh[81]), .C1(Inst_bSbox_AND_M50_U1_n9), .C2(Fresh[83]), .A(
        new_AGEMA_signal_3398), .ZN(Inst_bSbox_AND_M50_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M50_U1_U2 ( .A1(new_AGEMA_signal_3001), .A2(
        Fresh[82]), .B1(Fresh[80]), .B2(Inst_bSbox_AND_M50_U1_n9), .ZN(
        Inst_bSbox_AND_M50_U1_n11) );
  INV_X1 Inst_bSbox_AND_M50_U1_U1 ( .A(new_AGEMA_signal_3001), .ZN(
        Inst_bSbox_AND_M50_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M50_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3398), .CK(clk), .Q(Inst_bSbox_AND_M50_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M50_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3001), .CK(clk), .Q(Inst_bSbox_AND_M50_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M50_U1_Step1_ins_U9 ( .A(Fresh[83]), .B(
        Inst_bSbox_AND_M50_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M50_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M50_U1_Step1_ins_U8 ( .A1(Inst_bSbox_M38), .A2(
        Inst_bSbox_T9), .ZN(Inst_bSbox_AND_M50_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M50_U1_Step1_ins_U7 ( .A(Fresh[82]), .B(
        Inst_bSbox_AND_M50_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M50_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M50_U1_Step1_ins_U6 ( .A1(Inst_bSbox_T9), .A2(
        Inst_bSbox_AND_M50_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M50_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M50_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M50_U1_Step1_ins_n14), .B(Fresh[81]), .ZN(
        Inst_bSbox_AND_M50_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M50_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M50_U1_Step1_ins_n15), .A2(Inst_bSbox_T9), .ZN(
        Inst_bSbox_AND_M50_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M50_U1_Step1_ins_U3 ( .A(Inst_bSbox_M38), .ZN(
        Inst_bSbox_AND_M50_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M50_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M50_U1_Step1_ins_n13), .B(Fresh[80]), .ZN(
        Inst_bSbox_AND_M50_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M50_U1_Step1_ins_U1 ( .A1(Inst_bSbox_T9), .A2(
        Inst_bSbox_M38), .ZN(Inst_bSbox_AND_M50_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M50_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M50_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M50_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M50_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M50_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M50_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M50_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M50_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M50_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M50_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M50_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M50_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M50_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M50_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M50_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M50_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3407) );
  OAI221_X1 Inst_bSbox_AND_M50_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M50_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M50_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M50_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M50_U1_Step1_reg[3]), .A(
        Inst_bSbox_AND_M50_U1_in1_reg[1]), .ZN(
        Inst_bSbox_AND_M50_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M50_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M50_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M50_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M50_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M50_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M50_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M50_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M50_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M50_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M50_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M50_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M50), 
        .QN() );
  OAI21_X1 Inst_bSbox_AND_M51_U1_U4 ( .B1(new_AGEMA_signal_3397), .B2(
        Inst_bSbox_AND_M51_U1_n11), .A(Inst_bSbox_AND_M51_U1_n10), .ZN(
        Inst_bSbox_AND_M51_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M51_U1_U3 ( .B1(new_AGEMA_signal_3035), .B2(
        Fresh[85]), .C1(Inst_bSbox_AND_M51_U1_n9), .C2(Fresh[87]), .A(
        new_AGEMA_signal_3397), .ZN(Inst_bSbox_AND_M51_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M51_U1_U2 ( .A1(new_AGEMA_signal_3035), .A2(
        Fresh[86]), .B1(Fresh[84]), .B2(Inst_bSbox_AND_M51_U1_n9), .ZN(
        Inst_bSbox_AND_M51_U1_n11) );
  INV_X1 Inst_bSbox_AND_M51_U1_U1 ( .A(new_AGEMA_signal_3035), .ZN(
        Inst_bSbox_AND_M51_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M51_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3397), .CK(clk), .Q(Inst_bSbox_AND_M51_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M51_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3035), .CK(clk), .Q(Inst_bSbox_AND_M51_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M51_U1_Step1_ins_U9 ( .A(Fresh[87]), .B(
        Inst_bSbox_AND_M51_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M51_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M51_U1_Step1_ins_U8 ( .A1(Inst_bSbox_M37), .A2(
        Inst_bSbox_T17), .ZN(Inst_bSbox_AND_M51_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M51_U1_Step1_ins_U7 ( .A(Fresh[86]), .B(
        Inst_bSbox_AND_M51_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M51_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M51_U1_Step1_ins_U6 ( .A1(Inst_bSbox_T17), .A2(
        Inst_bSbox_AND_M51_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M51_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M51_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M51_U1_Step1_ins_n14), .B(Fresh[85]), .ZN(
        Inst_bSbox_AND_M51_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M51_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M51_U1_Step1_ins_n15), .A2(Inst_bSbox_T17), .ZN(
        Inst_bSbox_AND_M51_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M51_U1_Step1_ins_U3 ( .A(Inst_bSbox_M37), .ZN(
        Inst_bSbox_AND_M51_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M51_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M51_U1_Step1_ins_n13), .B(Fresh[84]), .ZN(
        Inst_bSbox_AND_M51_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M51_U1_Step1_ins_U1 ( .A1(Inst_bSbox_T17), .A2(
        Inst_bSbox_M37), .ZN(Inst_bSbox_AND_M51_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M51_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M51_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M51_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M51_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M51_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M51_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M51_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M51_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M51_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M51_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M51_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M51_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M51_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M51_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M51_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M51_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3408) );
  OAI221_X1 Inst_bSbox_AND_M51_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M51_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M51_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M51_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M51_U1_Step1_reg[3]), .A(
        Inst_bSbox_AND_M51_U1_in1_reg[1]), .ZN(
        Inst_bSbox_AND_M51_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M51_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M51_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M51_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M51_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M51_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M51_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M51_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M51_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M51_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M51_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M51_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M51), 
        .QN() );
  OAI21_X1 Inst_bSbox_AND_M52_U1_U4 ( .B1(new_AGEMA_signal_3402), .B2(
        Inst_bSbox_AND_M52_U1_n11), .A(Inst_bSbox_AND_M52_U1_n10), .ZN(
        Inst_bSbox_AND_M52_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M52_U1_U3 ( .B1(new_AGEMA_signal_3003), .B2(
        Fresh[89]), .C1(Inst_bSbox_AND_M52_U1_n9), .C2(Fresh[91]), .A(
        new_AGEMA_signal_3402), .ZN(Inst_bSbox_AND_M52_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M52_U1_U2 ( .A1(new_AGEMA_signal_3003), .A2(
        Fresh[90]), .B1(Fresh[88]), .B2(Inst_bSbox_AND_M52_U1_n9), .ZN(
        Inst_bSbox_AND_M52_U1_n11) );
  INV_X1 Inst_bSbox_AND_M52_U1_U1 ( .A(new_AGEMA_signal_3003), .ZN(
        Inst_bSbox_AND_M52_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M52_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3402), .CK(clk), .Q(Inst_bSbox_AND_M52_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M52_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3003), .CK(clk), .Q(Inst_bSbox_AND_M52_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M52_U1_Step1_ins_U9 ( .A(Fresh[91]), .B(
        Inst_bSbox_AND_M52_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M52_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M52_U1_Step1_ins_U8 ( .A1(Inst_bSbox_M42), .A2(
        Inst_bSbox_T15), .ZN(Inst_bSbox_AND_M52_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M52_U1_Step1_ins_U7 ( .A(Fresh[90]), .B(
        Inst_bSbox_AND_M52_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M52_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M52_U1_Step1_ins_U6 ( .A1(Inst_bSbox_T15), .A2(
        Inst_bSbox_AND_M52_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M52_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M52_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M52_U1_Step1_ins_n14), .B(Fresh[89]), .ZN(
        Inst_bSbox_AND_M52_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M52_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M52_U1_Step1_ins_n15), .A2(Inst_bSbox_T15), .ZN(
        Inst_bSbox_AND_M52_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M52_U1_Step1_ins_U3 ( .A(Inst_bSbox_M42), .ZN(
        Inst_bSbox_AND_M52_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M52_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M52_U1_Step1_ins_n13), .B(Fresh[88]), .ZN(
        Inst_bSbox_AND_M52_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M52_U1_Step1_ins_U1 ( .A1(Inst_bSbox_T15), .A2(
        Inst_bSbox_M42), .ZN(Inst_bSbox_AND_M52_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M52_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M52_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M52_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M52_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M52_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M52_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M52_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M52_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M52_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M52_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M52_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M52_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M52_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M52_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M52_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M52_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3416) );
  OAI221_X1 Inst_bSbox_AND_M52_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M52_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M52_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M52_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M52_U1_Step1_reg[3]), .A(
        Inst_bSbox_AND_M52_U1_in1_reg[1]), .ZN(
        Inst_bSbox_AND_M52_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M52_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M52_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M52_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M52_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M52_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M52_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M52_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M52_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M52_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M52_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M52_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M52), 
        .QN() );
  OAI21_X1 Inst_bSbox_AND_M53_U1_U4 ( .B1(new_AGEMA_signal_3413), .B2(
        Inst_bSbox_AND_M53_U1_n11), .A(Inst_bSbox_AND_M53_U1_n10), .ZN(
        Inst_bSbox_AND_M53_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M53_U1_U3 ( .B1(new_AGEMA_signal_3007), .B2(
        Fresh[93]), .C1(Inst_bSbox_AND_M53_U1_n9), .C2(Fresh[95]), .A(
        new_AGEMA_signal_3413), .ZN(Inst_bSbox_AND_M53_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M53_U1_U2 ( .A1(new_AGEMA_signal_3007), .A2(
        Fresh[94]), .B1(Fresh[92]), .B2(Inst_bSbox_AND_M53_U1_n9), .ZN(
        Inst_bSbox_AND_M53_U1_n11) );
  INV_X1 Inst_bSbox_AND_M53_U1_U1 ( .A(new_AGEMA_signal_3007), .ZN(
        Inst_bSbox_AND_M53_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M53_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3413), .CK(clk), .Q(Inst_bSbox_AND_M53_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M53_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3007), .CK(clk), .Q(Inst_bSbox_AND_M53_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M53_U1_Step1_ins_U9 ( .A(Fresh[95]), .B(
        Inst_bSbox_AND_M53_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M53_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M53_U1_Step1_ins_U8 ( .A1(Inst_bSbox_M45), .A2(
        Inst_bSbox_T27), .ZN(Inst_bSbox_AND_M53_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M53_U1_Step1_ins_U7 ( .A(Fresh[94]), .B(
        Inst_bSbox_AND_M53_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M53_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M53_U1_Step1_ins_U6 ( .A1(Inst_bSbox_T27), .A2(
        Inst_bSbox_AND_M53_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M53_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M53_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M53_U1_Step1_ins_n14), .B(Fresh[93]), .ZN(
        Inst_bSbox_AND_M53_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M53_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M53_U1_Step1_ins_n15), .A2(Inst_bSbox_T27), .ZN(
        Inst_bSbox_AND_M53_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M53_U1_Step1_ins_U3 ( .A(Inst_bSbox_M45), .ZN(
        Inst_bSbox_AND_M53_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M53_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M53_U1_Step1_ins_n13), .B(Fresh[92]), .ZN(
        Inst_bSbox_AND_M53_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M53_U1_Step1_ins_U1 ( .A1(Inst_bSbox_T27), .A2(
        Inst_bSbox_M45), .ZN(Inst_bSbox_AND_M53_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M53_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M53_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M53_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M53_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M53_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M53_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M53_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M53_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M53_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M53_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M53_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M53_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M53_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M53_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M53_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M53_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3425) );
  OAI221_X1 Inst_bSbox_AND_M53_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M53_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M53_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M53_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M53_U1_Step1_reg[3]), .A(
        Inst_bSbox_AND_M53_U1_in1_reg[1]), .ZN(
        Inst_bSbox_AND_M53_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M53_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M53_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M53_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M53_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M53_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M53_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M53_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M53_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M53_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M53_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M53_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M53), 
        .QN() );
  OAI21_X1 Inst_bSbox_AND_M54_U1_U4 ( .B1(new_AGEMA_signal_3401), .B2(
        Inst_bSbox_AND_M54_U1_n11), .A(Inst_bSbox_AND_M54_U1_n10), .ZN(
        Inst_bSbox_AND_M54_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M54_U1_U3 ( .B1(new_AGEMA_signal_3033), .B2(
        Fresh[97]), .C1(Inst_bSbox_AND_M54_U1_n9), .C2(Fresh[99]), .A(
        new_AGEMA_signal_3401), .ZN(Inst_bSbox_AND_M54_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M54_U1_U2 ( .A1(new_AGEMA_signal_3033), .A2(
        Fresh[98]), .B1(Fresh[96]), .B2(Inst_bSbox_AND_M54_U1_n9), .ZN(
        Inst_bSbox_AND_M54_U1_n11) );
  INV_X1 Inst_bSbox_AND_M54_U1_U1 ( .A(new_AGEMA_signal_3033), .ZN(
        Inst_bSbox_AND_M54_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M54_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3401), .CK(clk), .Q(Inst_bSbox_AND_M54_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M54_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3033), .CK(clk), .Q(Inst_bSbox_AND_M54_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M54_U1_Step1_ins_U9 ( .A(Fresh[99]), .B(
        Inst_bSbox_AND_M54_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M54_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M54_U1_Step1_ins_U8 ( .A1(Inst_bSbox_M41), .A2(
        Inst_bSbox_T10), .ZN(Inst_bSbox_AND_M54_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M54_U1_Step1_ins_U7 ( .A(Fresh[98]), .B(
        Inst_bSbox_AND_M54_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M54_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M54_U1_Step1_ins_U6 ( .A1(Inst_bSbox_T10), .A2(
        Inst_bSbox_AND_M54_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M54_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M54_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M54_U1_Step1_ins_n14), .B(Fresh[97]), .ZN(
        Inst_bSbox_AND_M54_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M54_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M54_U1_Step1_ins_n15), .A2(Inst_bSbox_T10), .ZN(
        Inst_bSbox_AND_M54_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M54_U1_Step1_ins_U3 ( .A(Inst_bSbox_M41), .ZN(
        Inst_bSbox_AND_M54_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M54_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M54_U1_Step1_ins_n13), .B(Fresh[96]), .ZN(
        Inst_bSbox_AND_M54_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M54_U1_Step1_ins_U1 ( .A1(Inst_bSbox_T10), .A2(
        Inst_bSbox_M41), .ZN(Inst_bSbox_AND_M54_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M54_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M54_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M54_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M54_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M54_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M54_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M54_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M54_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M54_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M54_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M54_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M54_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M54_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M54_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M54_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M54_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3417) );
  OAI221_X1 Inst_bSbox_AND_M54_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M54_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M54_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M54_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M54_U1_Step1_reg[3]), .A(
        Inst_bSbox_AND_M54_U1_in1_reg[1]), .ZN(
        Inst_bSbox_AND_M54_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M54_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M54_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M54_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M54_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M54_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M54_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M54_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M54_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M54_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M54_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M54_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M54), 
        .QN() );
  OAI21_X1 Inst_bSbox_AND_M55_U1_U4 ( .B1(new_AGEMA_signal_3404), .B2(
        Inst_bSbox_AND_M55_U1_n11), .A(Inst_bSbox_AND_M55_U1_n10), .ZN(
        Inst_bSbox_AND_M55_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M55_U1_U3 ( .B1(new_AGEMA_signal_3002), .B2(
        Fresh[101]), .C1(Inst_bSbox_AND_M55_U1_n9), .C2(Fresh[103]), .A(
        new_AGEMA_signal_3404), .ZN(Inst_bSbox_AND_M55_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M55_U1_U2 ( .A1(new_AGEMA_signal_3002), .A2(
        Fresh[102]), .B1(Fresh[100]), .B2(Inst_bSbox_AND_M55_U1_n9), .ZN(
        Inst_bSbox_AND_M55_U1_n11) );
  INV_X1 Inst_bSbox_AND_M55_U1_U1 ( .A(new_AGEMA_signal_3002), .ZN(
        Inst_bSbox_AND_M55_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M55_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3404), .CK(clk), .Q(Inst_bSbox_AND_M55_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M55_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3002), .CK(clk), .Q(Inst_bSbox_AND_M55_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M55_U1_Step1_ins_U9 ( .A(Fresh[103]), .B(
        Inst_bSbox_AND_M55_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M55_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M55_U1_Step1_ins_U8 ( .A1(Inst_bSbox_M44), .A2(
        Inst_bSbox_T13), .ZN(Inst_bSbox_AND_M55_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M55_U1_Step1_ins_U7 ( .A(Fresh[102]), .B(
        Inst_bSbox_AND_M55_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M55_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M55_U1_Step1_ins_U6 ( .A1(Inst_bSbox_T13), .A2(
        Inst_bSbox_AND_M55_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M55_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M55_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M55_U1_Step1_ins_n14), .B(Fresh[101]), .ZN(
        Inst_bSbox_AND_M55_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M55_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M55_U1_Step1_ins_n15), .A2(Inst_bSbox_T13), .ZN(
        Inst_bSbox_AND_M55_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M55_U1_Step1_ins_U3 ( .A(Inst_bSbox_M44), .ZN(
        Inst_bSbox_AND_M55_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M55_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M55_U1_Step1_ins_n13), .B(Fresh[100]), .ZN(
        Inst_bSbox_AND_M55_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M55_U1_Step1_ins_U1 ( .A1(Inst_bSbox_T13), .A2(
        Inst_bSbox_M44), .ZN(Inst_bSbox_AND_M55_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M55_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M55_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M55_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M55_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M55_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M55_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M55_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M55_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M55_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M55_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M55_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M55_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M55_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M55_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M55_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M55_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3418) );
  OAI221_X1 Inst_bSbox_AND_M55_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M55_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M55_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M55_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M55_U1_Step1_reg[3]), .A(
        Inst_bSbox_AND_M55_U1_in1_reg[1]), .ZN(
        Inst_bSbox_AND_M55_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M55_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M55_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M55_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M55_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M55_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M55_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M55_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M55_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M55_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M55_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M55_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M55), 
        .QN() );
  OAI21_X1 Inst_bSbox_AND_M56_U1_U4 ( .B1(new_AGEMA_signal_3400), .B2(
        Inst_bSbox_AND_M56_U1_n11), .A(Inst_bSbox_AND_M56_U1_n10), .ZN(
        Inst_bSbox_AND_M56_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M56_U1_U3 ( .B1(new_AGEMA_signal_3037), .B2(
        Fresh[105]), .C1(Inst_bSbox_AND_M56_U1_n9), .C2(Fresh[107]), .A(
        new_AGEMA_signal_3400), .ZN(Inst_bSbox_AND_M56_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M56_U1_U2 ( .A1(new_AGEMA_signal_3037), .A2(
        Fresh[106]), .B1(Fresh[104]), .B2(Inst_bSbox_AND_M56_U1_n9), .ZN(
        Inst_bSbox_AND_M56_U1_n11) );
  INV_X1 Inst_bSbox_AND_M56_U1_U1 ( .A(new_AGEMA_signal_3037), .ZN(
        Inst_bSbox_AND_M56_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M56_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3400), .CK(clk), .Q(Inst_bSbox_AND_M56_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M56_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3037), .CK(clk), .Q(Inst_bSbox_AND_M56_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M56_U1_Step1_ins_U9 ( .A(Fresh[107]), .B(
        Inst_bSbox_AND_M56_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M56_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M56_U1_Step1_ins_U8 ( .A1(Inst_bSbox_M40), .A2(
        Inst_bSbox_T23), .ZN(Inst_bSbox_AND_M56_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M56_U1_Step1_ins_U7 ( .A(Fresh[106]), .B(
        Inst_bSbox_AND_M56_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M56_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M56_U1_Step1_ins_U6 ( .A1(Inst_bSbox_T23), .A2(
        Inst_bSbox_AND_M56_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M56_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M56_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M56_U1_Step1_ins_n14), .B(Fresh[105]), .ZN(
        Inst_bSbox_AND_M56_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M56_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M56_U1_Step1_ins_n15), .A2(Inst_bSbox_T23), .ZN(
        Inst_bSbox_AND_M56_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M56_U1_Step1_ins_U3 ( .A(Inst_bSbox_M40), .ZN(
        Inst_bSbox_AND_M56_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M56_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M56_U1_Step1_ins_n13), .B(Fresh[104]), .ZN(
        Inst_bSbox_AND_M56_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M56_U1_Step1_ins_U1 ( .A1(Inst_bSbox_T23), .A2(
        Inst_bSbox_M40), .ZN(Inst_bSbox_AND_M56_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M56_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M56_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M56_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M56_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M56_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M56_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M56_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M56_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M56_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M56_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M56_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M56_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M56_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M56_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M56_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M56_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3409) );
  OAI221_X1 Inst_bSbox_AND_M56_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M56_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M56_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M56_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M56_U1_Step1_reg[3]), .A(
        Inst_bSbox_AND_M56_U1_in1_reg[1]), .ZN(
        Inst_bSbox_AND_M56_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M56_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M56_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M56_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M56_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M56_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M56_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M56_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M56_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M56_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M56_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M56_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M56), 
        .QN() );
  OAI21_X1 Inst_bSbox_AND_M57_U1_U4 ( .B1(new_AGEMA_signal_3399), .B2(
        Inst_bSbox_AND_M57_U1_n11), .A(Inst_bSbox_AND_M57_U1_n10), .ZN(
        Inst_bSbox_AND_M57_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M57_U1_U3 ( .B1(new_AGEMA_signal_3005), .B2(
        Fresh[109]), .C1(Inst_bSbox_AND_M57_U1_n9), .C2(Fresh[111]), .A(
        new_AGEMA_signal_3399), .ZN(Inst_bSbox_AND_M57_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M57_U1_U2 ( .A1(new_AGEMA_signal_3005), .A2(
        Fresh[110]), .B1(Fresh[108]), .B2(Inst_bSbox_AND_M57_U1_n9), .ZN(
        Inst_bSbox_AND_M57_U1_n11) );
  INV_X1 Inst_bSbox_AND_M57_U1_U1 ( .A(new_AGEMA_signal_3005), .ZN(
        Inst_bSbox_AND_M57_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M57_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3399), .CK(clk), .Q(Inst_bSbox_AND_M57_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M57_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3005), .CK(clk), .Q(Inst_bSbox_AND_M57_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M57_U1_Step1_ins_U9 ( .A(Fresh[111]), .B(
        Inst_bSbox_AND_M57_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M57_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M57_U1_Step1_ins_U8 ( .A1(Inst_bSbox_M39), .A2(
        Inst_bSbox_T19), .ZN(Inst_bSbox_AND_M57_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M57_U1_Step1_ins_U7 ( .A(Fresh[110]), .B(
        Inst_bSbox_AND_M57_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M57_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M57_U1_Step1_ins_U6 ( .A1(Inst_bSbox_T19), .A2(
        Inst_bSbox_AND_M57_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M57_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M57_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M57_U1_Step1_ins_n14), .B(Fresh[109]), .ZN(
        Inst_bSbox_AND_M57_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M57_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M57_U1_Step1_ins_n15), .A2(Inst_bSbox_T19), .ZN(
        Inst_bSbox_AND_M57_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M57_U1_Step1_ins_U3 ( .A(Inst_bSbox_M39), .ZN(
        Inst_bSbox_AND_M57_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M57_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M57_U1_Step1_ins_n13), .B(Fresh[108]), .ZN(
        Inst_bSbox_AND_M57_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M57_U1_Step1_ins_U1 ( .A1(Inst_bSbox_T19), .A2(
        Inst_bSbox_M39), .ZN(Inst_bSbox_AND_M57_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M57_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M57_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M57_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M57_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M57_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M57_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M57_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M57_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M57_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M57_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M57_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M57_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M57_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M57_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M57_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M57_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3410) );
  OAI221_X1 Inst_bSbox_AND_M57_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M57_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M57_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M57_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M57_U1_Step1_reg[3]), .A(
        Inst_bSbox_AND_M57_U1_in1_reg[1]), .ZN(
        Inst_bSbox_AND_M57_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M57_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M57_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M57_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M57_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M57_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M57_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M57_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M57_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M57_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M57_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M57_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M57), 
        .QN() );
  OAI21_X1 Inst_bSbox_AND_M58_U1_U4 ( .B1(new_AGEMA_signal_3403), .B2(
        Inst_bSbox_AND_M58_U1_n11), .A(Inst_bSbox_AND_M58_U1_n10), .ZN(
        Inst_bSbox_AND_M58_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M58_U1_U3 ( .B1(new_AGEMA_signal_2852), .B2(
        Fresh[113]), .C1(Inst_bSbox_AND_M58_U1_n9), .C2(Fresh[115]), .A(
        new_AGEMA_signal_3403), .ZN(Inst_bSbox_AND_M58_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M58_U1_U2 ( .A1(new_AGEMA_signal_2852), .A2(
        Fresh[114]), .B1(Fresh[112]), .B2(Inst_bSbox_AND_M58_U1_n9), .ZN(
        Inst_bSbox_AND_M58_U1_n11) );
  INV_X1 Inst_bSbox_AND_M58_U1_U1 ( .A(new_AGEMA_signal_2852), .ZN(
        Inst_bSbox_AND_M58_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M58_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3403), .CK(clk), .Q(Inst_bSbox_AND_M58_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M58_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_2852), .CK(clk), .Q(Inst_bSbox_AND_M58_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M58_U1_Step1_ins_U9 ( .A(Fresh[115]), .B(
        Inst_bSbox_AND_M58_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M58_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M58_U1_Step1_ins_U8 ( .A1(Inst_bSbox_M43), .A2(
        Inst_bSbox_T3), .ZN(Inst_bSbox_AND_M58_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M58_U1_Step1_ins_U7 ( .A(Fresh[114]), .B(
        Inst_bSbox_AND_M58_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M58_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M58_U1_Step1_ins_U6 ( .A1(Inst_bSbox_T3), .A2(
        Inst_bSbox_AND_M58_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M58_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M58_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M58_U1_Step1_ins_n14), .B(Fresh[113]), .ZN(
        Inst_bSbox_AND_M58_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M58_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M58_U1_Step1_ins_n15), .A2(Inst_bSbox_T3), .ZN(
        Inst_bSbox_AND_M58_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M58_U1_Step1_ins_U3 ( .A(Inst_bSbox_M43), .ZN(
        Inst_bSbox_AND_M58_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M58_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M58_U1_Step1_ins_n13), .B(Fresh[112]), .ZN(
        Inst_bSbox_AND_M58_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M58_U1_Step1_ins_U1 ( .A1(Inst_bSbox_T3), .A2(
        Inst_bSbox_M43), .ZN(Inst_bSbox_AND_M58_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M58_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M58_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M58_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M58_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M58_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M58_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M58_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M58_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M58_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M58_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M58_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M58_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M58_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M58_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M58_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M58_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3419) );
  OAI221_X1 Inst_bSbox_AND_M58_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M58_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M58_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M58_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M58_U1_Step1_reg[3]), .A(
        Inst_bSbox_AND_M58_U1_in1_reg[1]), .ZN(
        Inst_bSbox_AND_M58_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M58_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M58_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M58_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M58_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M58_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M58_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M58_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M58_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M58_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M58_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M58_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M58), 
        .QN() );
  OAI21_X1 Inst_bSbox_AND_M59_U1_U4 ( .B1(new_AGEMA_signal_3398), .B2(
        Inst_bSbox_AND_M59_U1_n11), .A(Inst_bSbox_AND_M59_U1_n10), .ZN(
        Inst_bSbox_AND_M59_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M59_U1_U3 ( .B1(new_AGEMA_signal_3006), .B2(
        Fresh[117]), .C1(Inst_bSbox_AND_M59_U1_n9), .C2(Fresh[119]), .A(
        new_AGEMA_signal_3398), .ZN(Inst_bSbox_AND_M59_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M59_U1_U2 ( .A1(new_AGEMA_signal_3006), .A2(
        Fresh[118]), .B1(Fresh[116]), .B2(Inst_bSbox_AND_M59_U1_n9), .ZN(
        Inst_bSbox_AND_M59_U1_n11) );
  INV_X1 Inst_bSbox_AND_M59_U1_U1 ( .A(new_AGEMA_signal_3006), .ZN(
        Inst_bSbox_AND_M59_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M59_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3398), .CK(clk), .Q(Inst_bSbox_AND_M59_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M59_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3006), .CK(clk), .Q(Inst_bSbox_AND_M59_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M59_U1_Step1_ins_U9 ( .A(Fresh[119]), .B(
        Inst_bSbox_AND_M59_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M59_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M59_U1_Step1_ins_U8 ( .A1(Inst_bSbox_M38), .A2(
        Inst_bSbox_T22), .ZN(Inst_bSbox_AND_M59_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M59_U1_Step1_ins_U7 ( .A(Fresh[118]), .B(
        Inst_bSbox_AND_M59_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M59_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M59_U1_Step1_ins_U6 ( .A1(Inst_bSbox_T22), .A2(
        Inst_bSbox_AND_M59_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M59_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M59_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M59_U1_Step1_ins_n14), .B(Fresh[117]), .ZN(
        Inst_bSbox_AND_M59_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M59_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M59_U1_Step1_ins_n15), .A2(Inst_bSbox_T22), .ZN(
        Inst_bSbox_AND_M59_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M59_U1_Step1_ins_U3 ( .A(Inst_bSbox_M38), .ZN(
        Inst_bSbox_AND_M59_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M59_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M59_U1_Step1_ins_n13), .B(Fresh[116]), .ZN(
        Inst_bSbox_AND_M59_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M59_U1_Step1_ins_U1 ( .A1(Inst_bSbox_T22), .A2(
        Inst_bSbox_M38), .ZN(Inst_bSbox_AND_M59_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M59_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M59_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M59_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M59_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M59_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M59_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M59_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M59_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M59_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M59_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M59_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M59_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M59_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M59_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M59_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M59_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3411) );
  OAI221_X1 Inst_bSbox_AND_M59_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M59_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M59_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M59_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M59_U1_Step1_reg[3]), .A(
        Inst_bSbox_AND_M59_U1_in1_reg[1]), .ZN(
        Inst_bSbox_AND_M59_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M59_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M59_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M59_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M59_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M59_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M59_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M59_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M59_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M59_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M59_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M59_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M59), 
        .QN() );
  OAI21_X1 Inst_bSbox_AND_M60_U1_U4 ( .B1(new_AGEMA_signal_3397), .B2(
        Inst_bSbox_AND_M60_U1_n11), .A(Inst_bSbox_AND_M60_U1_n10), .ZN(
        Inst_bSbox_AND_M60_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M60_U1_U3 ( .B1(new_AGEMA_signal_3036), .B2(
        Fresh[121]), .C1(Inst_bSbox_AND_M60_U1_n9), .C2(Fresh[123]), .A(
        new_AGEMA_signal_3397), .ZN(Inst_bSbox_AND_M60_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M60_U1_U2 ( .A1(new_AGEMA_signal_3036), .A2(
        Fresh[122]), .B1(Fresh[120]), .B2(Inst_bSbox_AND_M60_U1_n9), .ZN(
        Inst_bSbox_AND_M60_U1_n11) );
  INV_X1 Inst_bSbox_AND_M60_U1_U1 ( .A(new_AGEMA_signal_3036), .ZN(
        Inst_bSbox_AND_M60_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M60_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3397), .CK(clk), .Q(Inst_bSbox_AND_M60_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M60_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_3036), .CK(clk), .Q(Inst_bSbox_AND_M60_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M60_U1_Step1_ins_U9 ( .A(Fresh[123]), .B(
        Inst_bSbox_AND_M60_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M60_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M60_U1_Step1_ins_U8 ( .A1(Inst_bSbox_M37), .A2(
        Inst_bSbox_T20), .ZN(Inst_bSbox_AND_M60_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M60_U1_Step1_ins_U7 ( .A(Fresh[122]), .B(
        Inst_bSbox_AND_M60_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M60_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M60_U1_Step1_ins_U6 ( .A1(Inst_bSbox_T20), .A2(
        Inst_bSbox_AND_M60_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M60_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M60_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M60_U1_Step1_ins_n14), .B(Fresh[121]), .ZN(
        Inst_bSbox_AND_M60_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M60_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M60_U1_Step1_ins_n15), .A2(Inst_bSbox_T20), .ZN(
        Inst_bSbox_AND_M60_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M60_U1_Step1_ins_U3 ( .A(Inst_bSbox_M37), .ZN(
        Inst_bSbox_AND_M60_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M60_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M60_U1_Step1_ins_n13), .B(Fresh[120]), .ZN(
        Inst_bSbox_AND_M60_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M60_U1_Step1_ins_U1 ( .A1(Inst_bSbox_T20), .A2(
        Inst_bSbox_M37), .ZN(Inst_bSbox_AND_M60_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M60_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M60_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M60_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M60_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M60_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M60_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M60_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M60_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M60_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M60_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M60_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M60_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M60_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M60_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M60_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M60_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3412) );
  OAI221_X1 Inst_bSbox_AND_M60_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M60_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M60_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M60_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M60_U1_Step1_reg[3]), .A(
        Inst_bSbox_AND_M60_U1_in1_reg[1]), .ZN(
        Inst_bSbox_AND_M60_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M60_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M60_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M60_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M60_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M60_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M60_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M60_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M60_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M60_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M60_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M60_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M60), 
        .QN() );
  OAI21_X1 Inst_bSbox_AND_M61_U1_U4 ( .B1(new_AGEMA_signal_3402), .B2(
        Inst_bSbox_AND_M61_U1_n11), .A(Inst_bSbox_AND_M61_U1_n10), .ZN(
        Inst_bSbox_AND_M61_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M61_U1_U3 ( .B1(new_AGEMA_signal_2850), .B2(
        Fresh[125]), .C1(Inst_bSbox_AND_M61_U1_n9), .C2(Fresh[127]), .A(
        new_AGEMA_signal_3402), .ZN(Inst_bSbox_AND_M61_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M61_U1_U2 ( .A1(new_AGEMA_signal_2850), .A2(
        Fresh[126]), .B1(Fresh[124]), .B2(Inst_bSbox_AND_M61_U1_n9), .ZN(
        Inst_bSbox_AND_M61_U1_n11) );
  INV_X1 Inst_bSbox_AND_M61_U1_U1 ( .A(new_AGEMA_signal_2850), .ZN(
        Inst_bSbox_AND_M61_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M61_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3402), .CK(clk), .Q(Inst_bSbox_AND_M61_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M61_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_2850), .CK(clk), .Q(Inst_bSbox_AND_M61_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M61_U1_Step1_ins_U9 ( .A(Fresh[127]), .B(
        Inst_bSbox_AND_M61_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M61_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M61_U1_Step1_ins_U8 ( .A1(Inst_bSbox_M42), .A2(
        Inst_bSbox_T1), .ZN(Inst_bSbox_AND_M61_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M61_U1_Step1_ins_U7 ( .A(Fresh[126]), .B(
        Inst_bSbox_AND_M61_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M61_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M61_U1_Step1_ins_U6 ( .A1(Inst_bSbox_T1), .A2(
        Inst_bSbox_AND_M61_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M61_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M61_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M61_U1_Step1_ins_n14), .B(Fresh[125]), .ZN(
        Inst_bSbox_AND_M61_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M61_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M61_U1_Step1_ins_n15), .A2(Inst_bSbox_T1), .ZN(
        Inst_bSbox_AND_M61_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M61_U1_Step1_ins_U3 ( .A(Inst_bSbox_M42), .ZN(
        Inst_bSbox_AND_M61_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M61_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M61_U1_Step1_ins_n13), .B(Fresh[124]), .ZN(
        Inst_bSbox_AND_M61_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M61_U1_Step1_ins_U1 ( .A1(Inst_bSbox_T1), .A2(
        Inst_bSbox_M42), .ZN(Inst_bSbox_AND_M61_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M61_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M61_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M61_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M61_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M61_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M61_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M61_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M61_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M61_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M61_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M61_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M61_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M61_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M61_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M61_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M61_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3420) );
  OAI221_X1 Inst_bSbox_AND_M61_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M61_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M61_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M61_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M61_U1_Step1_reg[3]), .A(
        Inst_bSbox_AND_M61_U1_in1_reg[1]), .ZN(
        Inst_bSbox_AND_M61_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M61_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M61_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M61_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M61_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M61_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M61_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M61_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M61_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M61_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M61_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M61_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M61), 
        .QN() );
  OAI21_X1 Inst_bSbox_AND_M62_U1_U4 ( .B1(new_AGEMA_signal_3413), .B2(
        Inst_bSbox_AND_M62_U1_n11), .A(Inst_bSbox_AND_M62_U1_n10), .ZN(
        Inst_bSbox_AND_M62_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M62_U1_U3 ( .B1(new_AGEMA_signal_2853), .B2(
        Fresh[129]), .C1(Inst_bSbox_AND_M62_U1_n9), .C2(Fresh[131]), .A(
        new_AGEMA_signal_3413), .ZN(Inst_bSbox_AND_M62_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M62_U1_U2 ( .A1(new_AGEMA_signal_2853), .A2(
        Fresh[130]), .B1(Fresh[128]), .B2(Inst_bSbox_AND_M62_U1_n9), .ZN(
        Inst_bSbox_AND_M62_U1_n11) );
  INV_X1 Inst_bSbox_AND_M62_U1_U1 ( .A(new_AGEMA_signal_2853), .ZN(
        Inst_bSbox_AND_M62_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M62_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3413), .CK(clk), .Q(Inst_bSbox_AND_M62_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M62_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_2853), .CK(clk), .Q(Inst_bSbox_AND_M62_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M62_U1_Step1_ins_U9 ( .A(Fresh[131]), .B(
        Inst_bSbox_AND_M62_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M62_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M62_U1_Step1_ins_U8 ( .A1(Inst_bSbox_M45), .A2(
        Inst_bSbox_T4), .ZN(Inst_bSbox_AND_M62_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M62_U1_Step1_ins_U7 ( .A(Fresh[130]), .B(
        Inst_bSbox_AND_M62_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M62_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M62_U1_Step1_ins_U6 ( .A1(Inst_bSbox_T4), .A2(
        Inst_bSbox_AND_M62_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M62_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M62_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M62_U1_Step1_ins_n14), .B(Fresh[129]), .ZN(
        Inst_bSbox_AND_M62_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M62_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M62_U1_Step1_ins_n15), .A2(Inst_bSbox_T4), .ZN(
        Inst_bSbox_AND_M62_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M62_U1_Step1_ins_U3 ( .A(Inst_bSbox_M45), .ZN(
        Inst_bSbox_AND_M62_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M62_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M62_U1_Step1_ins_n13), .B(Fresh[128]), .ZN(
        Inst_bSbox_AND_M62_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M62_U1_Step1_ins_U1 ( .A1(Inst_bSbox_T4), .A2(
        Inst_bSbox_M45), .ZN(Inst_bSbox_AND_M62_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M62_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M62_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M62_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M62_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M62_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M62_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M62_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M62_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M62_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M62_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M62_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M62_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M62_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M62_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M62_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M62_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3426) );
  OAI221_X1 Inst_bSbox_AND_M62_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M62_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M62_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M62_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M62_U1_Step1_reg[3]), .A(
        Inst_bSbox_AND_M62_U1_in1_reg[1]), .ZN(
        Inst_bSbox_AND_M62_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M62_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M62_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M62_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M62_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M62_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M62_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M62_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M62_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M62_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M62_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M62_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M62), 
        .QN() );
  OAI21_X1 Inst_bSbox_AND_M63_U1_U4 ( .B1(new_AGEMA_signal_3401), .B2(
        Inst_bSbox_AND_M63_U1_n11), .A(Inst_bSbox_AND_M63_U1_n10), .ZN(
        Inst_bSbox_AND_M63_U1_out0_mid_0_) );
  OAI221_X1 Inst_bSbox_AND_M63_U1_U3 ( .B1(new_AGEMA_signal_2851), .B2(
        Fresh[133]), .C1(Inst_bSbox_AND_M63_U1_n9), .C2(Fresh[135]), .A(
        new_AGEMA_signal_3401), .ZN(Inst_bSbox_AND_M63_U1_n10) );
  AOI22_X1 Inst_bSbox_AND_M63_U1_U2 ( .A1(new_AGEMA_signal_2851), .A2(
        Fresh[134]), .B1(Fresh[132]), .B2(Inst_bSbox_AND_M63_U1_n9), .ZN(
        Inst_bSbox_AND_M63_U1_n11) );
  INV_X1 Inst_bSbox_AND_M63_U1_U1 ( .A(new_AGEMA_signal_2851), .ZN(
        Inst_bSbox_AND_M63_U1_n9) );
  DFF_X1 Inst_bSbox_AND_M63_U1_reg_ins1_0_s_current_state_reg ( .D(
        new_AGEMA_signal_3401), .CK(clk), .Q(Inst_bSbox_AND_M63_U1_in1_reg[0]), 
        .QN() );
  DFF_X1 Inst_bSbox_AND_M63_U1_reg_ins1_1_s_current_state_reg ( .D(
        new_AGEMA_signal_2851), .CK(clk), .Q(Inst_bSbox_AND_M63_U1_in1_reg[1]), 
        .QN() );
  XOR2_X1 Inst_bSbox_AND_M63_U1_Step1_ins_U9 ( .A(Fresh[135]), .B(
        Inst_bSbox_AND_M63_U1_Step1_ins_n17), .Z(
        Inst_bSbox_AND_M63_U1_Step1_ins_Step1[3]) );
  NOR2_X1 Inst_bSbox_AND_M63_U1_Step1_ins_U8 ( .A1(Inst_bSbox_M41), .A2(
        Inst_bSbox_T2), .ZN(Inst_bSbox_AND_M63_U1_Step1_ins_n17) );
  XOR2_X1 Inst_bSbox_AND_M63_U1_Step1_ins_U7 ( .A(Fresh[134]), .B(
        Inst_bSbox_AND_M63_U1_Step1_ins_n16), .Z(
        Inst_bSbox_AND_M63_U1_Step1_ins_Step1[2]) );
  NOR2_X1 Inst_bSbox_AND_M63_U1_Step1_ins_U6 ( .A1(Inst_bSbox_T2), .A2(
        Inst_bSbox_AND_M63_U1_Step1_ins_n15), .ZN(
        Inst_bSbox_AND_M63_U1_Step1_ins_n16) );
  XNOR2_X1 Inst_bSbox_AND_M63_U1_Step1_ins_U5 ( .A(
        Inst_bSbox_AND_M63_U1_Step1_ins_n14), .B(Fresh[133]), .ZN(
        Inst_bSbox_AND_M63_U1_Step1_ins_Step1[1]) );
  NAND2_X1 Inst_bSbox_AND_M63_U1_Step1_ins_U4 ( .A1(
        Inst_bSbox_AND_M63_U1_Step1_ins_n15), .A2(Inst_bSbox_T2), .ZN(
        Inst_bSbox_AND_M63_U1_Step1_ins_n14) );
  INV_X1 Inst_bSbox_AND_M63_U1_Step1_ins_U3 ( .A(Inst_bSbox_M41), .ZN(
        Inst_bSbox_AND_M63_U1_Step1_ins_n15) );
  XNOR2_X1 Inst_bSbox_AND_M63_U1_Step1_ins_U2 ( .A(
        Inst_bSbox_AND_M63_U1_Step1_ins_n13), .B(Fresh[132]), .ZN(
        Inst_bSbox_AND_M63_U1_Step1_ins_Step1[0]) );
  NAND2_X1 Inst_bSbox_AND_M63_U1_Step1_ins_U1 ( .A1(Inst_bSbox_T2), .A2(
        Inst_bSbox_M41), .ZN(Inst_bSbox_AND_M63_U1_Step1_ins_n13) );
  DFF_X1 Inst_bSbox_AND_M63_U1_Step1_ins_reg_ins_0_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M63_U1_Step1_ins_Step1[0]), .CK(clk), .Q(
        Inst_bSbox_AND_M63_U1_Step1_reg[0]), .QN() );
  DFF_X1 Inst_bSbox_AND_M63_U1_Step1_ins_reg_ins_0_1_s_current_state_reg ( .D(
        Inst_bSbox_AND_M63_U1_Step1_ins_Step1[1]), .CK(clk), .Q(
        Inst_bSbox_AND_M63_U1_Step1_reg[1]), .QN() );
  DFF_X1 Inst_bSbox_AND_M63_U1_Step1_ins_reg_ins_0_2_s_current_state_reg ( .D(
        Inst_bSbox_AND_M63_U1_Step1_ins_Step1[2]), .CK(clk), .Q(
        Inst_bSbox_AND_M63_U1_Step1_reg[2]), .QN() );
  DFF_X1 Inst_bSbox_AND_M63_U1_Step1_ins_reg_ins_0_3_s_current_state_reg ( .D(
        Inst_bSbox_AND_M63_U1_Step1_ins_Step1[3]), .CK(clk), .Q(
        Inst_bSbox_AND_M63_U1_Step1_reg[3]), .QN() );
  OAI21_X1 Inst_bSbox_AND_M63_U1_Step2_inst_U4 ( .B1(
        Inst_bSbox_AND_M63_U1_in1_reg[1]), .B2(
        Inst_bSbox_AND_M63_U1_Step2_inst_n11), .A(
        Inst_bSbox_AND_M63_U1_Step2_inst_n10), .ZN(new_AGEMA_signal_3421) );
  OAI221_X1 Inst_bSbox_AND_M63_U1_Step2_inst_U3 ( .B1(
        Inst_bSbox_AND_M63_U1_in1_reg[0]), .B2(
        Inst_bSbox_AND_M63_U1_Step1_reg[2]), .C1(
        Inst_bSbox_AND_M63_U1_Step2_inst_n9), .C2(
        Inst_bSbox_AND_M63_U1_Step1_reg[3]), .A(
        Inst_bSbox_AND_M63_U1_in1_reg[1]), .ZN(
        Inst_bSbox_AND_M63_U1_Step2_inst_n10) );
  AOI22_X1 Inst_bSbox_AND_M63_U1_Step2_inst_U2 ( .A1(
        Inst_bSbox_AND_M63_U1_in1_reg[0]), .A2(
        Inst_bSbox_AND_M63_U1_Step1_reg[1]), .B1(
        Inst_bSbox_AND_M63_U1_Step1_reg[0]), .B2(
        Inst_bSbox_AND_M63_U1_Step2_inst_n9), .ZN(
        Inst_bSbox_AND_M63_U1_Step2_inst_n11) );
  INV_X1 Inst_bSbox_AND_M63_U1_Step2_inst_U1 ( .A(
        Inst_bSbox_AND_M63_U1_in1_reg[0]), .ZN(
        Inst_bSbox_AND_M63_U1_Step2_inst_n9) );
  DFF_X1 Inst_bSbox_AND_M63_U1_reg_out0_ins2_0_s_current_state_reg ( .D(
        Inst_bSbox_AND_M63_U1_out0_mid_0_), .CK(clk), .Q(Inst_bSbox_M63), 
        .QN() );
  XOR2_X1 Inst_bSbox_XOR_L0_U1_Ins_0_U1 ( .A(Inst_bSbox_M61), .B(
        Inst_bSbox_M62), .Z(Inst_bSbox_L0) );
  XOR2_X1 Inst_bSbox_XOR_L0_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3420), .B(
        new_AGEMA_signal_3426), .Z(new_AGEMA_signal_3435) );
  XOR2_X1 Inst_bSbox_XOR_L1_U1_Ins_0_U1 ( .A(Inst_bSbox_M50), .B(
        Inst_bSbox_M56), .Z(Inst_bSbox_L1) );
  XOR2_X1 Inst_bSbox_XOR_L1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3407), .B(
        new_AGEMA_signal_3409), .Z(new_AGEMA_signal_3422) );
  XOR2_X1 Inst_bSbox_XOR_L2_U1_Ins_0_U1 ( .A(Inst_bSbox_M46), .B(
        Inst_bSbox_M48), .Z(Inst_bSbox_L2) );
  XOR2_X1 Inst_bSbox_XOR_L2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3414), .B(
        new_AGEMA_signal_3406), .Z(new_AGEMA_signal_3427) );
  XOR2_X1 Inst_bSbox_XOR_L3_U1_Ins_0_U1 ( .A(Inst_bSbox_M47), .B(
        Inst_bSbox_M55), .Z(Inst_bSbox_L3) );
  XOR2_X1 Inst_bSbox_XOR_L3_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3405), .B(
        new_AGEMA_signal_3418), .Z(new_AGEMA_signal_3428) );
  XOR2_X1 Inst_bSbox_XOR_L4_U1_Ins_0_U1 ( .A(Inst_bSbox_M54), .B(
        Inst_bSbox_M58), .Z(Inst_bSbox_L4) );
  XOR2_X1 Inst_bSbox_XOR_L4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3417), .B(
        new_AGEMA_signal_3419), .Z(new_AGEMA_signal_3429) );
  XOR2_X1 Inst_bSbox_XOR_L5_U1_Ins_0_U1 ( .A(Inst_bSbox_M49), .B(
        Inst_bSbox_M61), .Z(Inst_bSbox_L5) );
  XOR2_X1 Inst_bSbox_XOR_L5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3415), .B(
        new_AGEMA_signal_3420), .Z(new_AGEMA_signal_3430) );
  XOR2_X1 Inst_bSbox_XOR_L6_U1_Ins_0_U1 ( .A(Inst_bSbox_M62), .B(Inst_bSbox_L5), .Z(Inst_bSbox_L6) );
  XOR2_X1 Inst_bSbox_XOR_L6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3426), .B(
        new_AGEMA_signal_3430), .Z(new_AGEMA_signal_3436) );
  XOR2_X1 Inst_bSbox_XOR_L7_U1_Ins_0_U1 ( .A(Inst_bSbox_M46), .B(Inst_bSbox_L3), .Z(Inst_bSbox_L7) );
  XOR2_X1 Inst_bSbox_XOR_L7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3414), .B(
        new_AGEMA_signal_3428), .Z(new_AGEMA_signal_3437) );
  XOR2_X1 Inst_bSbox_XOR_L8_U1_Ins_0_U1 ( .A(Inst_bSbox_M51), .B(
        Inst_bSbox_M59), .Z(Inst_bSbox_L8) );
  XOR2_X1 Inst_bSbox_XOR_L8_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3408), .B(
        new_AGEMA_signal_3411), .Z(new_AGEMA_signal_3423) );
  XOR2_X1 Inst_bSbox_XOR_L9_U1_Ins_0_U1 ( .A(Inst_bSbox_M52), .B(
        Inst_bSbox_M53), .Z(Inst_bSbox_L9) );
  XOR2_X1 Inst_bSbox_XOR_L9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3416), .B(
        new_AGEMA_signal_3425), .Z(new_AGEMA_signal_3438) );
  XOR2_X1 Inst_bSbox_XOR_L10_U1_Ins_0_U1 ( .A(Inst_bSbox_M53), .B(
        Inst_bSbox_L4), .Z(Inst_bSbox_L10) );
  XOR2_X1 Inst_bSbox_XOR_L10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3425), .B(
        new_AGEMA_signal_3429), .Z(new_AGEMA_signal_3439) );
  XOR2_X1 Inst_bSbox_XOR_L11_U1_Ins_0_U1 ( .A(Inst_bSbox_M60), .B(
        Inst_bSbox_L2), .Z(Inst_bSbox_L11) );
  XOR2_X1 Inst_bSbox_XOR_L11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3412), .B(
        new_AGEMA_signal_3427), .Z(new_AGEMA_signal_3440) );
  XOR2_X1 Inst_bSbox_XOR_L12_U1_Ins_0_U1 ( .A(Inst_bSbox_M48), .B(
        Inst_bSbox_M51), .Z(Inst_bSbox_L12) );
  XOR2_X1 Inst_bSbox_XOR_L12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3406), .B(
        new_AGEMA_signal_3408), .Z(new_AGEMA_signal_3424) );
  XOR2_X1 Inst_bSbox_XOR_L13_U1_Ins_0_U1 ( .A(Inst_bSbox_M50), .B(
        Inst_bSbox_L0), .Z(Inst_bSbox_L13) );
  XOR2_X1 Inst_bSbox_XOR_L13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3407), .B(
        new_AGEMA_signal_3435), .Z(new_AGEMA_signal_3444) );
  XOR2_X1 Inst_bSbox_XOR_L14_U1_Ins_0_U1 ( .A(Inst_bSbox_M52), .B(
        Inst_bSbox_M61), .Z(Inst_bSbox_L14) );
  XOR2_X1 Inst_bSbox_XOR_L14_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3416), .B(
        new_AGEMA_signal_3420), .Z(new_AGEMA_signal_3431) );
  XOR2_X1 Inst_bSbox_XOR_L15_U1_Ins_0_U1 ( .A(Inst_bSbox_M55), .B(
        Inst_bSbox_L1), .Z(Inst_bSbox_L15) );
  XOR2_X1 Inst_bSbox_XOR_L15_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3418), .B(
        new_AGEMA_signal_3422), .Z(new_AGEMA_signal_3432) );
  XOR2_X1 Inst_bSbox_XOR_L16_U1_Ins_0_U1 ( .A(Inst_bSbox_M56), .B(
        Inst_bSbox_L0), .Z(Inst_bSbox_L16) );
  XOR2_X1 Inst_bSbox_XOR_L16_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3409), .B(
        new_AGEMA_signal_3435), .Z(new_AGEMA_signal_3445) );
  XOR2_X1 Inst_bSbox_XOR_L17_U1_Ins_0_U1 ( .A(Inst_bSbox_M57), .B(
        Inst_bSbox_L1), .Z(Inst_bSbox_L17) );
  XOR2_X1 Inst_bSbox_XOR_L17_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3410), .B(
        new_AGEMA_signal_3422), .Z(new_AGEMA_signal_3433) );
  XOR2_X1 Inst_bSbox_XOR_L18_U1_Ins_0_U1 ( .A(Inst_bSbox_M58), .B(
        Inst_bSbox_L8), .Z(Inst_bSbox_L18) );
  XOR2_X1 Inst_bSbox_XOR_L18_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3419), .B(
        new_AGEMA_signal_3423), .Z(new_AGEMA_signal_3434) );
  XOR2_X1 Inst_bSbox_XOR_L19_U1_Ins_0_U1 ( .A(Inst_bSbox_M63), .B(
        Inst_bSbox_L4), .Z(Inst_bSbox_L19) );
  XOR2_X1 Inst_bSbox_XOR_L19_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3421), .B(
        new_AGEMA_signal_3429), .Z(new_AGEMA_signal_3441) );
  XOR2_X1 Inst_bSbox_XOR_L20_U1_Ins_0_U1 ( .A(Inst_bSbox_L0), .B(Inst_bSbox_L1), .Z(Inst_bSbox_L20) );
  XOR2_X1 Inst_bSbox_XOR_L20_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3435), .B(
        new_AGEMA_signal_3422), .Z(new_AGEMA_signal_3446) );
  XOR2_X1 Inst_bSbox_XOR_L21_U1_Ins_0_U1 ( .A(Inst_bSbox_L1), .B(Inst_bSbox_L7), .Z(Inst_bSbox_L21) );
  XOR2_X1 Inst_bSbox_XOR_L21_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3422), .B(
        new_AGEMA_signal_3437), .Z(new_AGEMA_signal_3447) );
  XOR2_X1 Inst_bSbox_XOR_L22_U1_Ins_0_U1 ( .A(Inst_bSbox_L3), .B(
        Inst_bSbox_L12), .Z(Inst_bSbox_L22) );
  XOR2_X1 Inst_bSbox_XOR_L22_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3428), .B(
        new_AGEMA_signal_3424), .Z(new_AGEMA_signal_3442) );
  XOR2_X1 Inst_bSbox_XOR_L23_U1_Ins_0_U1 ( .A(Inst_bSbox_L18), .B(
        Inst_bSbox_L2), .Z(Inst_bSbox_L23) );
  XOR2_X1 Inst_bSbox_XOR_L23_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3434), .B(
        new_AGEMA_signal_3427), .Z(new_AGEMA_signal_3443) );
  XOR2_X1 Inst_bSbox_XOR_L24_U1_Ins_0_U1 ( .A(Inst_bSbox_L15), .B(
        Inst_bSbox_L9), .Z(Inst_bSbox_L24) );
  XOR2_X1 Inst_bSbox_XOR_L24_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3432), .B(
        new_AGEMA_signal_3438), .Z(new_AGEMA_signal_3448) );
  XOR2_X1 Inst_bSbox_XOR_L25_U1_Ins_0_U1 ( .A(Inst_bSbox_L6), .B(
        Inst_bSbox_L10), .Z(Inst_bSbox_L25) );
  XOR2_X1 Inst_bSbox_XOR_L25_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3436), .B(
        new_AGEMA_signal_3439), .Z(new_AGEMA_signal_3449) );
  XOR2_X1 Inst_bSbox_XOR_L26_U1_Ins_0_U1 ( .A(Inst_bSbox_L7), .B(Inst_bSbox_L9), .Z(Inst_bSbox_L26) );
  XOR2_X1 Inst_bSbox_XOR_L26_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3437), .B(
        new_AGEMA_signal_3438), .Z(new_AGEMA_signal_3450) );
  XOR2_X1 Inst_bSbox_XOR_L27_U1_Ins_0_U1 ( .A(Inst_bSbox_L8), .B(
        Inst_bSbox_L10), .Z(Inst_bSbox_L27) );
  XOR2_X1 Inst_bSbox_XOR_L27_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3423), .B(
        new_AGEMA_signal_3439), .Z(new_AGEMA_signal_3451) );
  XOR2_X1 Inst_bSbox_XOR_L28_U1_Ins_0_U1 ( .A(Inst_bSbox_L11), .B(
        Inst_bSbox_L14), .Z(Inst_bSbox_L28) );
  XOR2_X1 Inst_bSbox_XOR_L28_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3440), .B(
        new_AGEMA_signal_3431), .Z(new_AGEMA_signal_3452) );
  XOR2_X1 Inst_bSbox_XOR_L29_U1_Ins_0_U1 ( .A(Inst_bSbox_L11), .B(
        Inst_bSbox_L17), .Z(Inst_bSbox_L29) );
  XOR2_X1 Inst_bSbox_XOR_L29_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3440), .B(
        new_AGEMA_signal_3433), .Z(new_AGEMA_signal_3453) );
  XOR2_X1 Inst_bSbox_XOR_S0_U1_Ins_0_U1 ( .A(Inst_bSbox_L6), .B(Inst_bSbox_L24), .Z(SboxOut[7]) );
  XOR2_X1 Inst_bSbox_XOR_S0_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3436), .B(
        new_AGEMA_signal_3448), .Z(new_AGEMA_signal_3457) );
  XNOR2_X1 Inst_bSbox_XOR_S1_U1_Ins0_U1 ( .A(Inst_bSbox_L16), .B(
        Inst_bSbox_L26), .ZN(SboxOut[6]) );
  XOR2_X1 Inst_bSbox_XOR_S1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3445), .B(
        new_AGEMA_signal_3450), .Z(new_AGEMA_signal_3458) );
  XNOR2_X1 Inst_bSbox_XOR_S2_U1_Ins0_U1 ( .A(Inst_bSbox_L19), .B(
        Inst_bSbox_L28), .ZN(SboxOut[5]) );
  XOR2_X1 Inst_bSbox_XOR_S2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3441), .B(
        new_AGEMA_signal_3452), .Z(new_AGEMA_signal_3459) );
  XOR2_X1 Inst_bSbox_XOR_S3_U1_Ins_0_U1 ( .A(Inst_bSbox_L6), .B(Inst_bSbox_L21), .Z(SboxOut[4]) );
  XOR2_X1 Inst_bSbox_XOR_S3_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3436), .B(
        new_AGEMA_signal_3447), .Z(new_AGEMA_signal_3460) );
  XOR2_X1 Inst_bSbox_XOR_S4_U1_Ins_0_U1 ( .A(Inst_bSbox_L20), .B(
        Inst_bSbox_L22), .Z(SboxOut[3]) );
  XOR2_X1 Inst_bSbox_XOR_S4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3446), .B(
        new_AGEMA_signal_3442), .Z(new_AGEMA_signal_3461) );
  XOR2_X1 Inst_bSbox_XOR_S5_U1_Ins_0_U1 ( .A(Inst_bSbox_L25), .B(
        Inst_bSbox_L29), .Z(SboxOut[2]) );
  XOR2_X1 Inst_bSbox_XOR_S5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3449), .B(
        new_AGEMA_signal_3453), .Z(new_AGEMA_signal_3462) );
  XNOR2_X1 Inst_bSbox_XOR_S6_U1_Ins0_U1 ( .A(Inst_bSbox_L13), .B(
        Inst_bSbox_L27), .ZN(SboxOut[1]) );
  XOR2_X1 Inst_bSbox_XOR_S6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3444), .B(
        new_AGEMA_signal_3451), .Z(new_AGEMA_signal_3463) );
  XNOR2_X1 Inst_bSbox_XOR_S7_U1_Ins0_U1 ( .A(Inst_bSbox_L6), .B(Inst_bSbox_L23), .ZN(SboxOut[0]) );
  XOR2_X1 Inst_bSbox_XOR_S7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3436), .B(
        new_AGEMA_signal_3443), .Z(new_AGEMA_signal_3454) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S00reg_gff_1_SFF_0_QD), .CK(clk_gated), .Q(
        ciphertext_s0[120]), .QN() );
  DFF_X1 stateArray_S00reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3126), .CK(clk_gated), .Q(ciphertext_s1[120]), 
        .QN() );
  DFF_X1 stateArray_S00reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S00reg_gff_1_SFF_1_QD), .CK(clk_gated), .Q(
        ciphertext_s0[121]), .QN() );
  DFF_X1 stateArray_S00reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3127), .CK(clk_gated), .Q(ciphertext_s1[121]), 
        .QN() );
  DFF_X1 stateArray_S00reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S00reg_gff_1_SFF_2_QD), .CK(clk_gated), .Q(
        ciphertext_s0[122]), .QN() );
  DFF_X1 stateArray_S00reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3128), .CK(clk_gated), .Q(ciphertext_s1[122]), 
        .QN() );
  DFF_X1 stateArray_S00reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S00reg_gff_1_SFF_3_QD), .CK(clk_gated), .Q(
        ciphertext_s0[123]), .QN() );
  DFF_X1 stateArray_S00reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3129), .CK(clk_gated), .Q(ciphertext_s1[123]), 
        .QN() );
  DFF_X1 stateArray_S00reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S00reg_gff_1_SFF_4_QD), .CK(clk_gated), .Q(
        ciphertext_s0[124]), .QN() );
  DFF_X1 stateArray_S00reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3130), .CK(clk_gated), .Q(ciphertext_s1[124]), 
        .QN() );
  DFF_X1 stateArray_S00reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S00reg_gff_1_SFF_5_QD), .CK(clk_gated), .Q(
        ciphertext_s0[125]), .QN() );
  DFF_X1 stateArray_S00reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3131), .CK(clk_gated), .Q(ciphertext_s1[125]), 
        .QN() );
  DFF_X1 stateArray_S00reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S00reg_gff_1_SFF_6_QD), .CK(clk_gated), .Q(
        ciphertext_s0[126]), .QN() );
  DFF_X1 stateArray_S00reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3132), .CK(clk_gated), .Q(ciphertext_s1[126]), 
        .QN() );
  DFF_X1 stateArray_S00reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S00reg_gff_1_SFF_7_QD), .CK(clk_gated), .Q(
        ciphertext_s0[127]), .QN() );
  DFF_X1 stateArray_S00reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3133), .CK(clk_gated), .Q(ciphertext_s1[127]), 
        .QN() );
  DFF_X1 stateArray_S01reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S01reg_gff_1_SFF_0_QD), .CK(clk_gated), .Q(
        ciphertext_s0[112]), .QN() );
  DFF_X1 stateArray_S01reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3134), .CK(clk_gated), .Q(ciphertext_s1[112]), 
        .QN() );
  DFF_X1 stateArray_S01reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S01reg_gff_1_SFF_1_QD), .CK(clk_gated), .Q(
        ciphertext_s0[113]), .QN() );
  DFF_X1 stateArray_S01reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3135), .CK(clk_gated), .Q(ciphertext_s1[113]), 
        .QN() );
  DFF_X1 stateArray_S01reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S01reg_gff_1_SFF_2_QD), .CK(clk_gated), .Q(
        ciphertext_s0[114]), .QN() );
  DFF_X1 stateArray_S01reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3136), .CK(clk_gated), .Q(ciphertext_s1[114]), 
        .QN() );
  DFF_X1 stateArray_S01reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S01reg_gff_1_SFF_3_QD), .CK(clk_gated), .Q(
        ciphertext_s0[115]), .QN() );
  DFF_X1 stateArray_S01reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3137), .CK(clk_gated), .Q(ciphertext_s1[115]), 
        .QN() );
  DFF_X1 stateArray_S01reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S01reg_gff_1_SFF_4_QD), .CK(clk_gated), .Q(
        ciphertext_s0[116]), .QN() );
  DFF_X1 stateArray_S01reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3138), .CK(clk_gated), .Q(ciphertext_s1[116]), 
        .QN() );
  DFF_X1 stateArray_S01reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S01reg_gff_1_SFF_5_QD), .CK(clk_gated), .Q(
        ciphertext_s0[117]), .QN() );
  DFF_X1 stateArray_S01reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3139), .CK(clk_gated), .Q(ciphertext_s1[117]), 
        .QN() );
  DFF_X1 stateArray_S01reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S01reg_gff_1_SFF_6_QD), .CK(clk_gated), .Q(
        ciphertext_s0[118]), .QN() );
  DFF_X1 stateArray_S01reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3140), .CK(clk_gated), .Q(ciphertext_s1[118]), 
        .QN() );
  DFF_X1 stateArray_S01reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S01reg_gff_1_SFF_7_QD), .CK(clk_gated), .Q(
        ciphertext_s0[119]), .QN() );
  DFF_X1 stateArray_S01reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3141), .CK(clk_gated), .Q(ciphertext_s1[119]), 
        .QN() );
  DFF_X1 stateArray_S02reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S02reg_gff_1_SFF_0_QD), .CK(clk_gated), .Q(
        ciphertext_s0[104]), .QN() );
  DFF_X1 stateArray_S02reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3142), .CK(clk_gated), .Q(ciphertext_s1[104]), 
        .QN() );
  DFF_X1 stateArray_S02reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S02reg_gff_1_SFF_1_QD), .CK(clk_gated), .Q(
        ciphertext_s0[105]), .QN() );
  DFF_X1 stateArray_S02reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3143), .CK(clk_gated), .Q(ciphertext_s1[105]), 
        .QN() );
  DFF_X1 stateArray_S02reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S02reg_gff_1_SFF_2_QD), .CK(clk_gated), .Q(
        ciphertext_s0[106]), .QN() );
  DFF_X1 stateArray_S02reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3144), .CK(clk_gated), .Q(ciphertext_s1[106]), 
        .QN() );
  DFF_X1 stateArray_S02reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S02reg_gff_1_SFF_3_QD), .CK(clk_gated), .Q(
        ciphertext_s0[107]), .QN() );
  DFF_X1 stateArray_S02reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3145), .CK(clk_gated), .Q(ciphertext_s1[107]), 
        .QN() );
  DFF_X1 stateArray_S02reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S02reg_gff_1_SFF_4_QD), .CK(clk_gated), .Q(
        ciphertext_s0[108]), .QN() );
  DFF_X1 stateArray_S02reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3146), .CK(clk_gated), .Q(ciphertext_s1[108]), 
        .QN() );
  DFF_X1 stateArray_S02reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S02reg_gff_1_SFF_5_QD), .CK(clk_gated), .Q(
        ciphertext_s0[109]), .QN() );
  DFF_X1 stateArray_S02reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3147), .CK(clk_gated), .Q(ciphertext_s1[109]), 
        .QN() );
  DFF_X1 stateArray_S02reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S02reg_gff_1_SFF_6_QD), .CK(clk_gated), .Q(
        ciphertext_s0[110]), .QN() );
  DFF_X1 stateArray_S02reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3148), .CK(clk_gated), .Q(ciphertext_s1[110]), 
        .QN() );
  DFF_X1 stateArray_S02reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S02reg_gff_1_SFF_7_QD), .CK(clk_gated), .Q(
        ciphertext_s0[111]), .QN() );
  DFF_X1 stateArray_S02reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3149), .CK(clk_gated), .Q(ciphertext_s1[111]), 
        .QN() );
  DFF_X1 stateArray_S03reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S03reg_gff_1_SFF_0_QD), .CK(clk_gated), .Q(
        ciphertext_s0[96]), .QN() );
  DFF_X1 stateArray_S03reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3150), .CK(clk_gated), .Q(ciphertext_s1[96]), 
        .QN() );
  DFF_X1 stateArray_S03reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S03reg_gff_1_SFF_1_QD), .CK(clk_gated), .Q(
        ciphertext_s0[97]), .QN() );
  DFF_X1 stateArray_S03reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3151), .CK(clk_gated), .Q(ciphertext_s1[97]), 
        .QN() );
  DFF_X1 stateArray_S03reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S03reg_gff_1_SFF_2_QD), .CK(clk_gated), .Q(
        ciphertext_s0[98]), .QN() );
  DFF_X1 stateArray_S03reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3152), .CK(clk_gated), .Q(ciphertext_s1[98]), 
        .QN() );
  DFF_X1 stateArray_S03reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S03reg_gff_1_SFF_3_QD), .CK(clk_gated), .Q(
        ciphertext_s0[99]), .QN() );
  DFF_X1 stateArray_S03reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3153), .CK(clk_gated), .Q(ciphertext_s1[99]), 
        .QN() );
  DFF_X1 stateArray_S03reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S03reg_gff_1_SFF_4_QD), .CK(clk_gated), .Q(
        ciphertext_s0[100]), .QN() );
  DFF_X1 stateArray_S03reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3154), .CK(clk_gated), .Q(ciphertext_s1[100]), 
        .QN() );
  DFF_X1 stateArray_S03reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S03reg_gff_1_SFF_5_QD), .CK(clk_gated), .Q(
        ciphertext_s0[101]), .QN() );
  DFF_X1 stateArray_S03reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3155), .CK(clk_gated), .Q(ciphertext_s1[101]), 
        .QN() );
  DFF_X1 stateArray_S03reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S03reg_gff_1_SFF_6_QD), .CK(clk_gated), .Q(
        ciphertext_s0[102]), .QN() );
  DFF_X1 stateArray_S03reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3156), .CK(clk_gated), .Q(ciphertext_s1[102]), 
        .QN() );
  DFF_X1 stateArray_S03reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S03reg_gff_1_SFF_7_QD), .CK(clk_gated), .Q(
        ciphertext_s0[103]), .QN() );
  DFF_X1 stateArray_S03reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3157), .CK(clk_gated), .Q(ciphertext_s1[103]), 
        .QN() );
  DFF_X1 stateArray_S10reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S10reg_gff_1_SFF_0_QD), .CK(clk_gated), .Q(
        ciphertext_s0[88]), .QN() );
  DFF_X1 stateArray_S10reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3158), .CK(clk_gated), .Q(ciphertext_s1[88]), 
        .QN() );
  DFF_X1 stateArray_S10reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S10reg_gff_1_SFF_1_QD), .CK(clk_gated), .Q(
        ciphertext_s0[89]), .QN() );
  DFF_X1 stateArray_S10reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3159), .CK(clk_gated), .Q(ciphertext_s1[89]), 
        .QN() );
  DFF_X1 stateArray_S10reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S10reg_gff_1_SFF_2_QD), .CK(clk_gated), .Q(
        ciphertext_s0[90]), .QN() );
  DFF_X1 stateArray_S10reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3160), .CK(clk_gated), .Q(ciphertext_s1[90]), 
        .QN() );
  DFF_X1 stateArray_S10reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S10reg_gff_1_SFF_3_QD), .CK(clk_gated), .Q(
        ciphertext_s0[91]), .QN() );
  DFF_X1 stateArray_S10reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3161), .CK(clk_gated), .Q(ciphertext_s1[91]), 
        .QN() );
  DFF_X1 stateArray_S10reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S10reg_gff_1_SFF_4_QD), .CK(clk_gated), .Q(
        ciphertext_s0[92]), .QN() );
  DFF_X1 stateArray_S10reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3162), .CK(clk_gated), .Q(ciphertext_s1[92]), 
        .QN() );
  DFF_X1 stateArray_S10reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S10reg_gff_1_SFF_5_QD), .CK(clk_gated), .Q(
        ciphertext_s0[93]), .QN() );
  DFF_X1 stateArray_S10reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3163), .CK(clk_gated), .Q(ciphertext_s1[93]), 
        .QN() );
  DFF_X1 stateArray_S10reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S10reg_gff_1_SFF_6_QD), .CK(clk_gated), .Q(
        ciphertext_s0[94]), .QN() );
  DFF_X1 stateArray_S10reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3164), .CK(clk_gated), .Q(ciphertext_s1[94]), 
        .QN() );
  DFF_X1 stateArray_S10reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S10reg_gff_1_SFF_7_QD), .CK(clk_gated), .Q(
        ciphertext_s0[95]), .QN() );
  DFF_X1 stateArray_S10reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3165), .CK(clk_gated), .Q(ciphertext_s1[95]), 
        .QN() );
  DFF_X1 stateArray_S11reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S11reg_gff_1_SFF_0_QD), .CK(clk_gated), .Q(
        ciphertext_s0[80]), .QN() );
  DFF_X1 stateArray_S11reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3166), .CK(clk_gated), .Q(ciphertext_s1[80]), 
        .QN() );
  DFF_X1 stateArray_S11reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S11reg_gff_1_SFF_1_QD), .CK(clk_gated), .Q(
        ciphertext_s0[81]), .QN() );
  DFF_X1 stateArray_S11reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3167), .CK(clk_gated), .Q(ciphertext_s1[81]), 
        .QN() );
  DFF_X1 stateArray_S11reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S11reg_gff_1_SFF_2_QD), .CK(clk_gated), .Q(
        ciphertext_s0[82]), .QN() );
  DFF_X1 stateArray_S11reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3168), .CK(clk_gated), .Q(ciphertext_s1[82]), 
        .QN() );
  DFF_X1 stateArray_S11reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S11reg_gff_1_SFF_3_QD), .CK(clk_gated), .Q(
        ciphertext_s0[83]), .QN() );
  DFF_X1 stateArray_S11reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3169), .CK(clk_gated), .Q(ciphertext_s1[83]), 
        .QN() );
  DFF_X1 stateArray_S11reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S11reg_gff_1_SFF_4_QD), .CK(clk_gated), .Q(
        ciphertext_s0[84]), .QN() );
  DFF_X1 stateArray_S11reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3170), .CK(clk_gated), .Q(ciphertext_s1[84]), 
        .QN() );
  DFF_X1 stateArray_S11reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S11reg_gff_1_SFF_5_QD), .CK(clk_gated), .Q(
        ciphertext_s0[85]), .QN() );
  DFF_X1 stateArray_S11reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3171), .CK(clk_gated), .Q(ciphertext_s1[85]), 
        .QN() );
  DFF_X1 stateArray_S11reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S11reg_gff_1_SFF_6_QD), .CK(clk_gated), .Q(
        ciphertext_s0[86]), .QN() );
  DFF_X1 stateArray_S11reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3172), .CK(clk_gated), .Q(ciphertext_s1[86]), 
        .QN() );
  DFF_X1 stateArray_S11reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S11reg_gff_1_SFF_7_QD), .CK(clk_gated), .Q(
        ciphertext_s0[87]), .QN() );
  DFF_X1 stateArray_S11reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3173), .CK(clk_gated), .Q(ciphertext_s1[87]), 
        .QN() );
  DFF_X1 stateArray_S12reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S12reg_gff_1_SFF_0_QD), .CK(clk_gated), .Q(
        ciphertext_s0[72]), .QN() );
  DFF_X1 stateArray_S12reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3174), .CK(clk_gated), .Q(ciphertext_s1[72]), 
        .QN() );
  DFF_X1 stateArray_S12reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S12reg_gff_1_SFF_1_QD), .CK(clk_gated), .Q(
        ciphertext_s0[73]), .QN() );
  DFF_X1 stateArray_S12reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3175), .CK(clk_gated), .Q(ciphertext_s1[73]), 
        .QN() );
  DFF_X1 stateArray_S12reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S12reg_gff_1_SFF_2_QD), .CK(clk_gated), .Q(
        ciphertext_s0[74]), .QN() );
  DFF_X1 stateArray_S12reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3176), .CK(clk_gated), .Q(ciphertext_s1[74]), 
        .QN() );
  DFF_X1 stateArray_S12reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S12reg_gff_1_SFF_3_QD), .CK(clk_gated), .Q(
        ciphertext_s0[75]), .QN() );
  DFF_X1 stateArray_S12reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3177), .CK(clk_gated), .Q(ciphertext_s1[75]), 
        .QN() );
  DFF_X1 stateArray_S12reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S12reg_gff_1_SFF_4_QD), .CK(clk_gated), .Q(
        ciphertext_s0[76]), .QN() );
  DFF_X1 stateArray_S12reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3178), .CK(clk_gated), .Q(ciphertext_s1[76]), 
        .QN() );
  DFF_X1 stateArray_S12reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S12reg_gff_1_SFF_5_QD), .CK(clk_gated), .Q(
        ciphertext_s0[77]), .QN() );
  DFF_X1 stateArray_S12reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3179), .CK(clk_gated), .Q(ciphertext_s1[77]), 
        .QN() );
  DFF_X1 stateArray_S12reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S12reg_gff_1_SFF_6_QD), .CK(clk_gated), .Q(
        ciphertext_s0[78]), .QN() );
  DFF_X1 stateArray_S12reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3180), .CK(clk_gated), .Q(ciphertext_s1[78]), 
        .QN() );
  DFF_X1 stateArray_S12reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S12reg_gff_1_SFF_7_QD), .CK(clk_gated), .Q(
        ciphertext_s0[79]), .QN() );
  DFF_X1 stateArray_S12reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3181), .CK(clk_gated), .Q(ciphertext_s1[79]), 
        .QN() );
  DFF_X1 stateArray_S13reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S13reg_gff_1_SFF_0_QD), .CK(clk_gated), .Q(
        ciphertext_s0[64]), .QN() );
  DFF_X1 stateArray_S13reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3182), .CK(clk_gated), .Q(ciphertext_s1[64]), 
        .QN() );
  DFF_X1 stateArray_S13reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S13reg_gff_1_SFF_1_QD), .CK(clk_gated), .Q(
        ciphertext_s0[65]), .QN() );
  DFF_X1 stateArray_S13reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3183), .CK(clk_gated), .Q(ciphertext_s1[65]), 
        .QN() );
  DFF_X1 stateArray_S13reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S13reg_gff_1_SFF_2_QD), .CK(clk_gated), .Q(
        ciphertext_s0[66]), .QN() );
  DFF_X1 stateArray_S13reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3184), .CK(clk_gated), .Q(ciphertext_s1[66]), 
        .QN() );
  DFF_X1 stateArray_S13reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S13reg_gff_1_SFF_3_QD), .CK(clk_gated), .Q(
        ciphertext_s0[67]), .QN() );
  DFF_X1 stateArray_S13reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3185), .CK(clk_gated), .Q(ciphertext_s1[67]), 
        .QN() );
  DFF_X1 stateArray_S13reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S13reg_gff_1_SFF_4_QD), .CK(clk_gated), .Q(
        ciphertext_s0[68]), .QN() );
  DFF_X1 stateArray_S13reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3186), .CK(clk_gated), .Q(ciphertext_s1[68]), 
        .QN() );
  DFF_X1 stateArray_S13reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S13reg_gff_1_SFF_5_QD), .CK(clk_gated), .Q(
        ciphertext_s0[69]), .QN() );
  DFF_X1 stateArray_S13reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3187), .CK(clk_gated), .Q(ciphertext_s1[69]), 
        .QN() );
  DFF_X1 stateArray_S13reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S13reg_gff_1_SFF_6_QD), .CK(clk_gated), .Q(
        ciphertext_s0[70]), .QN() );
  DFF_X1 stateArray_S13reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3188), .CK(clk_gated), .Q(ciphertext_s1[70]), 
        .QN() );
  DFF_X1 stateArray_S13reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S13reg_gff_1_SFF_7_QD), .CK(clk_gated), .Q(
        ciphertext_s0[71]), .QN() );
  DFF_X1 stateArray_S13reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3189), .CK(clk_gated), .Q(ciphertext_s1[71]), 
        .QN() );
  DFF_X1 stateArray_S20reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S20reg_gff_1_SFF_0_QD), .CK(clk_gated), .Q(
        ciphertext_s0[56]), .QN() );
  DFF_X1 stateArray_S20reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3190), .CK(clk_gated), .Q(ciphertext_s1[56]), 
        .QN() );
  DFF_X1 stateArray_S20reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S20reg_gff_1_SFF_1_QD), .CK(clk_gated), .Q(
        ciphertext_s0[57]), .QN() );
  DFF_X1 stateArray_S20reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3191), .CK(clk_gated), .Q(ciphertext_s1[57]), 
        .QN() );
  DFF_X1 stateArray_S20reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S20reg_gff_1_SFF_2_QD), .CK(clk_gated), .Q(
        ciphertext_s0[58]), .QN() );
  DFF_X1 stateArray_S20reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3192), .CK(clk_gated), .Q(ciphertext_s1[58]), 
        .QN() );
  DFF_X1 stateArray_S20reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S20reg_gff_1_SFF_3_QD), .CK(clk_gated), .Q(
        ciphertext_s0[59]), .QN() );
  DFF_X1 stateArray_S20reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3193), .CK(clk_gated), .Q(ciphertext_s1[59]), 
        .QN() );
  DFF_X1 stateArray_S20reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S20reg_gff_1_SFF_4_QD), .CK(clk_gated), .Q(
        ciphertext_s0[60]), .QN() );
  DFF_X1 stateArray_S20reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3194), .CK(clk_gated), .Q(ciphertext_s1[60]), 
        .QN() );
  DFF_X1 stateArray_S20reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S20reg_gff_1_SFF_5_QD), .CK(clk_gated), .Q(
        ciphertext_s0[61]), .QN() );
  DFF_X1 stateArray_S20reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3195), .CK(clk_gated), .Q(ciphertext_s1[61]), 
        .QN() );
  DFF_X1 stateArray_S20reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S20reg_gff_1_SFF_6_QD), .CK(clk_gated), .Q(
        ciphertext_s0[62]), .QN() );
  DFF_X1 stateArray_S20reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3196), .CK(clk_gated), .Q(ciphertext_s1[62]), 
        .QN() );
  DFF_X1 stateArray_S20reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S20reg_gff_1_SFF_7_QD), .CK(clk_gated), .Q(
        ciphertext_s0[63]), .QN() );
  DFF_X1 stateArray_S20reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3197), .CK(clk_gated), .Q(ciphertext_s1[63]), 
        .QN() );
  DFF_X1 stateArray_S21reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S21reg_gff_1_SFF_0_QD), .CK(clk_gated), .Q(
        ciphertext_s0[48]), .QN() );
  DFF_X1 stateArray_S21reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3198), .CK(clk_gated), .Q(ciphertext_s1[48]), 
        .QN() );
  DFF_X1 stateArray_S21reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S21reg_gff_1_SFF_1_QD), .CK(clk_gated), .Q(
        ciphertext_s0[49]), .QN() );
  DFF_X1 stateArray_S21reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3199), .CK(clk_gated), .Q(ciphertext_s1[49]), 
        .QN() );
  DFF_X1 stateArray_S21reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S21reg_gff_1_SFF_2_QD), .CK(clk_gated), .Q(
        ciphertext_s0[50]), .QN() );
  DFF_X1 stateArray_S21reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3200), .CK(clk_gated), .Q(ciphertext_s1[50]), 
        .QN() );
  DFF_X1 stateArray_S21reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S21reg_gff_1_SFF_3_QD), .CK(clk_gated), .Q(
        ciphertext_s0[51]), .QN() );
  DFF_X1 stateArray_S21reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3201), .CK(clk_gated), .Q(ciphertext_s1[51]), 
        .QN() );
  DFF_X1 stateArray_S21reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S21reg_gff_1_SFF_4_QD), .CK(clk_gated), .Q(
        ciphertext_s0[52]), .QN() );
  DFF_X1 stateArray_S21reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3202), .CK(clk_gated), .Q(ciphertext_s1[52]), 
        .QN() );
  DFF_X1 stateArray_S21reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S21reg_gff_1_SFF_5_QD), .CK(clk_gated), .Q(
        ciphertext_s0[53]), .QN() );
  DFF_X1 stateArray_S21reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3203), .CK(clk_gated), .Q(ciphertext_s1[53]), 
        .QN() );
  DFF_X1 stateArray_S21reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S21reg_gff_1_SFF_6_QD), .CK(clk_gated), .Q(
        ciphertext_s0[54]), .QN() );
  DFF_X1 stateArray_S21reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3204), .CK(clk_gated), .Q(ciphertext_s1[54]), 
        .QN() );
  DFF_X1 stateArray_S21reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S21reg_gff_1_SFF_7_QD), .CK(clk_gated), .Q(
        ciphertext_s0[55]), .QN() );
  DFF_X1 stateArray_S21reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3205), .CK(clk_gated), .Q(ciphertext_s1[55]), 
        .QN() );
  DFF_X1 stateArray_S22reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S22reg_gff_1_SFF_0_QD), .CK(clk_gated), .Q(
        ciphertext_s0[40]), .QN() );
  DFF_X1 stateArray_S22reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3206), .CK(clk_gated), .Q(ciphertext_s1[40]), 
        .QN() );
  DFF_X1 stateArray_S22reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S22reg_gff_1_SFF_1_QD), .CK(clk_gated), .Q(
        ciphertext_s0[41]), .QN() );
  DFF_X1 stateArray_S22reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3207), .CK(clk_gated), .Q(ciphertext_s1[41]), 
        .QN() );
  DFF_X1 stateArray_S22reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S22reg_gff_1_SFF_2_QD), .CK(clk_gated), .Q(
        ciphertext_s0[42]), .QN() );
  DFF_X1 stateArray_S22reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3208), .CK(clk_gated), .Q(ciphertext_s1[42]), 
        .QN() );
  DFF_X1 stateArray_S22reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S22reg_gff_1_SFF_3_QD), .CK(clk_gated), .Q(
        ciphertext_s0[43]), .QN() );
  DFF_X1 stateArray_S22reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3209), .CK(clk_gated), .Q(ciphertext_s1[43]), 
        .QN() );
  DFF_X1 stateArray_S22reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S22reg_gff_1_SFF_4_QD), .CK(clk_gated), .Q(
        ciphertext_s0[44]), .QN() );
  DFF_X1 stateArray_S22reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3210), .CK(clk_gated), .Q(ciphertext_s1[44]), 
        .QN() );
  DFF_X1 stateArray_S22reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S22reg_gff_1_SFF_5_QD), .CK(clk_gated), .Q(
        ciphertext_s0[45]), .QN() );
  DFF_X1 stateArray_S22reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3211), .CK(clk_gated), .Q(ciphertext_s1[45]), 
        .QN() );
  DFF_X1 stateArray_S22reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S22reg_gff_1_SFF_6_QD), .CK(clk_gated), .Q(
        ciphertext_s0[46]), .QN() );
  DFF_X1 stateArray_S22reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3212), .CK(clk_gated), .Q(ciphertext_s1[46]), 
        .QN() );
  DFF_X1 stateArray_S22reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S22reg_gff_1_SFF_7_QD), .CK(clk_gated), .Q(
        ciphertext_s0[47]), .QN() );
  DFF_X1 stateArray_S22reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3213), .CK(clk_gated), .Q(ciphertext_s1[47]), 
        .QN() );
  DFF_X1 stateArray_S23reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S23reg_gff_1_SFF_0_QD), .CK(clk_gated), .Q(
        ciphertext_s0[32]), .QN() );
  DFF_X1 stateArray_S23reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3214), .CK(clk_gated), .Q(ciphertext_s1[32]), 
        .QN() );
  DFF_X1 stateArray_S23reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S23reg_gff_1_SFF_1_QD), .CK(clk_gated), .Q(
        ciphertext_s0[33]), .QN() );
  DFF_X1 stateArray_S23reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3215), .CK(clk_gated), .Q(ciphertext_s1[33]), 
        .QN() );
  DFF_X1 stateArray_S23reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S23reg_gff_1_SFF_2_QD), .CK(clk_gated), .Q(
        ciphertext_s0[34]), .QN() );
  DFF_X1 stateArray_S23reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3216), .CK(clk_gated), .Q(ciphertext_s1[34]), 
        .QN() );
  DFF_X1 stateArray_S23reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S23reg_gff_1_SFF_3_QD), .CK(clk_gated), .Q(
        ciphertext_s0[35]), .QN() );
  DFF_X1 stateArray_S23reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3217), .CK(clk_gated), .Q(ciphertext_s1[35]), 
        .QN() );
  DFF_X1 stateArray_S23reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S23reg_gff_1_SFF_4_QD), .CK(clk_gated), .Q(
        ciphertext_s0[36]), .QN() );
  DFF_X1 stateArray_S23reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3218), .CK(clk_gated), .Q(ciphertext_s1[36]), 
        .QN() );
  DFF_X1 stateArray_S23reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S23reg_gff_1_SFF_5_QD), .CK(clk_gated), .Q(
        ciphertext_s0[37]), .QN() );
  DFF_X1 stateArray_S23reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3219), .CK(clk_gated), .Q(ciphertext_s1[37]), 
        .QN() );
  DFF_X1 stateArray_S23reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S23reg_gff_1_SFF_6_QD), .CK(clk_gated), .Q(
        ciphertext_s0[38]), .QN() );
  DFF_X1 stateArray_S23reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3220), .CK(clk_gated), .Q(ciphertext_s1[38]), 
        .QN() );
  DFF_X1 stateArray_S23reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S23reg_gff_1_SFF_7_QD), .CK(clk_gated), .Q(
        ciphertext_s0[39]), .QN() );
  DFF_X1 stateArray_S23reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3221), .CK(clk_gated), .Q(ciphertext_s1[39]), 
        .QN() );
  DFF_X1 stateArray_S30reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S30reg_gff_1_SFF_0_QD), .CK(clk_gated), .Q(
        ciphertext_s0[24]), .QN() );
  DFF_X1 stateArray_S30reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3222), .CK(clk_gated), .Q(ciphertext_s1[24]), 
        .QN() );
  DFF_X1 stateArray_S30reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S30reg_gff_1_SFF_1_QD), .CK(clk_gated), .Q(
        ciphertext_s0[25]), .QN() );
  DFF_X1 stateArray_S30reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3223), .CK(clk_gated), .Q(ciphertext_s1[25]), 
        .QN() );
  DFF_X1 stateArray_S30reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S30reg_gff_1_SFF_2_QD), .CK(clk_gated), .Q(
        ciphertext_s0[26]), .QN() );
  DFF_X1 stateArray_S30reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3224), .CK(clk_gated), .Q(ciphertext_s1[26]), 
        .QN() );
  DFF_X1 stateArray_S30reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S30reg_gff_1_SFF_3_QD), .CK(clk_gated), .Q(
        ciphertext_s0[27]), .QN() );
  DFF_X1 stateArray_S30reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3225), .CK(clk_gated), .Q(ciphertext_s1[27]), 
        .QN() );
  DFF_X1 stateArray_S30reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S30reg_gff_1_SFF_4_QD), .CK(clk_gated), .Q(
        ciphertext_s0[28]), .QN() );
  DFF_X1 stateArray_S30reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3226), .CK(clk_gated), .Q(ciphertext_s1[28]), 
        .QN() );
  DFF_X1 stateArray_S30reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S30reg_gff_1_SFF_5_QD), .CK(clk_gated), .Q(
        ciphertext_s0[29]), .QN() );
  DFF_X1 stateArray_S30reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3227), .CK(clk_gated), .Q(ciphertext_s1[29]), 
        .QN() );
  DFF_X1 stateArray_S30reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S30reg_gff_1_SFF_6_QD), .CK(clk_gated), .Q(
        ciphertext_s0[30]), .QN() );
  DFF_X1 stateArray_S30reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3228), .CK(clk_gated), .Q(ciphertext_s1[30]), 
        .QN() );
  DFF_X1 stateArray_S30reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S30reg_gff_1_SFF_7_QD), .CK(clk_gated), .Q(
        ciphertext_s0[31]), .QN() );
  DFF_X1 stateArray_S30reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3229), .CK(clk_gated), .Q(ciphertext_s1[31]), 
        .QN() );
  DFF_X1 stateArray_S31reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S31reg_gff_1_SFF_0_QD), .CK(clk_gated), .Q(
        ciphertext_s0[16]), .QN() );
  DFF_X1 stateArray_S31reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3230), .CK(clk_gated), .Q(ciphertext_s1[16]), 
        .QN() );
  DFF_X1 stateArray_S31reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S31reg_gff_1_SFF_1_QD), .CK(clk_gated), .Q(
        ciphertext_s0[17]), .QN() );
  DFF_X1 stateArray_S31reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3231), .CK(clk_gated), .Q(ciphertext_s1[17]), 
        .QN() );
  DFF_X1 stateArray_S31reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S31reg_gff_1_SFF_2_QD), .CK(clk_gated), .Q(
        ciphertext_s0[18]), .QN() );
  DFF_X1 stateArray_S31reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3232), .CK(clk_gated), .Q(ciphertext_s1[18]), 
        .QN() );
  DFF_X1 stateArray_S31reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S31reg_gff_1_SFF_3_QD), .CK(clk_gated), .Q(
        ciphertext_s0[19]), .QN() );
  DFF_X1 stateArray_S31reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3233), .CK(clk_gated), .Q(ciphertext_s1[19]), 
        .QN() );
  DFF_X1 stateArray_S31reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S31reg_gff_1_SFF_4_QD), .CK(clk_gated), .Q(
        ciphertext_s0[20]), .QN() );
  DFF_X1 stateArray_S31reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3234), .CK(clk_gated), .Q(ciphertext_s1[20]), 
        .QN() );
  DFF_X1 stateArray_S31reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S31reg_gff_1_SFF_5_QD), .CK(clk_gated), .Q(
        ciphertext_s0[21]), .QN() );
  DFF_X1 stateArray_S31reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3235), .CK(clk_gated), .Q(ciphertext_s1[21]), 
        .QN() );
  DFF_X1 stateArray_S31reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S31reg_gff_1_SFF_6_QD), .CK(clk_gated), .Q(
        ciphertext_s0[22]), .QN() );
  DFF_X1 stateArray_S31reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3236), .CK(clk_gated), .Q(ciphertext_s1[22]), 
        .QN() );
  DFF_X1 stateArray_S31reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S31reg_gff_1_SFF_7_QD), .CK(clk_gated), .Q(
        ciphertext_s0[23]), .QN() );
  DFF_X1 stateArray_S31reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3237), .CK(clk_gated), .Q(ciphertext_s1[23]), 
        .QN() );
  DFF_X1 stateArray_S32reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S32reg_gff_1_SFF_0_QD), .CK(clk_gated), .Q(
        ciphertext_s0[8]), .QN() );
  DFF_X1 stateArray_S32reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3238), .CK(clk_gated), .Q(ciphertext_s1[8]), .QN()
         );
  DFF_X1 stateArray_S32reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S32reg_gff_1_SFF_1_QD), .CK(clk_gated), .Q(
        ciphertext_s0[9]), .QN() );
  DFF_X1 stateArray_S32reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3239), .CK(clk_gated), .Q(ciphertext_s1[9]), .QN()
         );
  DFF_X1 stateArray_S32reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S32reg_gff_1_SFF_2_QD), .CK(clk_gated), .Q(
        ciphertext_s0[10]), .QN() );
  DFF_X1 stateArray_S32reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3240), .CK(clk_gated), .Q(ciphertext_s1[10]), 
        .QN() );
  DFF_X1 stateArray_S32reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S32reg_gff_1_SFF_3_QD), .CK(clk_gated), .Q(
        ciphertext_s0[11]), .QN() );
  DFF_X1 stateArray_S32reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3241), .CK(clk_gated), .Q(ciphertext_s1[11]), 
        .QN() );
  DFF_X1 stateArray_S32reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S32reg_gff_1_SFF_4_QD), .CK(clk_gated), .Q(
        ciphertext_s0[12]), .QN() );
  DFF_X1 stateArray_S32reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3242), .CK(clk_gated), .Q(ciphertext_s1[12]), 
        .QN() );
  DFF_X1 stateArray_S32reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S32reg_gff_1_SFF_5_QD), .CK(clk_gated), .Q(
        ciphertext_s0[13]), .QN() );
  DFF_X1 stateArray_S32reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3243), .CK(clk_gated), .Q(ciphertext_s1[13]), 
        .QN() );
  DFF_X1 stateArray_S32reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S32reg_gff_1_SFF_6_QD), .CK(clk_gated), .Q(
        ciphertext_s0[14]), .QN() );
  DFF_X1 stateArray_S32reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3244), .CK(clk_gated), .Q(ciphertext_s1[14]), 
        .QN() );
  DFF_X1 stateArray_S32reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S32reg_gff_1_SFF_7_QD), .CK(clk_gated), .Q(
        ciphertext_s0[15]), .QN() );
  DFF_X1 stateArray_S32reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3245), .CK(clk_gated), .Q(ciphertext_s1[15]), 
        .QN() );
  DFF_X1 stateArray_S33reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S33reg_gff_1_SFF_0_QD), .CK(clk_gated), .Q(
        ciphertext_s0[0]), .QN() );
  DFF_X1 stateArray_S33reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3497), .CK(clk_gated), .Q(ciphertext_s1[0]), .QN()
         );
  DFF_X1 stateArray_S33reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S33reg_gff_1_SFF_1_QD), .CK(clk_gated), .Q(
        ciphertext_s0[1]), .QN() );
  DFF_X1 stateArray_S33reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3520), .CK(clk_gated), .Q(ciphertext_s1[1]), .QN()
         );
  DFF_X1 stateArray_S33reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S33reg_gff_1_SFF_2_QD), .CK(clk_gated), .Q(
        ciphertext_s0[2]), .QN() );
  DFF_X1 stateArray_S33reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3521), .CK(clk_gated), .Q(ciphertext_s1[2]), .QN()
         );
  DFF_X1 stateArray_S33reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S33reg_gff_1_SFF_3_QD), .CK(clk_gated), .Q(
        ciphertext_s0[3]), .QN() );
  DFF_X1 stateArray_S33reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3522), .CK(clk_gated), .Q(ciphertext_s1[3]), .QN()
         );
  DFF_X1 stateArray_S33reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S33reg_gff_1_SFF_4_QD), .CK(clk_gated), .Q(
        ciphertext_s0[4]), .QN() );
  DFF_X1 stateArray_S33reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3523), .CK(clk_gated), .Q(ciphertext_s1[4]), .QN()
         );
  DFF_X1 stateArray_S33reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S33reg_gff_1_SFF_5_QD), .CK(clk_gated), .Q(
        ciphertext_s0[5]), .QN() );
  DFF_X1 stateArray_S33reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3524), .CK(clk_gated), .Q(ciphertext_s1[5]), .QN()
         );
  DFF_X1 stateArray_S33reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S33reg_gff_1_SFF_6_QD), .CK(clk_gated), .Q(
        ciphertext_s0[6]), .QN() );
  DFF_X1 stateArray_S33reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3525), .CK(clk_gated), .Q(ciphertext_s1[6]), .QN()
         );
  DFF_X1 stateArray_S33reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(stateArray_S33reg_gff_1_SFF_7_QD), .CK(clk_gated), .Q(
        ciphertext_s0[7]), .QN() );
  DFF_X1 stateArray_S33reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3526), .CK(clk_gated), .Q(ciphertext_s1[7]), .QN()
         );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S00reg_gff_1_SFF_0_n5), .CK(clk_gated), .Q(keyStateIn[0]), 
        .QN() );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3375), .CK(clk_gated), .Q(new_AGEMA_signal_1983), 
        .QN() );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S00reg_gff_1_SFF_1_n6), .CK(clk_gated), .Q(keyStateIn[1]), 
        .QN() );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3376), .CK(clk_gated), .Q(new_AGEMA_signal_1986), 
        .QN() );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S00reg_gff_1_SFF_2_n6), .CK(clk_gated), .Q(keyStateIn[2]), 
        .QN() );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3377), .CK(clk_gated), .Q(new_AGEMA_signal_1989), 
        .QN() );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S00reg_gff_1_SFF_3_n6), .CK(clk_gated), .Q(keyStateIn[3]), 
        .QN() );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3378), .CK(clk_gated), .Q(new_AGEMA_signal_1992), 
        .QN() );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S00reg_gff_1_SFF_4_n6), .CK(clk_gated), .Q(keyStateIn[4]), 
        .QN() );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3379), .CK(clk_gated), .Q(new_AGEMA_signal_1995), 
        .QN() );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S00reg_gff_1_SFF_5_n6), .CK(clk_gated), .Q(keyStateIn[5]), 
        .QN() );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3380), .CK(clk_gated), .Q(new_AGEMA_signal_1998), 
        .QN() );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S00reg_gff_1_SFF_6_n6), .CK(clk_gated), .Q(keyStateIn[6]), 
        .QN() );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3381), .CK(clk_gated), .Q(new_AGEMA_signal_2001), 
        .QN() );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S00reg_gff_1_SFF_7_n6), .CK(clk_gated), .Q(keyStateIn[7]), 
        .QN() );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3382), .CK(clk_gated), .Q(new_AGEMA_signal_2004), 
        .QN() );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S01reg_gff_1_SFF_0_n6), .CK(clk_gated), .Q(
        KeyArray_outS01ser_0_), .QN() );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3275), .CK(clk_gated), .Q(new_AGEMA_signal_2020), 
        .QN() );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S01reg_gff_1_SFF_1_n6), .CK(clk_gated), .Q(
        KeyArray_outS01ser_1_), .QN() );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3276), .CK(clk_gated), .Q(new_AGEMA_signal_2018), 
        .QN() );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S01reg_gff_1_SFF_2_n6), .CK(clk_gated), .Q(
        KeyArray_outS01ser_2_), .QN() );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3277), .CK(clk_gated), .Q(new_AGEMA_signal_2016), 
        .QN() );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S01reg_gff_1_SFF_3_n6), .CK(clk_gated), .Q(
        KeyArray_outS01ser_3_), .QN() );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3278), .CK(clk_gated), .Q(new_AGEMA_signal_2014), 
        .QN() );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S01reg_gff_1_SFF_4_n6), .CK(clk_gated), .Q(
        KeyArray_outS01ser_4_), .QN() );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3279), .CK(clk_gated), .Q(new_AGEMA_signal_2012), 
        .QN() );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S01reg_gff_1_SFF_5_n6), .CK(clk_gated), .Q(
        KeyArray_outS01ser_5_), .QN() );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3280), .CK(clk_gated), .Q(new_AGEMA_signal_2010), 
        .QN() );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S01reg_gff_1_SFF_6_n6), .CK(clk_gated), .Q(
        KeyArray_outS01ser_6_), .QN() );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3281), .CK(clk_gated), .Q(new_AGEMA_signal_2008), 
        .QN() );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S01reg_gff_1_SFF_7_n6), .CK(clk_gated), .Q(
        KeyArray_outS01ser_7_), .QN() );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3282), .CK(clk_gated), .Q(new_AGEMA_signal_2006), 
        .QN() );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S02reg_gff_1_SFF_0_n6), .CK(clk_gated), .Q(
        KeyArray_outS02ser[0]), .QN() );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3283), .CK(clk_gated), .Q(new_AGEMA_signal_2443), 
        .QN() );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S02reg_gff_1_SFF_1_n6), .CK(clk_gated), .Q(
        KeyArray_outS02ser[1]), .QN() );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3284), .CK(clk_gated), .Q(new_AGEMA_signal_2446), 
        .QN() );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S02reg_gff_1_SFF_2_n6), .CK(clk_gated), .Q(
        KeyArray_outS02ser[2]), .QN() );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3285), .CK(clk_gated), .Q(new_AGEMA_signal_2449), 
        .QN() );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S02reg_gff_1_SFF_3_n6), .CK(clk_gated), .Q(
        KeyArray_outS02ser[3]), .QN() );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3286), .CK(clk_gated), .Q(new_AGEMA_signal_2452), 
        .QN() );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S02reg_gff_1_SFF_4_n6), .CK(clk_gated), .Q(
        KeyArray_outS02ser[4]), .QN() );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3287), .CK(clk_gated), .Q(new_AGEMA_signal_2455), 
        .QN() );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S02reg_gff_1_SFF_5_n6), .CK(clk_gated), .Q(
        KeyArray_outS02ser[5]), .QN() );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3288), .CK(clk_gated), .Q(new_AGEMA_signal_2458), 
        .QN() );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S02reg_gff_1_SFF_6_n6), .CK(clk_gated), .Q(
        KeyArray_outS02ser[6]), .QN() );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3289), .CK(clk_gated), .Q(new_AGEMA_signal_2461), 
        .QN() );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S02reg_gff_1_SFF_7_n6), .CK(clk_gated), .Q(
        KeyArray_outS02ser[7]), .QN() );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3290), .CK(clk_gated), .Q(new_AGEMA_signal_2464), 
        .QN() );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S03reg_gff_1_SFF_0_n6), .CK(clk_gated), .Q(
        KeyArray_outS03ser[0]), .QN() );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3291), .CK(clk_gated), .Q(new_AGEMA_signal_2467), 
        .QN() );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S03reg_gff_1_SFF_1_n6), .CK(clk_gated), .Q(
        KeyArray_outS03ser[1]), .QN() );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3292), .CK(clk_gated), .Q(new_AGEMA_signal_2470), 
        .QN() );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S03reg_gff_1_SFF_2_n6), .CK(clk_gated), .Q(
        KeyArray_outS03ser[2]), .QN() );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3293), .CK(clk_gated), .Q(new_AGEMA_signal_2473), 
        .QN() );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S03reg_gff_1_SFF_3_n6), .CK(clk_gated), .Q(
        KeyArray_outS03ser[3]), .QN() );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3294), .CK(clk_gated), .Q(new_AGEMA_signal_2476), 
        .QN() );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S03reg_gff_1_SFF_4_n6), .CK(clk_gated), .Q(
        KeyArray_outS03ser[4]), .QN() );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3295), .CK(clk_gated), .Q(new_AGEMA_signal_2479), 
        .QN() );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S03reg_gff_1_SFF_5_n5), .CK(clk_gated), .Q(
        KeyArray_outS03ser[5]), .QN() );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3296), .CK(clk_gated), .Q(new_AGEMA_signal_2482), 
        .QN() );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S03reg_gff_1_SFF_6_n5), .CK(clk_gated), .Q(
        KeyArray_outS03ser[6]), .QN() );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3297), .CK(clk_gated), .Q(new_AGEMA_signal_2485), 
        .QN() );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S03reg_gff_1_SFF_7_n5), .CK(clk_gated), .Q(
        KeyArray_outS03ser[7]), .QN() );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3298), .CK(clk_gated), .Q(new_AGEMA_signal_2488), 
        .QN() );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S10reg_gff_1_SFF_0_n5), .CK(clk_gated), .Q(
        KeyArray_outS10ser[0]), .QN() );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3299), .CK(clk_gated), .Q(new_AGEMA_signal_2491), 
        .QN() );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S10reg_gff_1_SFF_1_n5), .CK(clk_gated), .Q(
        KeyArray_outS10ser[1]), .QN() );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3300), .CK(clk_gated), .Q(new_AGEMA_signal_2494), 
        .QN() );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S10reg_gff_1_SFF_2_n5), .CK(clk_gated), .Q(
        KeyArray_outS10ser[2]), .QN() );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3301), .CK(clk_gated), .Q(new_AGEMA_signal_2497), 
        .QN() );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S10reg_gff_1_SFF_3_n5), .CK(clk_gated), .Q(
        KeyArray_outS10ser[3]), .QN() );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3302), .CK(clk_gated), .Q(new_AGEMA_signal_2500), 
        .QN() );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S10reg_gff_1_SFF_4_n5), .CK(clk_gated), .Q(
        KeyArray_outS10ser[4]), .QN() );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3303), .CK(clk_gated), .Q(new_AGEMA_signal_2503), 
        .QN() );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S10reg_gff_1_SFF_5_n5), .CK(clk_gated), .Q(
        KeyArray_outS10ser[5]), .QN() );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3304), .CK(clk_gated), .Q(new_AGEMA_signal_2506), 
        .QN() );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S10reg_gff_1_SFF_6_n5), .CK(clk_gated), .Q(
        KeyArray_outS10ser[6]), .QN() );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3305), .CK(clk_gated), .Q(new_AGEMA_signal_2509), 
        .QN() );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S10reg_gff_1_SFF_7_n5), .CK(clk_gated), .Q(
        KeyArray_outS10ser[7]), .QN() );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3306), .CK(clk_gated), .Q(new_AGEMA_signal_2512), 
        .QN() );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S11reg_gff_1_SFF_0_n6), .CK(clk_gated), .Q(
        KeyArray_outS11ser[0]), .QN() );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3307), .CK(clk_gated), .Q(new_AGEMA_signal_2515), 
        .QN() );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S11reg_gff_1_SFF_1_n6), .CK(clk_gated), .Q(
        KeyArray_outS11ser[1]), .QN() );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3308), .CK(clk_gated), .Q(new_AGEMA_signal_2518), 
        .QN() );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S11reg_gff_1_SFF_2_n6), .CK(clk_gated), .Q(
        KeyArray_outS11ser[2]), .QN() );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3309), .CK(clk_gated), .Q(new_AGEMA_signal_2521), 
        .QN() );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S11reg_gff_1_SFF_3_n6), .CK(clk_gated), .Q(
        KeyArray_outS11ser[3]), .QN() );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3310), .CK(clk_gated), .Q(new_AGEMA_signal_2524), 
        .QN() );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S11reg_gff_1_SFF_4_n6), .CK(clk_gated), .Q(
        KeyArray_outS11ser[4]), .QN() );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3311), .CK(clk_gated), .Q(new_AGEMA_signal_2527), 
        .QN() );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S11reg_gff_1_SFF_5_n6), .CK(clk_gated), .Q(
        KeyArray_outS11ser[5]), .QN() );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3312), .CK(clk_gated), .Q(new_AGEMA_signal_2530), 
        .QN() );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S11reg_gff_1_SFF_6_n6), .CK(clk_gated), .Q(
        KeyArray_outS11ser[6]), .QN() );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3313), .CK(clk_gated), .Q(new_AGEMA_signal_2533), 
        .QN() );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S11reg_gff_1_SFF_7_n6), .CK(clk_gated), .Q(
        KeyArray_outS11ser[7]), .QN() );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3314), .CK(clk_gated), .Q(new_AGEMA_signal_2536), 
        .QN() );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S12reg_gff_1_SFF_0_n6), .CK(clk_gated), .Q(
        KeyArray_outS12ser[0]), .QN() );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3093), .CK(clk_gated), .Q(new_AGEMA_signal_2539), 
        .QN() );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S12reg_gff_1_SFF_1_n6), .CK(clk_gated), .Q(
        KeyArray_outS12ser[1]), .QN() );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3094), .CK(clk_gated), .Q(new_AGEMA_signal_2542), 
        .QN() );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S12reg_gff_1_SFF_2_n6), .CK(clk_gated), .Q(
        KeyArray_outS12ser[2]), .QN() );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3095), .CK(clk_gated), .Q(new_AGEMA_signal_2545), 
        .QN() );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S12reg_gff_1_SFF_3_n6), .CK(clk_gated), .Q(
        KeyArray_outS12ser[3]), .QN() );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3096), .CK(clk_gated), .Q(new_AGEMA_signal_2548), 
        .QN() );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S12reg_gff_1_SFF_4_n6), .CK(clk_gated), .Q(
        KeyArray_outS12ser[4]), .QN() );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3097), .CK(clk_gated), .Q(new_AGEMA_signal_2551), 
        .QN() );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S12reg_gff_1_SFF_5_n6), .CK(clk_gated), .Q(
        KeyArray_outS12ser[5]), .QN() );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3098), .CK(clk_gated), .Q(new_AGEMA_signal_2554), 
        .QN() );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S12reg_gff_1_SFF_6_n6), .CK(clk_gated), .Q(
        KeyArray_outS12ser[6]), .QN() );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3099), .CK(clk_gated), .Q(new_AGEMA_signal_2557), 
        .QN() );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S12reg_gff_1_SFF_7_n6), .CK(clk_gated), .Q(
        KeyArray_outS12ser[7]), .QN() );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3100), .CK(clk_gated), .Q(new_AGEMA_signal_2560), 
        .QN() );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S13reg_gff_1_SFF_0_n6), .CK(clk_gated), .Q(keySBIn[0]), 
        .QN() );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3101), .CK(clk_gated), .Q(new_AGEMA_signal_2563), 
        .QN() );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S13reg_gff_1_SFF_1_n6), .CK(clk_gated), .Q(keySBIn[1]), 
        .QN() );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3102), .CK(clk_gated), .Q(new_AGEMA_signal_2566), 
        .QN() );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S13reg_gff_1_SFF_2_n6), .CK(clk_gated), .Q(keySBIn[2]), 
        .QN() );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3103), .CK(clk_gated), .Q(new_AGEMA_signal_2569), 
        .QN() );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S13reg_gff_1_SFF_3_n6), .CK(clk_gated), .Q(keySBIn[3]), 
        .QN() );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3104), .CK(clk_gated), .Q(new_AGEMA_signal_2572), 
        .QN() );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S13reg_gff_1_SFF_4_n6), .CK(clk_gated), .Q(keySBIn[4]), 
        .QN() );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3105), .CK(clk_gated), .Q(new_AGEMA_signal_2575), 
        .QN() );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S13reg_gff_1_SFF_5_n5), .CK(clk_gated), .Q(keySBIn[5]), 
        .QN() );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3106), .CK(clk_gated), .Q(new_AGEMA_signal_2578), 
        .QN() );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S13reg_gff_1_SFF_6_n5), .CK(clk_gated), .Q(keySBIn[6]), 
        .QN() );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3107), .CK(clk_gated), .Q(new_AGEMA_signal_2581), 
        .QN() );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S13reg_gff_1_SFF_7_n5), .CK(clk_gated), .Q(keySBIn[7]), 
        .QN() );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3108), .CK(clk_gated), .Q(new_AGEMA_signal_2584), 
        .QN() );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S20reg_gff_1_SFF_0_n5), .CK(clk_gated), .Q(
        KeyArray_outS20ser[0]), .QN() );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3315), .CK(clk_gated), .Q(new_AGEMA_signal_2587), 
        .QN() );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S20reg_gff_1_SFF_1_n5), .CK(clk_gated), .Q(
        KeyArray_outS20ser[1]), .QN() );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3316), .CK(clk_gated), .Q(new_AGEMA_signal_2590), 
        .QN() );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S20reg_gff_1_SFF_2_n5), .CK(clk_gated), .Q(
        KeyArray_outS20ser[2]), .QN() );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3317), .CK(clk_gated), .Q(new_AGEMA_signal_2593), 
        .QN() );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S20reg_gff_1_SFF_3_n5), .CK(clk_gated), .Q(
        KeyArray_outS20ser[3]), .QN() );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3318), .CK(clk_gated), .Q(new_AGEMA_signal_2596), 
        .QN() );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S20reg_gff_1_SFF_4_n5), .CK(clk_gated), .Q(
        KeyArray_outS20ser[4]), .QN() );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3319), .CK(clk_gated), .Q(new_AGEMA_signal_2599), 
        .QN() );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S20reg_gff_1_SFF_5_n5), .CK(clk_gated), .Q(
        KeyArray_outS20ser[5]), .QN() );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3320), .CK(clk_gated), .Q(new_AGEMA_signal_2602), 
        .QN() );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S20reg_gff_1_SFF_6_n5), .CK(clk_gated), .Q(
        KeyArray_outS20ser[6]), .QN() );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3321), .CK(clk_gated), .Q(new_AGEMA_signal_2605), 
        .QN() );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S20reg_gff_1_SFF_7_n5), .CK(clk_gated), .Q(
        KeyArray_outS20ser[7]), .QN() );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3322), .CK(clk_gated), .Q(new_AGEMA_signal_2608), 
        .QN() );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S21reg_gff_1_SFF_0_n6), .CK(clk_gated), .Q(
        KeyArray_outS21ser[0]), .QN() );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3323), .CK(clk_gated), .Q(new_AGEMA_signal_2611), 
        .QN() );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S21reg_gff_1_SFF_1_n6), .CK(clk_gated), .Q(
        KeyArray_outS21ser[1]), .QN() );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3324), .CK(clk_gated), .Q(new_AGEMA_signal_2614), 
        .QN() );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S21reg_gff_1_SFF_2_n6), .CK(clk_gated), .Q(
        KeyArray_outS21ser[2]), .QN() );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3325), .CK(clk_gated), .Q(new_AGEMA_signal_2617), 
        .QN() );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S21reg_gff_1_SFF_3_n6), .CK(clk_gated), .Q(
        KeyArray_outS21ser[3]), .QN() );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3326), .CK(clk_gated), .Q(new_AGEMA_signal_2620), 
        .QN() );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S21reg_gff_1_SFF_4_n6), .CK(clk_gated), .Q(
        KeyArray_outS21ser[4]), .QN() );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3327), .CK(clk_gated), .Q(new_AGEMA_signal_2623), 
        .QN() );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S21reg_gff_1_SFF_5_n6), .CK(clk_gated), .Q(
        KeyArray_outS21ser[5]), .QN() );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3328), .CK(clk_gated), .Q(new_AGEMA_signal_2626), 
        .QN() );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S21reg_gff_1_SFF_6_n6), .CK(clk_gated), .Q(
        KeyArray_outS21ser[6]), .QN() );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3329), .CK(clk_gated), .Q(new_AGEMA_signal_2629), 
        .QN() );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S21reg_gff_1_SFF_7_n6), .CK(clk_gated), .Q(
        KeyArray_outS21ser[7]), .QN() );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3330), .CK(clk_gated), .Q(new_AGEMA_signal_2632), 
        .QN() );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S22reg_gff_1_SFF_0_n6), .CK(clk_gated), .Q(
        KeyArray_outS22ser[0]), .QN() );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3331), .CK(clk_gated), .Q(new_AGEMA_signal_2635), 
        .QN() );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S22reg_gff_1_SFF_1_n6), .CK(clk_gated), .Q(
        KeyArray_outS22ser[1]), .QN() );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3332), .CK(clk_gated), .Q(new_AGEMA_signal_2638), 
        .QN() );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S22reg_gff_1_SFF_2_n6), .CK(clk_gated), .Q(
        KeyArray_outS22ser[2]), .QN() );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3333), .CK(clk_gated), .Q(new_AGEMA_signal_2641), 
        .QN() );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S22reg_gff_1_SFF_3_n6), .CK(clk_gated), .Q(
        KeyArray_outS22ser[3]), .QN() );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3334), .CK(clk_gated), .Q(new_AGEMA_signal_2644), 
        .QN() );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S22reg_gff_1_SFF_4_n6), .CK(clk_gated), .Q(
        KeyArray_outS22ser[4]), .QN() );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3335), .CK(clk_gated), .Q(new_AGEMA_signal_2647), 
        .QN() );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S22reg_gff_1_SFF_5_n6), .CK(clk_gated), .Q(
        KeyArray_outS22ser[5]), .QN() );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3336), .CK(clk_gated), .Q(new_AGEMA_signal_2650), 
        .QN() );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S22reg_gff_1_SFF_6_n6), .CK(clk_gated), .Q(
        KeyArray_outS22ser[6]), .QN() );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3337), .CK(clk_gated), .Q(new_AGEMA_signal_2653), 
        .QN() );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S22reg_gff_1_SFF_7_n6), .CK(clk_gated), .Q(
        KeyArray_outS22ser[7]), .QN() );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3338), .CK(clk_gated), .Q(new_AGEMA_signal_2656), 
        .QN() );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S23reg_gff_1_SFF_0_n6), .CK(clk_gated), .Q(
        KeyArray_outS23ser[0]), .QN() );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3339), .CK(clk_gated), .Q(new_AGEMA_signal_2659), 
        .QN() );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S23reg_gff_1_SFF_1_n6), .CK(clk_gated), .Q(
        KeyArray_outS23ser[1]), .QN() );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3340), .CK(clk_gated), .Q(new_AGEMA_signal_2662), 
        .QN() );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S23reg_gff_1_SFF_2_n6), .CK(clk_gated), .Q(
        KeyArray_outS23ser[2]), .QN() );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3341), .CK(clk_gated), .Q(new_AGEMA_signal_2665), 
        .QN() );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S23reg_gff_1_SFF_3_n6), .CK(clk_gated), .Q(
        KeyArray_outS23ser[3]), .QN() );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3342), .CK(clk_gated), .Q(new_AGEMA_signal_2668), 
        .QN() );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S23reg_gff_1_SFF_4_n6), .CK(clk_gated), .Q(
        KeyArray_outS23ser[4]), .QN() );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3343), .CK(clk_gated), .Q(new_AGEMA_signal_2671), 
        .QN() );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S23reg_gff_1_SFF_5_n5), .CK(clk_gated), .Q(
        KeyArray_outS23ser[5]), .QN() );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3344), .CK(clk_gated), .Q(new_AGEMA_signal_2674), 
        .QN() );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S23reg_gff_1_SFF_6_n5), .CK(clk_gated), .Q(
        KeyArray_outS23ser[6]), .QN() );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3345), .CK(clk_gated), .Q(new_AGEMA_signal_2677), 
        .QN() );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S23reg_gff_1_SFF_7_n5), .CK(clk_gated), .Q(
        KeyArray_outS23ser[7]), .QN() );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3346), .CK(clk_gated), .Q(new_AGEMA_signal_2680), 
        .QN() );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S30reg_gff_1_SFF_0_n5), .CK(clk_gated), .Q(
        KeyArray_outS30ser[0]), .QN() );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3512), .CK(clk_gated), .Q(new_AGEMA_signal_2683), 
        .QN() );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S30reg_gff_1_SFF_1_n5), .CK(clk_gated), .Q(
        KeyArray_outS30ser[1]), .QN() );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3527), .CK(clk_gated), .Q(new_AGEMA_signal_2686), 
        .QN() );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S30reg_gff_1_SFF_2_n5), .CK(clk_gated), .Q(
        KeyArray_outS30ser[2]), .QN() );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3528), .CK(clk_gated), .Q(new_AGEMA_signal_2689), 
        .QN() );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S30reg_gff_1_SFF_3_n5), .CK(clk_gated), .Q(
        KeyArray_outS30ser[3]), .QN() );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3529), .CK(clk_gated), .Q(new_AGEMA_signal_2692), 
        .QN() );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S30reg_gff_1_SFF_4_n5), .CK(clk_gated), .Q(
        KeyArray_outS30ser[4]), .QN() );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3530), .CK(clk_gated), .Q(new_AGEMA_signal_2695), 
        .QN() );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S30reg_gff_1_SFF_5_n5), .CK(clk_gated), .Q(
        KeyArray_outS30ser[5]), .QN() );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3531), .CK(clk_gated), .Q(new_AGEMA_signal_2698), 
        .QN() );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S30reg_gff_1_SFF_6_n5), .CK(clk_gated), .Q(
        KeyArray_outS30ser[6]), .QN() );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3532), .CK(clk_gated), .Q(new_AGEMA_signal_2701), 
        .QN() );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S30reg_gff_1_SFF_7_n5), .CK(clk_gated), .Q(
        KeyArray_outS30ser[7]), .QN() );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3533), .CK(clk_gated), .Q(new_AGEMA_signal_2704), 
        .QN() );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S31reg_gff_1_SFF_0_n6), .CK(clk_gated), .Q(
        KeyArray_outS31ser[0]), .QN() );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3347), .CK(clk_gated), .Q(new_AGEMA_signal_2707), 
        .QN() );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S31reg_gff_1_SFF_1_n6), .CK(clk_gated), .Q(
        KeyArray_outS31ser[1]), .QN() );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3348), .CK(clk_gated), .Q(new_AGEMA_signal_2710), 
        .QN() );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S31reg_gff_1_SFF_2_n6), .CK(clk_gated), .Q(
        KeyArray_outS31ser[2]), .QN() );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3349), .CK(clk_gated), .Q(new_AGEMA_signal_2713), 
        .QN() );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S31reg_gff_1_SFF_3_n6), .CK(clk_gated), .Q(
        KeyArray_outS31ser[3]), .QN() );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3350), .CK(clk_gated), .Q(new_AGEMA_signal_2716), 
        .QN() );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S31reg_gff_1_SFF_4_n6), .CK(clk_gated), .Q(
        KeyArray_outS31ser[4]), .QN() );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3351), .CK(clk_gated), .Q(new_AGEMA_signal_2719), 
        .QN() );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S31reg_gff_1_SFF_5_n6), .CK(clk_gated), .Q(
        KeyArray_outS31ser[5]), .QN() );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3352), .CK(clk_gated), .Q(new_AGEMA_signal_2722), 
        .QN() );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S31reg_gff_1_SFF_6_n6), .CK(clk_gated), .Q(
        KeyArray_outS31ser[6]), .QN() );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3353), .CK(clk_gated), .Q(new_AGEMA_signal_2725), 
        .QN() );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S31reg_gff_1_SFF_7_n6), .CK(clk_gated), .Q(
        KeyArray_outS31ser[7]), .QN() );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3354), .CK(clk_gated), .Q(new_AGEMA_signal_2728), 
        .QN() );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S32reg_gff_1_SFF_0_n6), .CK(clk_gated), .Q(
        KeyArray_outS32ser[0]), .QN() );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3355), .CK(clk_gated), .Q(new_AGEMA_signal_2731), 
        .QN() );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S32reg_gff_1_SFF_1_n6), .CK(clk_gated), .Q(
        KeyArray_outS32ser[1]), .QN() );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3356), .CK(clk_gated), .Q(new_AGEMA_signal_2734), 
        .QN() );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S32reg_gff_1_SFF_2_n6), .CK(clk_gated), .Q(
        KeyArray_outS32ser[2]), .QN() );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3357), .CK(clk_gated), .Q(new_AGEMA_signal_2737), 
        .QN() );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S32reg_gff_1_SFF_3_n6), .CK(clk_gated), .Q(
        KeyArray_outS32ser[3]), .QN() );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3358), .CK(clk_gated), .Q(new_AGEMA_signal_2740), 
        .QN() );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S32reg_gff_1_SFF_4_n6), .CK(clk_gated), .Q(
        KeyArray_outS32ser[4]), .QN() );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3359), .CK(clk_gated), .Q(new_AGEMA_signal_2743), 
        .QN() );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S32reg_gff_1_SFF_5_n6), .CK(clk_gated), .Q(
        KeyArray_outS32ser[5]), .QN() );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3360), .CK(clk_gated), .Q(new_AGEMA_signal_2746), 
        .QN() );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S32reg_gff_1_SFF_6_n5), .CK(clk_gated), .Q(
        KeyArray_outS32ser[6]), .QN() );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3361), .CK(clk_gated), .Q(new_AGEMA_signal_2749), 
        .QN() );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S32reg_gff_1_SFF_7_n5), .CK(clk_gated), .Q(
        KeyArray_outS32ser[7]), .QN() );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3362), .CK(clk_gated), .Q(new_AGEMA_signal_2752), 
        .QN() );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S33reg_gff_1_SFF_0_n5), .CK(clk_gated), .Q(
        KeyArray_outS33ser[0]), .QN() );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_0_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3363), .CK(clk_gated), .Q(new_AGEMA_signal_2755), 
        .QN() );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S33reg_gff_1_SFF_1_n5), .CK(clk_gated), .Q(
        KeyArray_outS33ser[1]), .QN() );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_1_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3364), .CK(clk_gated), .Q(new_AGEMA_signal_2758), 
        .QN() );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S33reg_gff_1_SFF_2_n5), .CK(clk_gated), .Q(
        KeyArray_outS33ser[2]), .QN() );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_2_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3365), .CK(clk_gated), .Q(new_AGEMA_signal_2761), 
        .QN() );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S33reg_gff_1_SFF_3_n5), .CK(clk_gated), .Q(
        KeyArray_outS33ser[3]), .QN() );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_3_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3366), .CK(clk_gated), .Q(new_AGEMA_signal_2764), 
        .QN() );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S33reg_gff_1_SFF_4_n5), .CK(clk_gated), .Q(
        KeyArray_outS33ser[4]), .QN() );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_4_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3367), .CK(clk_gated), .Q(new_AGEMA_signal_2767), 
        .QN() );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S33reg_gff_1_SFF_5_n5), .CK(clk_gated), .Q(
        KeyArray_outS33ser[5]), .QN() );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_5_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3368), .CK(clk_gated), .Q(new_AGEMA_signal_2770), 
        .QN() );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S33reg_gff_1_SFF_6_n5), .CK(clk_gated), .Q(
        KeyArray_outS33ser[6]), .QN() );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_6_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3369), .CK(clk_gated), .Q(new_AGEMA_signal_2773), 
        .QN() );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_0_s_current_state_reg ( 
        .D(KeyArray_S33reg_gff_1_SFF_7_n5), .CK(clk_gated), .Q(
        KeyArray_outS33ser[7]), .QN() );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_7_Q_reg_FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3370), .CK(clk_gated), .Q(new_AGEMA_signal_2776), 
        .QN() );
endmodule

