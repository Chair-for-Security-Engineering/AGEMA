/* modified netlist. Source: module sbox in file Designs/AESSbox/optBP2/AGEMA/sbox.v */
/* 8 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 9 register stage(s) in total */

module sbox_HPC2_AIG_Pipeline_d4 (X_s0, clk, X_s1, X_s2, X_s3, X_s4, Fresh, Y_s0, Y_s1, Y_s2, Y_s3, Y_s4);
    input [7:0] X_s0 ;
    input clk ;
    input [7:0] X_s1 ;
    input [7:0] X_s2 ;
    input [7:0] X_s3 ;
    input [7:0] X_s4 ;
    input [339:0] Fresh ;
    output [7:0] Y_s0 ;
    output [7:0] Y_s1 ;
    output [7:0] Y_s2 ;
    output [7:0] Y_s3 ;
    output [7:0] Y_s4 ;
    wire signal_143 ;
    wire signal_144 ;
    wire signal_145 ;
    wire signal_146 ;
    wire signal_147 ;
    wire signal_148 ;
    wire signal_149 ;
    wire signal_150 ;
    wire signal_151 ;
    wire signal_152 ;
    wire signal_153 ;
    wire signal_154 ;
    wire signal_155 ;
    wire signal_156 ;
    wire signal_157 ;
    wire signal_158 ;
    wire signal_159 ;
    wire signal_160 ;
    wire signal_161 ;
    wire signal_162 ;
    wire signal_163 ;
    wire signal_164 ;
    wire signal_165 ;
    wire signal_166 ;
    wire signal_167 ;
    wire signal_168 ;
    wire signal_169 ;
    wire signal_170 ;
    wire signal_171 ;
    wire signal_172 ;
    wire signal_173 ;
    wire signal_174 ;
    wire signal_175 ;
    wire signal_176 ;
    wire signal_177 ;
    wire signal_178 ;
    wire signal_179 ;
    wire signal_180 ;
    wire signal_181 ;
    wire signal_182 ;
    wire signal_183 ;
    wire signal_184 ;
    wire signal_185 ;
    wire signal_186 ;
    wire signal_187 ;
    wire signal_188 ;
    wire signal_189 ;
    wire signal_190 ;
    wire signal_191 ;
    wire signal_192 ;
    wire signal_193 ;
    wire signal_194 ;
    wire signal_195 ;
    wire signal_196 ;
    wire signal_197 ;
    wire signal_198 ;
    wire signal_199 ;
    wire signal_200 ;
    wire signal_201 ;
    wire signal_202 ;
    wire signal_203 ;
    wire signal_204 ;
    wire signal_205 ;
    wire signal_206 ;
    wire signal_207 ;
    wire signal_208 ;
    wire signal_209 ;
    wire signal_210 ;
    wire signal_211 ;
    wire signal_212 ;
    wire signal_213 ;
    wire signal_214 ;
    wire signal_215 ;
    wire signal_216 ;
    wire signal_217 ;
    wire signal_218 ;
    wire signal_219 ;
    wire signal_220 ;
    wire signal_221 ;
    wire signal_222 ;
    wire signal_223 ;
    wire signal_224 ;
    wire signal_225 ;
    wire signal_226 ;
    wire signal_227 ;
    wire signal_228 ;
    wire signal_229 ;
    wire signal_230 ;
    wire signal_231 ;
    wire signal_232 ;
    wire signal_233 ;
    wire signal_234 ;
    wire signal_235 ;
    wire signal_236 ;
    wire signal_237 ;
    wire signal_238 ;
    wire signal_239 ;
    wire signal_240 ;
    wire signal_241 ;
    wire signal_242 ;
    wire signal_243 ;
    wire signal_244 ;
    wire signal_245 ;
    wire signal_246 ;
    wire signal_247 ;
    wire signal_248 ;
    wire signal_249 ;
    wire signal_250 ;
    wire signal_251 ;
    wire signal_252 ;
    wire signal_253 ;
    wire signal_254 ;
    wire signal_255 ;
    wire signal_256 ;
    wire signal_257 ;
    wire signal_258 ;
    wire signal_259 ;
    wire signal_260 ;
    wire signal_261 ;
    wire signal_262 ;
    wire signal_263 ;
    wire signal_264 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_285 ;
    wire signal_286 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_352 ;
    wire signal_353 ;
    wire signal_354 ;
    wire signal_355 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_359 ;
    wire signal_360 ;
    wire signal_361 ;
    wire signal_362 ;
    wire signal_363 ;
    wire signal_364 ;
    wire signal_365 ;
    wire signal_366 ;
    wire signal_367 ;
    wire signal_368 ;
    wire signal_369 ;
    wire signal_370 ;
    wire signal_371 ;
    wire signal_372 ;
    wire signal_373 ;
    wire signal_374 ;
    wire signal_375 ;
    wire signal_376 ;
    wire signal_377 ;
    wire signal_378 ;
    wire signal_379 ;
    wire signal_380 ;
    wire signal_381 ;
    wire signal_382 ;
    wire signal_383 ;
    wire signal_384 ;
    wire signal_385 ;
    wire signal_386 ;
    wire signal_387 ;
    wire signal_388 ;
    wire signal_389 ;
    wire signal_390 ;
    wire signal_391 ;
    wire signal_392 ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_415 ;
    wire signal_416 ;
    wire signal_417 ;
    wire signal_418 ;
    wire signal_419 ;
    wire signal_420 ;
    wire signal_421 ;
    wire signal_422 ;
    wire signal_423 ;
    wire signal_424 ;
    wire signal_425 ;
    wire signal_426 ;
    wire signal_427 ;
    wire signal_428 ;
    wire signal_429 ;
    wire signal_430 ;
    wire signal_431 ;
    wire signal_432 ;
    wire signal_433 ;
    wire signal_434 ;
    wire signal_435 ;
    wire signal_436 ;
    wire signal_437 ;
    wire signal_438 ;
    wire signal_439 ;
    wire signal_440 ;
    wire signal_441 ;
    wire signal_442 ;
    wire signal_443 ;
    wire signal_444 ;
    wire signal_445 ;
    wire signal_446 ;
    wire signal_447 ;
    wire signal_448 ;
    wire signal_449 ;
    wire signal_450 ;
    wire signal_451 ;
    wire signal_452 ;
    wire signal_453 ;
    wire signal_454 ;
    wire signal_455 ;
    wire signal_456 ;
    wire signal_457 ;
    wire signal_458 ;
    wire signal_459 ;
    wire signal_460 ;
    wire signal_461 ;
    wire signal_462 ;
    wire signal_463 ;
    wire signal_464 ;
    wire signal_465 ;
    wire signal_466 ;
    wire signal_467 ;
    wire signal_468 ;
    wire signal_469 ;
    wire signal_470 ;
    wire signal_471 ;
    wire signal_472 ;
    wire signal_473 ;
    wire signal_474 ;
    wire signal_475 ;
    wire signal_476 ;
    wire signal_477 ;
    wire signal_478 ;
    wire signal_479 ;
    wire signal_480 ;
    wire signal_481 ;
    wire signal_482 ;
    wire signal_483 ;
    wire signal_484 ;
    wire signal_485 ;
    wire signal_486 ;
    wire signal_487 ;
    wire signal_488 ;
    wire signal_489 ;
    wire signal_490 ;
    wire signal_491 ;
    wire signal_492 ;
    wire signal_493 ;
    wire signal_494 ;
    wire signal_495 ;
    wire signal_496 ;
    wire signal_497 ;
    wire signal_498 ;
    wire signal_499 ;
    wire signal_500 ;
    wire signal_501 ;
    wire signal_502 ;
    wire signal_503 ;
    wire signal_504 ;
    wire signal_505 ;
    wire signal_506 ;
    wire signal_507 ;
    wire signal_508 ;
    wire signal_509 ;
    wire signal_510 ;
    wire signal_511 ;
    wire signal_512 ;
    wire signal_513 ;
    wire signal_514 ;
    wire signal_515 ;
    wire signal_516 ;
    wire signal_517 ;
    wire signal_518 ;
    wire signal_519 ;
    wire signal_520 ;
    wire signal_521 ;
    wire signal_522 ;
    wire signal_523 ;
    wire signal_524 ;
    wire signal_525 ;
    wire signal_526 ;
    wire signal_527 ;
    wire signal_528 ;
    wire signal_529 ;
    wire signal_530 ;
    wire signal_531 ;
    wire signal_532 ;
    wire signal_533 ;
    wire signal_534 ;
    wire signal_535 ;
    wire signal_536 ;
    wire signal_537 ;
    wire signal_538 ;
    wire signal_539 ;
    wire signal_540 ;
    wire signal_541 ;
    wire signal_542 ;
    wire signal_543 ;
    wire signal_544 ;
    wire signal_545 ;
    wire signal_546 ;
    wire signal_547 ;
    wire signal_548 ;
    wire signal_549 ;
    wire signal_550 ;
    wire signal_551 ;
    wire signal_552 ;
    wire signal_553 ;
    wire signal_554 ;
    wire signal_555 ;
    wire signal_556 ;
    wire signal_557 ;
    wire signal_558 ;
    wire signal_559 ;
    wire signal_560 ;
    wire signal_561 ;
    wire signal_562 ;
    wire signal_563 ;
    wire signal_564 ;
    wire signal_565 ;
    wire signal_566 ;
    wire signal_567 ;
    wire signal_568 ;
    wire signal_569 ;
    wire signal_570 ;
    wire signal_571 ;
    wire signal_572 ;
    wire signal_573 ;
    wire signal_574 ;
    wire signal_575 ;
    wire signal_576 ;
    wire signal_577 ;
    wire signal_578 ;
    wire signal_579 ;
    wire signal_580 ;
    wire signal_581 ;
    wire signal_582 ;
    wire signal_583 ;
    wire signal_584 ;
    wire signal_585 ;
    wire signal_586 ;
    wire signal_587 ;
    wire signal_588 ;
    wire signal_589 ;
    wire signal_590 ;
    wire signal_591 ;
    wire signal_592 ;
    wire signal_593 ;
    wire signal_594 ;
    wire signal_595 ;
    wire signal_596 ;
    wire signal_597 ;
    wire signal_598 ;
    wire signal_599 ;
    wire signal_600 ;
    wire signal_601 ;
    wire signal_602 ;
    wire signal_603 ;
    wire signal_604 ;
    wire signal_605 ;
    wire signal_606 ;
    wire signal_607 ;
    wire signal_608 ;
    wire signal_609 ;
    wire signal_610 ;
    wire signal_611 ;
    wire signal_612 ;
    wire signal_613 ;
    wire signal_614 ;
    wire signal_615 ;
    wire signal_616 ;
    wire signal_617 ;
    wire signal_618 ;
    wire signal_619 ;
    wire signal_620 ;
    wire signal_621 ;
    wire signal_622 ;
    wire signal_623 ;
    wire signal_624 ;
    wire signal_625 ;
    wire signal_626 ;
    wire signal_627 ;
    wire signal_628 ;
    wire signal_629 ;
    wire signal_630 ;
    wire signal_631 ;
    wire signal_632 ;
    wire signal_633 ;
    wire signal_634 ;
    wire signal_635 ;
    wire signal_636 ;
    wire signal_637 ;
    wire signal_638 ;
    wire signal_639 ;
    wire signal_640 ;
    wire signal_641 ;
    wire signal_642 ;
    wire signal_643 ;
    wire signal_644 ;
    wire signal_645 ;
    wire signal_646 ;
    wire signal_647 ;
    wire signal_648 ;
    wire signal_649 ;
    wire signal_650 ;
    wire signal_651 ;
    wire signal_652 ;
    wire signal_653 ;
    wire signal_654 ;
    wire signal_655 ;
    wire signal_656 ;
    wire signal_657 ;
    wire signal_658 ;
    wire signal_659 ;
    wire signal_660 ;
    wire signal_661 ;
    wire signal_662 ;
    wire signal_663 ;
    wire signal_664 ;
    wire signal_665 ;
    wire signal_666 ;
    wire signal_667 ;
    wire signal_668 ;
    wire signal_669 ;
    wire signal_670 ;
    wire signal_671 ;
    wire signal_672 ;
    wire signal_673 ;
    wire signal_674 ;
    wire signal_675 ;
    wire signal_676 ;
    wire signal_677 ;
    wire signal_678 ;
    wire signal_679 ;
    wire signal_680 ;
    wire signal_681 ;
    wire signal_682 ;
    wire signal_683 ;
    wire signal_684 ;
    wire signal_685 ;
    wire signal_686 ;
    wire signal_687 ;
    wire signal_688 ;
    wire signal_689 ;
    wire signal_690 ;
    wire signal_691 ;
    wire signal_692 ;
    wire signal_693 ;
    wire signal_694 ;
    wire signal_695 ;
    wire signal_696 ;
    wire signal_697 ;
    wire signal_698 ;
    wire signal_699 ;
    wire signal_700 ;
    wire signal_701 ;
    wire signal_702 ;
    wire signal_703 ;
    wire signal_704 ;
    wire signal_705 ;
    wire signal_706 ;
    wire signal_707 ;
    wire signal_708 ;
    wire signal_709 ;
    wire signal_710 ;
    wire signal_711 ;
    wire signal_712 ;
    wire signal_713 ;
    wire signal_714 ;
    wire signal_715 ;
    wire signal_716 ;
    wire signal_717 ;
    wire signal_718 ;
    wire signal_719 ;
    wire signal_720 ;
    wire signal_721 ;
    wire signal_722 ;
    wire signal_723 ;
    wire signal_724 ;
    wire signal_725 ;
    wire signal_726 ;
    wire signal_727 ;
    wire signal_728 ;
    wire signal_729 ;
    wire signal_730 ;
    wire signal_731 ;
    wire signal_732 ;
    wire signal_733 ;
    wire signal_734 ;
    wire signal_735 ;
    wire signal_736 ;
    wire signal_737 ;
    wire signal_738 ;
    wire signal_739 ;
    wire signal_740 ;
    wire signal_741 ;
    wire signal_742 ;
    wire signal_743 ;
    wire signal_744 ;
    wire signal_745 ;
    wire signal_746 ;
    wire signal_747 ;
    wire signal_748 ;
    wire signal_749 ;
    wire signal_750 ;
    wire signal_751 ;
    wire signal_752 ;
    wire signal_753 ;
    wire signal_754 ;
    wire signal_755 ;
    wire signal_756 ;
    wire signal_757 ;
    wire signal_758 ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_768 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_771 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_774 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_777 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_780 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_783 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_786 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_789 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_792 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_809 ;
    wire signal_810 ;
    wire signal_811 ;
    wire signal_812 ;
    wire signal_813 ;
    wire signal_814 ;
    wire signal_815 ;
    wire signal_816 ;
    wire signal_817 ;
    wire signal_818 ;
    wire signal_819 ;
    wire signal_820 ;
    wire signal_821 ;
    wire signal_822 ;
    wire signal_823 ;
    wire signal_824 ;
    wire signal_825 ;
    wire signal_826 ;
    wire signal_827 ;
    wire signal_828 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_831 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_834 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1276 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1279 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1282 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1285 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1288 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1294 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1297 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1300 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1303 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1309 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1494 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1499 ;
    wire signal_1500 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1503 ;
    wire signal_1504 ;
    wire signal_1505 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1509 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1512 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1518 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1521 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1527 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1530 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1536 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1539 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1564 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1623 ;
    wire signal_1624 ;
    wire signal_1625 ;
    wire signal_1626 ;
    wire signal_1627 ;
    wire signal_1628 ;
    wire signal_1629 ;
    wire signal_1630 ;
    wire signal_1631 ;
    wire signal_1632 ;
    wire signal_1633 ;
    wire signal_1634 ;
    wire signal_1635 ;
    wire signal_1636 ;
    wire signal_1637 ;
    wire signal_1638 ;
    wire signal_1639 ;
    wire signal_1640 ;
    wire signal_1641 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1657 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1660 ;
    wire signal_1661 ;
    wire signal_1662 ;
    wire signal_1663 ;
    wire signal_1664 ;
    wire signal_1665 ;
    wire signal_1666 ;
    wire signal_1667 ;
    wire signal_1668 ;
    wire signal_1669 ;
    wire signal_1670 ;
    wire signal_1671 ;
    wire signal_1672 ;
    wire signal_1673 ;
    wire signal_1674 ;
    wire signal_1675 ;
    wire signal_1676 ;
    wire signal_1677 ;
    wire signal_1678 ;
    wire signal_1679 ;
    wire signal_1680 ;
    wire signal_1681 ;
    wire signal_1682 ;
    wire signal_1683 ;
    wire signal_1684 ;
    wire signal_1685 ;
    wire signal_1686 ;
    wire signal_1687 ;
    wire signal_1688 ;
    wire signal_1689 ;
    wire signal_1690 ;
    wire signal_1691 ;
    wire signal_1692 ;
    wire signal_1693 ;
    wire signal_1694 ;
    wire signal_1695 ;
    wire signal_1696 ;
    wire signal_1697 ;
    wire signal_1698 ;
    wire signal_1699 ;
    wire signal_1700 ;
    wire signal_1701 ;
    wire signal_1702 ;
    wire signal_1703 ;
    wire signal_1704 ;
    wire signal_1705 ;
    wire signal_1706 ;
    wire signal_1707 ;
    wire signal_1708 ;
    wire signal_1709 ;
    wire signal_1710 ;
    wire signal_1711 ;
    wire signal_1712 ;
    wire signal_1713 ;
    wire signal_1714 ;
    wire signal_1715 ;
    wire signal_1716 ;
    wire signal_1717 ;
    wire signal_1718 ;
    wire signal_1719 ;
    wire signal_1720 ;
    wire signal_1721 ;
    wire signal_1722 ;
    wire signal_1723 ;
    wire signal_1724 ;
    wire signal_1725 ;
    wire signal_1726 ;
    wire signal_1727 ;
    wire signal_1728 ;
    wire signal_1729 ;
    wire signal_1730 ;
    wire signal_1731 ;
    wire signal_1732 ;
    wire signal_1733 ;
    wire signal_1734 ;
    wire signal_1735 ;
    wire signal_1736 ;
    wire signal_1737 ;
    wire signal_1738 ;
    wire signal_1739 ;
    wire signal_1740 ;
    wire signal_1741 ;
    wire signal_1742 ;
    wire signal_1743 ;
    wire signal_1744 ;
    wire signal_1745 ;
    wire signal_1746 ;
    wire signal_1747 ;
    wire signal_1748 ;
    wire signal_1749 ;
    wire signal_1750 ;
    wire signal_1751 ;
    wire signal_1752 ;
    wire signal_1753 ;
    wire signal_1754 ;
    wire signal_1755 ;
    wire signal_1756 ;
    wire signal_1757 ;
    wire signal_1758 ;
    wire signal_1759 ;
    wire signal_1760 ;
    wire signal_1761 ;
    wire signal_1762 ;
    wire signal_1763 ;
    wire signal_1764 ;
    wire signal_1765 ;
    wire signal_1766 ;
    wire signal_1767 ;
    wire signal_1768 ;
    wire signal_1769 ;
    wire signal_1770 ;
    wire signal_1771 ;
    wire signal_1772 ;
    wire signal_1773 ;
    wire signal_1774 ;
    wire signal_1775 ;
    wire signal_1776 ;
    wire signal_1777 ;
    wire signal_1778 ;
    wire signal_1779 ;
    wire signal_1780 ;
    wire signal_1781 ;
    wire signal_1782 ;
    wire signal_1783 ;
    wire signal_1784 ;
    wire signal_1785 ;
    wire signal_1786 ;
    wire signal_1787 ;
    wire signal_1788 ;
    wire signal_1789 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1792 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1795 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1813 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1844 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1854 ;
    wire signal_1855 ;
    wire signal_1856 ;
    wire signal_1857 ;
    wire signal_1858 ;
    wire signal_1859 ;
    wire signal_1860 ;
    wire signal_1861 ;
    wire signal_1862 ;
    wire signal_1863 ;
    wire signal_1864 ;
    wire signal_1865 ;
    wire signal_1866 ;

    /* cells in depth 0 */
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_136 ( .a ({X_s4[7], X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .c ({signal_286, signal_285, signal_284, signal_283, signal_151}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_137 ( .a ({X_s4[7], X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .c ({signal_294, signal_293, signal_292, signal_291, signal_152}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_138 ( .a ({X_s4[7], X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .c ({signal_302, signal_301, signal_300, signal_299, signal_153}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_139 ( .a ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .c ({signal_306, signal_305, signal_304, signal_303, signal_154}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_140 ( .a ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .c ({signal_314, signal_313, signal_312, signal_311, signal_155}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_141 ( .a ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({X_s4[5], X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .c ({signal_326, signal_325, signal_324, signal_323, signal_156}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_142 ( .a ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .c ({signal_330, signal_329, signal_328, signal_327, signal_157}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_143 ( .a ({X_s4[5], X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .b ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .c ({signal_334, signal_333, signal_332, signal_331, signal_158}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_144 ( .a ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({X_s4[0], X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .c ({signal_342, signal_341, signal_340, signal_339, signal_159}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_145 ( .a ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({X_s4[0], X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .c ({signal_346, signal_345, signal_344, signal_343, signal_160}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_146 ( .a ({signal_286, signal_285, signal_284, signal_283, signal_151}), .b ({signal_314, signal_313, signal_312, signal_311, signal_155}), .c ({signal_350, signal_349, signal_348, signal_347, signal_161}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_147 ( .a ({X_s4[0], X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({signal_326, signal_325, signal_324, signal_323, signal_156}), .c ({signal_354, signal_353, signal_352, signal_351, signal_162}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_148 ( .a ({signal_302, signal_301, signal_300, signal_299, signal_153}), .b ({signal_306, signal_305, signal_304, signal_303, signal_154}), .c ({signal_358, signal_357, signal_356, signal_355, signal_163}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_149 ( .a ({signal_314, signal_313, signal_312, signal_311, signal_155}), .b ({signal_330, signal_329, signal_328, signal_327, signal_157}), .c ({signal_362, signal_361, signal_360, signal_359, signal_164}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_150 ( .a ({signal_314, signal_313, signal_312, signal_311, signal_155}), .b ({signal_334, signal_333, signal_332, signal_331, signal_158}), .c ({signal_366, signal_365, signal_364, signal_363, signal_165}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_151 ( .a ({signal_326, signal_325, signal_324, signal_323, signal_156}), .b ({signal_342, signal_341, signal_340, signal_339, signal_159}), .c ({signal_370, signal_369, signal_368, signal_367, signal_166}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_152 ( .a ({signal_326, signal_325, signal_324, signal_323, signal_156}), .b ({signal_346, signal_345, signal_344, signal_343, signal_160}), .c ({signal_374, signal_373, signal_372, signal_371, signal_167}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_153 ( .a ({signal_286, signal_285, signal_284, signal_283, signal_151}), .b ({signal_334, signal_333, signal_332, signal_331, signal_158}), .c ({signal_378, signal_377, signal_376, signal_375, signal_168}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_160 ( .a ({X_s4[0], X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({signal_350, signal_349, signal_348, signal_347, signal_161}), .c ({signal_406, signal_405, signal_404, signal_403, signal_175}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_161 ( .a ({signal_326, signal_325, signal_324, signal_323, signal_156}), .b ({signal_350, signal_349, signal_348, signal_347, signal_161}), .c ({signal_410, signal_409, signal_408, signal_407, signal_176}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_162 ( .a ({signal_330, signal_329, signal_328, signal_327, signal_157}), .b ({signal_350, signal_349, signal_348, signal_347, signal_161}), .c ({signal_414, signal_413, signal_412, signal_411, signal_177}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_163 ( .a ({signal_354, signal_353, signal_352, signal_351, signal_162}), .b ({signal_366, signal_365, signal_364, signal_363, signal_165}), .c ({signal_418, signal_417, signal_416, signal_415, signal_178}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_164 ( .a ({signal_286, signal_285, signal_284, signal_283, signal_151}), .b ({signal_370, signal_369, signal_368, signal_367, signal_166}), .c ({signal_422, signal_421, signal_420, signal_419, signal_179}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_165 ( .a ({signal_294, signal_293, signal_292, signal_291, signal_152}), .b ({signal_374, signal_373, signal_372, signal_371, signal_167}), .c ({signal_426, signal_425, signal_424, signal_423, signal_180}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_166 ( .a ({signal_302, signal_301, signal_300, signal_299, signal_153}), .b ({signal_366, signal_365, signal_364, signal_363, signal_165}), .c ({signal_430, signal_429, signal_428, signal_427, signal_181}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_170 ( .a ({signal_294, signal_293, signal_292, signal_291, signal_152}), .b ({signal_410, signal_409, signal_408, signal_407, signal_176}), .c ({signal_446, signal_445, signal_444, signal_443, signal_185}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_171 ( .a ({signal_418, signal_417, signal_416, signal_415, signal_178}), .b ({signal_422, signal_421, signal_420, signal_419, signal_179}), .c ({signal_450, signal_449, signal_448, signal_447, signal_186}) ) ;

    /* cells in depth 1 */
    buf_clk cell_268 ( .C (clk), .D (signal_177), .Q (signal_1207) ) ;
    buf_clk cell_270 ( .C (clk), .D (signal_411), .Q (signal_1209) ) ;
    buf_clk cell_272 ( .C (clk), .D (signal_412), .Q (signal_1211) ) ;
    buf_clk cell_274 ( .C (clk), .D (signal_413), .Q (signal_1213) ) ;
    buf_clk cell_276 ( .C (clk), .D (signal_414), .Q (signal_1215) ) ;
    buf_clk cell_278 ( .C (clk), .D (signal_181), .Q (signal_1217) ) ;
    buf_clk cell_280 ( .C (clk), .D (signal_427), .Q (signal_1219) ) ;
    buf_clk cell_282 ( .C (clk), .D (signal_428), .Q (signal_1221) ) ;
    buf_clk cell_284 ( .C (clk), .D (signal_429), .Q (signal_1223) ) ;
    buf_clk cell_286 ( .C (clk), .D (signal_430), .Q (signal_1225) ) ;
    buf_clk cell_288 ( .C (clk), .D (signal_185), .Q (signal_1227) ) ;
    buf_clk cell_290 ( .C (clk), .D (signal_443), .Q (signal_1229) ) ;
    buf_clk cell_292 ( .C (clk), .D (signal_444), .Q (signal_1231) ) ;
    buf_clk cell_294 ( .C (clk), .D (signal_445), .Q (signal_1233) ) ;
    buf_clk cell_296 ( .C (clk), .D (signal_446), .Q (signal_1235) ) ;
    buf_clk cell_298 ( .C (clk), .D (signal_186), .Q (signal_1237) ) ;
    buf_clk cell_300 ( .C (clk), .D (signal_447), .Q (signal_1239) ) ;
    buf_clk cell_302 ( .C (clk), .D (signal_448), .Q (signal_1241) ) ;
    buf_clk cell_304 ( .C (clk), .D (signal_449), .Q (signal_1243) ) ;
    buf_clk cell_306 ( .C (clk), .D (signal_450), .Q (signal_1245) ) ;
    buf_clk cell_388 ( .C (clk), .D (signal_175), .Q (signal_1327) ) ;
    buf_clk cell_394 ( .C (clk), .D (signal_403), .Q (signal_1333) ) ;
    buf_clk cell_400 ( .C (clk), .D (signal_404), .Q (signal_1339) ) ;
    buf_clk cell_406 ( .C (clk), .D (signal_405), .Q (signal_1345) ) ;
    buf_clk cell_412 ( .C (clk), .D (signal_406), .Q (signal_1351) ) ;
    buf_clk cell_418 ( .C (clk), .D (X_s0[0]), .Q (signal_1357) ) ;
    buf_clk cell_424 ( .C (clk), .D (X_s1[0]), .Q (signal_1363) ) ;
    buf_clk cell_430 ( .C (clk), .D (X_s2[0]), .Q (signal_1369) ) ;
    buf_clk cell_436 ( .C (clk), .D (X_s3[0]), .Q (signal_1375) ) ;
    buf_clk cell_442 ( .C (clk), .D (X_s4[0]), .Q (signal_1381) ) ;
    buf_clk cell_448 ( .C (clk), .D (signal_162), .Q (signal_1387) ) ;
    buf_clk cell_454 ( .C (clk), .D (signal_351), .Q (signal_1393) ) ;
    buf_clk cell_460 ( .C (clk), .D (signal_352), .Q (signal_1399) ) ;
    buf_clk cell_466 ( .C (clk), .D (signal_353), .Q (signal_1405) ) ;
    buf_clk cell_472 ( .C (clk), .D (signal_354), .Q (signal_1411) ) ;
    buf_clk cell_478 ( .C (clk), .D (signal_178), .Q (signal_1417) ) ;
    buf_clk cell_484 ( .C (clk), .D (signal_415), .Q (signal_1423) ) ;
    buf_clk cell_490 ( .C (clk), .D (signal_416), .Q (signal_1429) ) ;
    buf_clk cell_496 ( .C (clk), .D (signal_417), .Q (signal_1435) ) ;
    buf_clk cell_502 ( .C (clk), .D (signal_418), .Q (signal_1441) ) ;
    buf_clk cell_508 ( .C (clk), .D (signal_180), .Q (signal_1447) ) ;
    buf_clk cell_514 ( .C (clk), .D (signal_423), .Q (signal_1453) ) ;
    buf_clk cell_520 ( .C (clk), .D (signal_424), .Q (signal_1459) ) ;
    buf_clk cell_526 ( .C (clk), .D (signal_425), .Q (signal_1465) ) ;
    buf_clk cell_532 ( .C (clk), .D (signal_426), .Q (signal_1471) ) ;
    buf_clk cell_538 ( .C (clk), .D (signal_166), .Q (signal_1477) ) ;
    buf_clk cell_544 ( .C (clk), .D (signal_367), .Q (signal_1483) ) ;
    buf_clk cell_550 ( .C (clk), .D (signal_368), .Q (signal_1489) ) ;
    buf_clk cell_556 ( .C (clk), .D (signal_369), .Q (signal_1495) ) ;
    buf_clk cell_562 ( .C (clk), .D (signal_370), .Q (signal_1501) ) ;
    buf_clk cell_568 ( .C (clk), .D (signal_167), .Q (signal_1507) ) ;
    buf_clk cell_574 ( .C (clk), .D (signal_371), .Q (signal_1513) ) ;
    buf_clk cell_580 ( .C (clk), .D (signal_372), .Q (signal_1519) ) ;
    buf_clk cell_586 ( .C (clk), .D (signal_373), .Q (signal_1525) ) ;
    buf_clk cell_592 ( .C (clk), .D (signal_374), .Q (signal_1531) ) ;
    buf_clk cell_598 ( .C (clk), .D (signal_179), .Q (signal_1537) ) ;
    buf_clk cell_604 ( .C (clk), .D (signal_419), .Q (signal_1543) ) ;
    buf_clk cell_610 ( .C (clk), .D (signal_420), .Q (signal_1549) ) ;
    buf_clk cell_616 ( .C (clk), .D (signal_421), .Q (signal_1555) ) ;
    buf_clk cell_622 ( .C (clk), .D (signal_422), .Q (signal_1561) ) ;
    buf_clk cell_628 ( .C (clk), .D (signal_161), .Q (signal_1567) ) ;
    buf_clk cell_634 ( .C (clk), .D (signal_347), .Q (signal_1573) ) ;
    buf_clk cell_640 ( .C (clk), .D (signal_348), .Q (signal_1579) ) ;
    buf_clk cell_646 ( .C (clk), .D (signal_349), .Q (signal_1585) ) ;
    buf_clk cell_652 ( .C (clk), .D (signal_350), .Q (signal_1591) ) ;
    buf_clk cell_658 ( .C (clk), .D (signal_165), .Q (signal_1597) ) ;
    buf_clk cell_664 ( .C (clk), .D (signal_363), .Q (signal_1603) ) ;
    buf_clk cell_670 ( .C (clk), .D (signal_364), .Q (signal_1609) ) ;
    buf_clk cell_676 ( .C (clk), .D (signal_365), .Q (signal_1615) ) ;
    buf_clk cell_682 ( .C (clk), .D (signal_366), .Q (signal_1621) ) ;
    buf_clk cell_688 ( .C (clk), .D (signal_164), .Q (signal_1627) ) ;
    buf_clk cell_694 ( .C (clk), .D (signal_359), .Q (signal_1633) ) ;
    buf_clk cell_700 ( .C (clk), .D (signal_360), .Q (signal_1639) ) ;
    buf_clk cell_706 ( .C (clk), .D (signal_361), .Q (signal_1645) ) ;
    buf_clk cell_712 ( .C (clk), .D (signal_362), .Q (signal_1651) ) ;
    buf_clk cell_718 ( .C (clk), .D (signal_176), .Q (signal_1657) ) ;
    buf_clk cell_724 ( .C (clk), .D (signal_407), .Q (signal_1663) ) ;
    buf_clk cell_730 ( .C (clk), .D (signal_408), .Q (signal_1669) ) ;
    buf_clk cell_736 ( .C (clk), .D (signal_409), .Q (signal_1675) ) ;
    buf_clk cell_742 ( .C (clk), .D (signal_410), .Q (signal_1681) ) ;
    buf_clk cell_748 ( .C (clk), .D (signal_163), .Q (signal_1687) ) ;
    buf_clk cell_754 ( .C (clk), .D (signal_355), .Q (signal_1693) ) ;
    buf_clk cell_760 ( .C (clk), .D (signal_356), .Q (signal_1699) ) ;
    buf_clk cell_766 ( .C (clk), .D (signal_357), .Q (signal_1705) ) ;
    buf_clk cell_772 ( .C (clk), .D (signal_358), .Q (signal_1711) ) ;
    buf_clk cell_778 ( .C (clk), .D (signal_153), .Q (signal_1717) ) ;
    buf_clk cell_784 ( .C (clk), .D (signal_299), .Q (signal_1723) ) ;
    buf_clk cell_790 ( .C (clk), .D (signal_300), .Q (signal_1729) ) ;
    buf_clk cell_796 ( .C (clk), .D (signal_301), .Q (signal_1735) ) ;
    buf_clk cell_802 ( .C (clk), .D (signal_302), .Q (signal_1741) ) ;
    buf_clk cell_808 ( .C (clk), .D (signal_151), .Q (signal_1747) ) ;
    buf_clk cell_814 ( .C (clk), .D (signal_283), .Q (signal_1753) ) ;
    buf_clk cell_820 ( .C (clk), .D (signal_284), .Q (signal_1759) ) ;
    buf_clk cell_826 ( .C (clk), .D (signal_285), .Q (signal_1765) ) ;
    buf_clk cell_832 ( .C (clk), .D (signal_286), .Q (signal_1771) ) ;
    buf_clk cell_838 ( .C (clk), .D (signal_152), .Q (signal_1777) ) ;
    buf_clk cell_844 ( .C (clk), .D (signal_291), .Q (signal_1783) ) ;
    buf_clk cell_850 ( .C (clk), .D (signal_292), .Q (signal_1789) ) ;
    buf_clk cell_856 ( .C (clk), .D (signal_293), .Q (signal_1795) ) ;
    buf_clk cell_862 ( .C (clk), .D (signal_294), .Q (signal_1801) ) ;
    buf_clk cell_868 ( .C (clk), .D (signal_168), .Q (signal_1807) ) ;
    buf_clk cell_874 ( .C (clk), .D (signal_375), .Q (signal_1813) ) ;
    buf_clk cell_880 ( .C (clk), .D (signal_376), .Q (signal_1819) ) ;
    buf_clk cell_886 ( .C (clk), .D (signal_377), .Q (signal_1825) ) ;
    buf_clk cell_892 ( .C (clk), .D (signal_378), .Q (signal_1831) ) ;
    buf_clk cell_898 ( .C (clk), .D (signal_154), .Q (signal_1837) ) ;
    buf_clk cell_904 ( .C (clk), .D (signal_303), .Q (signal_1843) ) ;
    buf_clk cell_910 ( .C (clk), .D (signal_304), .Q (signal_1849) ) ;
    buf_clk cell_916 ( .C (clk), .D (signal_305), .Q (signal_1855) ) ;
    buf_clk cell_922 ( .C (clk), .D (signal_306), .Q (signal_1861) ) ;

    /* cells in depth 2 */
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_154 ( .a ({signal_350, signal_349, signal_348, signal_347, signal_161}), .b ({signal_358, signal_357, signal_356, signal_355, signal_163}), .clk (clk), .r ({Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({signal_382, signal_381, signal_380, signal_379, signal_169}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_155 ( .a ({X_s4[0], X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({signal_370, signal_369, signal_368, signal_367, signal_166}), .clk (clk), .r ({Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10]}), .c ({signal_386, signal_385, signal_384, signal_383, signal_170}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_156 ( .a ({signal_302, signal_301, signal_300, signal_299, signal_153}), .b ({signal_366, signal_365, signal_364, signal_363, signal_165}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20]}), .c ({signal_390, signal_389, signal_388, signal_387, signal_171}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_157 ( .a ({signal_354, signal_353, signal_352, signal_351, signal_162}), .b ({signal_374, signal_373, signal_372, signal_371, signal_167}), .clk (clk), .r ({Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({signal_394, signal_393, signal_392, signal_391, signal_172}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_158 ( .a ({signal_286, signal_285, signal_284, signal_283, signal_151}), .b ({signal_362, signal_361, signal_360, signal_359, signal_164}), .clk (clk), .r ({Fresh[49], Fresh[48], Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40]}), .c ({signal_398, signal_397, signal_396, signal_395, signal_173}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_159 ( .a ({signal_306, signal_305, signal_304, signal_303, signal_154}), .b ({signal_378, signal_377, signal_376, signal_375, signal_168}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50]}), .c ({signal_402, signal_401, signal_400, signal_399, signal_174}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_167 ( .a ({signal_406, signal_405, signal_404, signal_403, signal_175}), .b ({signal_426, signal_425, signal_424, signal_423, signal_180}), .clk (clk), .r ({Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({signal_434, signal_433, signal_432, signal_431, signal_182}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_168 ( .a ({signal_418, signal_417, signal_416, signal_415, signal_178}), .b ({signal_422, signal_421, signal_420, signal_419, signal_179}), .clk (clk), .r ({Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72], Fresh[71], Fresh[70]}), .c ({signal_438, signal_437, signal_436, signal_435, signal_183}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_169 ( .a ({signal_294, signal_293, signal_292, signal_291, signal_152}), .b ({signal_410, signal_409, signal_408, signal_407, signal_176}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84], Fresh[83], Fresh[82], Fresh[81], Fresh[80]}), .c ({signal_442, signal_441, signal_440, signal_439, signal_184}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_172 ( .a ({signal_1216, signal_1214, signal_1212, signal_1210, signal_1208}), .b ({signal_382, signal_381, signal_380, signal_379, signal_169}), .c ({signal_454, signal_453, signal_452, signal_451, signal_187}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_173 ( .a ({signal_382, signal_381, signal_380, signal_379, signal_169}), .b ({signal_386, signal_385, signal_384, signal_383, signal_170}), .c ({signal_458, signal_457, signal_456, signal_455, signal_188}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_174 ( .a ({signal_1226, signal_1224, signal_1222, signal_1220, signal_1218}), .b ({signal_390, signal_389, signal_388, signal_387, signal_171}), .c ({signal_462, signal_461, signal_460, signal_459, signal_189}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_175 ( .a ({signal_398, signal_397, signal_396, signal_395, signal_173}), .b ({signal_402, signal_401, signal_400, signal_399, signal_174}), .c ({signal_466, signal_465, signal_464, signal_463, signal_190}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_176 ( .a ({signal_390, signal_389, signal_388, signal_387, signal_171}), .b ({signal_438, signal_437, signal_436, signal_435, signal_183}), .c ({signal_470, signal_469, signal_468, signal_467, signal_191}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_177 ( .a ({signal_398, signal_397, signal_396, signal_395, signal_173}), .b ({signal_442, signal_441, signal_440, signal_439, signal_184}), .c ({signal_474, signal_473, signal_472, signal_471, signal_192}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_178 ( .a ({signal_434, signal_433, signal_432, signal_431, signal_182}), .b ({signal_454, signal_453, signal_452, signal_451, signal_187}), .c ({signal_478, signal_477, signal_476, signal_475, signal_193}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_179 ( .a ({signal_1236, signal_1234, signal_1232, signal_1230, signal_1228}), .b ({signal_458, signal_457, signal_456, signal_455, signal_188}), .c ({signal_482, signal_481, signal_480, signal_479, signal_194}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_180 ( .a ({signal_394, signal_393, signal_392, signal_391, signal_172}), .b ({signal_462, signal_461, signal_460, signal_459, signal_189}), .c ({signal_486, signal_485, signal_484, signal_483, signal_195}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_181 ( .a ({signal_470, signal_469, signal_468, signal_467, signal_191}), .b ({signal_474, signal_473, signal_472, signal_471, signal_192}), .c ({signal_490, signal_489, signal_488, signal_487, signal_196}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_182 ( .a ({signal_466, signal_465, signal_464, signal_463, signal_190}), .b ({signal_478, signal_477, signal_476, signal_475, signal_193}), .c ({signal_494, signal_493, signal_492, signal_491, signal_197}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_183 ( .a ({signal_474, signal_473, signal_472, signal_471, signal_192}), .b ({signal_482, signal_481, signal_480, signal_479, signal_194}), .c ({signal_498, signal_497, signal_496, signal_495, signal_198}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_184 ( .a ({signal_466, signal_465, signal_464, signal_463, signal_190}), .b ({signal_486, signal_485, signal_484, signal_483, signal_195}), .c ({signal_502, signal_501, signal_500, signal_499, signal_199}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_187 ( .a ({signal_1246, signal_1244, signal_1242, signal_1240, signal_1238}), .b ({signal_490, signal_489, signal_488, signal_487, signal_196}), .c ({signal_514, signal_513, signal_512, signal_511, signal_202}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_188 ( .a ({signal_494, signal_493, signal_492, signal_491, signal_197}), .b ({signal_498, signal_497, signal_496, signal_495, signal_198}), .c ({signal_518, signal_517, signal_516, signal_515, signal_203}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_190 ( .a ({signal_502, signal_501, signal_500, signal_499, signal_199}), .b ({signal_514, signal_513, signal_512, signal_511, signal_202}), .c ({signal_526, signal_525, signal_524, signal_523, signal_205}) ) ;
    buf_clk cell_269 ( .C (clk), .D (signal_1207), .Q (signal_1208) ) ;
    buf_clk cell_271 ( .C (clk), .D (signal_1209), .Q (signal_1210) ) ;
    buf_clk cell_273 ( .C (clk), .D (signal_1211), .Q (signal_1212) ) ;
    buf_clk cell_275 ( .C (clk), .D (signal_1213), .Q (signal_1214) ) ;
    buf_clk cell_277 ( .C (clk), .D (signal_1215), .Q (signal_1216) ) ;
    buf_clk cell_279 ( .C (clk), .D (signal_1217), .Q (signal_1218) ) ;
    buf_clk cell_281 ( .C (clk), .D (signal_1219), .Q (signal_1220) ) ;
    buf_clk cell_283 ( .C (clk), .D (signal_1221), .Q (signal_1222) ) ;
    buf_clk cell_285 ( .C (clk), .D (signal_1223), .Q (signal_1224) ) ;
    buf_clk cell_287 ( .C (clk), .D (signal_1225), .Q (signal_1226) ) ;
    buf_clk cell_289 ( .C (clk), .D (signal_1227), .Q (signal_1228) ) ;
    buf_clk cell_291 ( .C (clk), .D (signal_1229), .Q (signal_1230) ) ;
    buf_clk cell_293 ( .C (clk), .D (signal_1231), .Q (signal_1232) ) ;
    buf_clk cell_295 ( .C (clk), .D (signal_1233), .Q (signal_1234) ) ;
    buf_clk cell_297 ( .C (clk), .D (signal_1235), .Q (signal_1236) ) ;
    buf_clk cell_299 ( .C (clk), .D (signal_1237), .Q (signal_1238) ) ;
    buf_clk cell_301 ( .C (clk), .D (signal_1239), .Q (signal_1240) ) ;
    buf_clk cell_303 ( .C (clk), .D (signal_1241), .Q (signal_1242) ) ;
    buf_clk cell_305 ( .C (clk), .D (signal_1243), .Q (signal_1244) ) ;
    buf_clk cell_307 ( .C (clk), .D (signal_1245), .Q (signal_1246) ) ;
    buf_clk cell_389 ( .C (clk), .D (signal_1327), .Q (signal_1328) ) ;
    buf_clk cell_395 ( .C (clk), .D (signal_1333), .Q (signal_1334) ) ;
    buf_clk cell_401 ( .C (clk), .D (signal_1339), .Q (signal_1340) ) ;
    buf_clk cell_407 ( .C (clk), .D (signal_1345), .Q (signal_1346) ) ;
    buf_clk cell_413 ( .C (clk), .D (signal_1351), .Q (signal_1352) ) ;
    buf_clk cell_419 ( .C (clk), .D (signal_1357), .Q (signal_1358) ) ;
    buf_clk cell_425 ( .C (clk), .D (signal_1363), .Q (signal_1364) ) ;
    buf_clk cell_431 ( .C (clk), .D (signal_1369), .Q (signal_1370) ) ;
    buf_clk cell_437 ( .C (clk), .D (signal_1375), .Q (signal_1376) ) ;
    buf_clk cell_443 ( .C (clk), .D (signal_1381), .Q (signal_1382) ) ;
    buf_clk cell_449 ( .C (clk), .D (signal_1387), .Q (signal_1388) ) ;
    buf_clk cell_455 ( .C (clk), .D (signal_1393), .Q (signal_1394) ) ;
    buf_clk cell_461 ( .C (clk), .D (signal_1399), .Q (signal_1400) ) ;
    buf_clk cell_467 ( .C (clk), .D (signal_1405), .Q (signal_1406) ) ;
    buf_clk cell_473 ( .C (clk), .D (signal_1411), .Q (signal_1412) ) ;
    buf_clk cell_479 ( .C (clk), .D (signal_1417), .Q (signal_1418) ) ;
    buf_clk cell_485 ( .C (clk), .D (signal_1423), .Q (signal_1424) ) ;
    buf_clk cell_491 ( .C (clk), .D (signal_1429), .Q (signal_1430) ) ;
    buf_clk cell_497 ( .C (clk), .D (signal_1435), .Q (signal_1436) ) ;
    buf_clk cell_503 ( .C (clk), .D (signal_1441), .Q (signal_1442) ) ;
    buf_clk cell_509 ( .C (clk), .D (signal_1447), .Q (signal_1448) ) ;
    buf_clk cell_515 ( .C (clk), .D (signal_1453), .Q (signal_1454) ) ;
    buf_clk cell_521 ( .C (clk), .D (signal_1459), .Q (signal_1460) ) ;
    buf_clk cell_527 ( .C (clk), .D (signal_1465), .Q (signal_1466) ) ;
    buf_clk cell_533 ( .C (clk), .D (signal_1471), .Q (signal_1472) ) ;
    buf_clk cell_539 ( .C (clk), .D (signal_1477), .Q (signal_1478) ) ;
    buf_clk cell_545 ( .C (clk), .D (signal_1483), .Q (signal_1484) ) ;
    buf_clk cell_551 ( .C (clk), .D (signal_1489), .Q (signal_1490) ) ;
    buf_clk cell_557 ( .C (clk), .D (signal_1495), .Q (signal_1496) ) ;
    buf_clk cell_563 ( .C (clk), .D (signal_1501), .Q (signal_1502) ) ;
    buf_clk cell_569 ( .C (clk), .D (signal_1507), .Q (signal_1508) ) ;
    buf_clk cell_575 ( .C (clk), .D (signal_1513), .Q (signal_1514) ) ;
    buf_clk cell_581 ( .C (clk), .D (signal_1519), .Q (signal_1520) ) ;
    buf_clk cell_587 ( .C (clk), .D (signal_1525), .Q (signal_1526) ) ;
    buf_clk cell_593 ( .C (clk), .D (signal_1531), .Q (signal_1532) ) ;
    buf_clk cell_599 ( .C (clk), .D (signal_1537), .Q (signal_1538) ) ;
    buf_clk cell_605 ( .C (clk), .D (signal_1543), .Q (signal_1544) ) ;
    buf_clk cell_611 ( .C (clk), .D (signal_1549), .Q (signal_1550) ) ;
    buf_clk cell_617 ( .C (clk), .D (signal_1555), .Q (signal_1556) ) ;
    buf_clk cell_623 ( .C (clk), .D (signal_1561), .Q (signal_1562) ) ;
    buf_clk cell_629 ( .C (clk), .D (signal_1567), .Q (signal_1568) ) ;
    buf_clk cell_635 ( .C (clk), .D (signal_1573), .Q (signal_1574) ) ;
    buf_clk cell_641 ( .C (clk), .D (signal_1579), .Q (signal_1580) ) ;
    buf_clk cell_647 ( .C (clk), .D (signal_1585), .Q (signal_1586) ) ;
    buf_clk cell_653 ( .C (clk), .D (signal_1591), .Q (signal_1592) ) ;
    buf_clk cell_659 ( .C (clk), .D (signal_1597), .Q (signal_1598) ) ;
    buf_clk cell_665 ( .C (clk), .D (signal_1603), .Q (signal_1604) ) ;
    buf_clk cell_671 ( .C (clk), .D (signal_1609), .Q (signal_1610) ) ;
    buf_clk cell_677 ( .C (clk), .D (signal_1615), .Q (signal_1616) ) ;
    buf_clk cell_683 ( .C (clk), .D (signal_1621), .Q (signal_1622) ) ;
    buf_clk cell_689 ( .C (clk), .D (signal_1627), .Q (signal_1628) ) ;
    buf_clk cell_695 ( .C (clk), .D (signal_1633), .Q (signal_1634) ) ;
    buf_clk cell_701 ( .C (clk), .D (signal_1639), .Q (signal_1640) ) ;
    buf_clk cell_707 ( .C (clk), .D (signal_1645), .Q (signal_1646) ) ;
    buf_clk cell_713 ( .C (clk), .D (signal_1651), .Q (signal_1652) ) ;
    buf_clk cell_719 ( .C (clk), .D (signal_1657), .Q (signal_1658) ) ;
    buf_clk cell_725 ( .C (clk), .D (signal_1663), .Q (signal_1664) ) ;
    buf_clk cell_731 ( .C (clk), .D (signal_1669), .Q (signal_1670) ) ;
    buf_clk cell_737 ( .C (clk), .D (signal_1675), .Q (signal_1676) ) ;
    buf_clk cell_743 ( .C (clk), .D (signal_1681), .Q (signal_1682) ) ;
    buf_clk cell_749 ( .C (clk), .D (signal_1687), .Q (signal_1688) ) ;
    buf_clk cell_755 ( .C (clk), .D (signal_1693), .Q (signal_1694) ) ;
    buf_clk cell_761 ( .C (clk), .D (signal_1699), .Q (signal_1700) ) ;
    buf_clk cell_767 ( .C (clk), .D (signal_1705), .Q (signal_1706) ) ;
    buf_clk cell_773 ( .C (clk), .D (signal_1711), .Q (signal_1712) ) ;
    buf_clk cell_779 ( .C (clk), .D (signal_1717), .Q (signal_1718) ) ;
    buf_clk cell_785 ( .C (clk), .D (signal_1723), .Q (signal_1724) ) ;
    buf_clk cell_791 ( .C (clk), .D (signal_1729), .Q (signal_1730) ) ;
    buf_clk cell_797 ( .C (clk), .D (signal_1735), .Q (signal_1736) ) ;
    buf_clk cell_803 ( .C (clk), .D (signal_1741), .Q (signal_1742) ) ;
    buf_clk cell_809 ( .C (clk), .D (signal_1747), .Q (signal_1748) ) ;
    buf_clk cell_815 ( .C (clk), .D (signal_1753), .Q (signal_1754) ) ;
    buf_clk cell_821 ( .C (clk), .D (signal_1759), .Q (signal_1760) ) ;
    buf_clk cell_827 ( .C (clk), .D (signal_1765), .Q (signal_1766) ) ;
    buf_clk cell_833 ( .C (clk), .D (signal_1771), .Q (signal_1772) ) ;
    buf_clk cell_839 ( .C (clk), .D (signal_1777), .Q (signal_1778) ) ;
    buf_clk cell_845 ( .C (clk), .D (signal_1783), .Q (signal_1784) ) ;
    buf_clk cell_851 ( .C (clk), .D (signal_1789), .Q (signal_1790) ) ;
    buf_clk cell_857 ( .C (clk), .D (signal_1795), .Q (signal_1796) ) ;
    buf_clk cell_863 ( .C (clk), .D (signal_1801), .Q (signal_1802) ) ;
    buf_clk cell_869 ( .C (clk), .D (signal_1807), .Q (signal_1808) ) ;
    buf_clk cell_875 ( .C (clk), .D (signal_1813), .Q (signal_1814) ) ;
    buf_clk cell_881 ( .C (clk), .D (signal_1819), .Q (signal_1820) ) ;
    buf_clk cell_887 ( .C (clk), .D (signal_1825), .Q (signal_1826) ) ;
    buf_clk cell_893 ( .C (clk), .D (signal_1831), .Q (signal_1832) ) ;
    buf_clk cell_899 ( .C (clk), .D (signal_1837), .Q (signal_1838) ) ;
    buf_clk cell_905 ( .C (clk), .D (signal_1843), .Q (signal_1844) ) ;
    buf_clk cell_911 ( .C (clk), .D (signal_1849), .Q (signal_1850) ) ;
    buf_clk cell_917 ( .C (clk), .D (signal_1855), .Q (signal_1856) ) ;
    buf_clk cell_923 ( .C (clk), .D (signal_1861), .Q (signal_1862) ) ;

    /* cells in depth 3 */
    buf_clk cell_308 ( .C (clk), .D (signal_198), .Q (signal_1247) ) ;
    buf_clk cell_310 ( .C (clk), .D (signal_495), .Q (signal_1249) ) ;
    buf_clk cell_312 ( .C (clk), .D (signal_496), .Q (signal_1251) ) ;
    buf_clk cell_314 ( .C (clk), .D (signal_497), .Q (signal_1253) ) ;
    buf_clk cell_316 ( .C (clk), .D (signal_498), .Q (signal_1255) ) ;
    buf_clk cell_318 ( .C (clk), .D (signal_202), .Q (signal_1257) ) ;
    buf_clk cell_320 ( .C (clk), .D (signal_511), .Q (signal_1259) ) ;
    buf_clk cell_322 ( .C (clk), .D (signal_512), .Q (signal_1261) ) ;
    buf_clk cell_324 ( .C (clk), .D (signal_513), .Q (signal_1263) ) ;
    buf_clk cell_326 ( .C (clk), .D (signal_514), .Q (signal_1265) ) ;
    buf_clk cell_328 ( .C (clk), .D (signal_203), .Q (signal_1267) ) ;
    buf_clk cell_330 ( .C (clk), .D (signal_515), .Q (signal_1269) ) ;
    buf_clk cell_332 ( .C (clk), .D (signal_516), .Q (signal_1271) ) ;
    buf_clk cell_334 ( .C (clk), .D (signal_517), .Q (signal_1273) ) ;
    buf_clk cell_336 ( .C (clk), .D (signal_518), .Q (signal_1275) ) ;
    buf_clk cell_338 ( .C (clk), .D (signal_205), .Q (signal_1277) ) ;
    buf_clk cell_340 ( .C (clk), .D (signal_523), .Q (signal_1279) ) ;
    buf_clk cell_342 ( .C (clk), .D (signal_524), .Q (signal_1281) ) ;
    buf_clk cell_344 ( .C (clk), .D (signal_525), .Q (signal_1283) ) ;
    buf_clk cell_346 ( .C (clk), .D (signal_526), .Q (signal_1285) ) ;
    buf_clk cell_390 ( .C (clk), .D (signal_1328), .Q (signal_1329) ) ;
    buf_clk cell_396 ( .C (clk), .D (signal_1334), .Q (signal_1335) ) ;
    buf_clk cell_402 ( .C (clk), .D (signal_1340), .Q (signal_1341) ) ;
    buf_clk cell_408 ( .C (clk), .D (signal_1346), .Q (signal_1347) ) ;
    buf_clk cell_414 ( .C (clk), .D (signal_1352), .Q (signal_1353) ) ;
    buf_clk cell_420 ( .C (clk), .D (signal_1358), .Q (signal_1359) ) ;
    buf_clk cell_426 ( .C (clk), .D (signal_1364), .Q (signal_1365) ) ;
    buf_clk cell_432 ( .C (clk), .D (signal_1370), .Q (signal_1371) ) ;
    buf_clk cell_438 ( .C (clk), .D (signal_1376), .Q (signal_1377) ) ;
    buf_clk cell_444 ( .C (clk), .D (signal_1382), .Q (signal_1383) ) ;
    buf_clk cell_450 ( .C (clk), .D (signal_1388), .Q (signal_1389) ) ;
    buf_clk cell_456 ( .C (clk), .D (signal_1394), .Q (signal_1395) ) ;
    buf_clk cell_462 ( .C (clk), .D (signal_1400), .Q (signal_1401) ) ;
    buf_clk cell_468 ( .C (clk), .D (signal_1406), .Q (signal_1407) ) ;
    buf_clk cell_474 ( .C (clk), .D (signal_1412), .Q (signal_1413) ) ;
    buf_clk cell_480 ( .C (clk), .D (signal_1418), .Q (signal_1419) ) ;
    buf_clk cell_486 ( .C (clk), .D (signal_1424), .Q (signal_1425) ) ;
    buf_clk cell_492 ( .C (clk), .D (signal_1430), .Q (signal_1431) ) ;
    buf_clk cell_498 ( .C (clk), .D (signal_1436), .Q (signal_1437) ) ;
    buf_clk cell_504 ( .C (clk), .D (signal_1442), .Q (signal_1443) ) ;
    buf_clk cell_510 ( .C (clk), .D (signal_1448), .Q (signal_1449) ) ;
    buf_clk cell_516 ( .C (clk), .D (signal_1454), .Q (signal_1455) ) ;
    buf_clk cell_522 ( .C (clk), .D (signal_1460), .Q (signal_1461) ) ;
    buf_clk cell_528 ( .C (clk), .D (signal_1466), .Q (signal_1467) ) ;
    buf_clk cell_534 ( .C (clk), .D (signal_1472), .Q (signal_1473) ) ;
    buf_clk cell_540 ( .C (clk), .D (signal_1478), .Q (signal_1479) ) ;
    buf_clk cell_546 ( .C (clk), .D (signal_1484), .Q (signal_1485) ) ;
    buf_clk cell_552 ( .C (clk), .D (signal_1490), .Q (signal_1491) ) ;
    buf_clk cell_558 ( .C (clk), .D (signal_1496), .Q (signal_1497) ) ;
    buf_clk cell_564 ( .C (clk), .D (signal_1502), .Q (signal_1503) ) ;
    buf_clk cell_570 ( .C (clk), .D (signal_1508), .Q (signal_1509) ) ;
    buf_clk cell_576 ( .C (clk), .D (signal_1514), .Q (signal_1515) ) ;
    buf_clk cell_582 ( .C (clk), .D (signal_1520), .Q (signal_1521) ) ;
    buf_clk cell_588 ( .C (clk), .D (signal_1526), .Q (signal_1527) ) ;
    buf_clk cell_594 ( .C (clk), .D (signal_1532), .Q (signal_1533) ) ;
    buf_clk cell_600 ( .C (clk), .D (signal_1538), .Q (signal_1539) ) ;
    buf_clk cell_606 ( .C (clk), .D (signal_1544), .Q (signal_1545) ) ;
    buf_clk cell_612 ( .C (clk), .D (signal_1550), .Q (signal_1551) ) ;
    buf_clk cell_618 ( .C (clk), .D (signal_1556), .Q (signal_1557) ) ;
    buf_clk cell_624 ( .C (clk), .D (signal_1562), .Q (signal_1563) ) ;
    buf_clk cell_630 ( .C (clk), .D (signal_1568), .Q (signal_1569) ) ;
    buf_clk cell_636 ( .C (clk), .D (signal_1574), .Q (signal_1575) ) ;
    buf_clk cell_642 ( .C (clk), .D (signal_1580), .Q (signal_1581) ) ;
    buf_clk cell_648 ( .C (clk), .D (signal_1586), .Q (signal_1587) ) ;
    buf_clk cell_654 ( .C (clk), .D (signal_1592), .Q (signal_1593) ) ;
    buf_clk cell_660 ( .C (clk), .D (signal_1598), .Q (signal_1599) ) ;
    buf_clk cell_666 ( .C (clk), .D (signal_1604), .Q (signal_1605) ) ;
    buf_clk cell_672 ( .C (clk), .D (signal_1610), .Q (signal_1611) ) ;
    buf_clk cell_678 ( .C (clk), .D (signal_1616), .Q (signal_1617) ) ;
    buf_clk cell_684 ( .C (clk), .D (signal_1622), .Q (signal_1623) ) ;
    buf_clk cell_690 ( .C (clk), .D (signal_1628), .Q (signal_1629) ) ;
    buf_clk cell_696 ( .C (clk), .D (signal_1634), .Q (signal_1635) ) ;
    buf_clk cell_702 ( .C (clk), .D (signal_1640), .Q (signal_1641) ) ;
    buf_clk cell_708 ( .C (clk), .D (signal_1646), .Q (signal_1647) ) ;
    buf_clk cell_714 ( .C (clk), .D (signal_1652), .Q (signal_1653) ) ;
    buf_clk cell_720 ( .C (clk), .D (signal_1658), .Q (signal_1659) ) ;
    buf_clk cell_726 ( .C (clk), .D (signal_1664), .Q (signal_1665) ) ;
    buf_clk cell_732 ( .C (clk), .D (signal_1670), .Q (signal_1671) ) ;
    buf_clk cell_738 ( .C (clk), .D (signal_1676), .Q (signal_1677) ) ;
    buf_clk cell_744 ( .C (clk), .D (signal_1682), .Q (signal_1683) ) ;
    buf_clk cell_750 ( .C (clk), .D (signal_1688), .Q (signal_1689) ) ;
    buf_clk cell_756 ( .C (clk), .D (signal_1694), .Q (signal_1695) ) ;
    buf_clk cell_762 ( .C (clk), .D (signal_1700), .Q (signal_1701) ) ;
    buf_clk cell_768 ( .C (clk), .D (signal_1706), .Q (signal_1707) ) ;
    buf_clk cell_774 ( .C (clk), .D (signal_1712), .Q (signal_1713) ) ;
    buf_clk cell_780 ( .C (clk), .D (signal_1718), .Q (signal_1719) ) ;
    buf_clk cell_786 ( .C (clk), .D (signal_1724), .Q (signal_1725) ) ;
    buf_clk cell_792 ( .C (clk), .D (signal_1730), .Q (signal_1731) ) ;
    buf_clk cell_798 ( .C (clk), .D (signal_1736), .Q (signal_1737) ) ;
    buf_clk cell_804 ( .C (clk), .D (signal_1742), .Q (signal_1743) ) ;
    buf_clk cell_810 ( .C (clk), .D (signal_1748), .Q (signal_1749) ) ;
    buf_clk cell_816 ( .C (clk), .D (signal_1754), .Q (signal_1755) ) ;
    buf_clk cell_822 ( .C (clk), .D (signal_1760), .Q (signal_1761) ) ;
    buf_clk cell_828 ( .C (clk), .D (signal_1766), .Q (signal_1767) ) ;
    buf_clk cell_834 ( .C (clk), .D (signal_1772), .Q (signal_1773) ) ;
    buf_clk cell_840 ( .C (clk), .D (signal_1778), .Q (signal_1779) ) ;
    buf_clk cell_846 ( .C (clk), .D (signal_1784), .Q (signal_1785) ) ;
    buf_clk cell_852 ( .C (clk), .D (signal_1790), .Q (signal_1791) ) ;
    buf_clk cell_858 ( .C (clk), .D (signal_1796), .Q (signal_1797) ) ;
    buf_clk cell_864 ( .C (clk), .D (signal_1802), .Q (signal_1803) ) ;
    buf_clk cell_870 ( .C (clk), .D (signal_1808), .Q (signal_1809) ) ;
    buf_clk cell_876 ( .C (clk), .D (signal_1814), .Q (signal_1815) ) ;
    buf_clk cell_882 ( .C (clk), .D (signal_1820), .Q (signal_1821) ) ;
    buf_clk cell_888 ( .C (clk), .D (signal_1826), .Q (signal_1827) ) ;
    buf_clk cell_894 ( .C (clk), .D (signal_1832), .Q (signal_1833) ) ;
    buf_clk cell_900 ( .C (clk), .D (signal_1838), .Q (signal_1839) ) ;
    buf_clk cell_906 ( .C (clk), .D (signal_1844), .Q (signal_1845) ) ;
    buf_clk cell_912 ( .C (clk), .D (signal_1850), .Q (signal_1851) ) ;
    buf_clk cell_918 ( .C (clk), .D (signal_1856), .Q (signal_1857) ) ;
    buf_clk cell_924 ( .C (clk), .D (signal_1862), .Q (signal_1863) ) ;

    /* cells in depth 4 */
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_185 ( .a ({signal_494, signal_493, signal_492, signal_491, signal_197}), .b ({signal_502, signal_501, signal_500, signal_499, signal_199}), .clk (clk), .r ({Fresh[99], Fresh[98], Fresh[97], Fresh[96], Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({signal_506, signal_505, signal_504, signal_503, signal_200}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_186 ( .a ({signal_498, signal_497, signal_496, signal_495, signal_198}), .b ({signal_502, signal_501, signal_500, signal_499, signal_199}), .clk (clk), .r ({Fresh[109], Fresh[108], Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100]}), .c ({signal_510, signal_509, signal_508, signal_507, signal_201}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_189 ( .a ({signal_494, signal_493, signal_492, signal_491, signal_197}), .b ({signal_514, signal_513, signal_512, signal_511, signal_202}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114], Fresh[113], Fresh[112], Fresh[111], Fresh[110]}), .c ({signal_522, signal_521, signal_520, signal_519, signal_204}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_191 ( .a ({signal_1256, signal_1254, signal_1252, signal_1250, signal_1248}), .b ({signal_506, signal_505, signal_504, signal_503, signal_200}), .c ({signal_530, signal_529, signal_528, signal_527, signal_206}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_192 ( .a ({signal_1266, signal_1264, signal_1262, signal_1260, signal_1258}), .b ({signal_506, signal_505, signal_504, signal_503, signal_200}), .c ({signal_534, signal_533, signal_532, signal_531, signal_207}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_193 ( .a ({signal_506, signal_505, signal_504, signal_503, signal_200}), .b ({signal_1276, signal_1274, signal_1272, signal_1270, signal_1268}), .c ({signal_538, signal_537, signal_536, signal_535, signal_208}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_198 ( .a ({signal_506, signal_505, signal_504, signal_503, signal_200}), .b ({signal_1286, signal_1284, signal_1282, signal_1280, signal_1278}), .c ({signal_558, signal_557, signal_556, signal_555, signal_213}) ) ;
    buf_clk cell_309 ( .C (clk), .D (signal_1247), .Q (signal_1248) ) ;
    buf_clk cell_311 ( .C (clk), .D (signal_1249), .Q (signal_1250) ) ;
    buf_clk cell_313 ( .C (clk), .D (signal_1251), .Q (signal_1252) ) ;
    buf_clk cell_315 ( .C (clk), .D (signal_1253), .Q (signal_1254) ) ;
    buf_clk cell_317 ( .C (clk), .D (signal_1255), .Q (signal_1256) ) ;
    buf_clk cell_319 ( .C (clk), .D (signal_1257), .Q (signal_1258) ) ;
    buf_clk cell_321 ( .C (clk), .D (signal_1259), .Q (signal_1260) ) ;
    buf_clk cell_323 ( .C (clk), .D (signal_1261), .Q (signal_1262) ) ;
    buf_clk cell_325 ( .C (clk), .D (signal_1263), .Q (signal_1264) ) ;
    buf_clk cell_327 ( .C (clk), .D (signal_1265), .Q (signal_1266) ) ;
    buf_clk cell_329 ( .C (clk), .D (signal_1267), .Q (signal_1268) ) ;
    buf_clk cell_331 ( .C (clk), .D (signal_1269), .Q (signal_1270) ) ;
    buf_clk cell_333 ( .C (clk), .D (signal_1271), .Q (signal_1272) ) ;
    buf_clk cell_335 ( .C (clk), .D (signal_1273), .Q (signal_1274) ) ;
    buf_clk cell_337 ( .C (clk), .D (signal_1275), .Q (signal_1276) ) ;
    buf_clk cell_339 ( .C (clk), .D (signal_1277), .Q (signal_1278) ) ;
    buf_clk cell_341 ( .C (clk), .D (signal_1279), .Q (signal_1280) ) ;
    buf_clk cell_343 ( .C (clk), .D (signal_1281), .Q (signal_1282) ) ;
    buf_clk cell_345 ( .C (clk), .D (signal_1283), .Q (signal_1284) ) ;
    buf_clk cell_347 ( .C (clk), .D (signal_1285), .Q (signal_1286) ) ;
    buf_clk cell_391 ( .C (clk), .D (signal_1329), .Q (signal_1330) ) ;
    buf_clk cell_397 ( .C (clk), .D (signal_1335), .Q (signal_1336) ) ;
    buf_clk cell_403 ( .C (clk), .D (signal_1341), .Q (signal_1342) ) ;
    buf_clk cell_409 ( .C (clk), .D (signal_1347), .Q (signal_1348) ) ;
    buf_clk cell_415 ( .C (clk), .D (signal_1353), .Q (signal_1354) ) ;
    buf_clk cell_421 ( .C (clk), .D (signal_1359), .Q (signal_1360) ) ;
    buf_clk cell_427 ( .C (clk), .D (signal_1365), .Q (signal_1366) ) ;
    buf_clk cell_433 ( .C (clk), .D (signal_1371), .Q (signal_1372) ) ;
    buf_clk cell_439 ( .C (clk), .D (signal_1377), .Q (signal_1378) ) ;
    buf_clk cell_445 ( .C (clk), .D (signal_1383), .Q (signal_1384) ) ;
    buf_clk cell_451 ( .C (clk), .D (signal_1389), .Q (signal_1390) ) ;
    buf_clk cell_457 ( .C (clk), .D (signal_1395), .Q (signal_1396) ) ;
    buf_clk cell_463 ( .C (clk), .D (signal_1401), .Q (signal_1402) ) ;
    buf_clk cell_469 ( .C (clk), .D (signal_1407), .Q (signal_1408) ) ;
    buf_clk cell_475 ( .C (clk), .D (signal_1413), .Q (signal_1414) ) ;
    buf_clk cell_481 ( .C (clk), .D (signal_1419), .Q (signal_1420) ) ;
    buf_clk cell_487 ( .C (clk), .D (signal_1425), .Q (signal_1426) ) ;
    buf_clk cell_493 ( .C (clk), .D (signal_1431), .Q (signal_1432) ) ;
    buf_clk cell_499 ( .C (clk), .D (signal_1437), .Q (signal_1438) ) ;
    buf_clk cell_505 ( .C (clk), .D (signal_1443), .Q (signal_1444) ) ;
    buf_clk cell_511 ( .C (clk), .D (signal_1449), .Q (signal_1450) ) ;
    buf_clk cell_517 ( .C (clk), .D (signal_1455), .Q (signal_1456) ) ;
    buf_clk cell_523 ( .C (clk), .D (signal_1461), .Q (signal_1462) ) ;
    buf_clk cell_529 ( .C (clk), .D (signal_1467), .Q (signal_1468) ) ;
    buf_clk cell_535 ( .C (clk), .D (signal_1473), .Q (signal_1474) ) ;
    buf_clk cell_541 ( .C (clk), .D (signal_1479), .Q (signal_1480) ) ;
    buf_clk cell_547 ( .C (clk), .D (signal_1485), .Q (signal_1486) ) ;
    buf_clk cell_553 ( .C (clk), .D (signal_1491), .Q (signal_1492) ) ;
    buf_clk cell_559 ( .C (clk), .D (signal_1497), .Q (signal_1498) ) ;
    buf_clk cell_565 ( .C (clk), .D (signal_1503), .Q (signal_1504) ) ;
    buf_clk cell_571 ( .C (clk), .D (signal_1509), .Q (signal_1510) ) ;
    buf_clk cell_577 ( .C (clk), .D (signal_1515), .Q (signal_1516) ) ;
    buf_clk cell_583 ( .C (clk), .D (signal_1521), .Q (signal_1522) ) ;
    buf_clk cell_589 ( .C (clk), .D (signal_1527), .Q (signal_1528) ) ;
    buf_clk cell_595 ( .C (clk), .D (signal_1533), .Q (signal_1534) ) ;
    buf_clk cell_601 ( .C (clk), .D (signal_1539), .Q (signal_1540) ) ;
    buf_clk cell_607 ( .C (clk), .D (signal_1545), .Q (signal_1546) ) ;
    buf_clk cell_613 ( .C (clk), .D (signal_1551), .Q (signal_1552) ) ;
    buf_clk cell_619 ( .C (clk), .D (signal_1557), .Q (signal_1558) ) ;
    buf_clk cell_625 ( .C (clk), .D (signal_1563), .Q (signal_1564) ) ;
    buf_clk cell_631 ( .C (clk), .D (signal_1569), .Q (signal_1570) ) ;
    buf_clk cell_637 ( .C (clk), .D (signal_1575), .Q (signal_1576) ) ;
    buf_clk cell_643 ( .C (clk), .D (signal_1581), .Q (signal_1582) ) ;
    buf_clk cell_649 ( .C (clk), .D (signal_1587), .Q (signal_1588) ) ;
    buf_clk cell_655 ( .C (clk), .D (signal_1593), .Q (signal_1594) ) ;
    buf_clk cell_661 ( .C (clk), .D (signal_1599), .Q (signal_1600) ) ;
    buf_clk cell_667 ( .C (clk), .D (signal_1605), .Q (signal_1606) ) ;
    buf_clk cell_673 ( .C (clk), .D (signal_1611), .Q (signal_1612) ) ;
    buf_clk cell_679 ( .C (clk), .D (signal_1617), .Q (signal_1618) ) ;
    buf_clk cell_685 ( .C (clk), .D (signal_1623), .Q (signal_1624) ) ;
    buf_clk cell_691 ( .C (clk), .D (signal_1629), .Q (signal_1630) ) ;
    buf_clk cell_697 ( .C (clk), .D (signal_1635), .Q (signal_1636) ) ;
    buf_clk cell_703 ( .C (clk), .D (signal_1641), .Q (signal_1642) ) ;
    buf_clk cell_709 ( .C (clk), .D (signal_1647), .Q (signal_1648) ) ;
    buf_clk cell_715 ( .C (clk), .D (signal_1653), .Q (signal_1654) ) ;
    buf_clk cell_721 ( .C (clk), .D (signal_1659), .Q (signal_1660) ) ;
    buf_clk cell_727 ( .C (clk), .D (signal_1665), .Q (signal_1666) ) ;
    buf_clk cell_733 ( .C (clk), .D (signal_1671), .Q (signal_1672) ) ;
    buf_clk cell_739 ( .C (clk), .D (signal_1677), .Q (signal_1678) ) ;
    buf_clk cell_745 ( .C (clk), .D (signal_1683), .Q (signal_1684) ) ;
    buf_clk cell_751 ( .C (clk), .D (signal_1689), .Q (signal_1690) ) ;
    buf_clk cell_757 ( .C (clk), .D (signal_1695), .Q (signal_1696) ) ;
    buf_clk cell_763 ( .C (clk), .D (signal_1701), .Q (signal_1702) ) ;
    buf_clk cell_769 ( .C (clk), .D (signal_1707), .Q (signal_1708) ) ;
    buf_clk cell_775 ( .C (clk), .D (signal_1713), .Q (signal_1714) ) ;
    buf_clk cell_781 ( .C (clk), .D (signal_1719), .Q (signal_1720) ) ;
    buf_clk cell_787 ( .C (clk), .D (signal_1725), .Q (signal_1726) ) ;
    buf_clk cell_793 ( .C (clk), .D (signal_1731), .Q (signal_1732) ) ;
    buf_clk cell_799 ( .C (clk), .D (signal_1737), .Q (signal_1738) ) ;
    buf_clk cell_805 ( .C (clk), .D (signal_1743), .Q (signal_1744) ) ;
    buf_clk cell_811 ( .C (clk), .D (signal_1749), .Q (signal_1750) ) ;
    buf_clk cell_817 ( .C (clk), .D (signal_1755), .Q (signal_1756) ) ;
    buf_clk cell_823 ( .C (clk), .D (signal_1761), .Q (signal_1762) ) ;
    buf_clk cell_829 ( .C (clk), .D (signal_1767), .Q (signal_1768) ) ;
    buf_clk cell_835 ( .C (clk), .D (signal_1773), .Q (signal_1774) ) ;
    buf_clk cell_841 ( .C (clk), .D (signal_1779), .Q (signal_1780) ) ;
    buf_clk cell_847 ( .C (clk), .D (signal_1785), .Q (signal_1786) ) ;
    buf_clk cell_853 ( .C (clk), .D (signal_1791), .Q (signal_1792) ) ;
    buf_clk cell_859 ( .C (clk), .D (signal_1797), .Q (signal_1798) ) ;
    buf_clk cell_865 ( .C (clk), .D (signal_1803), .Q (signal_1804) ) ;
    buf_clk cell_871 ( .C (clk), .D (signal_1809), .Q (signal_1810) ) ;
    buf_clk cell_877 ( .C (clk), .D (signal_1815), .Q (signal_1816) ) ;
    buf_clk cell_883 ( .C (clk), .D (signal_1821), .Q (signal_1822) ) ;
    buf_clk cell_889 ( .C (clk), .D (signal_1827), .Q (signal_1828) ) ;
    buf_clk cell_895 ( .C (clk), .D (signal_1833), .Q (signal_1834) ) ;
    buf_clk cell_901 ( .C (clk), .D (signal_1839), .Q (signal_1840) ) ;
    buf_clk cell_907 ( .C (clk), .D (signal_1845), .Q (signal_1846) ) ;
    buf_clk cell_913 ( .C (clk), .D (signal_1851), .Q (signal_1852) ) ;
    buf_clk cell_919 ( .C (clk), .D (signal_1857), .Q (signal_1858) ) ;
    buf_clk cell_925 ( .C (clk), .D (signal_1863), .Q (signal_1864) ) ;

    /* cells in depth 5 */
    buf_clk cell_348 ( .C (clk), .D (signal_1248), .Q (signal_1287) ) ;
    buf_clk cell_350 ( .C (clk), .D (signal_1250), .Q (signal_1289) ) ;
    buf_clk cell_352 ( .C (clk), .D (signal_1252), .Q (signal_1291) ) ;
    buf_clk cell_354 ( .C (clk), .D (signal_1254), .Q (signal_1293) ) ;
    buf_clk cell_356 ( .C (clk), .D (signal_1256), .Q (signal_1295) ) ;
    buf_clk cell_358 ( .C (clk), .D (signal_208), .Q (signal_1297) ) ;
    buf_clk cell_360 ( .C (clk), .D (signal_535), .Q (signal_1299) ) ;
    buf_clk cell_362 ( .C (clk), .D (signal_536), .Q (signal_1301) ) ;
    buf_clk cell_364 ( .C (clk), .D (signal_537), .Q (signal_1303) ) ;
    buf_clk cell_366 ( .C (clk), .D (signal_538), .Q (signal_1305) ) ;
    buf_clk cell_368 ( .C (clk), .D (signal_1258), .Q (signal_1307) ) ;
    buf_clk cell_370 ( .C (clk), .D (signal_1260), .Q (signal_1309) ) ;
    buf_clk cell_372 ( .C (clk), .D (signal_1262), .Q (signal_1311) ) ;
    buf_clk cell_374 ( .C (clk), .D (signal_1264), .Q (signal_1313) ) ;
    buf_clk cell_376 ( .C (clk), .D (signal_1266), .Q (signal_1315) ) ;
    buf_clk cell_378 ( .C (clk), .D (signal_213), .Q (signal_1317) ) ;
    buf_clk cell_380 ( .C (clk), .D (signal_555), .Q (signal_1319) ) ;
    buf_clk cell_382 ( .C (clk), .D (signal_556), .Q (signal_1321) ) ;
    buf_clk cell_384 ( .C (clk), .D (signal_557), .Q (signal_1323) ) ;
    buf_clk cell_386 ( .C (clk), .D (signal_558), .Q (signal_1325) ) ;
    buf_clk cell_392 ( .C (clk), .D (signal_1330), .Q (signal_1331) ) ;
    buf_clk cell_398 ( .C (clk), .D (signal_1336), .Q (signal_1337) ) ;
    buf_clk cell_404 ( .C (clk), .D (signal_1342), .Q (signal_1343) ) ;
    buf_clk cell_410 ( .C (clk), .D (signal_1348), .Q (signal_1349) ) ;
    buf_clk cell_416 ( .C (clk), .D (signal_1354), .Q (signal_1355) ) ;
    buf_clk cell_422 ( .C (clk), .D (signal_1360), .Q (signal_1361) ) ;
    buf_clk cell_428 ( .C (clk), .D (signal_1366), .Q (signal_1367) ) ;
    buf_clk cell_434 ( .C (clk), .D (signal_1372), .Q (signal_1373) ) ;
    buf_clk cell_440 ( .C (clk), .D (signal_1378), .Q (signal_1379) ) ;
    buf_clk cell_446 ( .C (clk), .D (signal_1384), .Q (signal_1385) ) ;
    buf_clk cell_452 ( .C (clk), .D (signal_1390), .Q (signal_1391) ) ;
    buf_clk cell_458 ( .C (clk), .D (signal_1396), .Q (signal_1397) ) ;
    buf_clk cell_464 ( .C (clk), .D (signal_1402), .Q (signal_1403) ) ;
    buf_clk cell_470 ( .C (clk), .D (signal_1408), .Q (signal_1409) ) ;
    buf_clk cell_476 ( .C (clk), .D (signal_1414), .Q (signal_1415) ) ;
    buf_clk cell_482 ( .C (clk), .D (signal_1420), .Q (signal_1421) ) ;
    buf_clk cell_488 ( .C (clk), .D (signal_1426), .Q (signal_1427) ) ;
    buf_clk cell_494 ( .C (clk), .D (signal_1432), .Q (signal_1433) ) ;
    buf_clk cell_500 ( .C (clk), .D (signal_1438), .Q (signal_1439) ) ;
    buf_clk cell_506 ( .C (clk), .D (signal_1444), .Q (signal_1445) ) ;
    buf_clk cell_512 ( .C (clk), .D (signal_1450), .Q (signal_1451) ) ;
    buf_clk cell_518 ( .C (clk), .D (signal_1456), .Q (signal_1457) ) ;
    buf_clk cell_524 ( .C (clk), .D (signal_1462), .Q (signal_1463) ) ;
    buf_clk cell_530 ( .C (clk), .D (signal_1468), .Q (signal_1469) ) ;
    buf_clk cell_536 ( .C (clk), .D (signal_1474), .Q (signal_1475) ) ;
    buf_clk cell_542 ( .C (clk), .D (signal_1480), .Q (signal_1481) ) ;
    buf_clk cell_548 ( .C (clk), .D (signal_1486), .Q (signal_1487) ) ;
    buf_clk cell_554 ( .C (clk), .D (signal_1492), .Q (signal_1493) ) ;
    buf_clk cell_560 ( .C (clk), .D (signal_1498), .Q (signal_1499) ) ;
    buf_clk cell_566 ( .C (clk), .D (signal_1504), .Q (signal_1505) ) ;
    buf_clk cell_572 ( .C (clk), .D (signal_1510), .Q (signal_1511) ) ;
    buf_clk cell_578 ( .C (clk), .D (signal_1516), .Q (signal_1517) ) ;
    buf_clk cell_584 ( .C (clk), .D (signal_1522), .Q (signal_1523) ) ;
    buf_clk cell_590 ( .C (clk), .D (signal_1528), .Q (signal_1529) ) ;
    buf_clk cell_596 ( .C (clk), .D (signal_1534), .Q (signal_1535) ) ;
    buf_clk cell_602 ( .C (clk), .D (signal_1540), .Q (signal_1541) ) ;
    buf_clk cell_608 ( .C (clk), .D (signal_1546), .Q (signal_1547) ) ;
    buf_clk cell_614 ( .C (clk), .D (signal_1552), .Q (signal_1553) ) ;
    buf_clk cell_620 ( .C (clk), .D (signal_1558), .Q (signal_1559) ) ;
    buf_clk cell_626 ( .C (clk), .D (signal_1564), .Q (signal_1565) ) ;
    buf_clk cell_632 ( .C (clk), .D (signal_1570), .Q (signal_1571) ) ;
    buf_clk cell_638 ( .C (clk), .D (signal_1576), .Q (signal_1577) ) ;
    buf_clk cell_644 ( .C (clk), .D (signal_1582), .Q (signal_1583) ) ;
    buf_clk cell_650 ( .C (clk), .D (signal_1588), .Q (signal_1589) ) ;
    buf_clk cell_656 ( .C (clk), .D (signal_1594), .Q (signal_1595) ) ;
    buf_clk cell_662 ( .C (clk), .D (signal_1600), .Q (signal_1601) ) ;
    buf_clk cell_668 ( .C (clk), .D (signal_1606), .Q (signal_1607) ) ;
    buf_clk cell_674 ( .C (clk), .D (signal_1612), .Q (signal_1613) ) ;
    buf_clk cell_680 ( .C (clk), .D (signal_1618), .Q (signal_1619) ) ;
    buf_clk cell_686 ( .C (clk), .D (signal_1624), .Q (signal_1625) ) ;
    buf_clk cell_692 ( .C (clk), .D (signal_1630), .Q (signal_1631) ) ;
    buf_clk cell_698 ( .C (clk), .D (signal_1636), .Q (signal_1637) ) ;
    buf_clk cell_704 ( .C (clk), .D (signal_1642), .Q (signal_1643) ) ;
    buf_clk cell_710 ( .C (clk), .D (signal_1648), .Q (signal_1649) ) ;
    buf_clk cell_716 ( .C (clk), .D (signal_1654), .Q (signal_1655) ) ;
    buf_clk cell_722 ( .C (clk), .D (signal_1660), .Q (signal_1661) ) ;
    buf_clk cell_728 ( .C (clk), .D (signal_1666), .Q (signal_1667) ) ;
    buf_clk cell_734 ( .C (clk), .D (signal_1672), .Q (signal_1673) ) ;
    buf_clk cell_740 ( .C (clk), .D (signal_1678), .Q (signal_1679) ) ;
    buf_clk cell_746 ( .C (clk), .D (signal_1684), .Q (signal_1685) ) ;
    buf_clk cell_752 ( .C (clk), .D (signal_1690), .Q (signal_1691) ) ;
    buf_clk cell_758 ( .C (clk), .D (signal_1696), .Q (signal_1697) ) ;
    buf_clk cell_764 ( .C (clk), .D (signal_1702), .Q (signal_1703) ) ;
    buf_clk cell_770 ( .C (clk), .D (signal_1708), .Q (signal_1709) ) ;
    buf_clk cell_776 ( .C (clk), .D (signal_1714), .Q (signal_1715) ) ;
    buf_clk cell_782 ( .C (clk), .D (signal_1720), .Q (signal_1721) ) ;
    buf_clk cell_788 ( .C (clk), .D (signal_1726), .Q (signal_1727) ) ;
    buf_clk cell_794 ( .C (clk), .D (signal_1732), .Q (signal_1733) ) ;
    buf_clk cell_800 ( .C (clk), .D (signal_1738), .Q (signal_1739) ) ;
    buf_clk cell_806 ( .C (clk), .D (signal_1744), .Q (signal_1745) ) ;
    buf_clk cell_812 ( .C (clk), .D (signal_1750), .Q (signal_1751) ) ;
    buf_clk cell_818 ( .C (clk), .D (signal_1756), .Q (signal_1757) ) ;
    buf_clk cell_824 ( .C (clk), .D (signal_1762), .Q (signal_1763) ) ;
    buf_clk cell_830 ( .C (clk), .D (signal_1768), .Q (signal_1769) ) ;
    buf_clk cell_836 ( .C (clk), .D (signal_1774), .Q (signal_1775) ) ;
    buf_clk cell_842 ( .C (clk), .D (signal_1780), .Q (signal_1781) ) ;
    buf_clk cell_848 ( .C (clk), .D (signal_1786), .Q (signal_1787) ) ;
    buf_clk cell_854 ( .C (clk), .D (signal_1792), .Q (signal_1793) ) ;
    buf_clk cell_860 ( .C (clk), .D (signal_1798), .Q (signal_1799) ) ;
    buf_clk cell_866 ( .C (clk), .D (signal_1804), .Q (signal_1805) ) ;
    buf_clk cell_872 ( .C (clk), .D (signal_1810), .Q (signal_1811) ) ;
    buf_clk cell_878 ( .C (clk), .D (signal_1816), .Q (signal_1817) ) ;
    buf_clk cell_884 ( .C (clk), .D (signal_1822), .Q (signal_1823) ) ;
    buf_clk cell_890 ( .C (clk), .D (signal_1828), .Q (signal_1829) ) ;
    buf_clk cell_896 ( .C (clk), .D (signal_1834), .Q (signal_1835) ) ;
    buf_clk cell_902 ( .C (clk), .D (signal_1840), .Q (signal_1841) ) ;
    buf_clk cell_908 ( .C (clk), .D (signal_1846), .Q (signal_1847) ) ;
    buf_clk cell_914 ( .C (clk), .D (signal_1852), .Q (signal_1853) ) ;
    buf_clk cell_920 ( .C (clk), .D (signal_1858), .Q (signal_1859) ) ;
    buf_clk cell_926 ( .C (clk), .D (signal_1864), .Q (signal_1865) ) ;

    /* cells in depth 6 */
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_194 ( .a ({signal_1276, signal_1274, signal_1272, signal_1270, signal_1268}), .b ({signal_534, signal_533, signal_532, signal_531, signal_207}), .clk (clk), .r ({Fresh[129], Fresh[128], Fresh[127], Fresh[126], Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({signal_542, signal_541, signal_540, signal_539, signal_209}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_195 ( .a ({signal_1286, signal_1284, signal_1282, signal_1280, signal_1278}), .b ({signal_530, signal_529, signal_528, signal_527, signal_206}), .clk (clk), .r ({Fresh[139], Fresh[138], Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132], Fresh[131], Fresh[130]}), .c ({signal_546, signal_545, signal_544, signal_543, signal_210}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_196 ( .a ({signal_1276, signal_1274, signal_1272, signal_1270, signal_1268}), .b ({signal_522, signal_521, signal_520, signal_519, signal_204}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144], Fresh[143], Fresh[142], Fresh[141], Fresh[140]}), .c ({signal_550, signal_549, signal_548, signal_547, signal_211}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_197 ( .a ({signal_510, signal_509, signal_508, signal_507, signal_201}), .b ({signal_1286, signal_1284, signal_1282, signal_1280, signal_1278}), .clk (clk), .r ({Fresh[159], Fresh[158], Fresh[157], Fresh[156], Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .c ({signal_554, signal_553, signal_552, signal_551, signal_212}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_199 ( .a ({signal_1296, signal_1294, signal_1292, signal_1290, signal_1288}), .b ({signal_542, signal_541, signal_540, signal_539, signal_209}), .c ({signal_562, signal_561, signal_560, signal_559, signal_214}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_200 ( .a ({signal_1306, signal_1304, signal_1302, signal_1300, signal_1298}), .b ({signal_550, signal_549, signal_548, signal_547, signal_211}), .c ({signal_566, signal_565, signal_564, signal_563, signal_215}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_201 ( .a ({signal_1316, signal_1314, signal_1312, signal_1310, signal_1308}), .b ({signal_546, signal_545, signal_544, signal_543, signal_210}), .c ({signal_570, signal_569, signal_568, signal_567, signal_216}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_202 ( .a ({signal_554, signal_553, signal_552, signal_551, signal_212}), .b ({signal_1326, signal_1324, signal_1322, signal_1320, signal_1318}), .c ({signal_574, signal_573, signal_572, signal_571, signal_217}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_211 ( .a ({signal_566, signal_565, signal_564, signal_563, signal_215}), .b ({signal_574, signal_573, signal_572, signal_571, signal_217}), .c ({signal_610, signal_609, signal_608, signal_607, signal_226}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_212 ( .a ({signal_562, signal_561, signal_560, signal_559, signal_214}), .b ({signal_570, signal_569, signal_568, signal_567, signal_216}), .c ({signal_614, signal_613, signal_612, signal_611, signal_227}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_213 ( .a ({signal_562, signal_561, signal_560, signal_559, signal_214}), .b ({signal_566, signal_565, signal_564, signal_563, signal_215}), .c ({signal_618, signal_617, signal_616, signal_615, signal_228}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_214 ( .a ({signal_570, signal_569, signal_568, signal_567, signal_216}), .b ({signal_574, signal_573, signal_572, signal_571, signal_217}), .c ({signal_622, signal_621, signal_620, signal_619, signal_229}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_223 ( .a ({signal_610, signal_609, signal_608, signal_607, signal_226}), .b ({signal_614, signal_613, signal_612, signal_611, signal_227}), .c ({signal_658, signal_657, signal_656, signal_655, signal_238}) ) ;
    buf_clk cell_349 ( .C (clk), .D (signal_1287), .Q (signal_1288) ) ;
    buf_clk cell_351 ( .C (clk), .D (signal_1289), .Q (signal_1290) ) ;
    buf_clk cell_353 ( .C (clk), .D (signal_1291), .Q (signal_1292) ) ;
    buf_clk cell_355 ( .C (clk), .D (signal_1293), .Q (signal_1294) ) ;
    buf_clk cell_357 ( .C (clk), .D (signal_1295), .Q (signal_1296) ) ;
    buf_clk cell_359 ( .C (clk), .D (signal_1297), .Q (signal_1298) ) ;
    buf_clk cell_361 ( .C (clk), .D (signal_1299), .Q (signal_1300) ) ;
    buf_clk cell_363 ( .C (clk), .D (signal_1301), .Q (signal_1302) ) ;
    buf_clk cell_365 ( .C (clk), .D (signal_1303), .Q (signal_1304) ) ;
    buf_clk cell_367 ( .C (clk), .D (signal_1305), .Q (signal_1306) ) ;
    buf_clk cell_369 ( .C (clk), .D (signal_1307), .Q (signal_1308) ) ;
    buf_clk cell_371 ( .C (clk), .D (signal_1309), .Q (signal_1310) ) ;
    buf_clk cell_373 ( .C (clk), .D (signal_1311), .Q (signal_1312) ) ;
    buf_clk cell_375 ( .C (clk), .D (signal_1313), .Q (signal_1314) ) ;
    buf_clk cell_377 ( .C (clk), .D (signal_1315), .Q (signal_1316) ) ;
    buf_clk cell_379 ( .C (clk), .D (signal_1317), .Q (signal_1318) ) ;
    buf_clk cell_381 ( .C (clk), .D (signal_1319), .Q (signal_1320) ) ;
    buf_clk cell_383 ( .C (clk), .D (signal_1321), .Q (signal_1322) ) ;
    buf_clk cell_385 ( .C (clk), .D (signal_1323), .Q (signal_1324) ) ;
    buf_clk cell_387 ( .C (clk), .D (signal_1325), .Q (signal_1326) ) ;
    buf_clk cell_393 ( .C (clk), .D (signal_1331), .Q (signal_1332) ) ;
    buf_clk cell_399 ( .C (clk), .D (signal_1337), .Q (signal_1338) ) ;
    buf_clk cell_405 ( .C (clk), .D (signal_1343), .Q (signal_1344) ) ;
    buf_clk cell_411 ( .C (clk), .D (signal_1349), .Q (signal_1350) ) ;
    buf_clk cell_417 ( .C (clk), .D (signal_1355), .Q (signal_1356) ) ;
    buf_clk cell_423 ( .C (clk), .D (signal_1361), .Q (signal_1362) ) ;
    buf_clk cell_429 ( .C (clk), .D (signal_1367), .Q (signal_1368) ) ;
    buf_clk cell_435 ( .C (clk), .D (signal_1373), .Q (signal_1374) ) ;
    buf_clk cell_441 ( .C (clk), .D (signal_1379), .Q (signal_1380) ) ;
    buf_clk cell_447 ( .C (clk), .D (signal_1385), .Q (signal_1386) ) ;
    buf_clk cell_453 ( .C (clk), .D (signal_1391), .Q (signal_1392) ) ;
    buf_clk cell_459 ( .C (clk), .D (signal_1397), .Q (signal_1398) ) ;
    buf_clk cell_465 ( .C (clk), .D (signal_1403), .Q (signal_1404) ) ;
    buf_clk cell_471 ( .C (clk), .D (signal_1409), .Q (signal_1410) ) ;
    buf_clk cell_477 ( .C (clk), .D (signal_1415), .Q (signal_1416) ) ;
    buf_clk cell_483 ( .C (clk), .D (signal_1421), .Q (signal_1422) ) ;
    buf_clk cell_489 ( .C (clk), .D (signal_1427), .Q (signal_1428) ) ;
    buf_clk cell_495 ( .C (clk), .D (signal_1433), .Q (signal_1434) ) ;
    buf_clk cell_501 ( .C (clk), .D (signal_1439), .Q (signal_1440) ) ;
    buf_clk cell_507 ( .C (clk), .D (signal_1445), .Q (signal_1446) ) ;
    buf_clk cell_513 ( .C (clk), .D (signal_1451), .Q (signal_1452) ) ;
    buf_clk cell_519 ( .C (clk), .D (signal_1457), .Q (signal_1458) ) ;
    buf_clk cell_525 ( .C (clk), .D (signal_1463), .Q (signal_1464) ) ;
    buf_clk cell_531 ( .C (clk), .D (signal_1469), .Q (signal_1470) ) ;
    buf_clk cell_537 ( .C (clk), .D (signal_1475), .Q (signal_1476) ) ;
    buf_clk cell_543 ( .C (clk), .D (signal_1481), .Q (signal_1482) ) ;
    buf_clk cell_549 ( .C (clk), .D (signal_1487), .Q (signal_1488) ) ;
    buf_clk cell_555 ( .C (clk), .D (signal_1493), .Q (signal_1494) ) ;
    buf_clk cell_561 ( .C (clk), .D (signal_1499), .Q (signal_1500) ) ;
    buf_clk cell_567 ( .C (clk), .D (signal_1505), .Q (signal_1506) ) ;
    buf_clk cell_573 ( .C (clk), .D (signal_1511), .Q (signal_1512) ) ;
    buf_clk cell_579 ( .C (clk), .D (signal_1517), .Q (signal_1518) ) ;
    buf_clk cell_585 ( .C (clk), .D (signal_1523), .Q (signal_1524) ) ;
    buf_clk cell_591 ( .C (clk), .D (signal_1529), .Q (signal_1530) ) ;
    buf_clk cell_597 ( .C (clk), .D (signal_1535), .Q (signal_1536) ) ;
    buf_clk cell_603 ( .C (clk), .D (signal_1541), .Q (signal_1542) ) ;
    buf_clk cell_609 ( .C (clk), .D (signal_1547), .Q (signal_1548) ) ;
    buf_clk cell_615 ( .C (clk), .D (signal_1553), .Q (signal_1554) ) ;
    buf_clk cell_621 ( .C (clk), .D (signal_1559), .Q (signal_1560) ) ;
    buf_clk cell_627 ( .C (clk), .D (signal_1565), .Q (signal_1566) ) ;
    buf_clk cell_633 ( .C (clk), .D (signal_1571), .Q (signal_1572) ) ;
    buf_clk cell_639 ( .C (clk), .D (signal_1577), .Q (signal_1578) ) ;
    buf_clk cell_645 ( .C (clk), .D (signal_1583), .Q (signal_1584) ) ;
    buf_clk cell_651 ( .C (clk), .D (signal_1589), .Q (signal_1590) ) ;
    buf_clk cell_657 ( .C (clk), .D (signal_1595), .Q (signal_1596) ) ;
    buf_clk cell_663 ( .C (clk), .D (signal_1601), .Q (signal_1602) ) ;
    buf_clk cell_669 ( .C (clk), .D (signal_1607), .Q (signal_1608) ) ;
    buf_clk cell_675 ( .C (clk), .D (signal_1613), .Q (signal_1614) ) ;
    buf_clk cell_681 ( .C (clk), .D (signal_1619), .Q (signal_1620) ) ;
    buf_clk cell_687 ( .C (clk), .D (signal_1625), .Q (signal_1626) ) ;
    buf_clk cell_693 ( .C (clk), .D (signal_1631), .Q (signal_1632) ) ;
    buf_clk cell_699 ( .C (clk), .D (signal_1637), .Q (signal_1638) ) ;
    buf_clk cell_705 ( .C (clk), .D (signal_1643), .Q (signal_1644) ) ;
    buf_clk cell_711 ( .C (clk), .D (signal_1649), .Q (signal_1650) ) ;
    buf_clk cell_717 ( .C (clk), .D (signal_1655), .Q (signal_1656) ) ;
    buf_clk cell_723 ( .C (clk), .D (signal_1661), .Q (signal_1662) ) ;
    buf_clk cell_729 ( .C (clk), .D (signal_1667), .Q (signal_1668) ) ;
    buf_clk cell_735 ( .C (clk), .D (signal_1673), .Q (signal_1674) ) ;
    buf_clk cell_741 ( .C (clk), .D (signal_1679), .Q (signal_1680) ) ;
    buf_clk cell_747 ( .C (clk), .D (signal_1685), .Q (signal_1686) ) ;
    buf_clk cell_753 ( .C (clk), .D (signal_1691), .Q (signal_1692) ) ;
    buf_clk cell_759 ( .C (clk), .D (signal_1697), .Q (signal_1698) ) ;
    buf_clk cell_765 ( .C (clk), .D (signal_1703), .Q (signal_1704) ) ;
    buf_clk cell_771 ( .C (clk), .D (signal_1709), .Q (signal_1710) ) ;
    buf_clk cell_777 ( .C (clk), .D (signal_1715), .Q (signal_1716) ) ;
    buf_clk cell_783 ( .C (clk), .D (signal_1721), .Q (signal_1722) ) ;
    buf_clk cell_789 ( .C (clk), .D (signal_1727), .Q (signal_1728) ) ;
    buf_clk cell_795 ( .C (clk), .D (signal_1733), .Q (signal_1734) ) ;
    buf_clk cell_801 ( .C (clk), .D (signal_1739), .Q (signal_1740) ) ;
    buf_clk cell_807 ( .C (clk), .D (signal_1745), .Q (signal_1746) ) ;
    buf_clk cell_813 ( .C (clk), .D (signal_1751), .Q (signal_1752) ) ;
    buf_clk cell_819 ( .C (clk), .D (signal_1757), .Q (signal_1758) ) ;
    buf_clk cell_825 ( .C (clk), .D (signal_1763), .Q (signal_1764) ) ;
    buf_clk cell_831 ( .C (clk), .D (signal_1769), .Q (signal_1770) ) ;
    buf_clk cell_837 ( .C (clk), .D (signal_1775), .Q (signal_1776) ) ;
    buf_clk cell_843 ( .C (clk), .D (signal_1781), .Q (signal_1782) ) ;
    buf_clk cell_849 ( .C (clk), .D (signal_1787), .Q (signal_1788) ) ;
    buf_clk cell_855 ( .C (clk), .D (signal_1793), .Q (signal_1794) ) ;
    buf_clk cell_861 ( .C (clk), .D (signal_1799), .Q (signal_1800) ) ;
    buf_clk cell_867 ( .C (clk), .D (signal_1805), .Q (signal_1806) ) ;
    buf_clk cell_873 ( .C (clk), .D (signal_1811), .Q (signal_1812) ) ;
    buf_clk cell_879 ( .C (clk), .D (signal_1817), .Q (signal_1818) ) ;
    buf_clk cell_885 ( .C (clk), .D (signal_1823), .Q (signal_1824) ) ;
    buf_clk cell_891 ( .C (clk), .D (signal_1829), .Q (signal_1830) ) ;
    buf_clk cell_897 ( .C (clk), .D (signal_1835), .Q (signal_1836) ) ;
    buf_clk cell_903 ( .C (clk), .D (signal_1841), .Q (signal_1842) ) ;
    buf_clk cell_909 ( .C (clk), .D (signal_1847), .Q (signal_1848) ) ;
    buf_clk cell_915 ( .C (clk), .D (signal_1853), .Q (signal_1854) ) ;
    buf_clk cell_921 ( .C (clk), .D (signal_1859), .Q (signal_1860) ) ;
    buf_clk cell_927 ( .C (clk), .D (signal_1865), .Q (signal_1866) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_203 ( .a ({signal_1356, signal_1350, signal_1344, signal_1338, signal_1332}), .b ({signal_574, signal_573, signal_572, signal_571, signal_217}), .clk (clk), .r ({Fresh[169], Fresh[168], Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162], Fresh[161], Fresh[160]}), .c ({signal_578, signal_577, signal_576, signal_575, signal_218}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_204 ( .a ({signal_1386, signal_1380, signal_1374, signal_1368, signal_1362}), .b ({signal_570, signal_569, signal_568, signal_567, signal_216}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174], Fresh[173], Fresh[172], Fresh[171], Fresh[170]}), .c ({signal_582, signal_581, signal_580, signal_579, signal_219}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_205 ( .a ({signal_1416, signal_1410, signal_1404, signal_1398, signal_1392}), .b ({signal_566, signal_565, signal_564, signal_563, signal_215}), .clk (clk), .r ({Fresh[189], Fresh[188], Fresh[187], Fresh[186], Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({signal_586, signal_585, signal_584, signal_583, signal_220}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_206 ( .a ({signal_1446, signal_1440, signal_1434, signal_1428, signal_1422}), .b ({signal_562, signal_561, signal_560, signal_559, signal_214}), .clk (clk), .r ({Fresh[199], Fresh[198], Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192], Fresh[191], Fresh[190]}), .c ({signal_590, signal_589, signal_588, signal_587, signal_221}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_207 ( .a ({signal_1476, signal_1470, signal_1464, signal_1458, signal_1452}), .b ({signal_574, signal_573, signal_572, signal_571, signal_217}), .clk (clk), .r ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204], Fresh[203], Fresh[202], Fresh[201], Fresh[200]}), .c ({signal_594, signal_593, signal_592, signal_591, signal_222}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_208 ( .a ({signal_1506, signal_1500, signal_1494, signal_1488, signal_1482}), .b ({signal_570, signal_569, signal_568, signal_567, signal_216}), .clk (clk), .r ({Fresh[219], Fresh[218], Fresh[217], Fresh[216], Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .c ({signal_598, signal_597, signal_596, signal_595, signal_223}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_209 ( .a ({signal_1536, signal_1530, signal_1524, signal_1518, signal_1512}), .b ({signal_566, signal_565, signal_564, signal_563, signal_215}), .clk (clk), .r ({Fresh[229], Fresh[228], Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222], Fresh[221], Fresh[220]}), .c ({signal_602, signal_601, signal_600, signal_599, signal_224}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_210 ( .a ({signal_1566, signal_1560, signal_1554, signal_1548, signal_1542}), .b ({signal_562, signal_561, signal_560, signal_559, signal_214}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234], Fresh[233], Fresh[232], Fresh[231], Fresh[230]}), .c ({signal_606, signal_605, signal_604, signal_603, signal_225}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_215 ( .a ({signal_1596, signal_1590, signal_1584, signal_1578, signal_1572}), .b ({signal_622, signal_621, signal_620, signal_619, signal_229}), .clk (clk), .r ({Fresh[249], Fresh[248], Fresh[247], Fresh[246], Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .c ({signal_626, signal_625, signal_624, signal_623, signal_230}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_216 ( .a ({signal_1626, signal_1620, signal_1614, signal_1608, signal_1602}), .b ({signal_618, signal_617, signal_616, signal_615, signal_228}), .clk (clk), .r ({Fresh[259], Fresh[258], Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252], Fresh[251], Fresh[250]}), .c ({signal_630, signal_629, signal_628, signal_627, signal_231}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_217 ( .a ({signal_1656, signal_1650, signal_1644, signal_1638, signal_1632}), .b ({signal_614, signal_613, signal_612, signal_611, signal_227}), .clk (clk), .r ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264], Fresh[263], Fresh[262], Fresh[261], Fresh[260]}), .c ({signal_634, signal_633, signal_632, signal_631, signal_232}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_218 ( .a ({signal_1686, signal_1680, signal_1674, signal_1668, signal_1662}), .b ({signal_610, signal_609, signal_608, signal_607, signal_226}), .clk (clk), .r ({Fresh[279], Fresh[278], Fresh[277], Fresh[276], Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .c ({signal_638, signal_637, signal_636, signal_635, signal_233}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_219 ( .a ({signal_1716, signal_1710, signal_1704, signal_1698, signal_1692}), .b ({signal_622, signal_621, signal_620, signal_619, signal_229}), .clk (clk), .r ({Fresh[289], Fresh[288], Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282], Fresh[281], Fresh[280]}), .c ({signal_642, signal_641, signal_640, signal_639, signal_234}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_220 ( .a ({signal_1746, signal_1740, signal_1734, signal_1728, signal_1722}), .b ({signal_618, signal_617, signal_616, signal_615, signal_228}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294], Fresh[293], Fresh[292], Fresh[291], Fresh[290]}), .c ({signal_646, signal_645, signal_644, signal_643, signal_235}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_221 ( .a ({signal_1776, signal_1770, signal_1764, signal_1758, signal_1752}), .b ({signal_614, signal_613, signal_612, signal_611, signal_227}), .clk (clk), .r ({Fresh[309], Fresh[308], Fresh[307], Fresh[306], Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .c ({signal_650, signal_649, signal_648, signal_647, signal_236}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_222 ( .a ({signal_1806, signal_1800, signal_1794, signal_1788, signal_1782}), .b ({signal_610, signal_609, signal_608, signal_607, signal_226}), .clk (clk), .r ({Fresh[319], Fresh[318], Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312], Fresh[311], Fresh[310]}), .c ({signal_654, signal_653, signal_652, signal_651, signal_237}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_224 ( .a ({signal_586, signal_585, signal_584, signal_583, signal_220}), .b ({signal_594, signal_593, signal_592, signal_591, signal_222}), .c ({signal_662, signal_661, signal_660, signal_659, signal_239}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_225 ( .a ({signal_590, signal_589, signal_588, signal_587, signal_221}), .b ({signal_602, signal_601, signal_600, signal_599, signal_224}), .c ({signal_666, signal_665, signal_664, signal_663, signal_240}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_226 ( .a ({signal_582, signal_581, signal_580, signal_579, signal_219}), .b ({signal_590, signal_589, signal_588, signal_587, signal_221}), .c ({signal_670, signal_669, signal_668, signal_667, signal_241}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_227 ( .a ({signal_1836, signal_1830, signal_1824, signal_1818, signal_1812}), .b ({signal_658, signal_657, signal_656, signal_655, signal_238}), .clk (clk), .r ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324], Fresh[323], Fresh[322], Fresh[321], Fresh[320]}), .c ({signal_674, signal_673, signal_672, signal_671, signal_242}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_228 ( .a ({signal_1866, signal_1860, signal_1854, signal_1848, signal_1842}), .b ({signal_658, signal_657, signal_656, signal_655, signal_238}), .clk (clk), .r ({Fresh[339], Fresh[338], Fresh[337], Fresh[336], Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .c ({signal_678, signal_677, signal_676, signal_675, signal_243}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_229 ( .a ({signal_582, signal_581, signal_580, signal_579, signal_219}), .b ({signal_626, signal_625, signal_624, signal_623, signal_230}), .c ({signal_682, signal_681, signal_680, signal_679, signal_244}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_230 ( .a ({signal_578, signal_577, signal_576, signal_575, signal_218}), .b ({signal_642, signal_641, signal_640, signal_639, signal_234}), .c ({signal_686, signal_685, signal_684, signal_683, signal_245}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_231 ( .a ({signal_638, signal_637, signal_636, signal_635, signal_233}), .b ({signal_646, signal_645, signal_644, signal_643, signal_235}), .c ({signal_690, signal_689, signal_688, signal_687, signal_246}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_232 ( .a ({signal_630, signal_629, signal_628, signal_627, signal_231}), .b ({signal_650, signal_649, signal_648, signal_647, signal_236}), .c ({signal_694, signal_693, signal_692, signal_691, signal_247}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_233 ( .a ({signal_634, signal_633, signal_632, signal_631, signal_232}), .b ({signal_650, signal_649, signal_648, signal_647, signal_236}), .c ({signal_698, signal_697, signal_696, signal_695, signal_248}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_234 ( .a ({signal_642, signal_641, signal_640, signal_639, signal_234}), .b ({signal_662, signal_661, signal_660, signal_659, signal_239}), .c ({signal_702, signal_701, signal_700, signal_699, signal_249}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_235 ( .a ({signal_598, signal_597, signal_596, signal_595, signal_223}), .b ({signal_662, signal_661, signal_660, signal_659, signal_239}), .c ({signal_706, signal_705, signal_704, signal_703, signal_250}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_236 ( .a ({signal_646, signal_645, signal_644, signal_643, signal_235}), .b ({signal_666, signal_665, signal_664, signal_663, signal_240}), .c ({signal_710, signal_709, signal_708, signal_707, signal_251}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_237 ( .a ({signal_650, signal_649, signal_648, signal_647, signal_236}), .b ({signal_678, signal_677, signal_676, signal_675, signal_243}), .c ({signal_714, signal_713, signal_712, signal_711, signal_252}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_238 ( .a ({signal_678, signal_677, signal_676, signal_675, signal_243}), .b ({signal_694, signal_693, signal_692, signal_691, signal_247}), .c ({signal_718, signal_717, signal_716, signal_715, signal_253}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_239 ( .a ({signal_626, signal_625, signal_624, signal_623, signal_230}), .b ({signal_686, signal_685, signal_684, signal_683, signal_245}), .c ({signal_722, signal_721, signal_720, signal_719, signal_254}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_240 ( .a ({signal_634, signal_633, signal_632, signal_631, signal_232}), .b ({signal_674, signal_673, signal_672, signal_671, signal_242}), .c ({signal_726, signal_725, signal_724, signal_723, signal_255}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_241 ( .a ({signal_674, signal_673, signal_672, signal_671, signal_242}), .b ({signal_690, signal_689, signal_688, signal_687, signal_246}), .c ({signal_730, signal_729, signal_728, signal_727, signal_256}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_242 ( .a ({signal_606, signal_605, signal_604, signal_603, signal_225}), .b ({signal_682, signal_681, signal_680, signal_679, signal_244}), .c ({signal_734, signal_733, signal_732, signal_731, signal_257}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_243 ( .a ({signal_654, signal_653, signal_652, signal_651, signal_237}), .b ({signal_690, signal_689, signal_688, signal_687, signal_246}), .c ({signal_738, signal_737, signal_736, signal_735, signal_258}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_244 ( .a ({signal_670, signal_669, signal_668, signal_667, signal_241}), .b ({signal_686, signal_685, signal_684, signal_683, signal_245}), .c ({signal_742, signal_741, signal_740, signal_739, signal_259}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_245 ( .a ({signal_682, signal_681, signal_680, signal_679, signal_244}), .b ({signal_710, signal_709, signal_708, signal_707, signal_251}), .c ({signal_746, signal_745, signal_744, signal_743, signal_260}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_246 ( .a ({signal_586, signal_585, signal_584, signal_583, signal_220}), .b ({signal_714, signal_713, signal_712, signal_711, signal_252}), .c ({signal_750, signal_749, signal_748, signal_747, signal_261}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_247 ( .a ({signal_594, signal_593, signal_592, signal_591, signal_222}), .b ({signal_714, signal_713, signal_712, signal_711, signal_252}), .c ({signal_754, signal_753, signal_752, signal_751, signal_262}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_248 ( .a ({signal_662, signal_661, signal_660, signal_659, signal_239}), .b ({signal_714, signal_713, signal_712, signal_711, signal_252}), .c ({signal_758, signal_757, signal_756, signal_755, signal_263}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_249 ( .a ({signal_662, signal_661, signal_660, signal_659, signal_239}), .b ({signal_722, signal_721, signal_720, signal_719, signal_254}), .c ({signal_762, signal_761, signal_760, signal_759, signal_264}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_250 ( .a ({signal_702, signal_701, signal_700, signal_699, signal_249}), .b ({signal_726, signal_725, signal_724, signal_723, signal_255}), .c ({signal_766, signal_765, signal_764, signal_763, signal_265}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_251 ( .a ({signal_718, signal_717, signal_716, signal_715, signal_253}), .b ({signal_730, signal_729, signal_728, signal_727, signal_256}), .c ({signal_770, signal_769, signal_768, signal_767, signal_266}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_252 ( .a ({signal_722, signal_721, signal_720, signal_719, signal_254}), .b ({signal_726, signal_725, signal_724, signal_723, signal_255}), .c ({signal_774, signal_773, signal_772, signal_771, signal_267}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_253 ( .a ({signal_666, signal_665, signal_664, signal_663, signal_240}), .b ({signal_730, signal_729, signal_728, signal_727, signal_256}), .c ({signal_778, signal_777, signal_776, signal_775, signal_268}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_254 ( .a ({signal_698, signal_697, signal_696, signal_695, signal_248}), .b ({signal_734, signal_733, signal_732, signal_731, signal_257}), .c ({signal_782, signal_781, signal_780, signal_779, signal_269}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_255 ( .a ({signal_706, signal_705, signal_704, signal_703, signal_250}), .b ({signal_734, signal_733, signal_732, signal_731, signal_257}), .c ({signal_786, signal_785, signal_784, signal_783, signal_270}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_256 ( .a ({signal_718, signal_717, signal_716, signal_715, signal_253}), .b ({signal_746, signal_745, signal_744, signal_743, signal_260}), .c ({signal_790, signal_789, signal_788, signal_787, signal_271}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_257 ( .a ({signal_790, signal_789, signal_788, signal_787, signal_271}), .b ({signal_794, signal_793, signal_792, signal_791, signal_150}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_258 ( .a ({signal_718, signal_717, signal_716, signal_715, signal_253}), .b ({signal_766, signal_765, signal_764, signal_763, signal_265}), .c ({signal_798, signal_797, signal_796, signal_795, signal_143}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_259 ( .a ({signal_754, signal_753, signal_752, signal_751, signal_262}), .b ({signal_774, signal_773, signal_772, signal_771, signal_267}), .c ({signal_802, signal_801, signal_800, signal_799, signal_272}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_260 ( .a ({signal_738, signal_737, signal_736, signal_735, signal_258}), .b ({signal_782, signal_781, signal_780, signal_779, signal_269}), .c ({signal_806, signal_805, signal_804, signal_803, signal_273}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_261 ( .a ({signal_718, signal_717, signal_716, signal_715, signal_253}), .b ({signal_762, signal_761, signal_760, signal_759, signal_264}), .c ({signal_810, signal_809, signal_808, signal_807, signal_146}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_262 ( .a ({signal_742, signal_741, signal_740, signal_739, signal_259}), .b ({signal_758, signal_757, signal_756, signal_755, signal_263}), .c ({signal_814, signal_813, signal_812, signal_811, signal_147}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_263 ( .a ({signal_770, signal_769, signal_768, signal_767, signal_266}), .b ({signal_786, signal_785, signal_784, signal_783, signal_270}), .c ({signal_818, signal_817, signal_816, signal_815, signal_148}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_264 ( .a ({signal_750, signal_749, signal_748, signal_747, signal_261}), .b ({signal_778, signal_777, signal_776, signal_775, signal_268}), .c ({signal_822, signal_821, signal_820, signal_819, signal_274}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_265 ( .a ({signal_802, signal_801, signal_800, signal_799, signal_272}), .b ({signal_826, signal_825, signal_824, signal_823, signal_144}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_266 ( .a ({signal_806, signal_805, signal_804, signal_803, signal_273}), .b ({signal_830, signal_829, signal_828, signal_827, signal_145}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_267 ( .a ({signal_822, signal_821, signal_820, signal_819, signal_274}), .b ({signal_834, signal_833, signal_832, signal_831, signal_149}) ) ;

    /* register cells */
    reg_masked #(.security_order(4), .pipeline(1)) cell_0 ( .clk (clk), .D ({signal_798, signal_797, signal_796, signal_795, signal_143}), .Q ({Y_s4[7], Y_s3[7], Y_s2[7], Y_s1[7], Y_s0[7]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) cell_1 ( .clk (clk), .D ({signal_826, signal_825, signal_824, signal_823, signal_144}), .Q ({Y_s4[6], Y_s3[6], Y_s2[6], Y_s1[6], Y_s0[6]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) cell_2 ( .clk (clk), .D ({signal_830, signal_829, signal_828, signal_827, signal_145}), .Q ({Y_s4[5], Y_s3[5], Y_s2[5], Y_s1[5], Y_s0[5]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) cell_3 ( .clk (clk), .D ({signal_810, signal_809, signal_808, signal_807, signal_146}), .Q ({Y_s4[4], Y_s3[4], Y_s2[4], Y_s1[4], Y_s0[4]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) cell_4 ( .clk (clk), .D ({signal_814, signal_813, signal_812, signal_811, signal_147}), .Q ({Y_s4[3], Y_s3[3], Y_s2[3], Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) cell_5 ( .clk (clk), .D ({signal_818, signal_817, signal_816, signal_815, signal_148}), .Q ({Y_s4[2], Y_s3[2], Y_s2[2], Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) cell_6 ( .clk (clk), .D ({signal_834, signal_833, signal_832, signal_831, signal_149}), .Q ({Y_s4[1], Y_s3[1], Y_s2[1], Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) cell_7 ( .clk (clk), .D ({signal_794, signal_793, signal_792, signal_791, signal_150}), .Q ({Y_s4[0], Y_s3[0], Y_s2[0], Y_s1[0], Y_s0[0]}) ) ;
endmodule
