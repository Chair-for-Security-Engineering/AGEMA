/* modified netlist. Source: module sbox in file Designs/AESSbox/lookup/AGEMA/sbox.v */
/* 34 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 35 register stage(s) in total */

module sbox_HPC1_Pipeline_d3 (SI_s0, clk, SI_s1, SI_s2, SI_s3, Fresh, SO_s0, SO_s1, SO_s2, SO_s3);
    input [7:0] SI_s0 ;
    input clk ;
    input [7:0] SI_s1 ;
    input [7:0] SI_s2 ;
    input [7:0] SI_s3 ;
    input [8679:0] Fresh ;
    output [7:0] SO_s0 ;
    output [7:0] SO_s1 ;
    output [7:0] SO_s2 ;
    output [7:0] SO_s3 ;
    wire N169 ;
    wire N277 ;
    wire N379 ;
    wire N470 ;
    wire N563 ;
    wire N639 ;
    wire N723 ;
    wire N789 ;
    wire n1922 ;
    wire n1923 ;
    wire n1924 ;
    wire n1925 ;
    wire n1926 ;
    wire n1927 ;
    wire n1928 ;
    wire n1929 ;
    wire n1930 ;
    wire n1931 ;
    wire n1932 ;
    wire n1933 ;
    wire n1934 ;
    wire n1935 ;
    wire n1936 ;
    wire n1937 ;
    wire n1938 ;
    wire n1939 ;
    wire n1940 ;
    wire n1941 ;
    wire n1942 ;
    wire n1943 ;
    wire n1944 ;
    wire n1945 ;
    wire n1946 ;
    wire n1947 ;
    wire n1948 ;
    wire n1949 ;
    wire n1950 ;
    wire n1951 ;
    wire n1952 ;
    wire n1953 ;
    wire n1954 ;
    wire n1955 ;
    wire n1956 ;
    wire n1957 ;
    wire n1958 ;
    wire n1959 ;
    wire n1960 ;
    wire n1961 ;
    wire n1962 ;
    wire n1963 ;
    wire n1964 ;
    wire n1965 ;
    wire n1966 ;
    wire n1967 ;
    wire n1968 ;
    wire n1969 ;
    wire n1970 ;
    wire n1971 ;
    wire n1972 ;
    wire n1973 ;
    wire n1974 ;
    wire n1975 ;
    wire n1976 ;
    wire n1977 ;
    wire n1978 ;
    wire n1979 ;
    wire n1980 ;
    wire n1981 ;
    wire n1982 ;
    wire n1983 ;
    wire n1984 ;
    wire n1985 ;
    wire n1986 ;
    wire n1987 ;
    wire n1988 ;
    wire n1989 ;
    wire n1990 ;
    wire n1991 ;
    wire n1992 ;
    wire n1993 ;
    wire n1994 ;
    wire n1995 ;
    wire n1996 ;
    wire n1997 ;
    wire n1998 ;
    wire n1999 ;
    wire n2000 ;
    wire n2001 ;
    wire n2002 ;
    wire n2003 ;
    wire n2004 ;
    wire n2005 ;
    wire n2006 ;
    wire n2007 ;
    wire n2008 ;
    wire n2009 ;
    wire n2010 ;
    wire n2011 ;
    wire n2012 ;
    wire n2013 ;
    wire n2014 ;
    wire n2015 ;
    wire n2016 ;
    wire n2017 ;
    wire n2018 ;
    wire n2019 ;
    wire n2020 ;
    wire n2021 ;
    wire n2022 ;
    wire n2023 ;
    wire n2024 ;
    wire n2025 ;
    wire n2026 ;
    wire n2027 ;
    wire n2028 ;
    wire n2029 ;
    wire n2030 ;
    wire n2031 ;
    wire n2032 ;
    wire n2033 ;
    wire n2034 ;
    wire n2035 ;
    wire n2036 ;
    wire n2037 ;
    wire n2038 ;
    wire n2039 ;
    wire n2040 ;
    wire n2041 ;
    wire n2042 ;
    wire n2043 ;
    wire n2044 ;
    wire n2045 ;
    wire n2046 ;
    wire n2047 ;
    wire n2048 ;
    wire n2049 ;
    wire n2050 ;
    wire n2051 ;
    wire n2052 ;
    wire n2053 ;
    wire n2054 ;
    wire n2055 ;
    wire n2056 ;
    wire n2057 ;
    wire n2058 ;
    wire n2059 ;
    wire n2060 ;
    wire n2061 ;
    wire n2062 ;
    wire n2063 ;
    wire n2064 ;
    wire n2065 ;
    wire n2066 ;
    wire n2067 ;
    wire n2068 ;
    wire n2069 ;
    wire n2070 ;
    wire n2071 ;
    wire n2072 ;
    wire n2073 ;
    wire n2074 ;
    wire n2075 ;
    wire n2076 ;
    wire n2077 ;
    wire n2078 ;
    wire n2079 ;
    wire n2080 ;
    wire n2081 ;
    wire n2082 ;
    wire n2083 ;
    wire n2084 ;
    wire n2085 ;
    wire n2086 ;
    wire n2087 ;
    wire n2088 ;
    wire n2089 ;
    wire n2090 ;
    wire n2091 ;
    wire n2092 ;
    wire n2093 ;
    wire n2094 ;
    wire n2095 ;
    wire n2096 ;
    wire n2097 ;
    wire n2098 ;
    wire n2099 ;
    wire n2100 ;
    wire n2101 ;
    wire n2102 ;
    wire n2103 ;
    wire n2104 ;
    wire n2105 ;
    wire n2106 ;
    wire n2107 ;
    wire n2108 ;
    wire n2109 ;
    wire n2110 ;
    wire n2111 ;
    wire n2112 ;
    wire n2113 ;
    wire n2114 ;
    wire n2115 ;
    wire n2116 ;
    wire n2117 ;
    wire n2118 ;
    wire n2119 ;
    wire n2120 ;
    wire n2121 ;
    wire n2122 ;
    wire n2123 ;
    wire n2124 ;
    wire n2125 ;
    wire n2126 ;
    wire n2127 ;
    wire n2128 ;
    wire n2129 ;
    wire n2130 ;
    wire n2131 ;
    wire n2132 ;
    wire n2133 ;
    wire n2134 ;
    wire n2135 ;
    wire n2136 ;
    wire n2137 ;
    wire n2138 ;
    wire n2139 ;
    wire n2140 ;
    wire n2141 ;
    wire n2142 ;
    wire n2143 ;
    wire n2144 ;
    wire n2145 ;
    wire n2146 ;
    wire n2147 ;
    wire n2148 ;
    wire n2149 ;
    wire n2150 ;
    wire n2151 ;
    wire n2152 ;
    wire n2153 ;
    wire n2154 ;
    wire n2155 ;
    wire n2156 ;
    wire n2157 ;
    wire n2158 ;
    wire n2159 ;
    wire n2160 ;
    wire n2161 ;
    wire n2162 ;
    wire n2163 ;
    wire n2164 ;
    wire n2165 ;
    wire n2166 ;
    wire n2167 ;
    wire n2168 ;
    wire n2169 ;
    wire n2170 ;
    wire n2171 ;
    wire n2172 ;
    wire n2173 ;
    wire n2174 ;
    wire n2175 ;
    wire n2176 ;
    wire n2177 ;
    wire n2178 ;
    wire n2179 ;
    wire n2180 ;
    wire n2181 ;
    wire n2182 ;
    wire n2183 ;
    wire n2184 ;
    wire n2185 ;
    wire n2186 ;
    wire n2187 ;
    wire n2188 ;
    wire n2189 ;
    wire n2190 ;
    wire n2191 ;
    wire n2192 ;
    wire n2193 ;
    wire n2194 ;
    wire n2195 ;
    wire n2196 ;
    wire n2197 ;
    wire n2198 ;
    wire n2199 ;
    wire n2200 ;
    wire n2201 ;
    wire n2202 ;
    wire n2203 ;
    wire n2204 ;
    wire n2205 ;
    wire n2206 ;
    wire n2207 ;
    wire n2208 ;
    wire n2209 ;
    wire n2210 ;
    wire n2211 ;
    wire n2212 ;
    wire n2213 ;
    wire n2214 ;
    wire n2215 ;
    wire n2216 ;
    wire n2217 ;
    wire n2218 ;
    wire n2219 ;
    wire n2220 ;
    wire n2221 ;
    wire n2222 ;
    wire n2223 ;
    wire n2224 ;
    wire n2225 ;
    wire n2226 ;
    wire n2227 ;
    wire n2228 ;
    wire n2229 ;
    wire n2230 ;
    wire n2231 ;
    wire n2232 ;
    wire n2233 ;
    wire n2234 ;
    wire n2235 ;
    wire n2236 ;
    wire n2237 ;
    wire n2238 ;
    wire n2239 ;
    wire n2240 ;
    wire n2241 ;
    wire n2242 ;
    wire n2243 ;
    wire n2244 ;
    wire n2245 ;
    wire n2246 ;
    wire n2247 ;
    wire n2248 ;
    wire n2249 ;
    wire n2250 ;
    wire n2251 ;
    wire n2252 ;
    wire n2253 ;
    wire n2254 ;
    wire n2255 ;
    wire n2256 ;
    wire n2257 ;
    wire n2258 ;
    wire n2259 ;
    wire n2260 ;
    wire n2261 ;
    wire n2262 ;
    wire n2263 ;
    wire n2264 ;
    wire n2265 ;
    wire n2266 ;
    wire n2267 ;
    wire n2268 ;
    wire n2269 ;
    wire n2270 ;
    wire n2271 ;
    wire n2272 ;
    wire n2273 ;
    wire n2274 ;
    wire n2275 ;
    wire n2276 ;
    wire n2277 ;
    wire n2278 ;
    wire n2279 ;
    wire n2280 ;
    wire n2281 ;
    wire n2282 ;
    wire n2283 ;
    wire n2284 ;
    wire n2285 ;
    wire n2286 ;
    wire n2287 ;
    wire n2288 ;
    wire n2289 ;
    wire n2290 ;
    wire n2291 ;
    wire n2292 ;
    wire n2293 ;
    wire n2294 ;
    wire n2295 ;
    wire n2296 ;
    wire n2297 ;
    wire n2298 ;
    wire n2299 ;
    wire n2300 ;
    wire n2301 ;
    wire n2302 ;
    wire n2303 ;
    wire n2304 ;
    wire n2305 ;
    wire n2306 ;
    wire n2307 ;
    wire n2308 ;
    wire n2309 ;
    wire n2310 ;
    wire n2311 ;
    wire n2312 ;
    wire n2313 ;
    wire n2314 ;
    wire n2315 ;
    wire n2316 ;
    wire n2317 ;
    wire n2318 ;
    wire n2319 ;
    wire n2320 ;
    wire n2321 ;
    wire n2322 ;
    wire n2323 ;
    wire n2324 ;
    wire n2325 ;
    wire n2326 ;
    wire n2327 ;
    wire n2328 ;
    wire n2329 ;
    wire n2330 ;
    wire n2331 ;
    wire n2332 ;
    wire n2333 ;
    wire n2334 ;
    wire n2335 ;
    wire n2336 ;
    wire n2337 ;
    wire n2338 ;
    wire n2339 ;
    wire n2340 ;
    wire n2341 ;
    wire n2342 ;
    wire n2343 ;
    wire n2344 ;
    wire n2345 ;
    wire n2346 ;
    wire n2347 ;
    wire n2348 ;
    wire n2349 ;
    wire n2350 ;
    wire n2351 ;
    wire n2352 ;
    wire n2353 ;
    wire n2354 ;
    wire n2355 ;
    wire n2356 ;
    wire n2357 ;
    wire n2358 ;
    wire n2359 ;
    wire n2360 ;
    wire n2361 ;
    wire n2362 ;
    wire n2363 ;
    wire n2364 ;
    wire n2365 ;
    wire n2366 ;
    wire n2367 ;
    wire n2368 ;
    wire n2369 ;
    wire n2370 ;
    wire n2371 ;
    wire n2372 ;
    wire n2373 ;
    wire n2374 ;
    wire n2375 ;
    wire n2376 ;
    wire n2377 ;
    wire n2378 ;
    wire n2379 ;
    wire n2380 ;
    wire n2381 ;
    wire n2382 ;
    wire n2383 ;
    wire n2384 ;
    wire n2385 ;
    wire n2386 ;
    wire n2387 ;
    wire n2388 ;
    wire n2389 ;
    wire n2390 ;
    wire n2391 ;
    wire n2392 ;
    wire n2393 ;
    wire n2394 ;
    wire n2395 ;
    wire n2396 ;
    wire n2397 ;
    wire n2398 ;
    wire n2399 ;
    wire n2400 ;
    wire n2401 ;
    wire n2402 ;
    wire n2403 ;
    wire n2404 ;
    wire n2405 ;
    wire n2406 ;
    wire n2407 ;
    wire n2408 ;
    wire n2409 ;
    wire n2410 ;
    wire n2411 ;
    wire n2412 ;
    wire n2413 ;
    wire n2414 ;
    wire n2415 ;
    wire n2416 ;
    wire n2417 ;
    wire n2418 ;
    wire n2419 ;
    wire n2420 ;
    wire n2421 ;
    wire n2422 ;
    wire n2423 ;
    wire n2424 ;
    wire n2425 ;
    wire n2426 ;
    wire n2427 ;
    wire n2428 ;
    wire n2429 ;
    wire n2430 ;
    wire n2431 ;
    wire n2432 ;
    wire n2433 ;
    wire n2434 ;
    wire n2435 ;
    wire n2436 ;
    wire n2437 ;
    wire n2438 ;
    wire n2439 ;
    wire n2440 ;
    wire n2441 ;
    wire n2442 ;
    wire n2443 ;
    wire n2444 ;
    wire n2445 ;
    wire n2446 ;
    wire n2447 ;
    wire n2448 ;
    wire n2449 ;
    wire n2450 ;
    wire n2451 ;
    wire n2452 ;
    wire n2453 ;
    wire n2454 ;
    wire n2455 ;
    wire n2456 ;
    wire n2457 ;
    wire n2458 ;
    wire n2459 ;
    wire n2460 ;
    wire n2461 ;
    wire n2462 ;
    wire n2463 ;
    wire n2464 ;
    wire n2465 ;
    wire n2466 ;
    wire n2467 ;
    wire n2468 ;
    wire n2469 ;
    wire n2470 ;
    wire n2471 ;
    wire n2472 ;
    wire n2473 ;
    wire n2474 ;
    wire n2475 ;
    wire n2476 ;
    wire n2477 ;
    wire n2478 ;
    wire n2479 ;
    wire n2480 ;
    wire n2481 ;
    wire n2482 ;
    wire n2483 ;
    wire n2484 ;
    wire n2485 ;
    wire n2486 ;
    wire n2487 ;
    wire n2488 ;
    wire n2489 ;
    wire n2490 ;
    wire n2491 ;
    wire n2492 ;
    wire n2493 ;
    wire n2494 ;
    wire n2495 ;
    wire n2496 ;
    wire n2497 ;
    wire n2498 ;
    wire n2499 ;
    wire n2500 ;
    wire n2501 ;
    wire n2502 ;
    wire n2503 ;
    wire n2504 ;
    wire n2505 ;
    wire n2506 ;
    wire n2507 ;
    wire n2508 ;
    wire n2509 ;
    wire n2510 ;
    wire n2511 ;
    wire n2512 ;
    wire n2513 ;
    wire n2514 ;
    wire n2515 ;
    wire n2516 ;
    wire n2517 ;
    wire n2518 ;
    wire n2519 ;
    wire n2520 ;
    wire n2521 ;
    wire n2522 ;
    wire n2523 ;
    wire n2524 ;
    wire n2525 ;
    wire n2526 ;
    wire n2527 ;
    wire n2528 ;
    wire n2529 ;
    wire n2530 ;
    wire n2531 ;
    wire n2532 ;
    wire n2533 ;
    wire n2534 ;
    wire n2535 ;
    wire n2536 ;
    wire n2537 ;
    wire n2538 ;
    wire n2539 ;
    wire n2540 ;
    wire n2541 ;
    wire n2542 ;
    wire n2543 ;
    wire n2544 ;
    wire n2545 ;
    wire n2546 ;
    wire n2547 ;
    wire n2548 ;
    wire n2549 ;
    wire n2550 ;
    wire n2551 ;
    wire n2552 ;
    wire n2553 ;
    wire n2554 ;
    wire n2555 ;
    wire n2556 ;
    wire n2557 ;
    wire n2558 ;
    wire n2559 ;
    wire n2560 ;
    wire n2561 ;
    wire n2562 ;
    wire n2563 ;
    wire n2564 ;
    wire n2565 ;
    wire n2566 ;
    wire n2567 ;
    wire n2568 ;
    wire n2569 ;
    wire n2570 ;
    wire n2571 ;
    wire n2572 ;
    wire n2573 ;
    wire n2574 ;
    wire n2575 ;
    wire n2576 ;
    wire n2577 ;
    wire n2578 ;
    wire n2579 ;
    wire n2580 ;
    wire n2581 ;
    wire n2582 ;
    wire n2583 ;
    wire n2584 ;
    wire n2585 ;
    wire n2586 ;
    wire n2587 ;
    wire n2588 ;
    wire n2589 ;
    wire n2590 ;
    wire n2591 ;
    wire n2592 ;
    wire n2593 ;
    wire n2594 ;
    wire n2595 ;
    wire n2596 ;
    wire n2597 ;
    wire n2598 ;
    wire n2599 ;
    wire n2600 ;
    wire n2601 ;
    wire n2602 ;
    wire n2603 ;
    wire n2604 ;
    wire n2605 ;
    wire n2606 ;
    wire n2607 ;
    wire n2608 ;
    wire n2609 ;
    wire n2610 ;
    wire n2611 ;
    wire n2612 ;
    wire n2613 ;
    wire n2614 ;
    wire n2615 ;
    wire n2616 ;
    wire n2617 ;
    wire n2618 ;
    wire n2619 ;
    wire n2620 ;
    wire n2621 ;
    wire n2622 ;
    wire n2623 ;
    wire n2624 ;
    wire n2625 ;
    wire n2626 ;
    wire n2627 ;
    wire n2628 ;
    wire n2629 ;
    wire n2630 ;
    wire n2631 ;
    wire n2632 ;
    wire n2633 ;
    wire n2634 ;
    wire n2635 ;
    wire n2636 ;
    wire n2637 ;
    wire n2638 ;
    wire n2639 ;
    wire n2640 ;
    wire n2641 ;
    wire n2642 ;
    wire n2643 ;
    wire n2644 ;
    wire n2645 ;
    wire n2646 ;
    wire n2647 ;
    wire n2648 ;
    wire n2649 ;
    wire n2650 ;
    wire n2651 ;
    wire n2652 ;
    wire n2653 ;
    wire n2654 ;
    wire n2655 ;
    wire n2656 ;
    wire n2657 ;
    wire n2658 ;
    wire n2659 ;
    wire n2660 ;
    wire n2661 ;
    wire n2662 ;
    wire n2663 ;
    wire n2664 ;
    wire n2665 ;
    wire n2666 ;
    wire n2667 ;
    wire n2668 ;
    wire n2669 ;
    wire n2670 ;
    wire n2671 ;
    wire n2672 ;
    wire n2673 ;
    wire n2674 ;
    wire n2675 ;
    wire n2676 ;
    wire n2677 ;
    wire n2678 ;
    wire n2679 ;
    wire n2680 ;
    wire n2681 ;
    wire n2682 ;
    wire n2683 ;
    wire n2684 ;
    wire n2685 ;
    wire n2686 ;
    wire n2687 ;
    wire n2688 ;
    wire n2689 ;
    wire n2690 ;
    wire n2691 ;
    wire n2692 ;
    wire n2693 ;
    wire n2694 ;
    wire n2695 ;
    wire n2696 ;
    wire n2697 ;
    wire n2698 ;
    wire n2699 ;
    wire n2700 ;
    wire n2701 ;
    wire n2702 ;
    wire n2703 ;
    wire n2704 ;
    wire n2705 ;
    wire n2706 ;
    wire n2707 ;
    wire n2708 ;
    wire n2709 ;
    wire n2710 ;
    wire n2711 ;
    wire n2712 ;
    wire n2713 ;
    wire n2714 ;
    wire n2715 ;
    wire n2716 ;
    wire n2717 ;
    wire n2718 ;
    wire n2719 ;
    wire n2720 ;
    wire n2721 ;
    wire n2722 ;
    wire n2723 ;
    wire n2724 ;
    wire n2725 ;
    wire n2726 ;
    wire n2727 ;
    wire n2728 ;
    wire n2729 ;
    wire n2730 ;
    wire n2731 ;
    wire n2732 ;
    wire n2733 ;
    wire n2734 ;
    wire n2735 ;
    wire n2736 ;
    wire n2737 ;
    wire n2738 ;
    wire n2739 ;
    wire n2740 ;
    wire n2741 ;
    wire n2742 ;
    wire n2743 ;
    wire n2744 ;
    wire n2745 ;
    wire n2746 ;
    wire n2747 ;
    wire n2748 ;
    wire n2749 ;
    wire n2750 ;
    wire n2751 ;
    wire n2752 ;
    wire n2753 ;
    wire n2754 ;
    wire n2755 ;
    wire n2756 ;
    wire n2757 ;
    wire n2758 ;
    wire n2759 ;
    wire n2760 ;
    wire n2761 ;
    wire n2762 ;
    wire n2763 ;
    wire n2764 ;
    wire n2765 ;
    wire n2766 ;
    wire n2767 ;
    wire n2768 ;
    wire n2769 ;
    wire n2770 ;
    wire n2771 ;
    wire n2772 ;
    wire n2773 ;
    wire n2774 ;
    wire n2775 ;
    wire n2776 ;
    wire n2777 ;
    wire n2778 ;
    wire n2779 ;
    wire n2780 ;
    wire n2781 ;
    wire n2782 ;
    wire n2783 ;
    wire n2784 ;
    wire n2785 ;
    wire n2786 ;
    wire n2787 ;
    wire n2788 ;
    wire n2789 ;
    wire n2790 ;
    wire n2791 ;
    wire n2792 ;
    wire n2793 ;
    wire n2794 ;
    wire n2795 ;
    wire n2796 ;
    wire n2797 ;
    wire n2798 ;
    wire n2799 ;
    wire n2800 ;
    wire n2801 ;
    wire n2802 ;
    wire n2803 ;
    wire n2804 ;
    wire n2805 ;
    wire n2806 ;
    wire n2807 ;
    wire n2808 ;
    wire n2809 ;
    wire n2810 ;
    wire n2811 ;
    wire n2812 ;
    wire n2813 ;
    wire n2814 ;
    wire n2815 ;
    wire n2816 ;
    wire n2817 ;
    wire n2818 ;
    wire n2819 ;
    wire n2820 ;
    wire n2821 ;
    wire n2822 ;
    wire n2823 ;
    wire n2824 ;
    wire n2825 ;
    wire n2826 ;
    wire n2827 ;
    wire n2828 ;
    wire n2829 ;
    wire n2830 ;
    wire n2831 ;
    wire n2832 ;
    wire new_AGEMA_signal_945 ;
    wire new_AGEMA_signal_946 ;
    wire new_AGEMA_signal_947 ;
    wire new_AGEMA_signal_951 ;
    wire new_AGEMA_signal_952 ;
    wire new_AGEMA_signal_953 ;
    wire new_AGEMA_signal_957 ;
    wire new_AGEMA_signal_958 ;
    wire new_AGEMA_signal_959 ;
    wire new_AGEMA_signal_963 ;
    wire new_AGEMA_signal_964 ;
    wire new_AGEMA_signal_965 ;
    wire new_AGEMA_signal_969 ;
    wire new_AGEMA_signal_970 ;
    wire new_AGEMA_signal_971 ;
    wire new_AGEMA_signal_975 ;
    wire new_AGEMA_signal_976 ;
    wire new_AGEMA_signal_977 ;
    wire new_AGEMA_signal_981 ;
    wire new_AGEMA_signal_982 ;
    wire new_AGEMA_signal_983 ;
    wire new_AGEMA_signal_987 ;
    wire new_AGEMA_signal_988 ;
    wire new_AGEMA_signal_989 ;
    wire new_AGEMA_signal_990 ;
    wire new_AGEMA_signal_991 ;
    wire new_AGEMA_signal_992 ;
    wire new_AGEMA_signal_993 ;
    wire new_AGEMA_signal_994 ;
    wire new_AGEMA_signal_995 ;
    wire new_AGEMA_signal_996 ;
    wire new_AGEMA_signal_997 ;
    wire new_AGEMA_signal_998 ;
    wire new_AGEMA_signal_999 ;
    wire new_AGEMA_signal_1000 ;
    wire new_AGEMA_signal_1001 ;
    wire new_AGEMA_signal_1002 ;
    wire new_AGEMA_signal_1003 ;
    wire new_AGEMA_signal_1004 ;
    wire new_AGEMA_signal_1005 ;
    wire new_AGEMA_signal_1006 ;
    wire new_AGEMA_signal_1007 ;
    wire new_AGEMA_signal_1008 ;
    wire new_AGEMA_signal_1009 ;
    wire new_AGEMA_signal_1010 ;
    wire new_AGEMA_signal_1011 ;
    wire new_AGEMA_signal_1012 ;
    wire new_AGEMA_signal_1013 ;
    wire new_AGEMA_signal_1014 ;
    wire new_AGEMA_signal_1015 ;
    wire new_AGEMA_signal_1016 ;
    wire new_AGEMA_signal_1017 ;
    wire new_AGEMA_signal_1018 ;
    wire new_AGEMA_signal_1019 ;
    wire new_AGEMA_signal_1020 ;
    wire new_AGEMA_signal_1021 ;
    wire new_AGEMA_signal_1022 ;
    wire new_AGEMA_signal_1023 ;
    wire new_AGEMA_signal_1024 ;
    wire new_AGEMA_signal_1025 ;
    wire new_AGEMA_signal_1026 ;
    wire new_AGEMA_signal_1027 ;
    wire new_AGEMA_signal_1028 ;
    wire new_AGEMA_signal_1029 ;
    wire new_AGEMA_signal_1030 ;
    wire new_AGEMA_signal_1031 ;
    wire new_AGEMA_signal_1032 ;
    wire new_AGEMA_signal_1033 ;
    wire new_AGEMA_signal_1034 ;
    wire new_AGEMA_signal_1035 ;
    wire new_AGEMA_signal_1036 ;
    wire new_AGEMA_signal_1037 ;
    wire new_AGEMA_signal_1038 ;
    wire new_AGEMA_signal_1039 ;
    wire new_AGEMA_signal_1040 ;
    wire new_AGEMA_signal_1041 ;
    wire new_AGEMA_signal_1042 ;
    wire new_AGEMA_signal_1043 ;
    wire new_AGEMA_signal_1044 ;
    wire new_AGEMA_signal_1045 ;
    wire new_AGEMA_signal_1046 ;
    wire new_AGEMA_signal_1047 ;
    wire new_AGEMA_signal_1048 ;
    wire new_AGEMA_signal_1049 ;
    wire new_AGEMA_signal_1050 ;
    wire new_AGEMA_signal_1051 ;
    wire new_AGEMA_signal_1052 ;
    wire new_AGEMA_signal_1053 ;
    wire new_AGEMA_signal_1054 ;
    wire new_AGEMA_signal_1055 ;
    wire new_AGEMA_signal_1056 ;
    wire new_AGEMA_signal_1057 ;
    wire new_AGEMA_signal_1058 ;
    wire new_AGEMA_signal_1059 ;
    wire new_AGEMA_signal_1060 ;
    wire new_AGEMA_signal_1061 ;
    wire new_AGEMA_signal_1062 ;
    wire new_AGEMA_signal_1063 ;
    wire new_AGEMA_signal_1064 ;
    wire new_AGEMA_signal_1065 ;
    wire new_AGEMA_signal_1066 ;
    wire new_AGEMA_signal_1067 ;
    wire new_AGEMA_signal_1068 ;
    wire new_AGEMA_signal_1069 ;
    wire new_AGEMA_signal_1070 ;
    wire new_AGEMA_signal_1071 ;
    wire new_AGEMA_signal_1072 ;
    wire new_AGEMA_signal_1073 ;
    wire new_AGEMA_signal_1074 ;
    wire new_AGEMA_signal_1075 ;
    wire new_AGEMA_signal_1076 ;
    wire new_AGEMA_signal_1077 ;
    wire new_AGEMA_signal_1078 ;
    wire new_AGEMA_signal_1079 ;
    wire new_AGEMA_signal_1080 ;
    wire new_AGEMA_signal_1081 ;
    wire new_AGEMA_signal_1082 ;
    wire new_AGEMA_signal_1083 ;
    wire new_AGEMA_signal_1084 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1086 ;
    wire new_AGEMA_signal_1087 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1089 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1091 ;
    wire new_AGEMA_signal_1092 ;
    wire new_AGEMA_signal_1093 ;
    wire new_AGEMA_signal_1094 ;
    wire new_AGEMA_signal_1095 ;
    wire new_AGEMA_signal_1096 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1098 ;
    wire new_AGEMA_signal_1099 ;
    wire new_AGEMA_signal_1100 ;
    wire new_AGEMA_signal_1101 ;
    wire new_AGEMA_signal_1102 ;
    wire new_AGEMA_signal_1103 ;
    wire new_AGEMA_signal_1104 ;
    wire new_AGEMA_signal_1105 ;
    wire new_AGEMA_signal_1106 ;
    wire new_AGEMA_signal_1107 ;
    wire new_AGEMA_signal_1108 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1110 ;
    wire new_AGEMA_signal_1111 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1113 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1115 ;
    wire new_AGEMA_signal_1116 ;
    wire new_AGEMA_signal_1117 ;
    wire new_AGEMA_signal_1118 ;
    wire new_AGEMA_signal_1119 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1121 ;
    wire new_AGEMA_signal_1122 ;
    wire new_AGEMA_signal_1123 ;
    wire new_AGEMA_signal_1124 ;
    wire new_AGEMA_signal_1125 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1127 ;
    wire new_AGEMA_signal_1128 ;
    wire new_AGEMA_signal_1129 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1131 ;
    wire new_AGEMA_signal_1132 ;
    wire new_AGEMA_signal_1133 ;
    wire new_AGEMA_signal_1134 ;
    wire new_AGEMA_signal_1135 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1137 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1139 ;
    wire new_AGEMA_signal_1140 ;
    wire new_AGEMA_signal_1141 ;
    wire new_AGEMA_signal_1142 ;
    wire new_AGEMA_signal_1143 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1146 ;
    wire new_AGEMA_signal_1147 ;
    wire new_AGEMA_signal_1148 ;
    wire new_AGEMA_signal_1149 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1152 ;
    wire new_AGEMA_signal_1153 ;
    wire new_AGEMA_signal_1154 ;
    wire new_AGEMA_signal_1155 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1158 ;
    wire new_AGEMA_signal_1159 ;
    wire new_AGEMA_signal_1160 ;
    wire new_AGEMA_signal_1161 ;
    wire new_AGEMA_signal_1162 ;
    wire new_AGEMA_signal_1163 ;
    wire new_AGEMA_signal_1164 ;
    wire new_AGEMA_signal_1165 ;
    wire new_AGEMA_signal_1166 ;
    wire new_AGEMA_signal_1167 ;
    wire new_AGEMA_signal_1168 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1170 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1172 ;
    wire new_AGEMA_signal_1173 ;
    wire new_AGEMA_signal_1174 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1176 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1179 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1182 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1184 ;
    wire new_AGEMA_signal_1185 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1188 ;
    wire new_AGEMA_signal_1189 ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1192 ;
    wire new_AGEMA_signal_1193 ;
    wire new_AGEMA_signal_1194 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1196 ;
    wire new_AGEMA_signal_1197 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1200 ;
    wire new_AGEMA_signal_1201 ;
    wire new_AGEMA_signal_1202 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1206 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1208 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1211 ;
    wire new_AGEMA_signal_1212 ;
    wire new_AGEMA_signal_1213 ;
    wire new_AGEMA_signal_1214 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1217 ;
    wire new_AGEMA_signal_1218 ;
    wire new_AGEMA_signal_1219 ;
    wire new_AGEMA_signal_1220 ;
    wire new_AGEMA_signal_1221 ;
    wire new_AGEMA_signal_1222 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1224 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1227 ;
    wire new_AGEMA_signal_1228 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1230 ;
    wire new_AGEMA_signal_1231 ;
    wire new_AGEMA_signal_1232 ;
    wire new_AGEMA_signal_1233 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1236 ;
    wire new_AGEMA_signal_1237 ;
    wire new_AGEMA_signal_1238 ;
    wire new_AGEMA_signal_1239 ;
    wire new_AGEMA_signal_1240 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1242 ;
    wire new_AGEMA_signal_1243 ;
    wire new_AGEMA_signal_1244 ;
    wire new_AGEMA_signal_1245 ;
    wire new_AGEMA_signal_1246 ;
    wire new_AGEMA_signal_1247 ;
    wire new_AGEMA_signal_1248 ;
    wire new_AGEMA_signal_1249 ;
    wire new_AGEMA_signal_1250 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1252 ;
    wire new_AGEMA_signal_1253 ;
    wire new_AGEMA_signal_1254 ;
    wire new_AGEMA_signal_1255 ;
    wire new_AGEMA_signal_1256 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1259 ;
    wire new_AGEMA_signal_1260 ;
    wire new_AGEMA_signal_1261 ;
    wire new_AGEMA_signal_1262 ;
    wire new_AGEMA_signal_1263 ;
    wire new_AGEMA_signal_1264 ;
    wire new_AGEMA_signal_1265 ;
    wire new_AGEMA_signal_1266 ;
    wire new_AGEMA_signal_1267 ;
    wire new_AGEMA_signal_1268 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1270 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1272 ;
    wire new_AGEMA_signal_1273 ;
    wire new_AGEMA_signal_1274 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1276 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1278 ;
    wire new_AGEMA_signal_1279 ;
    wire new_AGEMA_signal_1280 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1282 ;
    wire new_AGEMA_signal_1283 ;
    wire new_AGEMA_signal_1284 ;
    wire new_AGEMA_signal_1285 ;
    wire new_AGEMA_signal_1286 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1288 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1291 ;
    wire new_AGEMA_signal_1292 ;
    wire new_AGEMA_signal_1293 ;
    wire new_AGEMA_signal_1294 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1296 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1300 ;
    wire new_AGEMA_signal_1301 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1304 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1308 ;
    wire new_AGEMA_signal_1309 ;
    wire new_AGEMA_signal_1310 ;
    wire new_AGEMA_signal_1311 ;
    wire new_AGEMA_signal_1312 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1316 ;
    wire new_AGEMA_signal_1317 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1320 ;
    wire new_AGEMA_signal_1321 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1326 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1344 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1352 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1364 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1381 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1400 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1412 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1441 ;
    wire new_AGEMA_signal_1442 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1444 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1456 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1459 ;
    wire new_AGEMA_signal_1460 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1465 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1471 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1474 ;
    wire new_AGEMA_signal_1475 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1483 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1492 ;
    wire new_AGEMA_signal_1493 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1501 ;
    wire new_AGEMA_signal_1502 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1510 ;
    wire new_AGEMA_signal_1511 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1519 ;
    wire new_AGEMA_signal_1520 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1522 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1528 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1547 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1555 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1559 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1563 ;
    wire new_AGEMA_signal_1564 ;
    wire new_AGEMA_signal_1565 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1573 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1579 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1581 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1583 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1591 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1593 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1599 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1609 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1619 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1627 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1645 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1653 ;
    wire new_AGEMA_signal_1654 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1663 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1699 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1701 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1789 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1799 ;
    wire new_AGEMA_signal_1800 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1835 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1870 ;
    wire new_AGEMA_signal_1871 ;
    wire new_AGEMA_signal_1872 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1880 ;
    wire new_AGEMA_signal_1881 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1888 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1896 ;
    wire new_AGEMA_signal_1897 ;
    wire new_AGEMA_signal_1898 ;
    wire new_AGEMA_signal_1899 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1906 ;
    wire new_AGEMA_signal_1907 ;
    wire new_AGEMA_signal_1908 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1914 ;
    wire new_AGEMA_signal_1915 ;
    wire new_AGEMA_signal_1916 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1923 ;
    wire new_AGEMA_signal_1924 ;
    wire new_AGEMA_signal_1925 ;
    wire new_AGEMA_signal_1926 ;
    wire new_AGEMA_signal_1927 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1931 ;
    wire new_AGEMA_signal_1932 ;
    wire new_AGEMA_signal_1933 ;
    wire new_AGEMA_signal_1934 ;
    wire new_AGEMA_signal_1935 ;
    wire new_AGEMA_signal_1936 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1938 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1940 ;
    wire new_AGEMA_signal_1941 ;
    wire new_AGEMA_signal_1942 ;
    wire new_AGEMA_signal_1943 ;
    wire new_AGEMA_signal_1944 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1947 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1949 ;
    wire new_AGEMA_signal_1950 ;
    wire new_AGEMA_signal_1951 ;
    wire new_AGEMA_signal_1952 ;
    wire new_AGEMA_signal_1953 ;
    wire new_AGEMA_signal_1954 ;
    wire new_AGEMA_signal_1955 ;
    wire new_AGEMA_signal_1956 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1958 ;
    wire new_AGEMA_signal_1959 ;
    wire new_AGEMA_signal_1960 ;
    wire new_AGEMA_signal_1961 ;
    wire new_AGEMA_signal_1962 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1967 ;
    wire new_AGEMA_signal_1968 ;
    wire new_AGEMA_signal_1969 ;
    wire new_AGEMA_signal_1970 ;
    wire new_AGEMA_signal_1971 ;
    wire new_AGEMA_signal_1972 ;
    wire new_AGEMA_signal_1973 ;
    wire new_AGEMA_signal_1974 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1976 ;
    wire new_AGEMA_signal_1977 ;
    wire new_AGEMA_signal_1978 ;
    wire new_AGEMA_signal_1979 ;
    wire new_AGEMA_signal_1980 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1985 ;
    wire new_AGEMA_signal_1986 ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1988 ;
    wire new_AGEMA_signal_1989 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1995 ;
    wire new_AGEMA_signal_1996 ;
    wire new_AGEMA_signal_1997 ;
    wire new_AGEMA_signal_1998 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2003 ;
    wire new_AGEMA_signal_2004 ;
    wire new_AGEMA_signal_2005 ;
    wire new_AGEMA_signal_2006 ;
    wire new_AGEMA_signal_2007 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2014 ;
    wire new_AGEMA_signal_2015 ;
    wire new_AGEMA_signal_2016 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2022 ;
    wire new_AGEMA_signal_2023 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2025 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2032 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2034 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2041 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2043 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2050 ;
    wire new_AGEMA_signal_2051 ;
    wire new_AGEMA_signal_2052 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2059 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2061 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2086 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2097 ;
    wire new_AGEMA_signal_2098 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2102 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2104 ;
    wire new_AGEMA_signal_2105 ;
    wire new_AGEMA_signal_2106 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2114 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2116 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2120 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2122 ;
    wire new_AGEMA_signal_2123 ;
    wire new_AGEMA_signal_2124 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2127 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2130 ;
    wire new_AGEMA_signal_2131 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2133 ;
    wire new_AGEMA_signal_2134 ;
    wire new_AGEMA_signal_2135 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2139 ;
    wire new_AGEMA_signal_2140 ;
    wire new_AGEMA_signal_2141 ;
    wire new_AGEMA_signal_2142 ;
    wire new_AGEMA_signal_2143 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2147 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2150 ;
    wire new_AGEMA_signal_2151 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2154 ;
    wire new_AGEMA_signal_2155 ;
    wire new_AGEMA_signal_2156 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2158 ;
    wire new_AGEMA_signal_2159 ;
    wire new_AGEMA_signal_2160 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2166 ;
    wire new_AGEMA_signal_2167 ;
    wire new_AGEMA_signal_2168 ;
    wire new_AGEMA_signal_2169 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2171 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2175 ;
    wire new_AGEMA_signal_2176 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2178 ;
    wire new_AGEMA_signal_2179 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2183 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2186 ;
    wire new_AGEMA_signal_2187 ;
    wire new_AGEMA_signal_2188 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2191 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2194 ;
    wire new_AGEMA_signal_2195 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2199 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2203 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2205 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2209 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2211 ;
    wire new_AGEMA_signal_2212 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2214 ;
    wire new_AGEMA_signal_2215 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2221 ;
    wire new_AGEMA_signal_2222 ;
    wire new_AGEMA_signal_2223 ;
    wire new_AGEMA_signal_2224 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2226 ;
    wire new_AGEMA_signal_2227 ;
    wire new_AGEMA_signal_2228 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2230 ;
    wire new_AGEMA_signal_2231 ;
    wire new_AGEMA_signal_2232 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2235 ;
    wire new_AGEMA_signal_2236 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2239 ;
    wire new_AGEMA_signal_2240 ;
    wire new_AGEMA_signal_2241 ;
    wire new_AGEMA_signal_2242 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2247 ;
    wire new_AGEMA_signal_2248 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2250 ;
    wire new_AGEMA_signal_2251 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2259 ;
    wire new_AGEMA_signal_2260 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2262 ;
    wire new_AGEMA_signal_2263 ;
    wire new_AGEMA_signal_2264 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2266 ;
    wire new_AGEMA_signal_2267 ;
    wire new_AGEMA_signal_2268 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2271 ;
    wire new_AGEMA_signal_2272 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2275 ;
    wire new_AGEMA_signal_2276 ;
    wire new_AGEMA_signal_2277 ;
    wire new_AGEMA_signal_2278 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2280 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2282 ;
    wire new_AGEMA_signal_2283 ;
    wire new_AGEMA_signal_2284 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2286 ;
    wire new_AGEMA_signal_2287 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2290 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2294 ;
    wire new_AGEMA_signal_2295 ;
    wire new_AGEMA_signal_2296 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2298 ;
    wire new_AGEMA_signal_2299 ;
    wire new_AGEMA_signal_2300 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2302 ;
    wire new_AGEMA_signal_2303 ;
    wire new_AGEMA_signal_2304 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2307 ;
    wire new_AGEMA_signal_2308 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2311 ;
    wire new_AGEMA_signal_2312 ;
    wire new_AGEMA_signal_2313 ;
    wire new_AGEMA_signal_2314 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2319 ;
    wire new_AGEMA_signal_2320 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2322 ;
    wire new_AGEMA_signal_2323 ;
    wire new_AGEMA_signal_2324 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2326 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2330 ;
    wire new_AGEMA_signal_2331 ;
    wire new_AGEMA_signal_2332 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2334 ;
    wire new_AGEMA_signal_2335 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2350 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2367 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2371 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2375 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2392 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2826 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2914 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2926 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2934 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2942 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2950 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2962 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2966 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2970 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2976 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2988 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2992 ;
    wire new_AGEMA_signal_2993 ;
    wire new_AGEMA_signal_2994 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2996 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3000 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3004 ;
    wire new_AGEMA_signal_3005 ;
    wire new_AGEMA_signal_3006 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3012 ;
    wire new_AGEMA_signal_3013 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3016 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3020 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3022 ;
    wire new_AGEMA_signal_3023 ;
    wire new_AGEMA_signal_3024 ;
    wire new_AGEMA_signal_3025 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3028 ;
    wire new_AGEMA_signal_3029 ;
    wire new_AGEMA_signal_3030 ;
    wire new_AGEMA_signal_3031 ;
    wire new_AGEMA_signal_3032 ;
    wire new_AGEMA_signal_3033 ;
    wire new_AGEMA_signal_3034 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3036 ;
    wire new_AGEMA_signal_3037 ;
    wire new_AGEMA_signal_3038 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3040 ;
    wire new_AGEMA_signal_3041 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3043 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3047 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3049 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3051 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3055 ;
    wire new_AGEMA_signal_3056 ;
    wire new_AGEMA_signal_3057 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3059 ;
    wire new_AGEMA_signal_3060 ;
    wire new_AGEMA_signal_3061 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3065 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3067 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3069 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3073 ;
    wire new_AGEMA_signal_3074 ;
    wire new_AGEMA_signal_3075 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3077 ;
    wire new_AGEMA_signal_3078 ;
    wire new_AGEMA_signal_3079 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3083 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3085 ;
    wire new_AGEMA_signal_3086 ;
    wire new_AGEMA_signal_3087 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3132 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3139 ;
    wire new_AGEMA_signal_3140 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3248 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3256 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3374 ;
    wire new_AGEMA_signal_3375 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3391 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3411 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3418 ;
    wire new_AGEMA_signal_3419 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3423 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3427 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3447 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3483 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3502 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3561 ;
    wire new_AGEMA_signal_3562 ;
    wire new_AGEMA_signal_3563 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3567 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3569 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3571 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3579 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3583 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3587 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3590 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3615 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3617 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3623 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3634 ;
    wire new_AGEMA_signal_3635 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3659 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_12427 ;
    wire new_AGEMA_signal_12428 ;
    wire new_AGEMA_signal_12429 ;
    wire new_AGEMA_signal_12430 ;
    wire new_AGEMA_signal_12431 ;
    wire new_AGEMA_signal_12432 ;
    wire new_AGEMA_signal_12433 ;
    wire new_AGEMA_signal_12434 ;
    wire new_AGEMA_signal_12435 ;
    wire new_AGEMA_signal_12436 ;
    wire new_AGEMA_signal_12437 ;
    wire new_AGEMA_signal_12438 ;
    wire new_AGEMA_signal_12439 ;
    wire new_AGEMA_signal_12440 ;
    wire new_AGEMA_signal_12441 ;
    wire new_AGEMA_signal_12442 ;
    wire new_AGEMA_signal_12443 ;
    wire new_AGEMA_signal_12444 ;
    wire new_AGEMA_signal_12445 ;
    wire new_AGEMA_signal_12446 ;
    wire new_AGEMA_signal_12447 ;
    wire new_AGEMA_signal_12448 ;
    wire new_AGEMA_signal_12449 ;
    wire new_AGEMA_signal_12450 ;
    wire new_AGEMA_signal_12451 ;
    wire new_AGEMA_signal_12452 ;
    wire new_AGEMA_signal_12453 ;
    wire new_AGEMA_signal_12454 ;
    wire new_AGEMA_signal_12455 ;
    wire new_AGEMA_signal_12456 ;
    wire new_AGEMA_signal_12457 ;
    wire new_AGEMA_signal_12458 ;
    wire new_AGEMA_signal_12459 ;
    wire new_AGEMA_signal_12460 ;
    wire new_AGEMA_signal_12461 ;
    wire new_AGEMA_signal_12462 ;
    wire new_AGEMA_signal_12463 ;
    wire new_AGEMA_signal_12464 ;
    wire new_AGEMA_signal_12465 ;
    wire new_AGEMA_signal_12466 ;
    wire new_AGEMA_signal_12467 ;
    wire new_AGEMA_signal_12468 ;
    wire new_AGEMA_signal_12469 ;
    wire new_AGEMA_signal_12470 ;
    wire new_AGEMA_signal_12471 ;
    wire new_AGEMA_signal_12472 ;
    wire new_AGEMA_signal_12473 ;
    wire new_AGEMA_signal_12474 ;
    wire new_AGEMA_signal_12475 ;
    wire new_AGEMA_signal_12476 ;
    wire new_AGEMA_signal_12477 ;
    wire new_AGEMA_signal_12478 ;
    wire new_AGEMA_signal_12479 ;
    wire new_AGEMA_signal_12480 ;
    wire new_AGEMA_signal_12481 ;
    wire new_AGEMA_signal_12482 ;
    wire new_AGEMA_signal_12483 ;
    wire new_AGEMA_signal_12484 ;
    wire new_AGEMA_signal_12485 ;
    wire new_AGEMA_signal_12486 ;
    wire new_AGEMA_signal_12487 ;
    wire new_AGEMA_signal_12488 ;
    wire new_AGEMA_signal_12489 ;
    wire new_AGEMA_signal_12490 ;
    wire new_AGEMA_signal_12491 ;
    wire new_AGEMA_signal_12492 ;
    wire new_AGEMA_signal_12493 ;
    wire new_AGEMA_signal_12494 ;
    wire new_AGEMA_signal_12495 ;
    wire new_AGEMA_signal_12496 ;
    wire new_AGEMA_signal_12497 ;
    wire new_AGEMA_signal_12498 ;
    wire new_AGEMA_signal_12499 ;
    wire new_AGEMA_signal_12500 ;
    wire new_AGEMA_signal_12501 ;
    wire new_AGEMA_signal_12502 ;
    wire new_AGEMA_signal_12503 ;
    wire new_AGEMA_signal_12504 ;
    wire new_AGEMA_signal_12505 ;
    wire new_AGEMA_signal_12506 ;
    wire new_AGEMA_signal_12507 ;
    wire new_AGEMA_signal_12508 ;
    wire new_AGEMA_signal_12509 ;
    wire new_AGEMA_signal_12510 ;
    wire new_AGEMA_signal_12511 ;
    wire new_AGEMA_signal_12512 ;
    wire new_AGEMA_signal_12513 ;
    wire new_AGEMA_signal_12514 ;
    wire new_AGEMA_signal_12515 ;
    wire new_AGEMA_signal_12516 ;
    wire new_AGEMA_signal_12517 ;
    wire new_AGEMA_signal_12518 ;
    wire new_AGEMA_signal_12519 ;
    wire new_AGEMA_signal_12520 ;
    wire new_AGEMA_signal_12521 ;
    wire new_AGEMA_signal_12522 ;
    wire new_AGEMA_signal_12523 ;
    wire new_AGEMA_signal_12524 ;
    wire new_AGEMA_signal_12525 ;
    wire new_AGEMA_signal_12526 ;
    wire new_AGEMA_signal_12527 ;
    wire new_AGEMA_signal_12528 ;
    wire new_AGEMA_signal_12529 ;
    wire new_AGEMA_signal_12530 ;
    wire new_AGEMA_signal_12531 ;
    wire new_AGEMA_signal_12532 ;
    wire new_AGEMA_signal_12533 ;
    wire new_AGEMA_signal_12534 ;
    wire new_AGEMA_signal_12535 ;
    wire new_AGEMA_signal_12536 ;
    wire new_AGEMA_signal_12537 ;
    wire new_AGEMA_signal_12538 ;
    wire new_AGEMA_signal_12539 ;
    wire new_AGEMA_signal_12540 ;
    wire new_AGEMA_signal_12541 ;
    wire new_AGEMA_signal_12542 ;
    wire new_AGEMA_signal_12543 ;
    wire new_AGEMA_signal_12544 ;
    wire new_AGEMA_signal_12545 ;
    wire new_AGEMA_signal_12546 ;
    wire new_AGEMA_signal_12547 ;
    wire new_AGEMA_signal_12548 ;
    wire new_AGEMA_signal_12549 ;
    wire new_AGEMA_signal_12550 ;
    wire new_AGEMA_signal_12551 ;
    wire new_AGEMA_signal_12552 ;
    wire new_AGEMA_signal_12553 ;
    wire new_AGEMA_signal_12554 ;
    wire new_AGEMA_signal_12555 ;
    wire new_AGEMA_signal_12556 ;
    wire new_AGEMA_signal_12557 ;
    wire new_AGEMA_signal_12558 ;
    wire new_AGEMA_signal_12559 ;
    wire new_AGEMA_signal_12560 ;
    wire new_AGEMA_signal_12561 ;
    wire new_AGEMA_signal_12562 ;
    wire new_AGEMA_signal_12563 ;
    wire new_AGEMA_signal_12564 ;
    wire new_AGEMA_signal_12565 ;
    wire new_AGEMA_signal_12566 ;
    wire new_AGEMA_signal_12567 ;
    wire new_AGEMA_signal_12568 ;
    wire new_AGEMA_signal_12569 ;
    wire new_AGEMA_signal_12570 ;
    wire new_AGEMA_signal_12571 ;
    wire new_AGEMA_signal_12572 ;
    wire new_AGEMA_signal_12573 ;
    wire new_AGEMA_signal_12574 ;
    wire new_AGEMA_signal_12575 ;
    wire new_AGEMA_signal_12576 ;
    wire new_AGEMA_signal_12577 ;
    wire new_AGEMA_signal_12578 ;
    wire new_AGEMA_signal_12579 ;
    wire new_AGEMA_signal_12580 ;
    wire new_AGEMA_signal_12581 ;
    wire new_AGEMA_signal_12582 ;
    wire new_AGEMA_signal_12583 ;
    wire new_AGEMA_signal_12584 ;
    wire new_AGEMA_signal_12585 ;
    wire new_AGEMA_signal_12586 ;
    wire new_AGEMA_signal_12587 ;
    wire new_AGEMA_signal_12588 ;
    wire new_AGEMA_signal_12589 ;
    wire new_AGEMA_signal_12590 ;
    wire new_AGEMA_signal_12591 ;
    wire new_AGEMA_signal_12592 ;
    wire new_AGEMA_signal_12593 ;
    wire new_AGEMA_signal_12594 ;
    wire new_AGEMA_signal_12595 ;
    wire new_AGEMA_signal_12596 ;
    wire new_AGEMA_signal_12597 ;
    wire new_AGEMA_signal_12598 ;
    wire new_AGEMA_signal_12599 ;
    wire new_AGEMA_signal_12600 ;
    wire new_AGEMA_signal_12601 ;
    wire new_AGEMA_signal_12602 ;
    wire new_AGEMA_signal_12603 ;
    wire new_AGEMA_signal_12604 ;
    wire new_AGEMA_signal_12605 ;
    wire new_AGEMA_signal_12606 ;
    wire new_AGEMA_signal_12607 ;
    wire new_AGEMA_signal_12608 ;
    wire new_AGEMA_signal_12609 ;
    wire new_AGEMA_signal_12610 ;
    wire new_AGEMA_signal_12611 ;
    wire new_AGEMA_signal_12612 ;
    wire new_AGEMA_signal_12613 ;
    wire new_AGEMA_signal_12614 ;
    wire new_AGEMA_signal_12615 ;
    wire new_AGEMA_signal_12616 ;
    wire new_AGEMA_signal_12617 ;
    wire new_AGEMA_signal_12618 ;
    wire new_AGEMA_signal_12619 ;
    wire new_AGEMA_signal_12620 ;
    wire new_AGEMA_signal_12621 ;
    wire new_AGEMA_signal_12622 ;
    wire new_AGEMA_signal_12623 ;
    wire new_AGEMA_signal_12624 ;
    wire new_AGEMA_signal_12625 ;
    wire new_AGEMA_signal_12626 ;
    wire new_AGEMA_signal_12627 ;
    wire new_AGEMA_signal_12628 ;
    wire new_AGEMA_signal_12629 ;
    wire new_AGEMA_signal_12630 ;
    wire new_AGEMA_signal_12631 ;
    wire new_AGEMA_signal_12632 ;
    wire new_AGEMA_signal_12633 ;
    wire new_AGEMA_signal_12634 ;
    wire new_AGEMA_signal_12635 ;
    wire new_AGEMA_signal_12636 ;
    wire new_AGEMA_signal_12637 ;
    wire new_AGEMA_signal_12638 ;
    wire new_AGEMA_signal_12639 ;
    wire new_AGEMA_signal_12640 ;
    wire new_AGEMA_signal_12641 ;
    wire new_AGEMA_signal_12642 ;
    wire new_AGEMA_signal_12643 ;
    wire new_AGEMA_signal_12644 ;
    wire new_AGEMA_signal_12645 ;
    wire new_AGEMA_signal_12646 ;
    wire new_AGEMA_signal_12647 ;
    wire new_AGEMA_signal_12648 ;
    wire new_AGEMA_signal_12649 ;
    wire new_AGEMA_signal_12650 ;
    wire new_AGEMA_signal_12651 ;
    wire new_AGEMA_signal_12652 ;
    wire new_AGEMA_signal_12653 ;
    wire new_AGEMA_signal_12654 ;
    wire new_AGEMA_signal_12655 ;
    wire new_AGEMA_signal_12656 ;
    wire new_AGEMA_signal_12657 ;
    wire new_AGEMA_signal_12658 ;
    wire new_AGEMA_signal_12659 ;
    wire new_AGEMA_signal_12660 ;
    wire new_AGEMA_signal_12661 ;
    wire new_AGEMA_signal_12662 ;
    wire new_AGEMA_signal_12663 ;
    wire new_AGEMA_signal_12664 ;
    wire new_AGEMA_signal_12665 ;
    wire new_AGEMA_signal_12666 ;
    wire new_AGEMA_signal_12667 ;
    wire new_AGEMA_signal_12668 ;
    wire new_AGEMA_signal_12669 ;
    wire new_AGEMA_signal_12670 ;
    wire new_AGEMA_signal_12671 ;
    wire new_AGEMA_signal_12672 ;
    wire new_AGEMA_signal_12673 ;
    wire new_AGEMA_signal_12674 ;
    wire new_AGEMA_signal_12675 ;
    wire new_AGEMA_signal_12676 ;
    wire new_AGEMA_signal_12677 ;
    wire new_AGEMA_signal_12678 ;
    wire new_AGEMA_signal_12679 ;
    wire new_AGEMA_signal_12680 ;
    wire new_AGEMA_signal_12681 ;
    wire new_AGEMA_signal_12682 ;
    wire new_AGEMA_signal_12683 ;
    wire new_AGEMA_signal_12684 ;
    wire new_AGEMA_signal_12685 ;
    wire new_AGEMA_signal_12686 ;
    wire new_AGEMA_signal_12687 ;
    wire new_AGEMA_signal_12688 ;
    wire new_AGEMA_signal_12689 ;
    wire new_AGEMA_signal_12690 ;
    wire new_AGEMA_signal_12691 ;
    wire new_AGEMA_signal_12692 ;
    wire new_AGEMA_signal_12693 ;
    wire new_AGEMA_signal_12694 ;
    wire new_AGEMA_signal_12695 ;
    wire new_AGEMA_signal_12696 ;
    wire new_AGEMA_signal_12697 ;
    wire new_AGEMA_signal_12698 ;
    wire new_AGEMA_signal_12699 ;
    wire new_AGEMA_signal_12700 ;
    wire new_AGEMA_signal_12701 ;
    wire new_AGEMA_signal_12702 ;
    wire new_AGEMA_signal_12703 ;
    wire new_AGEMA_signal_12704 ;
    wire new_AGEMA_signal_12705 ;
    wire new_AGEMA_signal_12706 ;
    wire new_AGEMA_signal_12707 ;
    wire new_AGEMA_signal_12708 ;
    wire new_AGEMA_signal_12709 ;
    wire new_AGEMA_signal_12710 ;
    wire new_AGEMA_signal_12711 ;
    wire new_AGEMA_signal_12712 ;
    wire new_AGEMA_signal_12713 ;
    wire new_AGEMA_signal_12714 ;
    wire new_AGEMA_signal_12715 ;
    wire new_AGEMA_signal_12716 ;
    wire new_AGEMA_signal_12717 ;
    wire new_AGEMA_signal_12718 ;
    wire new_AGEMA_signal_12719 ;
    wire new_AGEMA_signal_12720 ;
    wire new_AGEMA_signal_12721 ;
    wire new_AGEMA_signal_12722 ;
    wire new_AGEMA_signal_12723 ;
    wire new_AGEMA_signal_12724 ;
    wire new_AGEMA_signal_12725 ;
    wire new_AGEMA_signal_12726 ;
    wire new_AGEMA_signal_12727 ;
    wire new_AGEMA_signal_12728 ;
    wire new_AGEMA_signal_12729 ;
    wire new_AGEMA_signal_12730 ;
    wire new_AGEMA_signal_12731 ;
    wire new_AGEMA_signal_12732 ;
    wire new_AGEMA_signal_12733 ;
    wire new_AGEMA_signal_12734 ;
    wire new_AGEMA_signal_12735 ;
    wire new_AGEMA_signal_12736 ;
    wire new_AGEMA_signal_12737 ;
    wire new_AGEMA_signal_12738 ;
    wire new_AGEMA_signal_12739 ;
    wire new_AGEMA_signal_12740 ;
    wire new_AGEMA_signal_12741 ;
    wire new_AGEMA_signal_12742 ;
    wire new_AGEMA_signal_12743 ;
    wire new_AGEMA_signal_12744 ;
    wire new_AGEMA_signal_12745 ;
    wire new_AGEMA_signal_12746 ;
    wire new_AGEMA_signal_12747 ;
    wire new_AGEMA_signal_12748 ;
    wire new_AGEMA_signal_12749 ;
    wire new_AGEMA_signal_12750 ;
    wire new_AGEMA_signal_12751 ;
    wire new_AGEMA_signal_12752 ;
    wire new_AGEMA_signal_12753 ;
    wire new_AGEMA_signal_12754 ;
    wire new_AGEMA_signal_12755 ;
    wire new_AGEMA_signal_12756 ;
    wire new_AGEMA_signal_12757 ;
    wire new_AGEMA_signal_12758 ;
    wire new_AGEMA_signal_12759 ;
    wire new_AGEMA_signal_12760 ;
    wire new_AGEMA_signal_12761 ;
    wire new_AGEMA_signal_12762 ;
    wire new_AGEMA_signal_12763 ;
    wire new_AGEMA_signal_12764 ;
    wire new_AGEMA_signal_12765 ;
    wire new_AGEMA_signal_12766 ;
    wire new_AGEMA_signal_12767 ;
    wire new_AGEMA_signal_12768 ;
    wire new_AGEMA_signal_12769 ;
    wire new_AGEMA_signal_12770 ;
    wire new_AGEMA_signal_12771 ;
    wire new_AGEMA_signal_12772 ;
    wire new_AGEMA_signal_12773 ;
    wire new_AGEMA_signal_12774 ;
    wire new_AGEMA_signal_12775 ;
    wire new_AGEMA_signal_12776 ;
    wire new_AGEMA_signal_12777 ;
    wire new_AGEMA_signal_12778 ;
    wire new_AGEMA_signal_12779 ;
    wire new_AGEMA_signal_12780 ;
    wire new_AGEMA_signal_12781 ;
    wire new_AGEMA_signal_12782 ;
    wire new_AGEMA_signal_12783 ;
    wire new_AGEMA_signal_12784 ;
    wire new_AGEMA_signal_12785 ;
    wire new_AGEMA_signal_12786 ;
    wire new_AGEMA_signal_12787 ;
    wire new_AGEMA_signal_12788 ;
    wire new_AGEMA_signal_12789 ;
    wire new_AGEMA_signal_12790 ;
    wire new_AGEMA_signal_12791 ;
    wire new_AGEMA_signal_12792 ;
    wire new_AGEMA_signal_12793 ;
    wire new_AGEMA_signal_12794 ;
    wire new_AGEMA_signal_12795 ;
    wire new_AGEMA_signal_12796 ;
    wire new_AGEMA_signal_12797 ;
    wire new_AGEMA_signal_12798 ;
    wire new_AGEMA_signal_12799 ;
    wire new_AGEMA_signal_12800 ;
    wire new_AGEMA_signal_12801 ;
    wire new_AGEMA_signal_12802 ;
    wire new_AGEMA_signal_12803 ;
    wire new_AGEMA_signal_12804 ;
    wire new_AGEMA_signal_12805 ;
    wire new_AGEMA_signal_12806 ;
    wire new_AGEMA_signal_12807 ;
    wire new_AGEMA_signal_12808 ;
    wire new_AGEMA_signal_12809 ;
    wire new_AGEMA_signal_12810 ;
    wire new_AGEMA_signal_12811 ;
    wire new_AGEMA_signal_12812 ;
    wire new_AGEMA_signal_12813 ;
    wire new_AGEMA_signal_12814 ;
    wire new_AGEMA_signal_12815 ;
    wire new_AGEMA_signal_12816 ;
    wire new_AGEMA_signal_12817 ;
    wire new_AGEMA_signal_12818 ;
    wire new_AGEMA_signal_12819 ;
    wire new_AGEMA_signal_12820 ;
    wire new_AGEMA_signal_12821 ;
    wire new_AGEMA_signal_12822 ;
    wire new_AGEMA_signal_12823 ;
    wire new_AGEMA_signal_12824 ;
    wire new_AGEMA_signal_12825 ;
    wire new_AGEMA_signal_12826 ;
    wire new_AGEMA_signal_12827 ;
    wire new_AGEMA_signal_12828 ;
    wire new_AGEMA_signal_12829 ;
    wire new_AGEMA_signal_12830 ;
    wire new_AGEMA_signal_12831 ;
    wire new_AGEMA_signal_12832 ;
    wire new_AGEMA_signal_12833 ;
    wire new_AGEMA_signal_12834 ;
    wire new_AGEMA_signal_12835 ;
    wire new_AGEMA_signal_12836 ;
    wire new_AGEMA_signal_12837 ;
    wire new_AGEMA_signal_12838 ;
    wire new_AGEMA_signal_12839 ;
    wire new_AGEMA_signal_12840 ;
    wire new_AGEMA_signal_12841 ;
    wire new_AGEMA_signal_12842 ;
    wire new_AGEMA_signal_12843 ;
    wire new_AGEMA_signal_12844 ;
    wire new_AGEMA_signal_12845 ;
    wire new_AGEMA_signal_12846 ;
    wire new_AGEMA_signal_12847 ;
    wire new_AGEMA_signal_12848 ;
    wire new_AGEMA_signal_12849 ;
    wire new_AGEMA_signal_12850 ;
    wire new_AGEMA_signal_12851 ;
    wire new_AGEMA_signal_12852 ;
    wire new_AGEMA_signal_12853 ;
    wire new_AGEMA_signal_12854 ;
    wire new_AGEMA_signal_12855 ;
    wire new_AGEMA_signal_12856 ;
    wire new_AGEMA_signal_12857 ;
    wire new_AGEMA_signal_12858 ;
    wire new_AGEMA_signal_12859 ;
    wire new_AGEMA_signal_12860 ;
    wire new_AGEMA_signal_12861 ;
    wire new_AGEMA_signal_12862 ;
    wire new_AGEMA_signal_12863 ;
    wire new_AGEMA_signal_12864 ;
    wire new_AGEMA_signal_12865 ;
    wire new_AGEMA_signal_12866 ;
    wire new_AGEMA_signal_12867 ;
    wire new_AGEMA_signal_12868 ;
    wire new_AGEMA_signal_12869 ;
    wire new_AGEMA_signal_12870 ;
    wire new_AGEMA_signal_12871 ;
    wire new_AGEMA_signal_12872 ;
    wire new_AGEMA_signal_12873 ;
    wire new_AGEMA_signal_12874 ;
    wire new_AGEMA_signal_12875 ;
    wire new_AGEMA_signal_12876 ;
    wire new_AGEMA_signal_12877 ;
    wire new_AGEMA_signal_12878 ;
    wire new_AGEMA_signal_12879 ;
    wire new_AGEMA_signal_12880 ;
    wire new_AGEMA_signal_12881 ;
    wire new_AGEMA_signal_12882 ;
    wire new_AGEMA_signal_12883 ;
    wire new_AGEMA_signal_12884 ;
    wire new_AGEMA_signal_12885 ;
    wire new_AGEMA_signal_12886 ;
    wire new_AGEMA_signal_12887 ;
    wire new_AGEMA_signal_12888 ;
    wire new_AGEMA_signal_12889 ;
    wire new_AGEMA_signal_12890 ;
    wire new_AGEMA_signal_12891 ;
    wire new_AGEMA_signal_12892 ;
    wire new_AGEMA_signal_12893 ;
    wire new_AGEMA_signal_12894 ;
    wire new_AGEMA_signal_12895 ;
    wire new_AGEMA_signal_12896 ;
    wire new_AGEMA_signal_12897 ;
    wire new_AGEMA_signal_12898 ;
    wire new_AGEMA_signal_12899 ;
    wire new_AGEMA_signal_12900 ;
    wire new_AGEMA_signal_12901 ;
    wire new_AGEMA_signal_12902 ;
    wire new_AGEMA_signal_12903 ;
    wire new_AGEMA_signal_12904 ;
    wire new_AGEMA_signal_12905 ;
    wire new_AGEMA_signal_12906 ;
    wire new_AGEMA_signal_12907 ;
    wire new_AGEMA_signal_12908 ;
    wire new_AGEMA_signal_12909 ;
    wire new_AGEMA_signal_12910 ;
    wire new_AGEMA_signal_12911 ;
    wire new_AGEMA_signal_12912 ;
    wire new_AGEMA_signal_12913 ;
    wire new_AGEMA_signal_12914 ;
    wire new_AGEMA_signal_12915 ;
    wire new_AGEMA_signal_12916 ;
    wire new_AGEMA_signal_12917 ;
    wire new_AGEMA_signal_12918 ;
    wire new_AGEMA_signal_12919 ;
    wire new_AGEMA_signal_12920 ;
    wire new_AGEMA_signal_12921 ;
    wire new_AGEMA_signal_12922 ;
    wire new_AGEMA_signal_12923 ;
    wire new_AGEMA_signal_12924 ;
    wire new_AGEMA_signal_12925 ;
    wire new_AGEMA_signal_12926 ;
    wire new_AGEMA_signal_12927 ;
    wire new_AGEMA_signal_12928 ;
    wire new_AGEMA_signal_12929 ;
    wire new_AGEMA_signal_12930 ;
    wire new_AGEMA_signal_12931 ;
    wire new_AGEMA_signal_12932 ;
    wire new_AGEMA_signal_12933 ;
    wire new_AGEMA_signal_12934 ;
    wire new_AGEMA_signal_12935 ;
    wire new_AGEMA_signal_12936 ;
    wire new_AGEMA_signal_12937 ;
    wire new_AGEMA_signal_12938 ;
    wire new_AGEMA_signal_12939 ;
    wire new_AGEMA_signal_12940 ;
    wire new_AGEMA_signal_12941 ;
    wire new_AGEMA_signal_12942 ;
    wire new_AGEMA_signal_12943 ;
    wire new_AGEMA_signal_12944 ;
    wire new_AGEMA_signal_12945 ;
    wire new_AGEMA_signal_12946 ;
    wire new_AGEMA_signal_12947 ;
    wire new_AGEMA_signal_12948 ;
    wire new_AGEMA_signal_12949 ;
    wire new_AGEMA_signal_12950 ;
    wire new_AGEMA_signal_12951 ;
    wire new_AGEMA_signal_12952 ;
    wire new_AGEMA_signal_12953 ;
    wire new_AGEMA_signal_12954 ;
    wire new_AGEMA_signal_12955 ;
    wire new_AGEMA_signal_12956 ;
    wire new_AGEMA_signal_12957 ;
    wire new_AGEMA_signal_12958 ;
    wire new_AGEMA_signal_12959 ;
    wire new_AGEMA_signal_12960 ;
    wire new_AGEMA_signal_12961 ;
    wire new_AGEMA_signal_12962 ;
    wire new_AGEMA_signal_12963 ;
    wire new_AGEMA_signal_12964 ;
    wire new_AGEMA_signal_12965 ;
    wire new_AGEMA_signal_12966 ;
    wire new_AGEMA_signal_12967 ;
    wire new_AGEMA_signal_12968 ;
    wire new_AGEMA_signal_12969 ;
    wire new_AGEMA_signal_12970 ;
    wire new_AGEMA_signal_12971 ;
    wire new_AGEMA_signal_12972 ;
    wire new_AGEMA_signal_12973 ;
    wire new_AGEMA_signal_12974 ;
    wire new_AGEMA_signal_12975 ;
    wire new_AGEMA_signal_12976 ;
    wire new_AGEMA_signal_12977 ;
    wire new_AGEMA_signal_12978 ;
    wire new_AGEMA_signal_12979 ;
    wire new_AGEMA_signal_12980 ;
    wire new_AGEMA_signal_12981 ;
    wire new_AGEMA_signal_12982 ;
    wire new_AGEMA_signal_12983 ;
    wire new_AGEMA_signal_12984 ;
    wire new_AGEMA_signal_12985 ;
    wire new_AGEMA_signal_12986 ;
    wire new_AGEMA_signal_12987 ;
    wire new_AGEMA_signal_12988 ;
    wire new_AGEMA_signal_12989 ;
    wire new_AGEMA_signal_12990 ;
    wire new_AGEMA_signal_12991 ;
    wire new_AGEMA_signal_12992 ;
    wire new_AGEMA_signal_12993 ;
    wire new_AGEMA_signal_12994 ;
    wire new_AGEMA_signal_12995 ;
    wire new_AGEMA_signal_12996 ;
    wire new_AGEMA_signal_12997 ;
    wire new_AGEMA_signal_12998 ;
    wire new_AGEMA_signal_12999 ;
    wire new_AGEMA_signal_13000 ;
    wire new_AGEMA_signal_13001 ;
    wire new_AGEMA_signal_13002 ;
    wire new_AGEMA_signal_13003 ;
    wire new_AGEMA_signal_13004 ;
    wire new_AGEMA_signal_13005 ;
    wire new_AGEMA_signal_13006 ;
    wire new_AGEMA_signal_13007 ;
    wire new_AGEMA_signal_13008 ;
    wire new_AGEMA_signal_13009 ;
    wire new_AGEMA_signal_13010 ;
    wire new_AGEMA_signal_13011 ;
    wire new_AGEMA_signal_13012 ;
    wire new_AGEMA_signal_13013 ;
    wire new_AGEMA_signal_13014 ;
    wire new_AGEMA_signal_13015 ;
    wire new_AGEMA_signal_13016 ;
    wire new_AGEMA_signal_13017 ;
    wire new_AGEMA_signal_13018 ;
    wire new_AGEMA_signal_13019 ;
    wire new_AGEMA_signal_13020 ;
    wire new_AGEMA_signal_13021 ;
    wire new_AGEMA_signal_13022 ;
    wire new_AGEMA_signal_13023 ;
    wire new_AGEMA_signal_13024 ;
    wire new_AGEMA_signal_13025 ;
    wire new_AGEMA_signal_13026 ;
    wire new_AGEMA_signal_13027 ;
    wire new_AGEMA_signal_13028 ;
    wire new_AGEMA_signal_13029 ;
    wire new_AGEMA_signal_13030 ;
    wire new_AGEMA_signal_13031 ;
    wire new_AGEMA_signal_13032 ;
    wire new_AGEMA_signal_13033 ;
    wire new_AGEMA_signal_13034 ;
    wire new_AGEMA_signal_13035 ;
    wire new_AGEMA_signal_13036 ;
    wire new_AGEMA_signal_13037 ;
    wire new_AGEMA_signal_13038 ;
    wire new_AGEMA_signal_13039 ;
    wire new_AGEMA_signal_13040 ;
    wire new_AGEMA_signal_13041 ;
    wire new_AGEMA_signal_13042 ;
    wire new_AGEMA_signal_13043 ;
    wire new_AGEMA_signal_13044 ;
    wire new_AGEMA_signal_13045 ;
    wire new_AGEMA_signal_13046 ;
    wire new_AGEMA_signal_13047 ;
    wire new_AGEMA_signal_13048 ;
    wire new_AGEMA_signal_13049 ;
    wire new_AGEMA_signal_13050 ;
    wire new_AGEMA_signal_13051 ;
    wire new_AGEMA_signal_13052 ;
    wire new_AGEMA_signal_13053 ;
    wire new_AGEMA_signal_13054 ;
    wire new_AGEMA_signal_13055 ;
    wire new_AGEMA_signal_13056 ;
    wire new_AGEMA_signal_13057 ;
    wire new_AGEMA_signal_13058 ;
    wire new_AGEMA_signal_13059 ;
    wire new_AGEMA_signal_13060 ;
    wire new_AGEMA_signal_13061 ;
    wire new_AGEMA_signal_13062 ;
    wire new_AGEMA_signal_13063 ;
    wire new_AGEMA_signal_13064 ;
    wire new_AGEMA_signal_13065 ;
    wire new_AGEMA_signal_13066 ;
    wire new_AGEMA_signal_13067 ;
    wire new_AGEMA_signal_13068 ;
    wire new_AGEMA_signal_13069 ;
    wire new_AGEMA_signal_13070 ;
    wire new_AGEMA_signal_13071 ;
    wire new_AGEMA_signal_13072 ;
    wire new_AGEMA_signal_13073 ;
    wire new_AGEMA_signal_13074 ;
    wire new_AGEMA_signal_13075 ;
    wire new_AGEMA_signal_13076 ;
    wire new_AGEMA_signal_13077 ;
    wire new_AGEMA_signal_13078 ;
    wire new_AGEMA_signal_13079 ;
    wire new_AGEMA_signal_13080 ;
    wire new_AGEMA_signal_13081 ;
    wire new_AGEMA_signal_13082 ;
    wire new_AGEMA_signal_13083 ;
    wire new_AGEMA_signal_13084 ;
    wire new_AGEMA_signal_13085 ;
    wire new_AGEMA_signal_13086 ;
    wire new_AGEMA_signal_13087 ;
    wire new_AGEMA_signal_13088 ;
    wire new_AGEMA_signal_13089 ;
    wire new_AGEMA_signal_13090 ;
    wire new_AGEMA_signal_13091 ;
    wire new_AGEMA_signal_13092 ;
    wire new_AGEMA_signal_13093 ;
    wire new_AGEMA_signal_13094 ;
    wire new_AGEMA_signal_13095 ;
    wire new_AGEMA_signal_13096 ;
    wire new_AGEMA_signal_13097 ;
    wire new_AGEMA_signal_13098 ;
    wire new_AGEMA_signal_13099 ;
    wire new_AGEMA_signal_13100 ;
    wire new_AGEMA_signal_13101 ;
    wire new_AGEMA_signal_13102 ;
    wire new_AGEMA_signal_13103 ;
    wire new_AGEMA_signal_13104 ;
    wire new_AGEMA_signal_13105 ;
    wire new_AGEMA_signal_13106 ;
    wire new_AGEMA_signal_13107 ;
    wire new_AGEMA_signal_13108 ;
    wire new_AGEMA_signal_13109 ;
    wire new_AGEMA_signal_13110 ;
    wire new_AGEMA_signal_13111 ;
    wire new_AGEMA_signal_13112 ;
    wire new_AGEMA_signal_13113 ;
    wire new_AGEMA_signal_13114 ;
    wire new_AGEMA_signal_13115 ;
    wire new_AGEMA_signal_13116 ;
    wire new_AGEMA_signal_13117 ;
    wire new_AGEMA_signal_13118 ;
    wire new_AGEMA_signal_13119 ;
    wire new_AGEMA_signal_13120 ;
    wire new_AGEMA_signal_13121 ;
    wire new_AGEMA_signal_13122 ;
    wire new_AGEMA_signal_13123 ;
    wire new_AGEMA_signal_13124 ;
    wire new_AGEMA_signal_13125 ;
    wire new_AGEMA_signal_13126 ;
    wire new_AGEMA_signal_13127 ;
    wire new_AGEMA_signal_13128 ;
    wire new_AGEMA_signal_13129 ;
    wire new_AGEMA_signal_13130 ;
    wire new_AGEMA_signal_13131 ;
    wire new_AGEMA_signal_13132 ;
    wire new_AGEMA_signal_13133 ;
    wire new_AGEMA_signal_13134 ;
    wire new_AGEMA_signal_13135 ;
    wire new_AGEMA_signal_13136 ;
    wire new_AGEMA_signal_13137 ;
    wire new_AGEMA_signal_13138 ;
    wire new_AGEMA_signal_13139 ;
    wire new_AGEMA_signal_13140 ;
    wire new_AGEMA_signal_13141 ;
    wire new_AGEMA_signal_13142 ;
    wire new_AGEMA_signal_13143 ;
    wire new_AGEMA_signal_13144 ;
    wire new_AGEMA_signal_13145 ;
    wire new_AGEMA_signal_13146 ;
    wire new_AGEMA_signal_13147 ;
    wire new_AGEMA_signal_13148 ;
    wire new_AGEMA_signal_13149 ;
    wire new_AGEMA_signal_13150 ;
    wire new_AGEMA_signal_13151 ;
    wire new_AGEMA_signal_13152 ;
    wire new_AGEMA_signal_13153 ;
    wire new_AGEMA_signal_13154 ;
    wire new_AGEMA_signal_13155 ;
    wire new_AGEMA_signal_13156 ;
    wire new_AGEMA_signal_13157 ;
    wire new_AGEMA_signal_13158 ;
    wire new_AGEMA_signal_13159 ;
    wire new_AGEMA_signal_13160 ;
    wire new_AGEMA_signal_13161 ;
    wire new_AGEMA_signal_13162 ;
    wire new_AGEMA_signal_13163 ;
    wire new_AGEMA_signal_13164 ;
    wire new_AGEMA_signal_13165 ;
    wire new_AGEMA_signal_13166 ;
    wire new_AGEMA_signal_13167 ;
    wire new_AGEMA_signal_13168 ;
    wire new_AGEMA_signal_13169 ;
    wire new_AGEMA_signal_13170 ;
    wire new_AGEMA_signal_13171 ;
    wire new_AGEMA_signal_13172 ;
    wire new_AGEMA_signal_13173 ;
    wire new_AGEMA_signal_13174 ;
    wire new_AGEMA_signal_13175 ;
    wire new_AGEMA_signal_13176 ;
    wire new_AGEMA_signal_13177 ;
    wire new_AGEMA_signal_13178 ;
    wire new_AGEMA_signal_13179 ;
    wire new_AGEMA_signal_13180 ;
    wire new_AGEMA_signal_13181 ;
    wire new_AGEMA_signal_13182 ;
    wire new_AGEMA_signal_13183 ;
    wire new_AGEMA_signal_13184 ;
    wire new_AGEMA_signal_13185 ;
    wire new_AGEMA_signal_13186 ;
    wire new_AGEMA_signal_13187 ;
    wire new_AGEMA_signal_13188 ;
    wire new_AGEMA_signal_13189 ;
    wire new_AGEMA_signal_13190 ;
    wire new_AGEMA_signal_13191 ;
    wire new_AGEMA_signal_13192 ;
    wire new_AGEMA_signal_13193 ;
    wire new_AGEMA_signal_13194 ;
    wire new_AGEMA_signal_13195 ;
    wire new_AGEMA_signal_13196 ;
    wire new_AGEMA_signal_13197 ;
    wire new_AGEMA_signal_13198 ;
    wire new_AGEMA_signal_13199 ;
    wire new_AGEMA_signal_13200 ;
    wire new_AGEMA_signal_13201 ;
    wire new_AGEMA_signal_13202 ;
    wire new_AGEMA_signal_13203 ;
    wire new_AGEMA_signal_13204 ;
    wire new_AGEMA_signal_13205 ;
    wire new_AGEMA_signal_13206 ;
    wire new_AGEMA_signal_13207 ;
    wire new_AGEMA_signal_13208 ;
    wire new_AGEMA_signal_13209 ;
    wire new_AGEMA_signal_13210 ;
    wire new_AGEMA_signal_13211 ;
    wire new_AGEMA_signal_13212 ;
    wire new_AGEMA_signal_13213 ;
    wire new_AGEMA_signal_13214 ;
    wire new_AGEMA_signal_13215 ;
    wire new_AGEMA_signal_13216 ;
    wire new_AGEMA_signal_13217 ;
    wire new_AGEMA_signal_13218 ;
    wire new_AGEMA_signal_13219 ;
    wire new_AGEMA_signal_13220 ;
    wire new_AGEMA_signal_13221 ;
    wire new_AGEMA_signal_13222 ;
    wire new_AGEMA_signal_13223 ;
    wire new_AGEMA_signal_13224 ;
    wire new_AGEMA_signal_13225 ;
    wire new_AGEMA_signal_13226 ;
    wire new_AGEMA_signal_13227 ;
    wire new_AGEMA_signal_13228 ;
    wire new_AGEMA_signal_13229 ;
    wire new_AGEMA_signal_13230 ;
    wire new_AGEMA_signal_13231 ;
    wire new_AGEMA_signal_13232 ;
    wire new_AGEMA_signal_13233 ;
    wire new_AGEMA_signal_13234 ;
    wire new_AGEMA_signal_13235 ;
    wire new_AGEMA_signal_13236 ;
    wire new_AGEMA_signal_13237 ;
    wire new_AGEMA_signal_13238 ;
    wire new_AGEMA_signal_13239 ;
    wire new_AGEMA_signal_13240 ;
    wire new_AGEMA_signal_13241 ;
    wire new_AGEMA_signal_13242 ;
    wire new_AGEMA_signal_13243 ;
    wire new_AGEMA_signal_13244 ;
    wire new_AGEMA_signal_13245 ;
    wire new_AGEMA_signal_13246 ;
    wire new_AGEMA_signal_13247 ;
    wire new_AGEMA_signal_13248 ;
    wire new_AGEMA_signal_13249 ;
    wire new_AGEMA_signal_13250 ;
    wire new_AGEMA_signal_13251 ;
    wire new_AGEMA_signal_13252 ;
    wire new_AGEMA_signal_13253 ;
    wire new_AGEMA_signal_13254 ;
    wire new_AGEMA_signal_13255 ;
    wire new_AGEMA_signal_13256 ;
    wire new_AGEMA_signal_13257 ;
    wire new_AGEMA_signal_13258 ;
    wire new_AGEMA_signal_13259 ;
    wire new_AGEMA_signal_13260 ;
    wire new_AGEMA_signal_13261 ;
    wire new_AGEMA_signal_13262 ;
    wire new_AGEMA_signal_13263 ;
    wire new_AGEMA_signal_13264 ;
    wire new_AGEMA_signal_13265 ;
    wire new_AGEMA_signal_13266 ;
    wire new_AGEMA_signal_13267 ;
    wire new_AGEMA_signal_13268 ;
    wire new_AGEMA_signal_13269 ;
    wire new_AGEMA_signal_13270 ;
    wire new_AGEMA_signal_13271 ;
    wire new_AGEMA_signal_13272 ;
    wire new_AGEMA_signal_13273 ;
    wire new_AGEMA_signal_13274 ;
    wire new_AGEMA_signal_13275 ;
    wire new_AGEMA_signal_13276 ;
    wire new_AGEMA_signal_13277 ;
    wire new_AGEMA_signal_13278 ;
    wire new_AGEMA_signal_13279 ;
    wire new_AGEMA_signal_13280 ;
    wire new_AGEMA_signal_13281 ;
    wire new_AGEMA_signal_13282 ;
    wire new_AGEMA_signal_13283 ;
    wire new_AGEMA_signal_13284 ;
    wire new_AGEMA_signal_13285 ;
    wire new_AGEMA_signal_13286 ;
    wire new_AGEMA_signal_13287 ;
    wire new_AGEMA_signal_13288 ;
    wire new_AGEMA_signal_13289 ;
    wire new_AGEMA_signal_13290 ;
    wire new_AGEMA_signal_13291 ;
    wire new_AGEMA_signal_13292 ;
    wire new_AGEMA_signal_13293 ;
    wire new_AGEMA_signal_13294 ;
    wire new_AGEMA_signal_13295 ;
    wire new_AGEMA_signal_13296 ;
    wire new_AGEMA_signal_13297 ;
    wire new_AGEMA_signal_13298 ;
    wire new_AGEMA_signal_13299 ;
    wire new_AGEMA_signal_13300 ;
    wire new_AGEMA_signal_13301 ;
    wire new_AGEMA_signal_13302 ;
    wire new_AGEMA_signal_13303 ;
    wire new_AGEMA_signal_13304 ;
    wire new_AGEMA_signal_13305 ;
    wire new_AGEMA_signal_13306 ;
    wire new_AGEMA_signal_13307 ;
    wire new_AGEMA_signal_13308 ;
    wire new_AGEMA_signal_13309 ;
    wire new_AGEMA_signal_13310 ;
    wire new_AGEMA_signal_13311 ;
    wire new_AGEMA_signal_13312 ;
    wire new_AGEMA_signal_13313 ;
    wire new_AGEMA_signal_13314 ;
    wire new_AGEMA_signal_13315 ;
    wire new_AGEMA_signal_13316 ;
    wire new_AGEMA_signal_13317 ;
    wire new_AGEMA_signal_13318 ;
    wire new_AGEMA_signal_13319 ;
    wire new_AGEMA_signal_13320 ;
    wire new_AGEMA_signal_13321 ;
    wire new_AGEMA_signal_13322 ;
    wire new_AGEMA_signal_13323 ;
    wire new_AGEMA_signal_13324 ;
    wire new_AGEMA_signal_13325 ;
    wire new_AGEMA_signal_13326 ;
    wire new_AGEMA_signal_13327 ;
    wire new_AGEMA_signal_13328 ;
    wire new_AGEMA_signal_13329 ;
    wire new_AGEMA_signal_13330 ;
    wire new_AGEMA_signal_13331 ;
    wire new_AGEMA_signal_13332 ;
    wire new_AGEMA_signal_13333 ;
    wire new_AGEMA_signal_13334 ;
    wire new_AGEMA_signal_13335 ;
    wire new_AGEMA_signal_13336 ;
    wire new_AGEMA_signal_13337 ;
    wire new_AGEMA_signal_13338 ;
    wire new_AGEMA_signal_13339 ;
    wire new_AGEMA_signal_13340 ;
    wire new_AGEMA_signal_13341 ;
    wire new_AGEMA_signal_13342 ;
    wire new_AGEMA_signal_13343 ;
    wire new_AGEMA_signal_13344 ;
    wire new_AGEMA_signal_13345 ;
    wire new_AGEMA_signal_13346 ;
    wire new_AGEMA_signal_13347 ;
    wire new_AGEMA_signal_13348 ;
    wire new_AGEMA_signal_13349 ;
    wire new_AGEMA_signal_13350 ;
    wire new_AGEMA_signal_13351 ;
    wire new_AGEMA_signal_13352 ;
    wire new_AGEMA_signal_13353 ;
    wire new_AGEMA_signal_13354 ;
    wire new_AGEMA_signal_13355 ;
    wire new_AGEMA_signal_13356 ;
    wire new_AGEMA_signal_13357 ;
    wire new_AGEMA_signal_13358 ;
    wire new_AGEMA_signal_13359 ;
    wire new_AGEMA_signal_13360 ;
    wire new_AGEMA_signal_13361 ;
    wire new_AGEMA_signal_13362 ;
    wire new_AGEMA_signal_13363 ;
    wire new_AGEMA_signal_13364 ;
    wire new_AGEMA_signal_13365 ;
    wire new_AGEMA_signal_13366 ;
    wire new_AGEMA_signal_13367 ;
    wire new_AGEMA_signal_13368 ;
    wire new_AGEMA_signal_13369 ;
    wire new_AGEMA_signal_13370 ;
    wire new_AGEMA_signal_13371 ;
    wire new_AGEMA_signal_13372 ;
    wire new_AGEMA_signal_13373 ;
    wire new_AGEMA_signal_13374 ;
    wire new_AGEMA_signal_13375 ;
    wire new_AGEMA_signal_13376 ;
    wire new_AGEMA_signal_13377 ;
    wire new_AGEMA_signal_13378 ;
    wire new_AGEMA_signal_13379 ;
    wire new_AGEMA_signal_13380 ;
    wire new_AGEMA_signal_13381 ;
    wire new_AGEMA_signal_13382 ;
    wire new_AGEMA_signal_13383 ;
    wire new_AGEMA_signal_13384 ;
    wire new_AGEMA_signal_13385 ;
    wire new_AGEMA_signal_13386 ;
    wire new_AGEMA_signal_13387 ;
    wire new_AGEMA_signal_13388 ;
    wire new_AGEMA_signal_13389 ;
    wire new_AGEMA_signal_13390 ;
    wire new_AGEMA_signal_13391 ;
    wire new_AGEMA_signal_13392 ;
    wire new_AGEMA_signal_13393 ;
    wire new_AGEMA_signal_13394 ;
    wire new_AGEMA_signal_13395 ;
    wire new_AGEMA_signal_13396 ;
    wire new_AGEMA_signal_13397 ;
    wire new_AGEMA_signal_13398 ;
    wire new_AGEMA_signal_13399 ;
    wire new_AGEMA_signal_13400 ;
    wire new_AGEMA_signal_13401 ;
    wire new_AGEMA_signal_13402 ;
    wire new_AGEMA_signal_13403 ;
    wire new_AGEMA_signal_13404 ;
    wire new_AGEMA_signal_13405 ;
    wire new_AGEMA_signal_13406 ;
    wire new_AGEMA_signal_13407 ;
    wire new_AGEMA_signal_13408 ;
    wire new_AGEMA_signal_13409 ;
    wire new_AGEMA_signal_13410 ;
    wire new_AGEMA_signal_13411 ;
    wire new_AGEMA_signal_13412 ;
    wire new_AGEMA_signal_13413 ;
    wire new_AGEMA_signal_13414 ;
    wire new_AGEMA_signal_13415 ;
    wire new_AGEMA_signal_13416 ;
    wire new_AGEMA_signal_13417 ;
    wire new_AGEMA_signal_13418 ;
    wire new_AGEMA_signal_13419 ;
    wire new_AGEMA_signal_13420 ;
    wire new_AGEMA_signal_13421 ;
    wire new_AGEMA_signal_13422 ;
    wire new_AGEMA_signal_13423 ;
    wire new_AGEMA_signal_13424 ;
    wire new_AGEMA_signal_13425 ;
    wire new_AGEMA_signal_13426 ;
    wire new_AGEMA_signal_13427 ;
    wire new_AGEMA_signal_13428 ;
    wire new_AGEMA_signal_13429 ;
    wire new_AGEMA_signal_13430 ;
    wire new_AGEMA_signal_13431 ;
    wire new_AGEMA_signal_13432 ;
    wire new_AGEMA_signal_13433 ;
    wire new_AGEMA_signal_13434 ;
    wire new_AGEMA_signal_13435 ;
    wire new_AGEMA_signal_13436 ;
    wire new_AGEMA_signal_13437 ;
    wire new_AGEMA_signal_13438 ;
    wire new_AGEMA_signal_13439 ;
    wire new_AGEMA_signal_13440 ;
    wire new_AGEMA_signal_13441 ;
    wire new_AGEMA_signal_13442 ;
    wire new_AGEMA_signal_13443 ;
    wire new_AGEMA_signal_13444 ;
    wire new_AGEMA_signal_13445 ;
    wire new_AGEMA_signal_13446 ;
    wire new_AGEMA_signal_13447 ;
    wire new_AGEMA_signal_13448 ;
    wire new_AGEMA_signal_13449 ;
    wire new_AGEMA_signal_13450 ;
    wire new_AGEMA_signal_13451 ;
    wire new_AGEMA_signal_13452 ;
    wire new_AGEMA_signal_13453 ;
    wire new_AGEMA_signal_13454 ;
    wire new_AGEMA_signal_13455 ;
    wire new_AGEMA_signal_13456 ;
    wire new_AGEMA_signal_13457 ;
    wire new_AGEMA_signal_13458 ;
    wire new_AGEMA_signal_13459 ;
    wire new_AGEMA_signal_13460 ;
    wire new_AGEMA_signal_13461 ;
    wire new_AGEMA_signal_13462 ;
    wire new_AGEMA_signal_13463 ;
    wire new_AGEMA_signal_13464 ;
    wire new_AGEMA_signal_13465 ;
    wire new_AGEMA_signal_13466 ;
    wire new_AGEMA_signal_13467 ;
    wire new_AGEMA_signal_13468 ;
    wire new_AGEMA_signal_13469 ;
    wire new_AGEMA_signal_13470 ;
    wire new_AGEMA_signal_13471 ;
    wire new_AGEMA_signal_13472 ;
    wire new_AGEMA_signal_13473 ;
    wire new_AGEMA_signal_13474 ;
    wire new_AGEMA_signal_13475 ;
    wire new_AGEMA_signal_13476 ;
    wire new_AGEMA_signal_13477 ;
    wire new_AGEMA_signal_13478 ;
    wire new_AGEMA_signal_13479 ;
    wire new_AGEMA_signal_13480 ;
    wire new_AGEMA_signal_13481 ;
    wire new_AGEMA_signal_13482 ;
    wire new_AGEMA_signal_13483 ;
    wire new_AGEMA_signal_13484 ;
    wire new_AGEMA_signal_13485 ;
    wire new_AGEMA_signal_13486 ;
    wire new_AGEMA_signal_13487 ;
    wire new_AGEMA_signal_13488 ;
    wire new_AGEMA_signal_13489 ;
    wire new_AGEMA_signal_13490 ;
    wire new_AGEMA_signal_13491 ;
    wire new_AGEMA_signal_13492 ;
    wire new_AGEMA_signal_13493 ;
    wire new_AGEMA_signal_13494 ;
    wire new_AGEMA_signal_13495 ;
    wire new_AGEMA_signal_13496 ;
    wire new_AGEMA_signal_13497 ;
    wire new_AGEMA_signal_13498 ;
    wire new_AGEMA_signal_13499 ;
    wire new_AGEMA_signal_13500 ;
    wire new_AGEMA_signal_13501 ;
    wire new_AGEMA_signal_13502 ;
    wire new_AGEMA_signal_13503 ;
    wire new_AGEMA_signal_13504 ;
    wire new_AGEMA_signal_13505 ;
    wire new_AGEMA_signal_13506 ;
    wire new_AGEMA_signal_13507 ;
    wire new_AGEMA_signal_13508 ;
    wire new_AGEMA_signal_13509 ;
    wire new_AGEMA_signal_13510 ;
    wire new_AGEMA_signal_13511 ;
    wire new_AGEMA_signal_13512 ;
    wire new_AGEMA_signal_13513 ;
    wire new_AGEMA_signal_13514 ;
    wire new_AGEMA_signal_13515 ;
    wire new_AGEMA_signal_13516 ;
    wire new_AGEMA_signal_13517 ;
    wire new_AGEMA_signal_13518 ;
    wire new_AGEMA_signal_13519 ;
    wire new_AGEMA_signal_13520 ;
    wire new_AGEMA_signal_13521 ;
    wire new_AGEMA_signal_13522 ;
    wire new_AGEMA_signal_13523 ;
    wire new_AGEMA_signal_13524 ;
    wire new_AGEMA_signal_13525 ;
    wire new_AGEMA_signal_13526 ;
    wire new_AGEMA_signal_13527 ;
    wire new_AGEMA_signal_13528 ;
    wire new_AGEMA_signal_13529 ;
    wire new_AGEMA_signal_13530 ;
    wire new_AGEMA_signal_13531 ;
    wire new_AGEMA_signal_13532 ;
    wire new_AGEMA_signal_13533 ;
    wire new_AGEMA_signal_13534 ;
    wire new_AGEMA_signal_13535 ;
    wire new_AGEMA_signal_13536 ;
    wire new_AGEMA_signal_13537 ;
    wire new_AGEMA_signal_13538 ;
    wire new_AGEMA_signal_13539 ;
    wire new_AGEMA_signal_13540 ;
    wire new_AGEMA_signal_13541 ;
    wire new_AGEMA_signal_13542 ;
    wire new_AGEMA_signal_13543 ;
    wire new_AGEMA_signal_13544 ;
    wire new_AGEMA_signal_13545 ;
    wire new_AGEMA_signal_13546 ;
    wire new_AGEMA_signal_13547 ;
    wire new_AGEMA_signal_13548 ;
    wire new_AGEMA_signal_13549 ;
    wire new_AGEMA_signal_13550 ;
    wire new_AGEMA_signal_13551 ;
    wire new_AGEMA_signal_13552 ;
    wire new_AGEMA_signal_13553 ;
    wire new_AGEMA_signal_13554 ;
    wire new_AGEMA_signal_13555 ;
    wire new_AGEMA_signal_13556 ;
    wire new_AGEMA_signal_13557 ;
    wire new_AGEMA_signal_13558 ;
    wire new_AGEMA_signal_13559 ;
    wire new_AGEMA_signal_13560 ;
    wire new_AGEMA_signal_13561 ;
    wire new_AGEMA_signal_13562 ;
    wire new_AGEMA_signal_13563 ;
    wire new_AGEMA_signal_13564 ;
    wire new_AGEMA_signal_13565 ;
    wire new_AGEMA_signal_13566 ;
    wire new_AGEMA_signal_13567 ;
    wire new_AGEMA_signal_13568 ;
    wire new_AGEMA_signal_13569 ;
    wire new_AGEMA_signal_13570 ;
    wire new_AGEMA_signal_13571 ;
    wire new_AGEMA_signal_13572 ;
    wire new_AGEMA_signal_13573 ;
    wire new_AGEMA_signal_13574 ;
    wire new_AGEMA_signal_13575 ;
    wire new_AGEMA_signal_13576 ;
    wire new_AGEMA_signal_13577 ;
    wire new_AGEMA_signal_13578 ;
    wire new_AGEMA_signal_13579 ;
    wire new_AGEMA_signal_13580 ;
    wire new_AGEMA_signal_13581 ;
    wire new_AGEMA_signal_13582 ;
    wire new_AGEMA_signal_13583 ;
    wire new_AGEMA_signal_13584 ;
    wire new_AGEMA_signal_13585 ;
    wire new_AGEMA_signal_13586 ;
    wire new_AGEMA_signal_13587 ;
    wire new_AGEMA_signal_13588 ;
    wire new_AGEMA_signal_13589 ;
    wire new_AGEMA_signal_13590 ;
    wire new_AGEMA_signal_13591 ;
    wire new_AGEMA_signal_13592 ;
    wire new_AGEMA_signal_13593 ;
    wire new_AGEMA_signal_13594 ;
    wire new_AGEMA_signal_13595 ;
    wire new_AGEMA_signal_13596 ;
    wire new_AGEMA_signal_13597 ;
    wire new_AGEMA_signal_13598 ;
    wire new_AGEMA_signal_13599 ;
    wire new_AGEMA_signal_13600 ;
    wire new_AGEMA_signal_13601 ;
    wire new_AGEMA_signal_13602 ;
    wire new_AGEMA_signal_13603 ;
    wire new_AGEMA_signal_13604 ;
    wire new_AGEMA_signal_13605 ;
    wire new_AGEMA_signal_13606 ;
    wire new_AGEMA_signal_13607 ;
    wire new_AGEMA_signal_13608 ;
    wire new_AGEMA_signal_13609 ;
    wire new_AGEMA_signal_13610 ;
    wire new_AGEMA_signal_13611 ;
    wire new_AGEMA_signal_13612 ;
    wire new_AGEMA_signal_13613 ;
    wire new_AGEMA_signal_13614 ;
    wire new_AGEMA_signal_13615 ;
    wire new_AGEMA_signal_13616 ;
    wire new_AGEMA_signal_13617 ;
    wire new_AGEMA_signal_13618 ;
    wire new_AGEMA_signal_13619 ;
    wire new_AGEMA_signal_13620 ;
    wire new_AGEMA_signal_13621 ;
    wire new_AGEMA_signal_13622 ;
    wire new_AGEMA_signal_13623 ;
    wire new_AGEMA_signal_13624 ;
    wire new_AGEMA_signal_13625 ;
    wire new_AGEMA_signal_13626 ;
    wire new_AGEMA_signal_13627 ;
    wire new_AGEMA_signal_13628 ;
    wire new_AGEMA_signal_13629 ;
    wire new_AGEMA_signal_13630 ;
    wire new_AGEMA_signal_13631 ;
    wire new_AGEMA_signal_13632 ;
    wire new_AGEMA_signal_13633 ;
    wire new_AGEMA_signal_13634 ;
    wire new_AGEMA_signal_13635 ;
    wire new_AGEMA_signal_13636 ;
    wire new_AGEMA_signal_13637 ;
    wire new_AGEMA_signal_13638 ;
    wire new_AGEMA_signal_13639 ;
    wire new_AGEMA_signal_13640 ;
    wire new_AGEMA_signal_13641 ;
    wire new_AGEMA_signal_13642 ;
    wire new_AGEMA_signal_13643 ;
    wire new_AGEMA_signal_13644 ;
    wire new_AGEMA_signal_13645 ;
    wire new_AGEMA_signal_13646 ;
    wire new_AGEMA_signal_13647 ;
    wire new_AGEMA_signal_13648 ;
    wire new_AGEMA_signal_13649 ;
    wire new_AGEMA_signal_13650 ;
    wire new_AGEMA_signal_13651 ;
    wire new_AGEMA_signal_13652 ;
    wire new_AGEMA_signal_13653 ;
    wire new_AGEMA_signal_13654 ;
    wire new_AGEMA_signal_13655 ;
    wire new_AGEMA_signal_13656 ;
    wire new_AGEMA_signal_13657 ;
    wire new_AGEMA_signal_13658 ;
    wire new_AGEMA_signal_13659 ;
    wire new_AGEMA_signal_13660 ;
    wire new_AGEMA_signal_13661 ;
    wire new_AGEMA_signal_13662 ;
    wire new_AGEMA_signal_13663 ;
    wire new_AGEMA_signal_13664 ;
    wire new_AGEMA_signal_13665 ;
    wire new_AGEMA_signal_13666 ;
    wire new_AGEMA_signal_13667 ;
    wire new_AGEMA_signal_13668 ;
    wire new_AGEMA_signal_13669 ;
    wire new_AGEMA_signal_13670 ;
    wire new_AGEMA_signal_13671 ;
    wire new_AGEMA_signal_13672 ;
    wire new_AGEMA_signal_13673 ;
    wire new_AGEMA_signal_13674 ;
    wire new_AGEMA_signal_13675 ;
    wire new_AGEMA_signal_13676 ;
    wire new_AGEMA_signal_13677 ;
    wire new_AGEMA_signal_13678 ;
    wire new_AGEMA_signal_13679 ;
    wire new_AGEMA_signal_13680 ;
    wire new_AGEMA_signal_13681 ;
    wire new_AGEMA_signal_13682 ;
    wire new_AGEMA_signal_13683 ;
    wire new_AGEMA_signal_13684 ;
    wire new_AGEMA_signal_13685 ;
    wire new_AGEMA_signal_13686 ;
    wire new_AGEMA_signal_13687 ;
    wire new_AGEMA_signal_13688 ;
    wire new_AGEMA_signal_13689 ;
    wire new_AGEMA_signal_13690 ;
    wire new_AGEMA_signal_13691 ;
    wire new_AGEMA_signal_13692 ;
    wire new_AGEMA_signal_13693 ;
    wire new_AGEMA_signal_13694 ;
    wire new_AGEMA_signal_13695 ;
    wire new_AGEMA_signal_13696 ;
    wire new_AGEMA_signal_13697 ;
    wire new_AGEMA_signal_13698 ;
    wire new_AGEMA_signal_13699 ;
    wire new_AGEMA_signal_13700 ;
    wire new_AGEMA_signal_13701 ;
    wire new_AGEMA_signal_13702 ;
    wire new_AGEMA_signal_13703 ;
    wire new_AGEMA_signal_13704 ;
    wire new_AGEMA_signal_13705 ;
    wire new_AGEMA_signal_13706 ;
    wire new_AGEMA_signal_13707 ;
    wire new_AGEMA_signal_13708 ;
    wire new_AGEMA_signal_13709 ;
    wire new_AGEMA_signal_13710 ;
    wire new_AGEMA_signal_13711 ;
    wire new_AGEMA_signal_13712 ;
    wire new_AGEMA_signal_13713 ;
    wire new_AGEMA_signal_13714 ;
    wire new_AGEMA_signal_13715 ;
    wire new_AGEMA_signal_13716 ;
    wire new_AGEMA_signal_13717 ;
    wire new_AGEMA_signal_13718 ;
    wire new_AGEMA_signal_13719 ;
    wire new_AGEMA_signal_13720 ;
    wire new_AGEMA_signal_13721 ;
    wire new_AGEMA_signal_13722 ;
    wire new_AGEMA_signal_13723 ;
    wire new_AGEMA_signal_13724 ;
    wire new_AGEMA_signal_13725 ;
    wire new_AGEMA_signal_13726 ;
    wire new_AGEMA_signal_13727 ;
    wire new_AGEMA_signal_13728 ;
    wire new_AGEMA_signal_13729 ;
    wire new_AGEMA_signal_13730 ;
    wire new_AGEMA_signal_13731 ;
    wire new_AGEMA_signal_13732 ;
    wire new_AGEMA_signal_13733 ;
    wire new_AGEMA_signal_13734 ;
    wire new_AGEMA_signal_13735 ;
    wire new_AGEMA_signal_13736 ;
    wire new_AGEMA_signal_13737 ;
    wire new_AGEMA_signal_13738 ;
    wire new_AGEMA_signal_13739 ;
    wire new_AGEMA_signal_13740 ;
    wire new_AGEMA_signal_13741 ;
    wire new_AGEMA_signal_13742 ;
    wire new_AGEMA_signal_13743 ;
    wire new_AGEMA_signal_13744 ;
    wire new_AGEMA_signal_13745 ;
    wire new_AGEMA_signal_13746 ;
    wire new_AGEMA_signal_13747 ;
    wire new_AGEMA_signal_13748 ;
    wire new_AGEMA_signal_13749 ;
    wire new_AGEMA_signal_13750 ;
    wire new_AGEMA_signal_13751 ;
    wire new_AGEMA_signal_13752 ;
    wire new_AGEMA_signal_13753 ;
    wire new_AGEMA_signal_13754 ;
    wire new_AGEMA_signal_13755 ;
    wire new_AGEMA_signal_13756 ;
    wire new_AGEMA_signal_13757 ;
    wire new_AGEMA_signal_13758 ;
    wire new_AGEMA_signal_13759 ;
    wire new_AGEMA_signal_13760 ;
    wire new_AGEMA_signal_13761 ;
    wire new_AGEMA_signal_13762 ;
    wire new_AGEMA_signal_13763 ;
    wire new_AGEMA_signal_13764 ;
    wire new_AGEMA_signal_13765 ;
    wire new_AGEMA_signal_13766 ;
    wire new_AGEMA_signal_13767 ;
    wire new_AGEMA_signal_13768 ;
    wire new_AGEMA_signal_13769 ;
    wire new_AGEMA_signal_13770 ;
    wire new_AGEMA_signal_13771 ;
    wire new_AGEMA_signal_13772 ;
    wire new_AGEMA_signal_13773 ;
    wire new_AGEMA_signal_13774 ;
    wire new_AGEMA_signal_13775 ;
    wire new_AGEMA_signal_13776 ;
    wire new_AGEMA_signal_13777 ;
    wire new_AGEMA_signal_13778 ;
    wire new_AGEMA_signal_13779 ;
    wire new_AGEMA_signal_13780 ;
    wire new_AGEMA_signal_13781 ;
    wire new_AGEMA_signal_13782 ;
    wire new_AGEMA_signal_13783 ;
    wire new_AGEMA_signal_13784 ;
    wire new_AGEMA_signal_13785 ;
    wire new_AGEMA_signal_13786 ;
    wire new_AGEMA_signal_13787 ;
    wire new_AGEMA_signal_13788 ;
    wire new_AGEMA_signal_13789 ;
    wire new_AGEMA_signal_13790 ;
    wire new_AGEMA_signal_13791 ;
    wire new_AGEMA_signal_13792 ;
    wire new_AGEMA_signal_13793 ;
    wire new_AGEMA_signal_13794 ;
    wire new_AGEMA_signal_13795 ;
    wire new_AGEMA_signal_13796 ;
    wire new_AGEMA_signal_13797 ;
    wire new_AGEMA_signal_13798 ;
    wire new_AGEMA_signal_13799 ;
    wire new_AGEMA_signal_13800 ;
    wire new_AGEMA_signal_13801 ;
    wire new_AGEMA_signal_13802 ;
    wire new_AGEMA_signal_13803 ;
    wire new_AGEMA_signal_13804 ;
    wire new_AGEMA_signal_13805 ;
    wire new_AGEMA_signal_13806 ;
    wire new_AGEMA_signal_13807 ;
    wire new_AGEMA_signal_13808 ;
    wire new_AGEMA_signal_13809 ;
    wire new_AGEMA_signal_13810 ;
    wire new_AGEMA_signal_13811 ;
    wire new_AGEMA_signal_13812 ;
    wire new_AGEMA_signal_13813 ;
    wire new_AGEMA_signal_13814 ;
    wire new_AGEMA_signal_13815 ;
    wire new_AGEMA_signal_13816 ;
    wire new_AGEMA_signal_13817 ;
    wire new_AGEMA_signal_13818 ;
    wire new_AGEMA_signal_13819 ;
    wire new_AGEMA_signal_13820 ;
    wire new_AGEMA_signal_13821 ;
    wire new_AGEMA_signal_13822 ;
    wire new_AGEMA_signal_13823 ;
    wire new_AGEMA_signal_13824 ;
    wire new_AGEMA_signal_13825 ;
    wire new_AGEMA_signal_13826 ;
    wire new_AGEMA_signal_13827 ;
    wire new_AGEMA_signal_13828 ;
    wire new_AGEMA_signal_13829 ;
    wire new_AGEMA_signal_13830 ;
    wire new_AGEMA_signal_13831 ;
    wire new_AGEMA_signal_13832 ;
    wire new_AGEMA_signal_13833 ;
    wire new_AGEMA_signal_13834 ;
    wire new_AGEMA_signal_13835 ;
    wire new_AGEMA_signal_13836 ;
    wire new_AGEMA_signal_13837 ;
    wire new_AGEMA_signal_13838 ;
    wire new_AGEMA_signal_13839 ;
    wire new_AGEMA_signal_13840 ;
    wire new_AGEMA_signal_13841 ;
    wire new_AGEMA_signal_13842 ;
    wire new_AGEMA_signal_13843 ;
    wire new_AGEMA_signal_13844 ;
    wire new_AGEMA_signal_13845 ;
    wire new_AGEMA_signal_13846 ;
    wire new_AGEMA_signal_13847 ;
    wire new_AGEMA_signal_13848 ;
    wire new_AGEMA_signal_13849 ;
    wire new_AGEMA_signal_13850 ;
    wire new_AGEMA_signal_13851 ;
    wire new_AGEMA_signal_13852 ;
    wire new_AGEMA_signal_13853 ;
    wire new_AGEMA_signal_13854 ;
    wire new_AGEMA_signal_13855 ;
    wire new_AGEMA_signal_13856 ;
    wire new_AGEMA_signal_13857 ;
    wire new_AGEMA_signal_13858 ;
    wire new_AGEMA_signal_13859 ;
    wire new_AGEMA_signal_13860 ;
    wire new_AGEMA_signal_13861 ;
    wire new_AGEMA_signal_13862 ;
    wire new_AGEMA_signal_13863 ;
    wire new_AGEMA_signal_13864 ;
    wire new_AGEMA_signal_13865 ;
    wire new_AGEMA_signal_13866 ;
    wire new_AGEMA_signal_13867 ;
    wire new_AGEMA_signal_13868 ;
    wire new_AGEMA_signal_13869 ;
    wire new_AGEMA_signal_13870 ;
    wire new_AGEMA_signal_13871 ;
    wire new_AGEMA_signal_13872 ;
    wire new_AGEMA_signal_13873 ;
    wire new_AGEMA_signal_13874 ;
    wire new_AGEMA_signal_13875 ;
    wire new_AGEMA_signal_13876 ;
    wire new_AGEMA_signal_13877 ;
    wire new_AGEMA_signal_13878 ;
    wire new_AGEMA_signal_13879 ;
    wire new_AGEMA_signal_13880 ;
    wire new_AGEMA_signal_13881 ;
    wire new_AGEMA_signal_13882 ;
    wire new_AGEMA_signal_13883 ;
    wire new_AGEMA_signal_13884 ;
    wire new_AGEMA_signal_13885 ;
    wire new_AGEMA_signal_13886 ;
    wire new_AGEMA_signal_13887 ;
    wire new_AGEMA_signal_13888 ;
    wire new_AGEMA_signal_13889 ;
    wire new_AGEMA_signal_13890 ;
    wire new_AGEMA_signal_13891 ;
    wire new_AGEMA_signal_13892 ;
    wire new_AGEMA_signal_13893 ;
    wire new_AGEMA_signal_13894 ;
    wire new_AGEMA_signal_13895 ;
    wire new_AGEMA_signal_13896 ;
    wire new_AGEMA_signal_13897 ;
    wire new_AGEMA_signal_13898 ;
    wire new_AGEMA_signal_13899 ;
    wire new_AGEMA_signal_13900 ;
    wire new_AGEMA_signal_13901 ;
    wire new_AGEMA_signal_13902 ;
    wire new_AGEMA_signal_13903 ;
    wire new_AGEMA_signal_13904 ;
    wire new_AGEMA_signal_13905 ;
    wire new_AGEMA_signal_13906 ;
    wire new_AGEMA_signal_13907 ;
    wire new_AGEMA_signal_13908 ;
    wire new_AGEMA_signal_13909 ;
    wire new_AGEMA_signal_13910 ;
    wire new_AGEMA_signal_13911 ;
    wire new_AGEMA_signal_13912 ;
    wire new_AGEMA_signal_13913 ;
    wire new_AGEMA_signal_13914 ;
    wire new_AGEMA_signal_13915 ;
    wire new_AGEMA_signal_13916 ;
    wire new_AGEMA_signal_13917 ;
    wire new_AGEMA_signal_13918 ;
    wire new_AGEMA_signal_13919 ;
    wire new_AGEMA_signal_13920 ;
    wire new_AGEMA_signal_13921 ;
    wire new_AGEMA_signal_13922 ;
    wire new_AGEMA_signal_13923 ;
    wire new_AGEMA_signal_13924 ;
    wire new_AGEMA_signal_13925 ;
    wire new_AGEMA_signal_13926 ;
    wire new_AGEMA_signal_13927 ;
    wire new_AGEMA_signal_13928 ;
    wire new_AGEMA_signal_13929 ;
    wire new_AGEMA_signal_13930 ;
    wire new_AGEMA_signal_13931 ;
    wire new_AGEMA_signal_13932 ;
    wire new_AGEMA_signal_13933 ;
    wire new_AGEMA_signal_13934 ;
    wire new_AGEMA_signal_13935 ;
    wire new_AGEMA_signal_13936 ;
    wire new_AGEMA_signal_13937 ;
    wire new_AGEMA_signal_13938 ;
    wire new_AGEMA_signal_13939 ;
    wire new_AGEMA_signal_13940 ;
    wire new_AGEMA_signal_13941 ;
    wire new_AGEMA_signal_13942 ;
    wire new_AGEMA_signal_13943 ;
    wire new_AGEMA_signal_13944 ;
    wire new_AGEMA_signal_13945 ;
    wire new_AGEMA_signal_13946 ;
    wire new_AGEMA_signal_13947 ;
    wire new_AGEMA_signal_13948 ;
    wire new_AGEMA_signal_13949 ;
    wire new_AGEMA_signal_13950 ;
    wire new_AGEMA_signal_13951 ;
    wire new_AGEMA_signal_13952 ;
    wire new_AGEMA_signal_13953 ;
    wire new_AGEMA_signal_13954 ;
    wire new_AGEMA_signal_13955 ;
    wire new_AGEMA_signal_13956 ;
    wire new_AGEMA_signal_13957 ;
    wire new_AGEMA_signal_13958 ;
    wire new_AGEMA_signal_13959 ;
    wire new_AGEMA_signal_13960 ;
    wire new_AGEMA_signal_13961 ;
    wire new_AGEMA_signal_13962 ;
    wire new_AGEMA_signal_13963 ;
    wire new_AGEMA_signal_13964 ;
    wire new_AGEMA_signal_13965 ;
    wire new_AGEMA_signal_13966 ;
    wire new_AGEMA_signal_13967 ;
    wire new_AGEMA_signal_13968 ;
    wire new_AGEMA_signal_13969 ;
    wire new_AGEMA_signal_13970 ;
    wire new_AGEMA_signal_13971 ;
    wire new_AGEMA_signal_13972 ;
    wire new_AGEMA_signal_13973 ;
    wire new_AGEMA_signal_13974 ;
    wire new_AGEMA_signal_13975 ;
    wire new_AGEMA_signal_13976 ;
    wire new_AGEMA_signal_13977 ;
    wire new_AGEMA_signal_13978 ;
    wire new_AGEMA_signal_13979 ;
    wire new_AGEMA_signal_13980 ;
    wire new_AGEMA_signal_13981 ;
    wire new_AGEMA_signal_13982 ;
    wire new_AGEMA_signal_13983 ;
    wire new_AGEMA_signal_13984 ;
    wire new_AGEMA_signal_13985 ;
    wire new_AGEMA_signal_13986 ;
    wire new_AGEMA_signal_13987 ;
    wire new_AGEMA_signal_13988 ;
    wire new_AGEMA_signal_13989 ;
    wire new_AGEMA_signal_13990 ;
    wire new_AGEMA_signal_13991 ;
    wire new_AGEMA_signal_13992 ;
    wire new_AGEMA_signal_13993 ;
    wire new_AGEMA_signal_13994 ;
    wire new_AGEMA_signal_13995 ;
    wire new_AGEMA_signal_13996 ;
    wire new_AGEMA_signal_13997 ;
    wire new_AGEMA_signal_13998 ;
    wire new_AGEMA_signal_13999 ;
    wire new_AGEMA_signal_14000 ;
    wire new_AGEMA_signal_14001 ;
    wire new_AGEMA_signal_14002 ;
    wire new_AGEMA_signal_14003 ;
    wire new_AGEMA_signal_14004 ;
    wire new_AGEMA_signal_14005 ;
    wire new_AGEMA_signal_14006 ;
    wire new_AGEMA_signal_14007 ;
    wire new_AGEMA_signal_14008 ;
    wire new_AGEMA_signal_14009 ;
    wire new_AGEMA_signal_14010 ;
    wire new_AGEMA_signal_14011 ;
    wire new_AGEMA_signal_14012 ;
    wire new_AGEMA_signal_14013 ;
    wire new_AGEMA_signal_14014 ;
    wire new_AGEMA_signal_14015 ;
    wire new_AGEMA_signal_14016 ;
    wire new_AGEMA_signal_14017 ;
    wire new_AGEMA_signal_14018 ;
    wire new_AGEMA_signal_14019 ;
    wire new_AGEMA_signal_14020 ;
    wire new_AGEMA_signal_14021 ;
    wire new_AGEMA_signal_14022 ;
    wire new_AGEMA_signal_14023 ;
    wire new_AGEMA_signal_14024 ;
    wire new_AGEMA_signal_14025 ;
    wire new_AGEMA_signal_14026 ;
    wire new_AGEMA_signal_14027 ;
    wire new_AGEMA_signal_14028 ;
    wire new_AGEMA_signal_14029 ;
    wire new_AGEMA_signal_14030 ;
    wire new_AGEMA_signal_14031 ;
    wire new_AGEMA_signal_14032 ;
    wire new_AGEMA_signal_14033 ;
    wire new_AGEMA_signal_14034 ;
    wire new_AGEMA_signal_14035 ;
    wire new_AGEMA_signal_14036 ;
    wire new_AGEMA_signal_14037 ;
    wire new_AGEMA_signal_14038 ;
    wire new_AGEMA_signal_14039 ;
    wire new_AGEMA_signal_14040 ;
    wire new_AGEMA_signal_14041 ;
    wire new_AGEMA_signal_14042 ;
    wire new_AGEMA_signal_14043 ;
    wire new_AGEMA_signal_14044 ;
    wire new_AGEMA_signal_14045 ;
    wire new_AGEMA_signal_14046 ;
    wire new_AGEMA_signal_14047 ;
    wire new_AGEMA_signal_14048 ;
    wire new_AGEMA_signal_14049 ;
    wire new_AGEMA_signal_14050 ;
    wire new_AGEMA_signal_14051 ;
    wire new_AGEMA_signal_14052 ;
    wire new_AGEMA_signal_14053 ;
    wire new_AGEMA_signal_14054 ;
    wire new_AGEMA_signal_14055 ;
    wire new_AGEMA_signal_14056 ;
    wire new_AGEMA_signal_14057 ;
    wire new_AGEMA_signal_14058 ;
    wire new_AGEMA_signal_14059 ;
    wire new_AGEMA_signal_14060 ;
    wire new_AGEMA_signal_14061 ;
    wire new_AGEMA_signal_14062 ;
    wire new_AGEMA_signal_14063 ;
    wire new_AGEMA_signal_14064 ;
    wire new_AGEMA_signal_14065 ;
    wire new_AGEMA_signal_14066 ;
    wire new_AGEMA_signal_14067 ;
    wire new_AGEMA_signal_14068 ;
    wire new_AGEMA_signal_14069 ;
    wire new_AGEMA_signal_14070 ;
    wire new_AGEMA_signal_14071 ;
    wire new_AGEMA_signal_14072 ;
    wire new_AGEMA_signal_14073 ;
    wire new_AGEMA_signal_14074 ;
    wire new_AGEMA_signal_14075 ;
    wire new_AGEMA_signal_14076 ;
    wire new_AGEMA_signal_14077 ;
    wire new_AGEMA_signal_14078 ;
    wire new_AGEMA_signal_14079 ;
    wire new_AGEMA_signal_14080 ;
    wire new_AGEMA_signal_14081 ;
    wire new_AGEMA_signal_14082 ;
    wire new_AGEMA_signal_14083 ;
    wire new_AGEMA_signal_14084 ;
    wire new_AGEMA_signal_14085 ;
    wire new_AGEMA_signal_14086 ;
    wire new_AGEMA_signal_14087 ;
    wire new_AGEMA_signal_14088 ;
    wire new_AGEMA_signal_14089 ;
    wire new_AGEMA_signal_14090 ;
    wire new_AGEMA_signal_14091 ;
    wire new_AGEMA_signal_14092 ;
    wire new_AGEMA_signal_14093 ;
    wire new_AGEMA_signal_14094 ;
    wire new_AGEMA_signal_14095 ;
    wire new_AGEMA_signal_14096 ;
    wire new_AGEMA_signal_14097 ;
    wire new_AGEMA_signal_14098 ;
    wire new_AGEMA_signal_14099 ;
    wire new_AGEMA_signal_14100 ;
    wire new_AGEMA_signal_14101 ;
    wire new_AGEMA_signal_14102 ;
    wire new_AGEMA_signal_14103 ;
    wire new_AGEMA_signal_14104 ;
    wire new_AGEMA_signal_14105 ;
    wire new_AGEMA_signal_14106 ;
    wire new_AGEMA_signal_14107 ;
    wire new_AGEMA_signal_14108 ;
    wire new_AGEMA_signal_14109 ;
    wire new_AGEMA_signal_14110 ;
    wire new_AGEMA_signal_14111 ;
    wire new_AGEMA_signal_14112 ;
    wire new_AGEMA_signal_14113 ;
    wire new_AGEMA_signal_14114 ;
    wire new_AGEMA_signal_14115 ;
    wire new_AGEMA_signal_14116 ;
    wire new_AGEMA_signal_14117 ;
    wire new_AGEMA_signal_14118 ;
    wire new_AGEMA_signal_14119 ;
    wire new_AGEMA_signal_14120 ;
    wire new_AGEMA_signal_14121 ;
    wire new_AGEMA_signal_14122 ;
    wire new_AGEMA_signal_14123 ;
    wire new_AGEMA_signal_14124 ;
    wire new_AGEMA_signal_14125 ;
    wire new_AGEMA_signal_14126 ;
    wire new_AGEMA_signal_14127 ;
    wire new_AGEMA_signal_14128 ;
    wire new_AGEMA_signal_14129 ;
    wire new_AGEMA_signal_14130 ;
    wire new_AGEMA_signal_14131 ;
    wire new_AGEMA_signal_14132 ;
    wire new_AGEMA_signal_14133 ;
    wire new_AGEMA_signal_14134 ;
    wire new_AGEMA_signal_14135 ;
    wire new_AGEMA_signal_14136 ;
    wire new_AGEMA_signal_14137 ;
    wire new_AGEMA_signal_14138 ;
    wire new_AGEMA_signal_14139 ;
    wire new_AGEMA_signal_14140 ;
    wire new_AGEMA_signal_14141 ;
    wire new_AGEMA_signal_14142 ;
    wire new_AGEMA_signal_14143 ;
    wire new_AGEMA_signal_14144 ;
    wire new_AGEMA_signal_14145 ;
    wire new_AGEMA_signal_14146 ;
    wire new_AGEMA_signal_14147 ;
    wire new_AGEMA_signal_14148 ;
    wire new_AGEMA_signal_14149 ;
    wire new_AGEMA_signal_14150 ;
    wire new_AGEMA_signal_14151 ;
    wire new_AGEMA_signal_14152 ;
    wire new_AGEMA_signal_14153 ;
    wire new_AGEMA_signal_14154 ;
    wire new_AGEMA_signal_14155 ;
    wire new_AGEMA_signal_14156 ;
    wire new_AGEMA_signal_14157 ;
    wire new_AGEMA_signal_14158 ;
    wire new_AGEMA_signal_14159 ;
    wire new_AGEMA_signal_14160 ;
    wire new_AGEMA_signal_14161 ;
    wire new_AGEMA_signal_14162 ;
    wire new_AGEMA_signal_14163 ;
    wire new_AGEMA_signal_14164 ;
    wire new_AGEMA_signal_14165 ;
    wire new_AGEMA_signal_14166 ;
    wire new_AGEMA_signal_14167 ;
    wire new_AGEMA_signal_14168 ;
    wire new_AGEMA_signal_14169 ;
    wire new_AGEMA_signal_14170 ;
    wire new_AGEMA_signal_14171 ;
    wire new_AGEMA_signal_14172 ;
    wire new_AGEMA_signal_14173 ;
    wire new_AGEMA_signal_14174 ;
    wire new_AGEMA_signal_14175 ;
    wire new_AGEMA_signal_14176 ;
    wire new_AGEMA_signal_14177 ;
    wire new_AGEMA_signal_14178 ;
    wire new_AGEMA_signal_14179 ;
    wire new_AGEMA_signal_14180 ;
    wire new_AGEMA_signal_14181 ;
    wire new_AGEMA_signal_14182 ;
    wire new_AGEMA_signal_14183 ;
    wire new_AGEMA_signal_14184 ;
    wire new_AGEMA_signal_14185 ;
    wire new_AGEMA_signal_14186 ;
    wire new_AGEMA_signal_14187 ;
    wire new_AGEMA_signal_14188 ;
    wire new_AGEMA_signal_14189 ;
    wire new_AGEMA_signal_14190 ;
    wire new_AGEMA_signal_14191 ;
    wire new_AGEMA_signal_14192 ;
    wire new_AGEMA_signal_14193 ;
    wire new_AGEMA_signal_14194 ;
    wire new_AGEMA_signal_14195 ;
    wire new_AGEMA_signal_14196 ;
    wire new_AGEMA_signal_14197 ;
    wire new_AGEMA_signal_14198 ;
    wire new_AGEMA_signal_14199 ;
    wire new_AGEMA_signal_14200 ;
    wire new_AGEMA_signal_14201 ;
    wire new_AGEMA_signal_14202 ;
    wire new_AGEMA_signal_14203 ;
    wire new_AGEMA_signal_14204 ;
    wire new_AGEMA_signal_14205 ;
    wire new_AGEMA_signal_14206 ;
    wire new_AGEMA_signal_14207 ;
    wire new_AGEMA_signal_14208 ;
    wire new_AGEMA_signal_14209 ;
    wire new_AGEMA_signal_14210 ;
    wire new_AGEMA_signal_14211 ;
    wire new_AGEMA_signal_14212 ;
    wire new_AGEMA_signal_14213 ;
    wire new_AGEMA_signal_14214 ;
    wire new_AGEMA_signal_14215 ;
    wire new_AGEMA_signal_14216 ;
    wire new_AGEMA_signal_14217 ;
    wire new_AGEMA_signal_14218 ;
    wire new_AGEMA_signal_14219 ;
    wire new_AGEMA_signal_14220 ;
    wire new_AGEMA_signal_14221 ;
    wire new_AGEMA_signal_14222 ;
    wire new_AGEMA_signal_14223 ;
    wire new_AGEMA_signal_14224 ;
    wire new_AGEMA_signal_14225 ;
    wire new_AGEMA_signal_14226 ;
    wire new_AGEMA_signal_14227 ;
    wire new_AGEMA_signal_14228 ;
    wire new_AGEMA_signal_14229 ;
    wire new_AGEMA_signal_14230 ;
    wire new_AGEMA_signal_14231 ;
    wire new_AGEMA_signal_14232 ;
    wire new_AGEMA_signal_14233 ;
    wire new_AGEMA_signal_14234 ;
    wire new_AGEMA_signal_14235 ;
    wire new_AGEMA_signal_14236 ;
    wire new_AGEMA_signal_14237 ;
    wire new_AGEMA_signal_14238 ;
    wire new_AGEMA_signal_14239 ;
    wire new_AGEMA_signal_14240 ;
    wire new_AGEMA_signal_14241 ;
    wire new_AGEMA_signal_14242 ;
    wire new_AGEMA_signal_14243 ;
    wire new_AGEMA_signal_14244 ;
    wire new_AGEMA_signal_14245 ;
    wire new_AGEMA_signal_14246 ;
    wire new_AGEMA_signal_14247 ;
    wire new_AGEMA_signal_14248 ;
    wire new_AGEMA_signal_14249 ;
    wire new_AGEMA_signal_14250 ;
    wire new_AGEMA_signal_14251 ;
    wire new_AGEMA_signal_14252 ;
    wire new_AGEMA_signal_14253 ;
    wire new_AGEMA_signal_14254 ;
    wire new_AGEMA_signal_14255 ;
    wire new_AGEMA_signal_14256 ;
    wire new_AGEMA_signal_14257 ;
    wire new_AGEMA_signal_14258 ;
    wire new_AGEMA_signal_14259 ;
    wire new_AGEMA_signal_14260 ;
    wire new_AGEMA_signal_14261 ;
    wire new_AGEMA_signal_14262 ;
    wire new_AGEMA_signal_14263 ;
    wire new_AGEMA_signal_14264 ;
    wire new_AGEMA_signal_14265 ;
    wire new_AGEMA_signal_14266 ;
    wire new_AGEMA_signal_14267 ;
    wire new_AGEMA_signal_14268 ;
    wire new_AGEMA_signal_14269 ;
    wire new_AGEMA_signal_14270 ;
    wire new_AGEMA_signal_14271 ;
    wire new_AGEMA_signal_14272 ;
    wire new_AGEMA_signal_14273 ;
    wire new_AGEMA_signal_14274 ;
    wire new_AGEMA_signal_14275 ;
    wire new_AGEMA_signal_14276 ;
    wire new_AGEMA_signal_14277 ;
    wire new_AGEMA_signal_14278 ;
    wire new_AGEMA_signal_14279 ;
    wire new_AGEMA_signal_14280 ;
    wire new_AGEMA_signal_14281 ;
    wire new_AGEMA_signal_14282 ;
    wire new_AGEMA_signal_14283 ;
    wire new_AGEMA_signal_14284 ;
    wire new_AGEMA_signal_14285 ;
    wire new_AGEMA_signal_14286 ;
    wire new_AGEMA_signal_14287 ;
    wire new_AGEMA_signal_14288 ;
    wire new_AGEMA_signal_14289 ;
    wire new_AGEMA_signal_14290 ;
    wire new_AGEMA_signal_14291 ;
    wire new_AGEMA_signal_14292 ;
    wire new_AGEMA_signal_14293 ;
    wire new_AGEMA_signal_14294 ;
    wire new_AGEMA_signal_14295 ;
    wire new_AGEMA_signal_14296 ;
    wire new_AGEMA_signal_14297 ;
    wire new_AGEMA_signal_14298 ;
    wire new_AGEMA_signal_14299 ;
    wire new_AGEMA_signal_14300 ;
    wire new_AGEMA_signal_14301 ;
    wire new_AGEMA_signal_14302 ;
    wire new_AGEMA_signal_14303 ;
    wire new_AGEMA_signal_14304 ;
    wire new_AGEMA_signal_14305 ;
    wire new_AGEMA_signal_14306 ;
    wire new_AGEMA_signal_14307 ;
    wire new_AGEMA_signal_14308 ;
    wire new_AGEMA_signal_14309 ;
    wire new_AGEMA_signal_14310 ;
    wire new_AGEMA_signal_14311 ;
    wire new_AGEMA_signal_14312 ;
    wire new_AGEMA_signal_14313 ;
    wire new_AGEMA_signal_14314 ;
    wire new_AGEMA_signal_14315 ;
    wire new_AGEMA_signal_14316 ;
    wire new_AGEMA_signal_14317 ;
    wire new_AGEMA_signal_14318 ;
    wire new_AGEMA_signal_14319 ;
    wire new_AGEMA_signal_14320 ;
    wire new_AGEMA_signal_14321 ;
    wire new_AGEMA_signal_14322 ;
    wire new_AGEMA_signal_14323 ;
    wire new_AGEMA_signal_14324 ;
    wire new_AGEMA_signal_14325 ;
    wire new_AGEMA_signal_14326 ;
    wire new_AGEMA_signal_14327 ;
    wire new_AGEMA_signal_14328 ;
    wire new_AGEMA_signal_14329 ;
    wire new_AGEMA_signal_14330 ;
    wire new_AGEMA_signal_14331 ;
    wire new_AGEMA_signal_14332 ;
    wire new_AGEMA_signal_14333 ;
    wire new_AGEMA_signal_14334 ;
    wire new_AGEMA_signal_14335 ;
    wire new_AGEMA_signal_14336 ;
    wire new_AGEMA_signal_14337 ;
    wire new_AGEMA_signal_14338 ;
    wire new_AGEMA_signal_14339 ;
    wire new_AGEMA_signal_14340 ;
    wire new_AGEMA_signal_14341 ;
    wire new_AGEMA_signal_14342 ;
    wire new_AGEMA_signal_14343 ;
    wire new_AGEMA_signal_14344 ;
    wire new_AGEMA_signal_14345 ;
    wire new_AGEMA_signal_14346 ;
    wire new_AGEMA_signal_14347 ;
    wire new_AGEMA_signal_14348 ;
    wire new_AGEMA_signal_14349 ;
    wire new_AGEMA_signal_14350 ;
    wire new_AGEMA_signal_14351 ;
    wire new_AGEMA_signal_14352 ;
    wire new_AGEMA_signal_14353 ;
    wire new_AGEMA_signal_14354 ;
    wire new_AGEMA_signal_14355 ;
    wire new_AGEMA_signal_14356 ;
    wire new_AGEMA_signal_14357 ;
    wire new_AGEMA_signal_14358 ;
    wire new_AGEMA_signal_14359 ;
    wire new_AGEMA_signal_14360 ;
    wire new_AGEMA_signal_14361 ;
    wire new_AGEMA_signal_14362 ;
    wire new_AGEMA_signal_14363 ;
    wire new_AGEMA_signal_14364 ;
    wire new_AGEMA_signal_14365 ;
    wire new_AGEMA_signal_14366 ;
    wire new_AGEMA_signal_14367 ;
    wire new_AGEMA_signal_14368 ;
    wire new_AGEMA_signal_14369 ;
    wire new_AGEMA_signal_14370 ;
    wire new_AGEMA_signal_14371 ;
    wire new_AGEMA_signal_14372 ;
    wire new_AGEMA_signal_14373 ;
    wire new_AGEMA_signal_14374 ;
    wire new_AGEMA_signal_14375 ;
    wire new_AGEMA_signal_14376 ;
    wire new_AGEMA_signal_14377 ;
    wire new_AGEMA_signal_14378 ;
    wire new_AGEMA_signal_14379 ;
    wire new_AGEMA_signal_14380 ;
    wire new_AGEMA_signal_14381 ;
    wire new_AGEMA_signal_14382 ;
    wire new_AGEMA_signal_14383 ;
    wire new_AGEMA_signal_14384 ;
    wire new_AGEMA_signal_14385 ;
    wire new_AGEMA_signal_14386 ;
    wire new_AGEMA_signal_14387 ;
    wire new_AGEMA_signal_14388 ;
    wire new_AGEMA_signal_14389 ;
    wire new_AGEMA_signal_14390 ;
    wire new_AGEMA_signal_14391 ;
    wire new_AGEMA_signal_14392 ;
    wire new_AGEMA_signal_14393 ;
    wire new_AGEMA_signal_14394 ;
    wire new_AGEMA_signal_14395 ;
    wire new_AGEMA_signal_14396 ;
    wire new_AGEMA_signal_14397 ;
    wire new_AGEMA_signal_14398 ;
    wire new_AGEMA_signal_14399 ;
    wire new_AGEMA_signal_14400 ;
    wire new_AGEMA_signal_14401 ;
    wire new_AGEMA_signal_14402 ;
    wire new_AGEMA_signal_14403 ;
    wire new_AGEMA_signal_14404 ;
    wire new_AGEMA_signal_14405 ;
    wire new_AGEMA_signal_14406 ;
    wire new_AGEMA_signal_14407 ;
    wire new_AGEMA_signal_14408 ;
    wire new_AGEMA_signal_14409 ;
    wire new_AGEMA_signal_14410 ;
    wire new_AGEMA_signal_14411 ;
    wire new_AGEMA_signal_14412 ;
    wire new_AGEMA_signal_14413 ;
    wire new_AGEMA_signal_14414 ;
    wire new_AGEMA_signal_14415 ;
    wire new_AGEMA_signal_14416 ;
    wire new_AGEMA_signal_14417 ;
    wire new_AGEMA_signal_14418 ;
    wire new_AGEMA_signal_14419 ;
    wire new_AGEMA_signal_14420 ;
    wire new_AGEMA_signal_14421 ;
    wire new_AGEMA_signal_14422 ;
    wire new_AGEMA_signal_14423 ;
    wire new_AGEMA_signal_14424 ;
    wire new_AGEMA_signal_14425 ;
    wire new_AGEMA_signal_14426 ;
    wire new_AGEMA_signal_14427 ;
    wire new_AGEMA_signal_14428 ;
    wire new_AGEMA_signal_14429 ;
    wire new_AGEMA_signal_14430 ;
    wire new_AGEMA_signal_14431 ;
    wire new_AGEMA_signal_14432 ;
    wire new_AGEMA_signal_14433 ;
    wire new_AGEMA_signal_14434 ;
    wire new_AGEMA_signal_14435 ;
    wire new_AGEMA_signal_14436 ;
    wire new_AGEMA_signal_14437 ;
    wire new_AGEMA_signal_14438 ;
    wire new_AGEMA_signal_14439 ;
    wire new_AGEMA_signal_14440 ;
    wire new_AGEMA_signal_14441 ;
    wire new_AGEMA_signal_14442 ;
    wire new_AGEMA_signal_14443 ;
    wire new_AGEMA_signal_14444 ;
    wire new_AGEMA_signal_14445 ;
    wire new_AGEMA_signal_14446 ;
    wire new_AGEMA_signal_14447 ;
    wire new_AGEMA_signal_14448 ;
    wire new_AGEMA_signal_14449 ;
    wire new_AGEMA_signal_14450 ;
    wire new_AGEMA_signal_14451 ;
    wire new_AGEMA_signal_14452 ;
    wire new_AGEMA_signal_14453 ;
    wire new_AGEMA_signal_14454 ;
    wire new_AGEMA_signal_14455 ;
    wire new_AGEMA_signal_14456 ;
    wire new_AGEMA_signal_14457 ;
    wire new_AGEMA_signal_14458 ;
    wire new_AGEMA_signal_14459 ;
    wire new_AGEMA_signal_14460 ;
    wire new_AGEMA_signal_14461 ;
    wire new_AGEMA_signal_14462 ;
    wire new_AGEMA_signal_14463 ;
    wire new_AGEMA_signal_14464 ;
    wire new_AGEMA_signal_14465 ;
    wire new_AGEMA_signal_14466 ;
    wire new_AGEMA_signal_14467 ;
    wire new_AGEMA_signal_14468 ;
    wire new_AGEMA_signal_14469 ;
    wire new_AGEMA_signal_14470 ;
    wire new_AGEMA_signal_14471 ;
    wire new_AGEMA_signal_14472 ;
    wire new_AGEMA_signal_14473 ;
    wire new_AGEMA_signal_14474 ;
    wire new_AGEMA_signal_14475 ;
    wire new_AGEMA_signal_14476 ;
    wire new_AGEMA_signal_14477 ;
    wire new_AGEMA_signal_14478 ;
    wire new_AGEMA_signal_14479 ;
    wire new_AGEMA_signal_14480 ;
    wire new_AGEMA_signal_14481 ;
    wire new_AGEMA_signal_14482 ;
    wire new_AGEMA_signal_14483 ;
    wire new_AGEMA_signal_14484 ;
    wire new_AGEMA_signal_14485 ;
    wire new_AGEMA_signal_14486 ;
    wire new_AGEMA_signal_14487 ;
    wire new_AGEMA_signal_14488 ;
    wire new_AGEMA_signal_14489 ;
    wire new_AGEMA_signal_14490 ;
    wire new_AGEMA_signal_14491 ;
    wire new_AGEMA_signal_14492 ;
    wire new_AGEMA_signal_14493 ;
    wire new_AGEMA_signal_14494 ;
    wire new_AGEMA_signal_14495 ;
    wire new_AGEMA_signal_14496 ;
    wire new_AGEMA_signal_14497 ;
    wire new_AGEMA_signal_14498 ;
    wire new_AGEMA_signal_14499 ;
    wire new_AGEMA_signal_14500 ;
    wire new_AGEMA_signal_14501 ;
    wire new_AGEMA_signal_14502 ;
    wire new_AGEMA_signal_14503 ;
    wire new_AGEMA_signal_14504 ;
    wire new_AGEMA_signal_14505 ;
    wire new_AGEMA_signal_14506 ;
    wire new_AGEMA_signal_14507 ;
    wire new_AGEMA_signal_14508 ;
    wire new_AGEMA_signal_14509 ;
    wire new_AGEMA_signal_14510 ;
    wire new_AGEMA_signal_14511 ;
    wire new_AGEMA_signal_14512 ;
    wire new_AGEMA_signal_14513 ;
    wire new_AGEMA_signal_14514 ;
    wire new_AGEMA_signal_14515 ;
    wire new_AGEMA_signal_14516 ;
    wire new_AGEMA_signal_14517 ;
    wire new_AGEMA_signal_14518 ;
    wire new_AGEMA_signal_14519 ;
    wire new_AGEMA_signal_14520 ;
    wire new_AGEMA_signal_14521 ;
    wire new_AGEMA_signal_14522 ;
    wire new_AGEMA_signal_14523 ;
    wire new_AGEMA_signal_14524 ;
    wire new_AGEMA_signal_14525 ;
    wire new_AGEMA_signal_14526 ;
    wire new_AGEMA_signal_14527 ;
    wire new_AGEMA_signal_14528 ;
    wire new_AGEMA_signal_14529 ;
    wire new_AGEMA_signal_14530 ;
    wire new_AGEMA_signal_14531 ;
    wire new_AGEMA_signal_14532 ;
    wire new_AGEMA_signal_14533 ;
    wire new_AGEMA_signal_14534 ;
    wire new_AGEMA_signal_14535 ;
    wire new_AGEMA_signal_14536 ;
    wire new_AGEMA_signal_14537 ;
    wire new_AGEMA_signal_14538 ;
    wire new_AGEMA_signal_14539 ;
    wire new_AGEMA_signal_14540 ;
    wire new_AGEMA_signal_14541 ;
    wire new_AGEMA_signal_14542 ;
    wire new_AGEMA_signal_14543 ;
    wire new_AGEMA_signal_14544 ;
    wire new_AGEMA_signal_14545 ;
    wire new_AGEMA_signal_14546 ;
    wire new_AGEMA_signal_14547 ;
    wire new_AGEMA_signal_14548 ;
    wire new_AGEMA_signal_14549 ;
    wire new_AGEMA_signal_14550 ;
    wire new_AGEMA_signal_14551 ;
    wire new_AGEMA_signal_14552 ;
    wire new_AGEMA_signal_14553 ;
    wire new_AGEMA_signal_14554 ;
    wire new_AGEMA_signal_14555 ;
    wire new_AGEMA_signal_14556 ;
    wire new_AGEMA_signal_14557 ;
    wire new_AGEMA_signal_14558 ;
    wire new_AGEMA_signal_14559 ;
    wire new_AGEMA_signal_14560 ;
    wire new_AGEMA_signal_14561 ;
    wire new_AGEMA_signal_14562 ;
    wire new_AGEMA_signal_14563 ;
    wire new_AGEMA_signal_14564 ;
    wire new_AGEMA_signal_14565 ;
    wire new_AGEMA_signal_14566 ;
    wire new_AGEMA_signal_14567 ;
    wire new_AGEMA_signal_14568 ;
    wire new_AGEMA_signal_14569 ;
    wire new_AGEMA_signal_14570 ;
    wire new_AGEMA_signal_14571 ;
    wire new_AGEMA_signal_14572 ;
    wire new_AGEMA_signal_14573 ;
    wire new_AGEMA_signal_14574 ;
    wire new_AGEMA_signal_14575 ;
    wire new_AGEMA_signal_14576 ;
    wire new_AGEMA_signal_14577 ;
    wire new_AGEMA_signal_14578 ;
    wire new_AGEMA_signal_14579 ;
    wire new_AGEMA_signal_14580 ;
    wire new_AGEMA_signal_14581 ;
    wire new_AGEMA_signal_14582 ;
    wire new_AGEMA_signal_14583 ;
    wire new_AGEMA_signal_14584 ;
    wire new_AGEMA_signal_14585 ;
    wire new_AGEMA_signal_14586 ;
    wire new_AGEMA_signal_14587 ;
    wire new_AGEMA_signal_14588 ;
    wire new_AGEMA_signal_14589 ;
    wire new_AGEMA_signal_14590 ;
    wire new_AGEMA_signal_14591 ;
    wire new_AGEMA_signal_14592 ;
    wire new_AGEMA_signal_14593 ;
    wire new_AGEMA_signal_14594 ;
    wire new_AGEMA_signal_14595 ;
    wire new_AGEMA_signal_14596 ;
    wire new_AGEMA_signal_14597 ;
    wire new_AGEMA_signal_14598 ;
    wire new_AGEMA_signal_14599 ;
    wire new_AGEMA_signal_14600 ;
    wire new_AGEMA_signal_14601 ;
    wire new_AGEMA_signal_14602 ;
    wire new_AGEMA_signal_14603 ;
    wire new_AGEMA_signal_14604 ;
    wire new_AGEMA_signal_14605 ;
    wire new_AGEMA_signal_14606 ;
    wire new_AGEMA_signal_14607 ;
    wire new_AGEMA_signal_14608 ;
    wire new_AGEMA_signal_14609 ;
    wire new_AGEMA_signal_14610 ;
    wire new_AGEMA_signal_14611 ;
    wire new_AGEMA_signal_14612 ;
    wire new_AGEMA_signal_14613 ;
    wire new_AGEMA_signal_14614 ;
    wire new_AGEMA_signal_14615 ;
    wire new_AGEMA_signal_14616 ;
    wire new_AGEMA_signal_14617 ;
    wire new_AGEMA_signal_14618 ;
    wire new_AGEMA_signal_14619 ;
    wire new_AGEMA_signal_14620 ;
    wire new_AGEMA_signal_14621 ;
    wire new_AGEMA_signal_14622 ;
    wire new_AGEMA_signal_14623 ;
    wire new_AGEMA_signal_14624 ;
    wire new_AGEMA_signal_14625 ;
    wire new_AGEMA_signal_14626 ;
    wire new_AGEMA_signal_14627 ;
    wire new_AGEMA_signal_14628 ;
    wire new_AGEMA_signal_14629 ;
    wire new_AGEMA_signal_14630 ;
    wire new_AGEMA_signal_14631 ;
    wire new_AGEMA_signal_14632 ;
    wire new_AGEMA_signal_14633 ;
    wire new_AGEMA_signal_14634 ;
    wire new_AGEMA_signal_14635 ;
    wire new_AGEMA_signal_14636 ;
    wire new_AGEMA_signal_14637 ;
    wire new_AGEMA_signal_14638 ;
    wire new_AGEMA_signal_14639 ;
    wire new_AGEMA_signal_14640 ;
    wire new_AGEMA_signal_14641 ;
    wire new_AGEMA_signal_14642 ;
    wire new_AGEMA_signal_14643 ;
    wire new_AGEMA_signal_14644 ;
    wire new_AGEMA_signal_14645 ;
    wire new_AGEMA_signal_14646 ;
    wire new_AGEMA_signal_14647 ;
    wire new_AGEMA_signal_14648 ;
    wire new_AGEMA_signal_14649 ;
    wire new_AGEMA_signal_14650 ;
    wire new_AGEMA_signal_14651 ;
    wire new_AGEMA_signal_14652 ;
    wire new_AGEMA_signal_14653 ;
    wire new_AGEMA_signal_14654 ;
    wire new_AGEMA_signal_14655 ;
    wire new_AGEMA_signal_14656 ;
    wire new_AGEMA_signal_14657 ;
    wire new_AGEMA_signal_14658 ;
    wire new_AGEMA_signal_14659 ;
    wire new_AGEMA_signal_14660 ;
    wire new_AGEMA_signal_14661 ;
    wire new_AGEMA_signal_14662 ;
    wire new_AGEMA_signal_14663 ;
    wire new_AGEMA_signal_14664 ;
    wire new_AGEMA_signal_14665 ;
    wire new_AGEMA_signal_14666 ;
    wire new_AGEMA_signal_14667 ;
    wire new_AGEMA_signal_14668 ;
    wire new_AGEMA_signal_14669 ;
    wire new_AGEMA_signal_14670 ;
    wire new_AGEMA_signal_14671 ;
    wire new_AGEMA_signal_14672 ;
    wire new_AGEMA_signal_14673 ;
    wire new_AGEMA_signal_14674 ;
    wire new_AGEMA_signal_14675 ;
    wire new_AGEMA_signal_14676 ;
    wire new_AGEMA_signal_14677 ;
    wire new_AGEMA_signal_14678 ;
    wire new_AGEMA_signal_14679 ;
    wire new_AGEMA_signal_14680 ;
    wire new_AGEMA_signal_14681 ;
    wire new_AGEMA_signal_14682 ;
    wire new_AGEMA_signal_14683 ;
    wire new_AGEMA_signal_14684 ;
    wire new_AGEMA_signal_14685 ;
    wire new_AGEMA_signal_14686 ;
    wire new_AGEMA_signal_14687 ;
    wire new_AGEMA_signal_14688 ;
    wire new_AGEMA_signal_14689 ;
    wire new_AGEMA_signal_14690 ;
    wire new_AGEMA_signal_14691 ;
    wire new_AGEMA_signal_14692 ;
    wire new_AGEMA_signal_14693 ;
    wire new_AGEMA_signal_14694 ;
    wire new_AGEMA_signal_14695 ;
    wire new_AGEMA_signal_14696 ;
    wire new_AGEMA_signal_14697 ;
    wire new_AGEMA_signal_14698 ;
    wire new_AGEMA_signal_14699 ;
    wire new_AGEMA_signal_14700 ;
    wire new_AGEMA_signal_14701 ;
    wire new_AGEMA_signal_14702 ;
    wire new_AGEMA_signal_14703 ;
    wire new_AGEMA_signal_14704 ;
    wire new_AGEMA_signal_14705 ;
    wire new_AGEMA_signal_14706 ;
    wire new_AGEMA_signal_14707 ;
    wire new_AGEMA_signal_14708 ;
    wire new_AGEMA_signal_14709 ;
    wire new_AGEMA_signal_14710 ;
    wire new_AGEMA_signal_14711 ;
    wire new_AGEMA_signal_14712 ;
    wire new_AGEMA_signal_14713 ;
    wire new_AGEMA_signal_14714 ;
    wire new_AGEMA_signal_14715 ;
    wire new_AGEMA_signal_14716 ;
    wire new_AGEMA_signal_14717 ;
    wire new_AGEMA_signal_14718 ;
    wire new_AGEMA_signal_14719 ;
    wire new_AGEMA_signal_14720 ;
    wire new_AGEMA_signal_14721 ;
    wire new_AGEMA_signal_14722 ;
    wire new_AGEMA_signal_14723 ;
    wire new_AGEMA_signal_14724 ;
    wire new_AGEMA_signal_14725 ;
    wire new_AGEMA_signal_14726 ;
    wire new_AGEMA_signal_14727 ;
    wire new_AGEMA_signal_14728 ;
    wire new_AGEMA_signal_14729 ;
    wire new_AGEMA_signal_14730 ;
    wire new_AGEMA_signal_14731 ;
    wire new_AGEMA_signal_14732 ;
    wire new_AGEMA_signal_14733 ;
    wire new_AGEMA_signal_14734 ;
    wire new_AGEMA_signal_14735 ;
    wire new_AGEMA_signal_14736 ;
    wire new_AGEMA_signal_14737 ;
    wire new_AGEMA_signal_14738 ;
    wire new_AGEMA_signal_14739 ;
    wire new_AGEMA_signal_14740 ;
    wire new_AGEMA_signal_14741 ;
    wire new_AGEMA_signal_14742 ;
    wire new_AGEMA_signal_14743 ;
    wire new_AGEMA_signal_14744 ;
    wire new_AGEMA_signal_14745 ;
    wire new_AGEMA_signal_14746 ;
    wire new_AGEMA_signal_14747 ;
    wire new_AGEMA_signal_14748 ;
    wire new_AGEMA_signal_14749 ;
    wire new_AGEMA_signal_14750 ;
    wire new_AGEMA_signal_14751 ;
    wire new_AGEMA_signal_14752 ;
    wire new_AGEMA_signal_14753 ;
    wire new_AGEMA_signal_14754 ;
    wire new_AGEMA_signal_14755 ;
    wire new_AGEMA_signal_14756 ;
    wire new_AGEMA_signal_14757 ;
    wire new_AGEMA_signal_14758 ;
    wire new_AGEMA_signal_14759 ;
    wire new_AGEMA_signal_14760 ;
    wire new_AGEMA_signal_14761 ;
    wire new_AGEMA_signal_14762 ;
    wire new_AGEMA_signal_14763 ;
    wire new_AGEMA_signal_14764 ;
    wire new_AGEMA_signal_14765 ;
    wire new_AGEMA_signal_14766 ;
    wire new_AGEMA_signal_14767 ;
    wire new_AGEMA_signal_14768 ;
    wire new_AGEMA_signal_14769 ;
    wire new_AGEMA_signal_14770 ;
    wire new_AGEMA_signal_14771 ;
    wire new_AGEMA_signal_14772 ;
    wire new_AGEMA_signal_14773 ;
    wire new_AGEMA_signal_14774 ;
    wire new_AGEMA_signal_14775 ;
    wire new_AGEMA_signal_14776 ;
    wire new_AGEMA_signal_14777 ;
    wire new_AGEMA_signal_14778 ;
    wire new_AGEMA_signal_14779 ;
    wire new_AGEMA_signal_14780 ;
    wire new_AGEMA_signal_14781 ;
    wire new_AGEMA_signal_14782 ;
    wire new_AGEMA_signal_14783 ;
    wire new_AGEMA_signal_14784 ;
    wire new_AGEMA_signal_14785 ;
    wire new_AGEMA_signal_14786 ;
    wire new_AGEMA_signal_14787 ;
    wire new_AGEMA_signal_14788 ;
    wire new_AGEMA_signal_14789 ;
    wire new_AGEMA_signal_14790 ;
    wire new_AGEMA_signal_14791 ;
    wire new_AGEMA_signal_14792 ;
    wire new_AGEMA_signal_14793 ;
    wire new_AGEMA_signal_14794 ;
    wire new_AGEMA_signal_14795 ;
    wire new_AGEMA_signal_14796 ;
    wire new_AGEMA_signal_14797 ;
    wire new_AGEMA_signal_14798 ;
    wire new_AGEMA_signal_14799 ;
    wire new_AGEMA_signal_14800 ;
    wire new_AGEMA_signal_14801 ;
    wire new_AGEMA_signal_14802 ;
    wire new_AGEMA_signal_14803 ;
    wire new_AGEMA_signal_14804 ;
    wire new_AGEMA_signal_14805 ;
    wire new_AGEMA_signal_14806 ;
    wire new_AGEMA_signal_14807 ;
    wire new_AGEMA_signal_14808 ;
    wire new_AGEMA_signal_14809 ;
    wire new_AGEMA_signal_14810 ;
    wire new_AGEMA_signal_14811 ;
    wire new_AGEMA_signal_14812 ;
    wire new_AGEMA_signal_14813 ;
    wire new_AGEMA_signal_14814 ;
    wire new_AGEMA_signal_14815 ;
    wire new_AGEMA_signal_14816 ;
    wire new_AGEMA_signal_14817 ;
    wire new_AGEMA_signal_14818 ;
    wire new_AGEMA_signal_14819 ;
    wire new_AGEMA_signal_14820 ;
    wire new_AGEMA_signal_14821 ;
    wire new_AGEMA_signal_14822 ;
    wire new_AGEMA_signal_14823 ;
    wire new_AGEMA_signal_14824 ;
    wire new_AGEMA_signal_14825 ;
    wire new_AGEMA_signal_14826 ;
    wire new_AGEMA_signal_14827 ;
    wire new_AGEMA_signal_14828 ;
    wire new_AGEMA_signal_14829 ;
    wire new_AGEMA_signal_14830 ;
    wire new_AGEMA_signal_14831 ;
    wire new_AGEMA_signal_14832 ;
    wire new_AGEMA_signal_14833 ;
    wire new_AGEMA_signal_14834 ;
    wire new_AGEMA_signal_14835 ;
    wire new_AGEMA_signal_14836 ;
    wire new_AGEMA_signal_14837 ;
    wire new_AGEMA_signal_14838 ;
    wire new_AGEMA_signal_14839 ;
    wire new_AGEMA_signal_14840 ;
    wire new_AGEMA_signal_14841 ;
    wire new_AGEMA_signal_14842 ;
    wire new_AGEMA_signal_14843 ;
    wire new_AGEMA_signal_14844 ;
    wire new_AGEMA_signal_14845 ;
    wire new_AGEMA_signal_14846 ;
    wire new_AGEMA_signal_14847 ;
    wire new_AGEMA_signal_14848 ;
    wire new_AGEMA_signal_14849 ;
    wire new_AGEMA_signal_14850 ;
    wire new_AGEMA_signal_14851 ;
    wire new_AGEMA_signal_14852 ;
    wire new_AGEMA_signal_14853 ;
    wire new_AGEMA_signal_14854 ;
    wire new_AGEMA_signal_14855 ;
    wire new_AGEMA_signal_14856 ;
    wire new_AGEMA_signal_14857 ;
    wire new_AGEMA_signal_14858 ;
    wire new_AGEMA_signal_14859 ;
    wire new_AGEMA_signal_14860 ;
    wire new_AGEMA_signal_14861 ;
    wire new_AGEMA_signal_14862 ;
    wire new_AGEMA_signal_14863 ;
    wire new_AGEMA_signal_14864 ;
    wire new_AGEMA_signal_14865 ;
    wire new_AGEMA_signal_14866 ;
    wire new_AGEMA_signal_14867 ;
    wire new_AGEMA_signal_14868 ;
    wire new_AGEMA_signal_14869 ;
    wire new_AGEMA_signal_14870 ;
    wire new_AGEMA_signal_14871 ;
    wire new_AGEMA_signal_14872 ;
    wire new_AGEMA_signal_14873 ;
    wire new_AGEMA_signal_14874 ;
    wire new_AGEMA_signal_14875 ;
    wire new_AGEMA_signal_14876 ;
    wire new_AGEMA_signal_14877 ;
    wire new_AGEMA_signal_14878 ;
    wire new_AGEMA_signal_14879 ;
    wire new_AGEMA_signal_14880 ;
    wire new_AGEMA_signal_14881 ;
    wire new_AGEMA_signal_14882 ;
    wire new_AGEMA_signal_14883 ;
    wire new_AGEMA_signal_14884 ;
    wire new_AGEMA_signal_14885 ;
    wire new_AGEMA_signal_14886 ;
    wire new_AGEMA_signal_14887 ;
    wire new_AGEMA_signal_14888 ;
    wire new_AGEMA_signal_14889 ;
    wire new_AGEMA_signal_14890 ;
    wire new_AGEMA_signal_14891 ;
    wire new_AGEMA_signal_14892 ;
    wire new_AGEMA_signal_14893 ;
    wire new_AGEMA_signal_14894 ;
    wire new_AGEMA_signal_14895 ;
    wire new_AGEMA_signal_14896 ;
    wire new_AGEMA_signal_14897 ;
    wire new_AGEMA_signal_14898 ;
    wire new_AGEMA_signal_14899 ;
    wire new_AGEMA_signal_14900 ;
    wire new_AGEMA_signal_14901 ;
    wire new_AGEMA_signal_14902 ;
    wire new_AGEMA_signal_14903 ;
    wire new_AGEMA_signal_14904 ;
    wire new_AGEMA_signal_14905 ;
    wire new_AGEMA_signal_14906 ;
    wire new_AGEMA_signal_14907 ;
    wire new_AGEMA_signal_14908 ;
    wire new_AGEMA_signal_14909 ;
    wire new_AGEMA_signal_14910 ;
    wire new_AGEMA_signal_14911 ;
    wire new_AGEMA_signal_14912 ;
    wire new_AGEMA_signal_14913 ;
    wire new_AGEMA_signal_14914 ;
    wire new_AGEMA_signal_14915 ;
    wire new_AGEMA_signal_14916 ;
    wire new_AGEMA_signal_14917 ;
    wire new_AGEMA_signal_14918 ;
    wire new_AGEMA_signal_14919 ;
    wire new_AGEMA_signal_14920 ;
    wire new_AGEMA_signal_14921 ;
    wire new_AGEMA_signal_14922 ;
    wire new_AGEMA_signal_14923 ;
    wire new_AGEMA_signal_14924 ;
    wire new_AGEMA_signal_14925 ;
    wire new_AGEMA_signal_14926 ;
    wire new_AGEMA_signal_14927 ;
    wire new_AGEMA_signal_14928 ;
    wire new_AGEMA_signal_14929 ;
    wire new_AGEMA_signal_14930 ;
    wire new_AGEMA_signal_14931 ;
    wire new_AGEMA_signal_14932 ;
    wire new_AGEMA_signal_14933 ;
    wire new_AGEMA_signal_14934 ;
    wire new_AGEMA_signal_14935 ;
    wire new_AGEMA_signal_14936 ;
    wire new_AGEMA_signal_14937 ;
    wire new_AGEMA_signal_14938 ;
    wire new_AGEMA_signal_14939 ;
    wire new_AGEMA_signal_14940 ;
    wire new_AGEMA_signal_14941 ;
    wire new_AGEMA_signal_14942 ;
    wire new_AGEMA_signal_14943 ;
    wire new_AGEMA_signal_14944 ;
    wire new_AGEMA_signal_14945 ;
    wire new_AGEMA_signal_14946 ;
    wire new_AGEMA_signal_14947 ;
    wire new_AGEMA_signal_14948 ;
    wire new_AGEMA_signal_14949 ;
    wire new_AGEMA_signal_14950 ;
    wire new_AGEMA_signal_14951 ;
    wire new_AGEMA_signal_14952 ;
    wire new_AGEMA_signal_14953 ;
    wire new_AGEMA_signal_14954 ;
    wire new_AGEMA_signal_14955 ;
    wire new_AGEMA_signal_14956 ;
    wire new_AGEMA_signal_14957 ;
    wire new_AGEMA_signal_14958 ;
    wire new_AGEMA_signal_14959 ;
    wire new_AGEMA_signal_14960 ;
    wire new_AGEMA_signal_14961 ;
    wire new_AGEMA_signal_14962 ;
    wire new_AGEMA_signal_14963 ;
    wire new_AGEMA_signal_14964 ;
    wire new_AGEMA_signal_14965 ;
    wire new_AGEMA_signal_14966 ;
    wire new_AGEMA_signal_14967 ;
    wire new_AGEMA_signal_14968 ;
    wire new_AGEMA_signal_14969 ;
    wire new_AGEMA_signal_14970 ;
    wire new_AGEMA_signal_14971 ;
    wire new_AGEMA_signal_14972 ;
    wire new_AGEMA_signal_14973 ;
    wire new_AGEMA_signal_14974 ;
    wire new_AGEMA_signal_14975 ;
    wire new_AGEMA_signal_14976 ;
    wire new_AGEMA_signal_14977 ;
    wire new_AGEMA_signal_14978 ;
    wire new_AGEMA_signal_14979 ;
    wire new_AGEMA_signal_14980 ;
    wire new_AGEMA_signal_14981 ;
    wire new_AGEMA_signal_14982 ;
    wire new_AGEMA_signal_14983 ;
    wire new_AGEMA_signal_14984 ;
    wire new_AGEMA_signal_14985 ;
    wire new_AGEMA_signal_14986 ;
    wire new_AGEMA_signal_14987 ;
    wire new_AGEMA_signal_14988 ;
    wire new_AGEMA_signal_14989 ;
    wire new_AGEMA_signal_14990 ;
    wire new_AGEMA_signal_14991 ;
    wire new_AGEMA_signal_14992 ;
    wire new_AGEMA_signal_14993 ;
    wire new_AGEMA_signal_14994 ;
    wire new_AGEMA_signal_14995 ;
    wire new_AGEMA_signal_14996 ;
    wire new_AGEMA_signal_14997 ;
    wire new_AGEMA_signal_14998 ;
    wire new_AGEMA_signal_14999 ;
    wire new_AGEMA_signal_15000 ;
    wire new_AGEMA_signal_15001 ;
    wire new_AGEMA_signal_15002 ;
    wire new_AGEMA_signal_15003 ;
    wire new_AGEMA_signal_15004 ;
    wire new_AGEMA_signal_15005 ;
    wire new_AGEMA_signal_15006 ;
    wire new_AGEMA_signal_15007 ;
    wire new_AGEMA_signal_15008 ;
    wire new_AGEMA_signal_15009 ;
    wire new_AGEMA_signal_15010 ;
    wire new_AGEMA_signal_15011 ;
    wire new_AGEMA_signal_15012 ;
    wire new_AGEMA_signal_15013 ;
    wire new_AGEMA_signal_15014 ;
    wire new_AGEMA_signal_15015 ;
    wire new_AGEMA_signal_15016 ;
    wire new_AGEMA_signal_15017 ;
    wire new_AGEMA_signal_15018 ;
    wire new_AGEMA_signal_15019 ;
    wire new_AGEMA_signal_15020 ;
    wire new_AGEMA_signal_15021 ;
    wire new_AGEMA_signal_15022 ;
    wire new_AGEMA_signal_15023 ;
    wire new_AGEMA_signal_15024 ;
    wire new_AGEMA_signal_15025 ;
    wire new_AGEMA_signal_15026 ;
    wire new_AGEMA_signal_15027 ;
    wire new_AGEMA_signal_15028 ;
    wire new_AGEMA_signal_15029 ;
    wire new_AGEMA_signal_15030 ;
    wire new_AGEMA_signal_15031 ;
    wire new_AGEMA_signal_15032 ;
    wire new_AGEMA_signal_15033 ;
    wire new_AGEMA_signal_15034 ;
    wire new_AGEMA_signal_15035 ;
    wire new_AGEMA_signal_15036 ;
    wire new_AGEMA_signal_15037 ;
    wire new_AGEMA_signal_15038 ;
    wire new_AGEMA_signal_15039 ;
    wire new_AGEMA_signal_15040 ;
    wire new_AGEMA_signal_15041 ;
    wire new_AGEMA_signal_15042 ;
    wire new_AGEMA_signal_15043 ;
    wire new_AGEMA_signal_15044 ;
    wire new_AGEMA_signal_15045 ;
    wire new_AGEMA_signal_15046 ;
    wire new_AGEMA_signal_15047 ;
    wire new_AGEMA_signal_15048 ;
    wire new_AGEMA_signal_15049 ;
    wire new_AGEMA_signal_15050 ;
    wire new_AGEMA_signal_15051 ;
    wire new_AGEMA_signal_15052 ;
    wire new_AGEMA_signal_15053 ;
    wire new_AGEMA_signal_15054 ;
    wire new_AGEMA_signal_15055 ;
    wire new_AGEMA_signal_15056 ;
    wire new_AGEMA_signal_15057 ;
    wire new_AGEMA_signal_15058 ;
    wire new_AGEMA_signal_15059 ;
    wire new_AGEMA_signal_15060 ;
    wire new_AGEMA_signal_15061 ;
    wire new_AGEMA_signal_15062 ;
    wire new_AGEMA_signal_15063 ;
    wire new_AGEMA_signal_15064 ;
    wire new_AGEMA_signal_15065 ;
    wire new_AGEMA_signal_15066 ;
    wire new_AGEMA_signal_15067 ;
    wire new_AGEMA_signal_15068 ;
    wire new_AGEMA_signal_15069 ;
    wire new_AGEMA_signal_15070 ;
    wire new_AGEMA_signal_15071 ;
    wire new_AGEMA_signal_15072 ;
    wire new_AGEMA_signal_15073 ;
    wire new_AGEMA_signal_15074 ;
    wire new_AGEMA_signal_15075 ;
    wire new_AGEMA_signal_15076 ;
    wire new_AGEMA_signal_15077 ;
    wire new_AGEMA_signal_15078 ;
    wire new_AGEMA_signal_15079 ;
    wire new_AGEMA_signal_15080 ;
    wire new_AGEMA_signal_15081 ;
    wire new_AGEMA_signal_15082 ;
    wire new_AGEMA_signal_15083 ;
    wire new_AGEMA_signal_15084 ;
    wire new_AGEMA_signal_15085 ;
    wire new_AGEMA_signal_15086 ;
    wire new_AGEMA_signal_15087 ;
    wire new_AGEMA_signal_15088 ;
    wire new_AGEMA_signal_15089 ;
    wire new_AGEMA_signal_15090 ;
    wire new_AGEMA_signal_15091 ;
    wire new_AGEMA_signal_15092 ;
    wire new_AGEMA_signal_15093 ;
    wire new_AGEMA_signal_15094 ;
    wire new_AGEMA_signal_15095 ;
    wire new_AGEMA_signal_15096 ;
    wire new_AGEMA_signal_15097 ;
    wire new_AGEMA_signal_15098 ;
    wire new_AGEMA_signal_15099 ;
    wire new_AGEMA_signal_15100 ;
    wire new_AGEMA_signal_15101 ;
    wire new_AGEMA_signal_15102 ;
    wire new_AGEMA_signal_15103 ;
    wire new_AGEMA_signal_15104 ;
    wire new_AGEMA_signal_15105 ;
    wire new_AGEMA_signal_15106 ;
    wire new_AGEMA_signal_15107 ;
    wire new_AGEMA_signal_15108 ;
    wire new_AGEMA_signal_15109 ;
    wire new_AGEMA_signal_15110 ;
    wire new_AGEMA_signal_15111 ;
    wire new_AGEMA_signal_15112 ;
    wire new_AGEMA_signal_15113 ;
    wire new_AGEMA_signal_15114 ;
    wire new_AGEMA_signal_15115 ;
    wire new_AGEMA_signal_15116 ;
    wire new_AGEMA_signal_15117 ;
    wire new_AGEMA_signal_15118 ;
    wire new_AGEMA_signal_15119 ;
    wire new_AGEMA_signal_15120 ;
    wire new_AGEMA_signal_15121 ;
    wire new_AGEMA_signal_15122 ;
    wire new_AGEMA_signal_15123 ;
    wire new_AGEMA_signal_15124 ;
    wire new_AGEMA_signal_15125 ;
    wire new_AGEMA_signal_15126 ;
    wire new_AGEMA_signal_15127 ;
    wire new_AGEMA_signal_15128 ;
    wire new_AGEMA_signal_15129 ;
    wire new_AGEMA_signal_15130 ;
    wire new_AGEMA_signal_15131 ;
    wire new_AGEMA_signal_15132 ;
    wire new_AGEMA_signal_15133 ;
    wire new_AGEMA_signal_15134 ;
    wire new_AGEMA_signal_15135 ;
    wire new_AGEMA_signal_15136 ;
    wire new_AGEMA_signal_15137 ;
    wire new_AGEMA_signal_15138 ;
    wire new_AGEMA_signal_15139 ;
    wire new_AGEMA_signal_15140 ;
    wire new_AGEMA_signal_15141 ;
    wire new_AGEMA_signal_15142 ;
    wire new_AGEMA_signal_15143 ;
    wire new_AGEMA_signal_15144 ;
    wire new_AGEMA_signal_15145 ;
    wire new_AGEMA_signal_15146 ;
    wire new_AGEMA_signal_15147 ;
    wire new_AGEMA_signal_15148 ;
    wire new_AGEMA_signal_15149 ;
    wire new_AGEMA_signal_15150 ;
    wire new_AGEMA_signal_15151 ;
    wire new_AGEMA_signal_15152 ;
    wire new_AGEMA_signal_15153 ;
    wire new_AGEMA_signal_15154 ;
    wire new_AGEMA_signal_15155 ;
    wire new_AGEMA_signal_15156 ;
    wire new_AGEMA_signal_15157 ;
    wire new_AGEMA_signal_15158 ;
    wire new_AGEMA_signal_15159 ;
    wire new_AGEMA_signal_15160 ;
    wire new_AGEMA_signal_15161 ;
    wire new_AGEMA_signal_15162 ;
    wire new_AGEMA_signal_15163 ;
    wire new_AGEMA_signal_15164 ;
    wire new_AGEMA_signal_15165 ;
    wire new_AGEMA_signal_15166 ;
    wire new_AGEMA_signal_15167 ;
    wire new_AGEMA_signal_15168 ;
    wire new_AGEMA_signal_15169 ;
    wire new_AGEMA_signal_15170 ;
    wire new_AGEMA_signal_15171 ;
    wire new_AGEMA_signal_15172 ;
    wire new_AGEMA_signal_15173 ;
    wire new_AGEMA_signal_15174 ;
    wire new_AGEMA_signal_15175 ;
    wire new_AGEMA_signal_15176 ;
    wire new_AGEMA_signal_15177 ;
    wire new_AGEMA_signal_15178 ;
    wire new_AGEMA_signal_15179 ;
    wire new_AGEMA_signal_15180 ;
    wire new_AGEMA_signal_15181 ;
    wire new_AGEMA_signal_15182 ;
    wire new_AGEMA_signal_15183 ;
    wire new_AGEMA_signal_15184 ;
    wire new_AGEMA_signal_15185 ;
    wire new_AGEMA_signal_15186 ;
    wire new_AGEMA_signal_15187 ;
    wire new_AGEMA_signal_15188 ;
    wire new_AGEMA_signal_15189 ;
    wire new_AGEMA_signal_15190 ;
    wire new_AGEMA_signal_15191 ;
    wire new_AGEMA_signal_15192 ;
    wire new_AGEMA_signal_15193 ;
    wire new_AGEMA_signal_15194 ;
    wire new_AGEMA_signal_15195 ;
    wire new_AGEMA_signal_15196 ;
    wire new_AGEMA_signal_15197 ;
    wire new_AGEMA_signal_15198 ;
    wire new_AGEMA_signal_15199 ;
    wire new_AGEMA_signal_15200 ;
    wire new_AGEMA_signal_15201 ;
    wire new_AGEMA_signal_15202 ;
    wire new_AGEMA_signal_15203 ;
    wire new_AGEMA_signal_15204 ;
    wire new_AGEMA_signal_15205 ;
    wire new_AGEMA_signal_15206 ;
    wire new_AGEMA_signal_15207 ;
    wire new_AGEMA_signal_15208 ;
    wire new_AGEMA_signal_15209 ;
    wire new_AGEMA_signal_15210 ;
    wire new_AGEMA_signal_15211 ;
    wire new_AGEMA_signal_15212 ;
    wire new_AGEMA_signal_15213 ;
    wire new_AGEMA_signal_15214 ;
    wire new_AGEMA_signal_15215 ;
    wire new_AGEMA_signal_15216 ;
    wire new_AGEMA_signal_15217 ;
    wire new_AGEMA_signal_15218 ;
    wire new_AGEMA_signal_15219 ;
    wire new_AGEMA_signal_15220 ;
    wire new_AGEMA_signal_15221 ;
    wire new_AGEMA_signal_15222 ;
    wire new_AGEMA_signal_15223 ;
    wire new_AGEMA_signal_15224 ;
    wire new_AGEMA_signal_15225 ;
    wire new_AGEMA_signal_15226 ;
    wire new_AGEMA_signal_15227 ;
    wire new_AGEMA_signal_15228 ;
    wire new_AGEMA_signal_15229 ;
    wire new_AGEMA_signal_15230 ;
    wire new_AGEMA_signal_15231 ;
    wire new_AGEMA_signal_15232 ;
    wire new_AGEMA_signal_15233 ;
    wire new_AGEMA_signal_15234 ;
    wire new_AGEMA_signal_15235 ;
    wire new_AGEMA_signal_15236 ;
    wire new_AGEMA_signal_15237 ;
    wire new_AGEMA_signal_15238 ;
    wire new_AGEMA_signal_15239 ;
    wire new_AGEMA_signal_15240 ;
    wire new_AGEMA_signal_15241 ;
    wire new_AGEMA_signal_15242 ;
    wire new_AGEMA_signal_15243 ;
    wire new_AGEMA_signal_15244 ;
    wire new_AGEMA_signal_15245 ;
    wire new_AGEMA_signal_15246 ;
    wire new_AGEMA_signal_15247 ;
    wire new_AGEMA_signal_15248 ;
    wire new_AGEMA_signal_15249 ;
    wire new_AGEMA_signal_15250 ;
    wire new_AGEMA_signal_15251 ;
    wire new_AGEMA_signal_15252 ;
    wire new_AGEMA_signal_15253 ;
    wire new_AGEMA_signal_15254 ;
    wire new_AGEMA_signal_15255 ;
    wire new_AGEMA_signal_15256 ;
    wire new_AGEMA_signal_15257 ;
    wire new_AGEMA_signal_15258 ;
    wire new_AGEMA_signal_15259 ;
    wire new_AGEMA_signal_15260 ;
    wire new_AGEMA_signal_15261 ;
    wire new_AGEMA_signal_15262 ;
    wire new_AGEMA_signal_15263 ;
    wire new_AGEMA_signal_15264 ;
    wire new_AGEMA_signal_15265 ;
    wire new_AGEMA_signal_15266 ;
    wire new_AGEMA_signal_15267 ;
    wire new_AGEMA_signal_15268 ;
    wire new_AGEMA_signal_15269 ;
    wire new_AGEMA_signal_15270 ;
    wire new_AGEMA_signal_15271 ;
    wire new_AGEMA_signal_15272 ;
    wire new_AGEMA_signal_15273 ;
    wire new_AGEMA_signal_15274 ;
    wire new_AGEMA_signal_15275 ;
    wire new_AGEMA_signal_15276 ;
    wire new_AGEMA_signal_15277 ;
    wire new_AGEMA_signal_15278 ;
    wire new_AGEMA_signal_15279 ;
    wire new_AGEMA_signal_15280 ;
    wire new_AGEMA_signal_15281 ;
    wire new_AGEMA_signal_15282 ;
    wire new_AGEMA_signal_15283 ;
    wire new_AGEMA_signal_15284 ;
    wire new_AGEMA_signal_15285 ;
    wire new_AGEMA_signal_15286 ;
    wire new_AGEMA_signal_15287 ;
    wire new_AGEMA_signal_15288 ;
    wire new_AGEMA_signal_15289 ;
    wire new_AGEMA_signal_15290 ;
    wire new_AGEMA_signal_15291 ;
    wire new_AGEMA_signal_15292 ;
    wire new_AGEMA_signal_15293 ;
    wire new_AGEMA_signal_15294 ;
    wire new_AGEMA_signal_15295 ;
    wire new_AGEMA_signal_15296 ;
    wire new_AGEMA_signal_15297 ;
    wire new_AGEMA_signal_15298 ;
    wire new_AGEMA_signal_15299 ;
    wire new_AGEMA_signal_15300 ;
    wire new_AGEMA_signal_15301 ;
    wire new_AGEMA_signal_15302 ;
    wire new_AGEMA_signal_15303 ;
    wire new_AGEMA_signal_15304 ;
    wire new_AGEMA_signal_15305 ;
    wire new_AGEMA_signal_15306 ;
    wire new_AGEMA_signal_15307 ;
    wire new_AGEMA_signal_15308 ;
    wire new_AGEMA_signal_15309 ;
    wire new_AGEMA_signal_15310 ;
    wire new_AGEMA_signal_15311 ;
    wire new_AGEMA_signal_15312 ;
    wire new_AGEMA_signal_15313 ;
    wire new_AGEMA_signal_15314 ;
    wire new_AGEMA_signal_15315 ;
    wire new_AGEMA_signal_15316 ;
    wire new_AGEMA_signal_15317 ;
    wire new_AGEMA_signal_15318 ;
    wire new_AGEMA_signal_15319 ;
    wire new_AGEMA_signal_15320 ;
    wire new_AGEMA_signal_15321 ;
    wire new_AGEMA_signal_15322 ;
    wire new_AGEMA_signal_15323 ;
    wire new_AGEMA_signal_15324 ;
    wire new_AGEMA_signal_15325 ;
    wire new_AGEMA_signal_15326 ;
    wire new_AGEMA_signal_15327 ;
    wire new_AGEMA_signal_15328 ;
    wire new_AGEMA_signal_15329 ;
    wire new_AGEMA_signal_15330 ;
    wire new_AGEMA_signal_15331 ;
    wire new_AGEMA_signal_15332 ;
    wire new_AGEMA_signal_15333 ;
    wire new_AGEMA_signal_15334 ;
    wire new_AGEMA_signal_15335 ;
    wire new_AGEMA_signal_15336 ;
    wire new_AGEMA_signal_15337 ;
    wire new_AGEMA_signal_15338 ;
    wire new_AGEMA_signal_15339 ;
    wire new_AGEMA_signal_15340 ;
    wire new_AGEMA_signal_15341 ;
    wire new_AGEMA_signal_15342 ;
    wire new_AGEMA_signal_15343 ;
    wire new_AGEMA_signal_15344 ;
    wire new_AGEMA_signal_15345 ;
    wire new_AGEMA_signal_15346 ;
    wire new_AGEMA_signal_15347 ;
    wire new_AGEMA_signal_15348 ;
    wire new_AGEMA_signal_15349 ;
    wire new_AGEMA_signal_15350 ;
    wire new_AGEMA_signal_15351 ;
    wire new_AGEMA_signal_15352 ;
    wire new_AGEMA_signal_15353 ;
    wire new_AGEMA_signal_15354 ;
    wire new_AGEMA_signal_15355 ;
    wire new_AGEMA_signal_15356 ;
    wire new_AGEMA_signal_15357 ;
    wire new_AGEMA_signal_15358 ;
    wire new_AGEMA_signal_15359 ;
    wire new_AGEMA_signal_15360 ;
    wire new_AGEMA_signal_15361 ;
    wire new_AGEMA_signal_15362 ;
    wire new_AGEMA_signal_15363 ;
    wire new_AGEMA_signal_15364 ;
    wire new_AGEMA_signal_15365 ;
    wire new_AGEMA_signal_15366 ;
    wire new_AGEMA_signal_15367 ;
    wire new_AGEMA_signal_15368 ;
    wire new_AGEMA_signal_15369 ;
    wire new_AGEMA_signal_15370 ;
    wire new_AGEMA_signal_15371 ;
    wire new_AGEMA_signal_15372 ;
    wire new_AGEMA_signal_15373 ;
    wire new_AGEMA_signal_15374 ;
    wire new_AGEMA_signal_15375 ;
    wire new_AGEMA_signal_15376 ;
    wire new_AGEMA_signal_15377 ;
    wire new_AGEMA_signal_15378 ;
    wire new_AGEMA_signal_15379 ;
    wire new_AGEMA_signal_15380 ;
    wire new_AGEMA_signal_15381 ;
    wire new_AGEMA_signal_15382 ;
    wire new_AGEMA_signal_15383 ;
    wire new_AGEMA_signal_15384 ;
    wire new_AGEMA_signal_15385 ;
    wire new_AGEMA_signal_15386 ;
    wire new_AGEMA_signal_15387 ;
    wire new_AGEMA_signal_15388 ;
    wire new_AGEMA_signal_15389 ;
    wire new_AGEMA_signal_15390 ;
    wire new_AGEMA_signal_15391 ;
    wire new_AGEMA_signal_15392 ;
    wire new_AGEMA_signal_15393 ;
    wire new_AGEMA_signal_15394 ;
    wire new_AGEMA_signal_15395 ;
    wire new_AGEMA_signal_15396 ;
    wire new_AGEMA_signal_15397 ;
    wire new_AGEMA_signal_15398 ;
    wire new_AGEMA_signal_15399 ;
    wire new_AGEMA_signal_15400 ;
    wire new_AGEMA_signal_15401 ;
    wire new_AGEMA_signal_15402 ;
    wire new_AGEMA_signal_15403 ;
    wire new_AGEMA_signal_15404 ;
    wire new_AGEMA_signal_15405 ;
    wire new_AGEMA_signal_15406 ;
    wire new_AGEMA_signal_15407 ;
    wire new_AGEMA_signal_15408 ;
    wire new_AGEMA_signal_15409 ;
    wire new_AGEMA_signal_15410 ;
    wire new_AGEMA_signal_15411 ;
    wire new_AGEMA_signal_15412 ;
    wire new_AGEMA_signal_15413 ;
    wire new_AGEMA_signal_15414 ;
    wire new_AGEMA_signal_15415 ;
    wire new_AGEMA_signal_15416 ;
    wire new_AGEMA_signal_15417 ;
    wire new_AGEMA_signal_15418 ;
    wire new_AGEMA_signal_15419 ;
    wire new_AGEMA_signal_15420 ;
    wire new_AGEMA_signal_15421 ;
    wire new_AGEMA_signal_15422 ;
    wire new_AGEMA_signal_15423 ;
    wire new_AGEMA_signal_15424 ;
    wire new_AGEMA_signal_15425 ;
    wire new_AGEMA_signal_15426 ;
    wire new_AGEMA_signal_15427 ;
    wire new_AGEMA_signal_15428 ;
    wire new_AGEMA_signal_15429 ;
    wire new_AGEMA_signal_15430 ;
    wire new_AGEMA_signal_15431 ;
    wire new_AGEMA_signal_15432 ;
    wire new_AGEMA_signal_15433 ;
    wire new_AGEMA_signal_15434 ;
    wire new_AGEMA_signal_15435 ;
    wire new_AGEMA_signal_15436 ;
    wire new_AGEMA_signal_15437 ;
    wire new_AGEMA_signal_15438 ;
    wire new_AGEMA_signal_15439 ;
    wire new_AGEMA_signal_15440 ;
    wire new_AGEMA_signal_15441 ;
    wire new_AGEMA_signal_15442 ;
    wire new_AGEMA_signal_15443 ;
    wire new_AGEMA_signal_15444 ;
    wire new_AGEMA_signal_15445 ;
    wire new_AGEMA_signal_15446 ;
    wire new_AGEMA_signal_15447 ;
    wire new_AGEMA_signal_15448 ;
    wire new_AGEMA_signal_15449 ;
    wire new_AGEMA_signal_15450 ;
    wire new_AGEMA_signal_15451 ;
    wire new_AGEMA_signal_15452 ;
    wire new_AGEMA_signal_15453 ;
    wire new_AGEMA_signal_15454 ;
    wire new_AGEMA_signal_15455 ;
    wire new_AGEMA_signal_15456 ;
    wire new_AGEMA_signal_15457 ;
    wire new_AGEMA_signal_15458 ;
    wire new_AGEMA_signal_15459 ;
    wire new_AGEMA_signal_15460 ;
    wire new_AGEMA_signal_15461 ;
    wire new_AGEMA_signal_15462 ;
    wire new_AGEMA_signal_15463 ;
    wire new_AGEMA_signal_15464 ;
    wire new_AGEMA_signal_15465 ;
    wire new_AGEMA_signal_15466 ;
    wire new_AGEMA_signal_15467 ;
    wire new_AGEMA_signal_15468 ;
    wire new_AGEMA_signal_15469 ;
    wire new_AGEMA_signal_15470 ;
    wire new_AGEMA_signal_15471 ;
    wire new_AGEMA_signal_15472 ;
    wire new_AGEMA_signal_15473 ;
    wire new_AGEMA_signal_15474 ;
    wire new_AGEMA_signal_15475 ;
    wire new_AGEMA_signal_15476 ;
    wire new_AGEMA_signal_15477 ;
    wire new_AGEMA_signal_15478 ;
    wire new_AGEMA_signal_15479 ;
    wire new_AGEMA_signal_15480 ;
    wire new_AGEMA_signal_15481 ;
    wire new_AGEMA_signal_15482 ;
    wire new_AGEMA_signal_15483 ;
    wire new_AGEMA_signal_15484 ;
    wire new_AGEMA_signal_15485 ;
    wire new_AGEMA_signal_15486 ;
    wire new_AGEMA_signal_15487 ;
    wire new_AGEMA_signal_15488 ;
    wire new_AGEMA_signal_15489 ;
    wire new_AGEMA_signal_15490 ;
    wire new_AGEMA_signal_15491 ;
    wire new_AGEMA_signal_15492 ;
    wire new_AGEMA_signal_15493 ;
    wire new_AGEMA_signal_15494 ;
    wire new_AGEMA_signal_15495 ;
    wire new_AGEMA_signal_15496 ;
    wire new_AGEMA_signal_15497 ;
    wire new_AGEMA_signal_15498 ;
    wire new_AGEMA_signal_15499 ;
    wire new_AGEMA_signal_15500 ;
    wire new_AGEMA_signal_15501 ;
    wire new_AGEMA_signal_15502 ;
    wire new_AGEMA_signal_15503 ;
    wire new_AGEMA_signal_15504 ;
    wire new_AGEMA_signal_15505 ;
    wire new_AGEMA_signal_15506 ;
    wire new_AGEMA_signal_15507 ;
    wire new_AGEMA_signal_15508 ;
    wire new_AGEMA_signal_15509 ;
    wire new_AGEMA_signal_15510 ;
    wire new_AGEMA_signal_15511 ;
    wire new_AGEMA_signal_15512 ;
    wire new_AGEMA_signal_15513 ;
    wire new_AGEMA_signal_15514 ;
    wire new_AGEMA_signal_15515 ;
    wire new_AGEMA_signal_15516 ;
    wire new_AGEMA_signal_15517 ;
    wire new_AGEMA_signal_15518 ;
    wire new_AGEMA_signal_15519 ;
    wire new_AGEMA_signal_15520 ;
    wire new_AGEMA_signal_15521 ;
    wire new_AGEMA_signal_15522 ;
    wire new_AGEMA_signal_15523 ;
    wire new_AGEMA_signal_15524 ;
    wire new_AGEMA_signal_15525 ;
    wire new_AGEMA_signal_15526 ;
    wire new_AGEMA_signal_15527 ;
    wire new_AGEMA_signal_15528 ;
    wire new_AGEMA_signal_15529 ;
    wire new_AGEMA_signal_15530 ;
    wire new_AGEMA_signal_15531 ;
    wire new_AGEMA_signal_15532 ;
    wire new_AGEMA_signal_15533 ;
    wire new_AGEMA_signal_15534 ;
    wire new_AGEMA_signal_15535 ;
    wire new_AGEMA_signal_15536 ;
    wire new_AGEMA_signal_15537 ;
    wire new_AGEMA_signal_15538 ;
    wire new_AGEMA_signal_15539 ;
    wire new_AGEMA_signal_15540 ;
    wire new_AGEMA_signal_15541 ;
    wire new_AGEMA_signal_15542 ;
    wire new_AGEMA_signal_15543 ;
    wire new_AGEMA_signal_15544 ;
    wire new_AGEMA_signal_15545 ;
    wire new_AGEMA_signal_15546 ;
    wire new_AGEMA_signal_15547 ;
    wire new_AGEMA_signal_15548 ;
    wire new_AGEMA_signal_15549 ;
    wire new_AGEMA_signal_15550 ;
    wire new_AGEMA_signal_15551 ;
    wire new_AGEMA_signal_15552 ;
    wire new_AGEMA_signal_15553 ;
    wire new_AGEMA_signal_15554 ;
    wire new_AGEMA_signal_15555 ;
    wire new_AGEMA_signal_15556 ;
    wire new_AGEMA_signal_15557 ;
    wire new_AGEMA_signal_15558 ;
    wire new_AGEMA_signal_15559 ;
    wire new_AGEMA_signal_15560 ;
    wire new_AGEMA_signal_15561 ;
    wire new_AGEMA_signal_15562 ;
    wire new_AGEMA_signal_15563 ;
    wire new_AGEMA_signal_15564 ;
    wire new_AGEMA_signal_15565 ;
    wire new_AGEMA_signal_15566 ;
    wire new_AGEMA_signal_15567 ;
    wire new_AGEMA_signal_15568 ;
    wire new_AGEMA_signal_15569 ;
    wire new_AGEMA_signal_15570 ;
    wire new_AGEMA_signal_15571 ;
    wire new_AGEMA_signal_15572 ;
    wire new_AGEMA_signal_15573 ;
    wire new_AGEMA_signal_15574 ;
    wire new_AGEMA_signal_15575 ;
    wire new_AGEMA_signal_15576 ;
    wire new_AGEMA_signal_15577 ;
    wire new_AGEMA_signal_15578 ;
    wire new_AGEMA_signal_15579 ;
    wire new_AGEMA_signal_15580 ;
    wire new_AGEMA_signal_15581 ;
    wire new_AGEMA_signal_15582 ;
    wire new_AGEMA_signal_15583 ;
    wire new_AGEMA_signal_15584 ;
    wire new_AGEMA_signal_15585 ;
    wire new_AGEMA_signal_15586 ;
    wire new_AGEMA_signal_15587 ;
    wire new_AGEMA_signal_15588 ;
    wire new_AGEMA_signal_15589 ;
    wire new_AGEMA_signal_15590 ;
    wire new_AGEMA_signal_15591 ;
    wire new_AGEMA_signal_15592 ;
    wire new_AGEMA_signal_15593 ;
    wire new_AGEMA_signal_15594 ;
    wire new_AGEMA_signal_15595 ;
    wire new_AGEMA_signal_15596 ;
    wire new_AGEMA_signal_15597 ;
    wire new_AGEMA_signal_15598 ;
    wire new_AGEMA_signal_15599 ;
    wire new_AGEMA_signal_15600 ;
    wire new_AGEMA_signal_15601 ;
    wire new_AGEMA_signal_15602 ;
    wire new_AGEMA_signal_15603 ;
    wire new_AGEMA_signal_15604 ;
    wire new_AGEMA_signal_15605 ;
    wire new_AGEMA_signal_15606 ;
    wire new_AGEMA_signal_15607 ;
    wire new_AGEMA_signal_15608 ;
    wire new_AGEMA_signal_15609 ;
    wire new_AGEMA_signal_15610 ;
    wire new_AGEMA_signal_15611 ;
    wire new_AGEMA_signal_15612 ;
    wire new_AGEMA_signal_15613 ;
    wire new_AGEMA_signal_15614 ;
    wire new_AGEMA_signal_15615 ;
    wire new_AGEMA_signal_15616 ;
    wire new_AGEMA_signal_15617 ;
    wire new_AGEMA_signal_15618 ;
    wire new_AGEMA_signal_15619 ;
    wire new_AGEMA_signal_15620 ;
    wire new_AGEMA_signal_15621 ;
    wire new_AGEMA_signal_15622 ;
    wire new_AGEMA_signal_15623 ;
    wire new_AGEMA_signal_15624 ;
    wire new_AGEMA_signal_15625 ;
    wire new_AGEMA_signal_15626 ;
    wire new_AGEMA_signal_15627 ;
    wire new_AGEMA_signal_15628 ;
    wire new_AGEMA_signal_15629 ;
    wire new_AGEMA_signal_15630 ;
    wire new_AGEMA_signal_15631 ;
    wire new_AGEMA_signal_15632 ;
    wire new_AGEMA_signal_15633 ;
    wire new_AGEMA_signal_15634 ;
    wire new_AGEMA_signal_15635 ;
    wire new_AGEMA_signal_15636 ;
    wire new_AGEMA_signal_15637 ;
    wire new_AGEMA_signal_15638 ;
    wire new_AGEMA_signal_15639 ;
    wire new_AGEMA_signal_15640 ;
    wire new_AGEMA_signal_15641 ;
    wire new_AGEMA_signal_15642 ;
    wire new_AGEMA_signal_15643 ;
    wire new_AGEMA_signal_15644 ;
    wire new_AGEMA_signal_15645 ;
    wire new_AGEMA_signal_15646 ;
    wire new_AGEMA_signal_15647 ;
    wire new_AGEMA_signal_15648 ;
    wire new_AGEMA_signal_15649 ;
    wire new_AGEMA_signal_15650 ;
    wire new_AGEMA_signal_15651 ;
    wire new_AGEMA_signal_15652 ;
    wire new_AGEMA_signal_15653 ;
    wire new_AGEMA_signal_15654 ;
    wire new_AGEMA_signal_15655 ;
    wire new_AGEMA_signal_15656 ;
    wire new_AGEMA_signal_15657 ;
    wire new_AGEMA_signal_15658 ;
    wire new_AGEMA_signal_15659 ;
    wire new_AGEMA_signal_15660 ;
    wire new_AGEMA_signal_15661 ;
    wire new_AGEMA_signal_15662 ;
    wire new_AGEMA_signal_15663 ;
    wire new_AGEMA_signal_15664 ;
    wire new_AGEMA_signal_15665 ;
    wire new_AGEMA_signal_15666 ;
    wire new_AGEMA_signal_15667 ;
    wire new_AGEMA_signal_15668 ;
    wire new_AGEMA_signal_15669 ;
    wire new_AGEMA_signal_15670 ;
    wire new_AGEMA_signal_15671 ;
    wire new_AGEMA_signal_15672 ;
    wire new_AGEMA_signal_15673 ;
    wire new_AGEMA_signal_15674 ;
    wire new_AGEMA_signal_15675 ;
    wire new_AGEMA_signal_15676 ;
    wire new_AGEMA_signal_15677 ;
    wire new_AGEMA_signal_15678 ;
    wire new_AGEMA_signal_15679 ;
    wire new_AGEMA_signal_15680 ;
    wire new_AGEMA_signal_15681 ;
    wire new_AGEMA_signal_15682 ;
    wire new_AGEMA_signal_15683 ;
    wire new_AGEMA_signal_15684 ;
    wire new_AGEMA_signal_15685 ;
    wire new_AGEMA_signal_15686 ;
    wire new_AGEMA_signal_15687 ;
    wire new_AGEMA_signal_15688 ;
    wire new_AGEMA_signal_15689 ;
    wire new_AGEMA_signal_15690 ;
    wire new_AGEMA_signal_15691 ;
    wire new_AGEMA_signal_15692 ;
    wire new_AGEMA_signal_15693 ;
    wire new_AGEMA_signal_15694 ;
    wire new_AGEMA_signal_15695 ;
    wire new_AGEMA_signal_15696 ;
    wire new_AGEMA_signal_15697 ;
    wire new_AGEMA_signal_15698 ;
    wire new_AGEMA_signal_15699 ;
    wire new_AGEMA_signal_15700 ;
    wire new_AGEMA_signal_15701 ;
    wire new_AGEMA_signal_15702 ;
    wire new_AGEMA_signal_15703 ;
    wire new_AGEMA_signal_15704 ;
    wire new_AGEMA_signal_15705 ;
    wire new_AGEMA_signal_15706 ;
    wire new_AGEMA_signal_15707 ;
    wire new_AGEMA_signal_15708 ;
    wire new_AGEMA_signal_15709 ;
    wire new_AGEMA_signal_15710 ;
    wire new_AGEMA_signal_15711 ;
    wire new_AGEMA_signal_15712 ;
    wire new_AGEMA_signal_15713 ;
    wire new_AGEMA_signal_15714 ;
    wire new_AGEMA_signal_15715 ;
    wire new_AGEMA_signal_15716 ;
    wire new_AGEMA_signal_15717 ;
    wire new_AGEMA_signal_15718 ;
    wire new_AGEMA_signal_15719 ;
    wire new_AGEMA_signal_15720 ;
    wire new_AGEMA_signal_15721 ;
    wire new_AGEMA_signal_15722 ;
    wire new_AGEMA_signal_15723 ;
    wire new_AGEMA_signal_15724 ;
    wire new_AGEMA_signal_15725 ;
    wire new_AGEMA_signal_15726 ;
    wire new_AGEMA_signal_15727 ;
    wire new_AGEMA_signal_15728 ;
    wire new_AGEMA_signal_15729 ;
    wire new_AGEMA_signal_15730 ;
    wire new_AGEMA_signal_15731 ;
    wire new_AGEMA_signal_15732 ;
    wire new_AGEMA_signal_15733 ;
    wire new_AGEMA_signal_15734 ;
    wire new_AGEMA_signal_15735 ;
    wire new_AGEMA_signal_15736 ;
    wire new_AGEMA_signal_15737 ;
    wire new_AGEMA_signal_15738 ;
    wire new_AGEMA_signal_15739 ;
    wire new_AGEMA_signal_15740 ;
    wire new_AGEMA_signal_15741 ;
    wire new_AGEMA_signal_15742 ;
    wire new_AGEMA_signal_15743 ;
    wire new_AGEMA_signal_15744 ;
    wire new_AGEMA_signal_15745 ;
    wire new_AGEMA_signal_15746 ;
    wire new_AGEMA_signal_15747 ;
    wire new_AGEMA_signal_15748 ;
    wire new_AGEMA_signal_15749 ;
    wire new_AGEMA_signal_15750 ;
    wire new_AGEMA_signal_15751 ;
    wire new_AGEMA_signal_15752 ;
    wire new_AGEMA_signal_15753 ;
    wire new_AGEMA_signal_15754 ;
    wire new_AGEMA_signal_15755 ;
    wire new_AGEMA_signal_15756 ;
    wire new_AGEMA_signal_15757 ;
    wire new_AGEMA_signal_15758 ;
    wire new_AGEMA_signal_15759 ;
    wire new_AGEMA_signal_15760 ;
    wire new_AGEMA_signal_15761 ;
    wire new_AGEMA_signal_15762 ;
    wire new_AGEMA_signal_15763 ;
    wire new_AGEMA_signal_15764 ;
    wire new_AGEMA_signal_15765 ;
    wire new_AGEMA_signal_15766 ;
    wire new_AGEMA_signal_15767 ;
    wire new_AGEMA_signal_15768 ;
    wire new_AGEMA_signal_15769 ;
    wire new_AGEMA_signal_15770 ;
    wire new_AGEMA_signal_15771 ;
    wire new_AGEMA_signal_15772 ;
    wire new_AGEMA_signal_15773 ;
    wire new_AGEMA_signal_15774 ;
    wire new_AGEMA_signal_15775 ;
    wire new_AGEMA_signal_15776 ;
    wire new_AGEMA_signal_15777 ;
    wire new_AGEMA_signal_15778 ;
    wire new_AGEMA_signal_15779 ;
    wire new_AGEMA_signal_15780 ;
    wire new_AGEMA_signal_15781 ;
    wire new_AGEMA_signal_15782 ;
    wire new_AGEMA_signal_15783 ;
    wire new_AGEMA_signal_15784 ;
    wire new_AGEMA_signal_15785 ;
    wire new_AGEMA_signal_15786 ;
    wire new_AGEMA_signal_15787 ;
    wire new_AGEMA_signal_15788 ;
    wire new_AGEMA_signal_15789 ;
    wire new_AGEMA_signal_15790 ;
    wire new_AGEMA_signal_15791 ;
    wire new_AGEMA_signal_15792 ;
    wire new_AGEMA_signal_15793 ;
    wire new_AGEMA_signal_15794 ;
    wire new_AGEMA_signal_15795 ;
    wire new_AGEMA_signal_15796 ;
    wire new_AGEMA_signal_15797 ;
    wire new_AGEMA_signal_15798 ;
    wire new_AGEMA_signal_15799 ;
    wire new_AGEMA_signal_15800 ;
    wire new_AGEMA_signal_15801 ;
    wire new_AGEMA_signal_15802 ;
    wire new_AGEMA_signal_15803 ;
    wire new_AGEMA_signal_15804 ;
    wire new_AGEMA_signal_15805 ;
    wire new_AGEMA_signal_15806 ;
    wire new_AGEMA_signal_15807 ;
    wire new_AGEMA_signal_15808 ;
    wire new_AGEMA_signal_15809 ;
    wire new_AGEMA_signal_15810 ;
    wire new_AGEMA_signal_15811 ;
    wire new_AGEMA_signal_15812 ;
    wire new_AGEMA_signal_15813 ;
    wire new_AGEMA_signal_15814 ;
    wire new_AGEMA_signal_15815 ;
    wire new_AGEMA_signal_15816 ;
    wire new_AGEMA_signal_15817 ;
    wire new_AGEMA_signal_15818 ;
    wire new_AGEMA_signal_15819 ;
    wire new_AGEMA_signal_15820 ;
    wire new_AGEMA_signal_15821 ;
    wire new_AGEMA_signal_15822 ;
    wire new_AGEMA_signal_15823 ;
    wire new_AGEMA_signal_15824 ;
    wire new_AGEMA_signal_15825 ;
    wire new_AGEMA_signal_15826 ;
    wire new_AGEMA_signal_15827 ;
    wire new_AGEMA_signal_15828 ;
    wire new_AGEMA_signal_15829 ;
    wire new_AGEMA_signal_15830 ;
    wire new_AGEMA_signal_15831 ;
    wire new_AGEMA_signal_15832 ;
    wire new_AGEMA_signal_15833 ;
    wire new_AGEMA_signal_15834 ;
    wire new_AGEMA_signal_15835 ;
    wire new_AGEMA_signal_15836 ;
    wire new_AGEMA_signal_15837 ;
    wire new_AGEMA_signal_15838 ;
    wire new_AGEMA_signal_15839 ;
    wire new_AGEMA_signal_15840 ;
    wire new_AGEMA_signal_15841 ;
    wire new_AGEMA_signal_15842 ;
    wire new_AGEMA_signal_15843 ;
    wire new_AGEMA_signal_15844 ;
    wire new_AGEMA_signal_15845 ;
    wire new_AGEMA_signal_15846 ;
    wire new_AGEMA_signal_15847 ;
    wire new_AGEMA_signal_15848 ;
    wire new_AGEMA_signal_15849 ;
    wire new_AGEMA_signal_15850 ;
    wire new_AGEMA_signal_15851 ;
    wire new_AGEMA_signal_15852 ;
    wire new_AGEMA_signal_15853 ;
    wire new_AGEMA_signal_15854 ;
    wire new_AGEMA_signal_15855 ;
    wire new_AGEMA_signal_15856 ;
    wire new_AGEMA_signal_15857 ;
    wire new_AGEMA_signal_15858 ;
    wire new_AGEMA_signal_15859 ;
    wire new_AGEMA_signal_15860 ;
    wire new_AGEMA_signal_15861 ;
    wire new_AGEMA_signal_15862 ;
    wire new_AGEMA_signal_15863 ;
    wire new_AGEMA_signal_15864 ;
    wire new_AGEMA_signal_15865 ;
    wire new_AGEMA_signal_15866 ;
    wire new_AGEMA_signal_15867 ;
    wire new_AGEMA_signal_15868 ;
    wire new_AGEMA_signal_15869 ;
    wire new_AGEMA_signal_15870 ;
    wire new_AGEMA_signal_15871 ;
    wire new_AGEMA_signal_15872 ;
    wire new_AGEMA_signal_15873 ;
    wire new_AGEMA_signal_15874 ;
    wire new_AGEMA_signal_15875 ;
    wire new_AGEMA_signal_15876 ;
    wire new_AGEMA_signal_15877 ;
    wire new_AGEMA_signal_15878 ;
    wire new_AGEMA_signal_15879 ;
    wire new_AGEMA_signal_15880 ;
    wire new_AGEMA_signal_15881 ;
    wire new_AGEMA_signal_15882 ;
    wire new_AGEMA_signal_15883 ;
    wire new_AGEMA_signal_15884 ;
    wire new_AGEMA_signal_15885 ;
    wire new_AGEMA_signal_15886 ;
    wire new_AGEMA_signal_15887 ;
    wire new_AGEMA_signal_15888 ;
    wire new_AGEMA_signal_15889 ;
    wire new_AGEMA_signal_15890 ;
    wire new_AGEMA_signal_15891 ;
    wire new_AGEMA_signal_15892 ;
    wire new_AGEMA_signal_15893 ;
    wire new_AGEMA_signal_15894 ;
    wire new_AGEMA_signal_15895 ;
    wire new_AGEMA_signal_15896 ;
    wire new_AGEMA_signal_15897 ;
    wire new_AGEMA_signal_15898 ;
    wire new_AGEMA_signal_15899 ;
    wire new_AGEMA_signal_15900 ;
    wire new_AGEMA_signal_15901 ;
    wire new_AGEMA_signal_15902 ;
    wire new_AGEMA_signal_15903 ;
    wire new_AGEMA_signal_15904 ;
    wire new_AGEMA_signal_15905 ;
    wire new_AGEMA_signal_15906 ;
    wire new_AGEMA_signal_15907 ;
    wire new_AGEMA_signal_15908 ;
    wire new_AGEMA_signal_15909 ;
    wire new_AGEMA_signal_15910 ;
    wire new_AGEMA_signal_15911 ;
    wire new_AGEMA_signal_15912 ;
    wire new_AGEMA_signal_15913 ;
    wire new_AGEMA_signal_15914 ;
    wire new_AGEMA_signal_15915 ;
    wire new_AGEMA_signal_15916 ;
    wire new_AGEMA_signal_15917 ;
    wire new_AGEMA_signal_15918 ;
    wire new_AGEMA_signal_15919 ;
    wire new_AGEMA_signal_15920 ;
    wire new_AGEMA_signal_15921 ;
    wire new_AGEMA_signal_15922 ;
    wire new_AGEMA_signal_15923 ;
    wire new_AGEMA_signal_15924 ;
    wire new_AGEMA_signal_15925 ;
    wire new_AGEMA_signal_15926 ;
    wire new_AGEMA_signal_15927 ;
    wire new_AGEMA_signal_15928 ;
    wire new_AGEMA_signal_15929 ;
    wire new_AGEMA_signal_15930 ;
    wire new_AGEMA_signal_15931 ;
    wire new_AGEMA_signal_15932 ;
    wire new_AGEMA_signal_15933 ;
    wire new_AGEMA_signal_15934 ;
    wire new_AGEMA_signal_15935 ;
    wire new_AGEMA_signal_15936 ;
    wire new_AGEMA_signal_15937 ;
    wire new_AGEMA_signal_15938 ;
    wire new_AGEMA_signal_15939 ;
    wire new_AGEMA_signal_15940 ;
    wire new_AGEMA_signal_15941 ;
    wire new_AGEMA_signal_15942 ;
    wire new_AGEMA_signal_15943 ;
    wire new_AGEMA_signal_15944 ;
    wire new_AGEMA_signal_15945 ;
    wire new_AGEMA_signal_15946 ;
    wire new_AGEMA_signal_15947 ;
    wire new_AGEMA_signal_15948 ;
    wire new_AGEMA_signal_15949 ;
    wire new_AGEMA_signal_15950 ;
    wire new_AGEMA_signal_15951 ;
    wire new_AGEMA_signal_15952 ;
    wire new_AGEMA_signal_15953 ;
    wire new_AGEMA_signal_15954 ;
    wire new_AGEMA_signal_15955 ;
    wire new_AGEMA_signal_15956 ;
    wire new_AGEMA_signal_15957 ;
    wire new_AGEMA_signal_15958 ;
    wire new_AGEMA_signal_15959 ;
    wire new_AGEMA_signal_15960 ;
    wire new_AGEMA_signal_15961 ;
    wire new_AGEMA_signal_15962 ;
    wire new_AGEMA_signal_15963 ;
    wire new_AGEMA_signal_15964 ;
    wire new_AGEMA_signal_15965 ;
    wire new_AGEMA_signal_15966 ;
    wire new_AGEMA_signal_15967 ;
    wire new_AGEMA_signal_15968 ;
    wire new_AGEMA_signal_15969 ;
    wire new_AGEMA_signal_15970 ;
    wire new_AGEMA_signal_15971 ;
    wire new_AGEMA_signal_15972 ;
    wire new_AGEMA_signal_15973 ;
    wire new_AGEMA_signal_15974 ;
    wire new_AGEMA_signal_15975 ;
    wire new_AGEMA_signal_15976 ;
    wire new_AGEMA_signal_15977 ;
    wire new_AGEMA_signal_15978 ;
    wire new_AGEMA_signal_15979 ;
    wire new_AGEMA_signal_15980 ;
    wire new_AGEMA_signal_15981 ;
    wire new_AGEMA_signal_15982 ;
    wire new_AGEMA_signal_15983 ;
    wire new_AGEMA_signal_15984 ;
    wire new_AGEMA_signal_15985 ;
    wire new_AGEMA_signal_15986 ;
    wire new_AGEMA_signal_15987 ;
    wire new_AGEMA_signal_15988 ;
    wire new_AGEMA_signal_15989 ;
    wire new_AGEMA_signal_15990 ;
    wire new_AGEMA_signal_15991 ;
    wire new_AGEMA_signal_15992 ;
    wire new_AGEMA_signal_15993 ;
    wire new_AGEMA_signal_15994 ;
    wire new_AGEMA_signal_15995 ;
    wire new_AGEMA_signal_15996 ;
    wire new_AGEMA_signal_15997 ;
    wire new_AGEMA_signal_15998 ;
    wire new_AGEMA_signal_15999 ;
    wire new_AGEMA_signal_16000 ;
    wire new_AGEMA_signal_16001 ;
    wire new_AGEMA_signal_16002 ;
    wire new_AGEMA_signal_16003 ;
    wire new_AGEMA_signal_16004 ;
    wire new_AGEMA_signal_16005 ;
    wire new_AGEMA_signal_16006 ;
    wire new_AGEMA_signal_16007 ;
    wire new_AGEMA_signal_16008 ;
    wire new_AGEMA_signal_16009 ;
    wire new_AGEMA_signal_16010 ;
    wire new_AGEMA_signal_16011 ;
    wire new_AGEMA_signal_16012 ;
    wire new_AGEMA_signal_16013 ;
    wire new_AGEMA_signal_16014 ;
    wire new_AGEMA_signal_16015 ;
    wire new_AGEMA_signal_16016 ;
    wire new_AGEMA_signal_16017 ;
    wire new_AGEMA_signal_16018 ;
    wire new_AGEMA_signal_16019 ;
    wire new_AGEMA_signal_16020 ;
    wire new_AGEMA_signal_16021 ;
    wire new_AGEMA_signal_16022 ;
    wire new_AGEMA_signal_16023 ;
    wire new_AGEMA_signal_16024 ;
    wire new_AGEMA_signal_16025 ;
    wire new_AGEMA_signal_16026 ;
    wire new_AGEMA_signal_16027 ;
    wire new_AGEMA_signal_16028 ;
    wire new_AGEMA_signal_16029 ;
    wire new_AGEMA_signal_16030 ;
    wire new_AGEMA_signal_16031 ;
    wire new_AGEMA_signal_16032 ;
    wire new_AGEMA_signal_16033 ;
    wire new_AGEMA_signal_16034 ;
    wire new_AGEMA_signal_16035 ;
    wire new_AGEMA_signal_16036 ;
    wire new_AGEMA_signal_16037 ;
    wire new_AGEMA_signal_16038 ;
    wire new_AGEMA_signal_16039 ;
    wire new_AGEMA_signal_16040 ;
    wire new_AGEMA_signal_16041 ;
    wire new_AGEMA_signal_16042 ;
    wire new_AGEMA_signal_16043 ;
    wire new_AGEMA_signal_16044 ;
    wire new_AGEMA_signal_16045 ;
    wire new_AGEMA_signal_16046 ;
    wire new_AGEMA_signal_16047 ;
    wire new_AGEMA_signal_16048 ;
    wire new_AGEMA_signal_16049 ;
    wire new_AGEMA_signal_16050 ;
    wire new_AGEMA_signal_16051 ;
    wire new_AGEMA_signal_16052 ;
    wire new_AGEMA_signal_16053 ;
    wire new_AGEMA_signal_16054 ;
    wire new_AGEMA_signal_16055 ;
    wire new_AGEMA_signal_16056 ;
    wire new_AGEMA_signal_16057 ;
    wire new_AGEMA_signal_16058 ;
    wire new_AGEMA_signal_16059 ;
    wire new_AGEMA_signal_16060 ;
    wire new_AGEMA_signal_16061 ;
    wire new_AGEMA_signal_16062 ;
    wire new_AGEMA_signal_16063 ;
    wire new_AGEMA_signal_16064 ;
    wire new_AGEMA_signal_16065 ;
    wire new_AGEMA_signal_16066 ;
    wire new_AGEMA_signal_16067 ;
    wire new_AGEMA_signal_16068 ;
    wire new_AGEMA_signal_16069 ;
    wire new_AGEMA_signal_16070 ;
    wire new_AGEMA_signal_16071 ;
    wire new_AGEMA_signal_16072 ;
    wire new_AGEMA_signal_16073 ;
    wire new_AGEMA_signal_16074 ;
    wire new_AGEMA_signal_16075 ;
    wire new_AGEMA_signal_16076 ;
    wire new_AGEMA_signal_16077 ;
    wire new_AGEMA_signal_16078 ;
    wire new_AGEMA_signal_16079 ;
    wire new_AGEMA_signal_16080 ;
    wire new_AGEMA_signal_16081 ;
    wire new_AGEMA_signal_16082 ;
    wire new_AGEMA_signal_16083 ;
    wire new_AGEMA_signal_16084 ;
    wire new_AGEMA_signal_16085 ;
    wire new_AGEMA_signal_16086 ;
    wire new_AGEMA_signal_16087 ;
    wire new_AGEMA_signal_16088 ;
    wire new_AGEMA_signal_16089 ;
    wire new_AGEMA_signal_16090 ;
    wire new_AGEMA_signal_16091 ;
    wire new_AGEMA_signal_16092 ;
    wire new_AGEMA_signal_16093 ;
    wire new_AGEMA_signal_16094 ;
    wire new_AGEMA_signal_16095 ;
    wire new_AGEMA_signal_16096 ;
    wire new_AGEMA_signal_16097 ;
    wire new_AGEMA_signal_16098 ;
    wire new_AGEMA_signal_16099 ;
    wire new_AGEMA_signal_16100 ;
    wire new_AGEMA_signal_16101 ;
    wire new_AGEMA_signal_16102 ;
    wire new_AGEMA_signal_16103 ;
    wire new_AGEMA_signal_16104 ;
    wire new_AGEMA_signal_16105 ;
    wire new_AGEMA_signal_16106 ;
    wire new_AGEMA_signal_16107 ;
    wire new_AGEMA_signal_16108 ;
    wire new_AGEMA_signal_16109 ;
    wire new_AGEMA_signal_16110 ;
    wire new_AGEMA_signal_16111 ;
    wire new_AGEMA_signal_16112 ;
    wire new_AGEMA_signal_16113 ;
    wire new_AGEMA_signal_16114 ;
    wire new_AGEMA_signal_16115 ;
    wire new_AGEMA_signal_16116 ;
    wire new_AGEMA_signal_16117 ;
    wire new_AGEMA_signal_16118 ;
    wire new_AGEMA_signal_16119 ;
    wire new_AGEMA_signal_16120 ;
    wire new_AGEMA_signal_16121 ;
    wire new_AGEMA_signal_16122 ;
    wire new_AGEMA_signal_16123 ;
    wire new_AGEMA_signal_16124 ;
    wire new_AGEMA_signal_16125 ;
    wire new_AGEMA_signal_16126 ;
    wire new_AGEMA_signal_16127 ;
    wire new_AGEMA_signal_16128 ;
    wire new_AGEMA_signal_16129 ;
    wire new_AGEMA_signal_16130 ;
    wire new_AGEMA_signal_16131 ;
    wire new_AGEMA_signal_16132 ;
    wire new_AGEMA_signal_16133 ;
    wire new_AGEMA_signal_16134 ;
    wire new_AGEMA_signal_16135 ;
    wire new_AGEMA_signal_16136 ;
    wire new_AGEMA_signal_16137 ;
    wire new_AGEMA_signal_16138 ;
    wire new_AGEMA_signal_16139 ;
    wire new_AGEMA_signal_16140 ;
    wire new_AGEMA_signal_16141 ;
    wire new_AGEMA_signal_16142 ;
    wire new_AGEMA_signal_16143 ;
    wire new_AGEMA_signal_16144 ;
    wire new_AGEMA_signal_16145 ;
    wire new_AGEMA_signal_16146 ;
    wire new_AGEMA_signal_16147 ;
    wire new_AGEMA_signal_16148 ;
    wire new_AGEMA_signal_16149 ;
    wire new_AGEMA_signal_16150 ;
    wire new_AGEMA_signal_16151 ;
    wire new_AGEMA_signal_16152 ;
    wire new_AGEMA_signal_16153 ;
    wire new_AGEMA_signal_16154 ;
    wire new_AGEMA_signal_16155 ;
    wire new_AGEMA_signal_16156 ;
    wire new_AGEMA_signal_16157 ;
    wire new_AGEMA_signal_16158 ;
    wire new_AGEMA_signal_16159 ;
    wire new_AGEMA_signal_16160 ;
    wire new_AGEMA_signal_16161 ;
    wire new_AGEMA_signal_16162 ;
    wire new_AGEMA_signal_16163 ;
    wire new_AGEMA_signal_16164 ;
    wire new_AGEMA_signal_16165 ;
    wire new_AGEMA_signal_16166 ;
    wire new_AGEMA_signal_16167 ;
    wire new_AGEMA_signal_16168 ;
    wire new_AGEMA_signal_16169 ;
    wire new_AGEMA_signal_16170 ;
    wire new_AGEMA_signal_16171 ;
    wire new_AGEMA_signal_16172 ;
    wire new_AGEMA_signal_16173 ;
    wire new_AGEMA_signal_16174 ;
    wire new_AGEMA_signal_16175 ;
    wire new_AGEMA_signal_16176 ;
    wire new_AGEMA_signal_16177 ;
    wire new_AGEMA_signal_16178 ;
    wire new_AGEMA_signal_16179 ;
    wire new_AGEMA_signal_16180 ;
    wire new_AGEMA_signal_16181 ;
    wire new_AGEMA_signal_16182 ;
    wire new_AGEMA_signal_16183 ;
    wire new_AGEMA_signal_16184 ;
    wire new_AGEMA_signal_16185 ;
    wire new_AGEMA_signal_16186 ;
    wire new_AGEMA_signal_16187 ;
    wire new_AGEMA_signal_16188 ;
    wire new_AGEMA_signal_16189 ;
    wire new_AGEMA_signal_16190 ;
    wire new_AGEMA_signal_16191 ;
    wire new_AGEMA_signal_16192 ;
    wire new_AGEMA_signal_16193 ;
    wire new_AGEMA_signal_16194 ;
    wire new_AGEMA_signal_16195 ;
    wire new_AGEMA_signal_16196 ;
    wire new_AGEMA_signal_16197 ;
    wire new_AGEMA_signal_16198 ;
    wire new_AGEMA_signal_16199 ;
    wire new_AGEMA_signal_16200 ;
    wire new_AGEMA_signal_16201 ;
    wire new_AGEMA_signal_16202 ;
    wire new_AGEMA_signal_16203 ;
    wire new_AGEMA_signal_16204 ;
    wire new_AGEMA_signal_16205 ;
    wire new_AGEMA_signal_16206 ;
    wire new_AGEMA_signal_16207 ;
    wire new_AGEMA_signal_16208 ;
    wire new_AGEMA_signal_16209 ;
    wire new_AGEMA_signal_16210 ;
    wire new_AGEMA_signal_16211 ;
    wire new_AGEMA_signal_16212 ;
    wire new_AGEMA_signal_16213 ;
    wire new_AGEMA_signal_16214 ;
    wire new_AGEMA_signal_16215 ;
    wire new_AGEMA_signal_16216 ;
    wire new_AGEMA_signal_16217 ;
    wire new_AGEMA_signal_16218 ;
    wire new_AGEMA_signal_16219 ;
    wire new_AGEMA_signal_16220 ;
    wire new_AGEMA_signal_16221 ;
    wire new_AGEMA_signal_16222 ;
    wire new_AGEMA_signal_16223 ;
    wire new_AGEMA_signal_16224 ;
    wire new_AGEMA_signal_16225 ;
    wire new_AGEMA_signal_16226 ;
    wire new_AGEMA_signal_16227 ;
    wire new_AGEMA_signal_16228 ;
    wire new_AGEMA_signal_16229 ;
    wire new_AGEMA_signal_16230 ;
    wire new_AGEMA_signal_16231 ;
    wire new_AGEMA_signal_16232 ;
    wire new_AGEMA_signal_16233 ;
    wire new_AGEMA_signal_16234 ;
    wire new_AGEMA_signal_16235 ;
    wire new_AGEMA_signal_16236 ;
    wire new_AGEMA_signal_16237 ;
    wire new_AGEMA_signal_16238 ;
    wire new_AGEMA_signal_16239 ;
    wire new_AGEMA_signal_16240 ;
    wire new_AGEMA_signal_16241 ;
    wire new_AGEMA_signal_16242 ;
    wire new_AGEMA_signal_16243 ;
    wire new_AGEMA_signal_16244 ;
    wire new_AGEMA_signal_16245 ;
    wire new_AGEMA_signal_16246 ;
    wire new_AGEMA_signal_16247 ;
    wire new_AGEMA_signal_16248 ;
    wire new_AGEMA_signal_16249 ;
    wire new_AGEMA_signal_16250 ;
    wire new_AGEMA_signal_16251 ;
    wire new_AGEMA_signal_16252 ;
    wire new_AGEMA_signal_16253 ;
    wire new_AGEMA_signal_16254 ;
    wire new_AGEMA_signal_16255 ;
    wire new_AGEMA_signal_16256 ;
    wire new_AGEMA_signal_16257 ;
    wire new_AGEMA_signal_16258 ;
    wire new_AGEMA_signal_16259 ;
    wire new_AGEMA_signal_16260 ;
    wire new_AGEMA_signal_16261 ;
    wire new_AGEMA_signal_16262 ;
    wire new_AGEMA_signal_16263 ;
    wire new_AGEMA_signal_16264 ;
    wire new_AGEMA_signal_16265 ;
    wire new_AGEMA_signal_16266 ;
    wire new_AGEMA_signal_16267 ;
    wire new_AGEMA_signal_16268 ;
    wire new_AGEMA_signal_16269 ;
    wire new_AGEMA_signal_16270 ;
    wire new_AGEMA_signal_16271 ;
    wire new_AGEMA_signal_16272 ;
    wire new_AGEMA_signal_16273 ;
    wire new_AGEMA_signal_16274 ;
    wire new_AGEMA_signal_16275 ;
    wire new_AGEMA_signal_16276 ;
    wire new_AGEMA_signal_16277 ;
    wire new_AGEMA_signal_16278 ;
    wire new_AGEMA_signal_16279 ;
    wire new_AGEMA_signal_16280 ;
    wire new_AGEMA_signal_16281 ;
    wire new_AGEMA_signal_16282 ;
    wire new_AGEMA_signal_16283 ;
    wire new_AGEMA_signal_16284 ;
    wire new_AGEMA_signal_16285 ;
    wire new_AGEMA_signal_16286 ;
    wire new_AGEMA_signal_16287 ;
    wire new_AGEMA_signal_16288 ;
    wire new_AGEMA_signal_16289 ;
    wire new_AGEMA_signal_16290 ;
    wire new_AGEMA_signal_16291 ;
    wire new_AGEMA_signal_16292 ;
    wire new_AGEMA_signal_16293 ;
    wire new_AGEMA_signal_16294 ;
    wire new_AGEMA_signal_16295 ;
    wire new_AGEMA_signal_16296 ;
    wire new_AGEMA_signal_16297 ;
    wire new_AGEMA_signal_16298 ;
    wire new_AGEMA_signal_16299 ;
    wire new_AGEMA_signal_16300 ;
    wire new_AGEMA_signal_16301 ;
    wire new_AGEMA_signal_16302 ;
    wire new_AGEMA_signal_16303 ;
    wire new_AGEMA_signal_16304 ;
    wire new_AGEMA_signal_16305 ;
    wire new_AGEMA_signal_16306 ;
    wire new_AGEMA_signal_16307 ;
    wire new_AGEMA_signal_16308 ;
    wire new_AGEMA_signal_16309 ;
    wire new_AGEMA_signal_16310 ;
    wire new_AGEMA_signal_16311 ;
    wire new_AGEMA_signal_16312 ;
    wire new_AGEMA_signal_16313 ;
    wire new_AGEMA_signal_16314 ;
    wire new_AGEMA_signal_16315 ;
    wire new_AGEMA_signal_16316 ;
    wire new_AGEMA_signal_16317 ;
    wire new_AGEMA_signal_16318 ;
    wire new_AGEMA_signal_16319 ;
    wire new_AGEMA_signal_16320 ;
    wire new_AGEMA_signal_16321 ;
    wire new_AGEMA_signal_16322 ;
    wire new_AGEMA_signal_16323 ;
    wire new_AGEMA_signal_16324 ;
    wire new_AGEMA_signal_16325 ;
    wire new_AGEMA_signal_16326 ;
    wire new_AGEMA_signal_16327 ;
    wire new_AGEMA_signal_16328 ;
    wire new_AGEMA_signal_16329 ;
    wire new_AGEMA_signal_16330 ;
    wire new_AGEMA_signal_16331 ;
    wire new_AGEMA_signal_16332 ;
    wire new_AGEMA_signal_16333 ;
    wire new_AGEMA_signal_16334 ;
    wire new_AGEMA_signal_16335 ;
    wire new_AGEMA_signal_16336 ;
    wire new_AGEMA_signal_16337 ;
    wire new_AGEMA_signal_16338 ;
    wire new_AGEMA_signal_16339 ;
    wire new_AGEMA_signal_16340 ;
    wire new_AGEMA_signal_16341 ;
    wire new_AGEMA_signal_16342 ;
    wire new_AGEMA_signal_16343 ;
    wire new_AGEMA_signal_16344 ;
    wire new_AGEMA_signal_16345 ;
    wire new_AGEMA_signal_16346 ;
    wire new_AGEMA_signal_16347 ;
    wire new_AGEMA_signal_16348 ;
    wire new_AGEMA_signal_16349 ;
    wire new_AGEMA_signal_16350 ;
    wire new_AGEMA_signal_16351 ;
    wire new_AGEMA_signal_16352 ;
    wire new_AGEMA_signal_16353 ;
    wire new_AGEMA_signal_16354 ;
    wire new_AGEMA_signal_16355 ;
    wire new_AGEMA_signal_16356 ;
    wire new_AGEMA_signal_16357 ;
    wire new_AGEMA_signal_16358 ;
    wire new_AGEMA_signal_16359 ;
    wire new_AGEMA_signal_16360 ;
    wire new_AGEMA_signal_16361 ;
    wire new_AGEMA_signal_16362 ;
    wire new_AGEMA_signal_16363 ;
    wire new_AGEMA_signal_16364 ;
    wire new_AGEMA_signal_16365 ;
    wire new_AGEMA_signal_16366 ;
    wire new_AGEMA_signal_16367 ;
    wire new_AGEMA_signal_16368 ;
    wire new_AGEMA_signal_16369 ;
    wire new_AGEMA_signal_16370 ;
    wire new_AGEMA_signal_16371 ;
    wire new_AGEMA_signal_16372 ;
    wire new_AGEMA_signal_16373 ;
    wire new_AGEMA_signal_16374 ;
    wire new_AGEMA_signal_16375 ;
    wire new_AGEMA_signal_16376 ;
    wire new_AGEMA_signal_16377 ;
    wire new_AGEMA_signal_16378 ;
    wire new_AGEMA_signal_16379 ;
    wire new_AGEMA_signal_16380 ;
    wire new_AGEMA_signal_16381 ;
    wire new_AGEMA_signal_16382 ;
    wire new_AGEMA_signal_16383 ;
    wire new_AGEMA_signal_16384 ;
    wire new_AGEMA_signal_16385 ;
    wire new_AGEMA_signal_16386 ;
    wire new_AGEMA_signal_16387 ;
    wire new_AGEMA_signal_16388 ;
    wire new_AGEMA_signal_16389 ;
    wire new_AGEMA_signal_16390 ;
    wire new_AGEMA_signal_16391 ;
    wire new_AGEMA_signal_16392 ;
    wire new_AGEMA_signal_16393 ;
    wire new_AGEMA_signal_16394 ;
    wire new_AGEMA_signal_16395 ;
    wire new_AGEMA_signal_16396 ;
    wire new_AGEMA_signal_16397 ;
    wire new_AGEMA_signal_16398 ;
    wire new_AGEMA_signal_16399 ;
    wire new_AGEMA_signal_16400 ;
    wire new_AGEMA_signal_16401 ;
    wire new_AGEMA_signal_16402 ;
    wire new_AGEMA_signal_16403 ;
    wire new_AGEMA_signal_16404 ;
    wire new_AGEMA_signal_16405 ;
    wire new_AGEMA_signal_16406 ;
    wire new_AGEMA_signal_16407 ;
    wire new_AGEMA_signal_16408 ;
    wire new_AGEMA_signal_16409 ;
    wire new_AGEMA_signal_16410 ;
    wire new_AGEMA_signal_16411 ;
    wire new_AGEMA_signal_16412 ;
    wire new_AGEMA_signal_16413 ;
    wire new_AGEMA_signal_16414 ;
    wire new_AGEMA_signal_16415 ;
    wire new_AGEMA_signal_16416 ;
    wire new_AGEMA_signal_16417 ;
    wire new_AGEMA_signal_16418 ;
    wire new_AGEMA_signal_16419 ;
    wire new_AGEMA_signal_16420 ;
    wire new_AGEMA_signal_16421 ;
    wire new_AGEMA_signal_16422 ;
    wire new_AGEMA_signal_16423 ;
    wire new_AGEMA_signal_16424 ;
    wire new_AGEMA_signal_16425 ;
    wire new_AGEMA_signal_16426 ;
    wire new_AGEMA_signal_16427 ;
    wire new_AGEMA_signal_16428 ;
    wire new_AGEMA_signal_16429 ;
    wire new_AGEMA_signal_16430 ;
    wire new_AGEMA_signal_16431 ;
    wire new_AGEMA_signal_16432 ;
    wire new_AGEMA_signal_16433 ;
    wire new_AGEMA_signal_16434 ;
    wire new_AGEMA_signal_16435 ;
    wire new_AGEMA_signal_16436 ;
    wire new_AGEMA_signal_16437 ;
    wire new_AGEMA_signal_16438 ;
    wire new_AGEMA_signal_16439 ;
    wire new_AGEMA_signal_16440 ;
    wire new_AGEMA_signal_16441 ;
    wire new_AGEMA_signal_16442 ;
    wire new_AGEMA_signal_16443 ;
    wire new_AGEMA_signal_16444 ;
    wire new_AGEMA_signal_16445 ;
    wire new_AGEMA_signal_16446 ;
    wire new_AGEMA_signal_16447 ;
    wire new_AGEMA_signal_16448 ;
    wire new_AGEMA_signal_16449 ;
    wire new_AGEMA_signal_16450 ;
    wire new_AGEMA_signal_16451 ;
    wire new_AGEMA_signal_16452 ;
    wire new_AGEMA_signal_16453 ;
    wire new_AGEMA_signal_16454 ;
    wire new_AGEMA_signal_16455 ;
    wire new_AGEMA_signal_16456 ;
    wire new_AGEMA_signal_16457 ;
    wire new_AGEMA_signal_16458 ;
    wire new_AGEMA_signal_16459 ;
    wire new_AGEMA_signal_16460 ;
    wire new_AGEMA_signal_16461 ;
    wire new_AGEMA_signal_16462 ;
    wire new_AGEMA_signal_16463 ;
    wire new_AGEMA_signal_16464 ;
    wire new_AGEMA_signal_16465 ;
    wire new_AGEMA_signal_16466 ;
    wire new_AGEMA_signal_16467 ;
    wire new_AGEMA_signal_16468 ;
    wire new_AGEMA_signal_16469 ;
    wire new_AGEMA_signal_16470 ;
    wire new_AGEMA_signal_16471 ;
    wire new_AGEMA_signal_16472 ;
    wire new_AGEMA_signal_16473 ;
    wire new_AGEMA_signal_16474 ;
    wire new_AGEMA_signal_16475 ;
    wire new_AGEMA_signal_16476 ;
    wire new_AGEMA_signal_16477 ;
    wire new_AGEMA_signal_16478 ;
    wire new_AGEMA_signal_16479 ;
    wire new_AGEMA_signal_16480 ;
    wire new_AGEMA_signal_16481 ;
    wire new_AGEMA_signal_16482 ;
    wire new_AGEMA_signal_16483 ;
    wire new_AGEMA_signal_16484 ;
    wire new_AGEMA_signal_16485 ;
    wire new_AGEMA_signal_16486 ;
    wire new_AGEMA_signal_16487 ;
    wire new_AGEMA_signal_16488 ;
    wire new_AGEMA_signal_16489 ;
    wire new_AGEMA_signal_16490 ;
    wire new_AGEMA_signal_16491 ;
    wire new_AGEMA_signal_16492 ;
    wire new_AGEMA_signal_16493 ;
    wire new_AGEMA_signal_16494 ;
    wire new_AGEMA_signal_16495 ;
    wire new_AGEMA_signal_16496 ;
    wire new_AGEMA_signal_16497 ;
    wire new_AGEMA_signal_16498 ;
    wire new_AGEMA_signal_16499 ;
    wire new_AGEMA_signal_16500 ;
    wire new_AGEMA_signal_16501 ;
    wire new_AGEMA_signal_16502 ;
    wire new_AGEMA_signal_16503 ;
    wire new_AGEMA_signal_16504 ;
    wire new_AGEMA_signal_16505 ;
    wire new_AGEMA_signal_16506 ;
    wire new_AGEMA_signal_16507 ;
    wire new_AGEMA_signal_16508 ;
    wire new_AGEMA_signal_16509 ;
    wire new_AGEMA_signal_16510 ;
    wire new_AGEMA_signal_16511 ;
    wire new_AGEMA_signal_16512 ;
    wire new_AGEMA_signal_16513 ;
    wire new_AGEMA_signal_16514 ;
    wire new_AGEMA_signal_16515 ;
    wire new_AGEMA_signal_16516 ;
    wire new_AGEMA_signal_16517 ;
    wire new_AGEMA_signal_16518 ;
    wire new_AGEMA_signal_16519 ;
    wire new_AGEMA_signal_16520 ;
    wire new_AGEMA_signal_16521 ;
    wire new_AGEMA_signal_16522 ;
    wire new_AGEMA_signal_16523 ;
    wire new_AGEMA_signal_16524 ;
    wire new_AGEMA_signal_16525 ;
    wire new_AGEMA_signal_16526 ;
    wire new_AGEMA_signal_16527 ;
    wire new_AGEMA_signal_16528 ;
    wire new_AGEMA_signal_16529 ;
    wire new_AGEMA_signal_16530 ;
    wire new_AGEMA_signal_16531 ;
    wire new_AGEMA_signal_16532 ;
    wire new_AGEMA_signal_16533 ;
    wire new_AGEMA_signal_16534 ;
    wire new_AGEMA_signal_16535 ;
    wire new_AGEMA_signal_16536 ;
    wire new_AGEMA_signal_16537 ;
    wire new_AGEMA_signal_16538 ;
    wire new_AGEMA_signal_16539 ;
    wire new_AGEMA_signal_16540 ;
    wire new_AGEMA_signal_16541 ;
    wire new_AGEMA_signal_16542 ;
    wire new_AGEMA_signal_16543 ;
    wire new_AGEMA_signal_16544 ;
    wire new_AGEMA_signal_16545 ;
    wire new_AGEMA_signal_16546 ;
    wire new_AGEMA_signal_16547 ;
    wire new_AGEMA_signal_16548 ;
    wire new_AGEMA_signal_16549 ;
    wire new_AGEMA_signal_16550 ;
    wire new_AGEMA_signal_16551 ;
    wire new_AGEMA_signal_16552 ;
    wire new_AGEMA_signal_16553 ;
    wire new_AGEMA_signal_16554 ;
    wire new_AGEMA_signal_16555 ;
    wire new_AGEMA_signal_16556 ;
    wire new_AGEMA_signal_16557 ;
    wire new_AGEMA_signal_16558 ;
    wire new_AGEMA_signal_16559 ;
    wire new_AGEMA_signal_16560 ;
    wire new_AGEMA_signal_16561 ;
    wire new_AGEMA_signal_16562 ;
    wire new_AGEMA_signal_16563 ;
    wire new_AGEMA_signal_16564 ;
    wire new_AGEMA_signal_16565 ;
    wire new_AGEMA_signal_16566 ;
    wire new_AGEMA_signal_16567 ;
    wire new_AGEMA_signal_16568 ;
    wire new_AGEMA_signal_16569 ;
    wire new_AGEMA_signal_16570 ;
    wire new_AGEMA_signal_16571 ;
    wire new_AGEMA_signal_16572 ;
    wire new_AGEMA_signal_16573 ;
    wire new_AGEMA_signal_16574 ;
    wire new_AGEMA_signal_16575 ;
    wire new_AGEMA_signal_16576 ;
    wire new_AGEMA_signal_16577 ;
    wire new_AGEMA_signal_16578 ;
    wire new_AGEMA_signal_16579 ;
    wire new_AGEMA_signal_16580 ;
    wire new_AGEMA_signal_16581 ;
    wire new_AGEMA_signal_16582 ;
    wire new_AGEMA_signal_16583 ;
    wire new_AGEMA_signal_16584 ;
    wire new_AGEMA_signal_16585 ;
    wire new_AGEMA_signal_16586 ;
    wire new_AGEMA_signal_16587 ;
    wire new_AGEMA_signal_16588 ;
    wire new_AGEMA_signal_16589 ;
    wire new_AGEMA_signal_16590 ;
    wire new_AGEMA_signal_16591 ;
    wire new_AGEMA_signal_16592 ;
    wire new_AGEMA_signal_16593 ;
    wire new_AGEMA_signal_16594 ;
    wire new_AGEMA_signal_16595 ;
    wire new_AGEMA_signal_16596 ;
    wire new_AGEMA_signal_16597 ;
    wire new_AGEMA_signal_16598 ;
    wire new_AGEMA_signal_16599 ;
    wire new_AGEMA_signal_16600 ;
    wire new_AGEMA_signal_16601 ;
    wire new_AGEMA_signal_16602 ;
    wire new_AGEMA_signal_16603 ;
    wire new_AGEMA_signal_16604 ;
    wire new_AGEMA_signal_16605 ;
    wire new_AGEMA_signal_16606 ;
    wire new_AGEMA_signal_16607 ;
    wire new_AGEMA_signal_16608 ;
    wire new_AGEMA_signal_16609 ;
    wire new_AGEMA_signal_16610 ;
    wire new_AGEMA_signal_16611 ;
    wire new_AGEMA_signal_16612 ;
    wire new_AGEMA_signal_16613 ;
    wire new_AGEMA_signal_16614 ;
    wire new_AGEMA_signal_16615 ;
    wire new_AGEMA_signal_16616 ;
    wire new_AGEMA_signal_16617 ;
    wire new_AGEMA_signal_16618 ;
    wire new_AGEMA_signal_16619 ;
    wire new_AGEMA_signal_16620 ;
    wire new_AGEMA_signal_16621 ;
    wire new_AGEMA_signal_16622 ;
    wire new_AGEMA_signal_16623 ;
    wire new_AGEMA_signal_16624 ;
    wire new_AGEMA_signal_16625 ;
    wire new_AGEMA_signal_16626 ;
    wire new_AGEMA_signal_16627 ;
    wire new_AGEMA_signal_16628 ;
    wire new_AGEMA_signal_16629 ;
    wire new_AGEMA_signal_16630 ;
    wire new_AGEMA_signal_16631 ;
    wire new_AGEMA_signal_16632 ;
    wire new_AGEMA_signal_16633 ;
    wire new_AGEMA_signal_16634 ;
    wire new_AGEMA_signal_16635 ;
    wire new_AGEMA_signal_16636 ;
    wire new_AGEMA_signal_16637 ;
    wire new_AGEMA_signal_16638 ;
    wire new_AGEMA_signal_16639 ;
    wire new_AGEMA_signal_16640 ;
    wire new_AGEMA_signal_16641 ;
    wire new_AGEMA_signal_16642 ;
    wire new_AGEMA_signal_16643 ;
    wire new_AGEMA_signal_16644 ;
    wire new_AGEMA_signal_16645 ;
    wire new_AGEMA_signal_16646 ;
    wire new_AGEMA_signal_16647 ;
    wire new_AGEMA_signal_16648 ;
    wire new_AGEMA_signal_16649 ;
    wire new_AGEMA_signal_16650 ;
    wire new_AGEMA_signal_16651 ;
    wire new_AGEMA_signal_16652 ;
    wire new_AGEMA_signal_16653 ;
    wire new_AGEMA_signal_16654 ;
    wire new_AGEMA_signal_16655 ;
    wire new_AGEMA_signal_16656 ;
    wire new_AGEMA_signal_16657 ;
    wire new_AGEMA_signal_16658 ;
    wire new_AGEMA_signal_16659 ;
    wire new_AGEMA_signal_16660 ;
    wire new_AGEMA_signal_16661 ;
    wire new_AGEMA_signal_16662 ;
    wire new_AGEMA_signal_16663 ;
    wire new_AGEMA_signal_16664 ;
    wire new_AGEMA_signal_16665 ;
    wire new_AGEMA_signal_16666 ;
    wire new_AGEMA_signal_16667 ;
    wire new_AGEMA_signal_16668 ;
    wire new_AGEMA_signal_16669 ;
    wire new_AGEMA_signal_16670 ;
    wire new_AGEMA_signal_16671 ;
    wire new_AGEMA_signal_16672 ;
    wire new_AGEMA_signal_16673 ;
    wire new_AGEMA_signal_16674 ;
    wire new_AGEMA_signal_16675 ;
    wire new_AGEMA_signal_16676 ;
    wire new_AGEMA_signal_16677 ;
    wire new_AGEMA_signal_16678 ;
    wire new_AGEMA_signal_16679 ;
    wire new_AGEMA_signal_16680 ;
    wire new_AGEMA_signal_16681 ;
    wire new_AGEMA_signal_16682 ;
    wire new_AGEMA_signal_16683 ;
    wire new_AGEMA_signal_16684 ;
    wire new_AGEMA_signal_16685 ;
    wire new_AGEMA_signal_16686 ;
    wire new_AGEMA_signal_16687 ;
    wire new_AGEMA_signal_16688 ;
    wire new_AGEMA_signal_16689 ;
    wire new_AGEMA_signal_16690 ;
    wire new_AGEMA_signal_16691 ;
    wire new_AGEMA_signal_16692 ;
    wire new_AGEMA_signal_16693 ;
    wire new_AGEMA_signal_16694 ;
    wire new_AGEMA_signal_16695 ;
    wire new_AGEMA_signal_16696 ;
    wire new_AGEMA_signal_16697 ;
    wire new_AGEMA_signal_16698 ;
    wire new_AGEMA_signal_16699 ;
    wire new_AGEMA_signal_16700 ;
    wire new_AGEMA_signal_16701 ;
    wire new_AGEMA_signal_16702 ;
    wire new_AGEMA_signal_16703 ;
    wire new_AGEMA_signal_16704 ;
    wire new_AGEMA_signal_16705 ;
    wire new_AGEMA_signal_16706 ;
    wire new_AGEMA_signal_16707 ;
    wire new_AGEMA_signal_16708 ;
    wire new_AGEMA_signal_16709 ;
    wire new_AGEMA_signal_16710 ;
    wire new_AGEMA_signal_16711 ;
    wire new_AGEMA_signal_16712 ;
    wire new_AGEMA_signal_16713 ;
    wire new_AGEMA_signal_16714 ;
    wire new_AGEMA_signal_16715 ;
    wire new_AGEMA_signal_16716 ;
    wire new_AGEMA_signal_16717 ;
    wire new_AGEMA_signal_16718 ;
    wire new_AGEMA_signal_16719 ;
    wire new_AGEMA_signal_16720 ;
    wire new_AGEMA_signal_16721 ;
    wire new_AGEMA_signal_16722 ;
    wire new_AGEMA_signal_16723 ;
    wire new_AGEMA_signal_16724 ;
    wire new_AGEMA_signal_16725 ;
    wire new_AGEMA_signal_16726 ;
    wire new_AGEMA_signal_16727 ;
    wire new_AGEMA_signal_16728 ;
    wire new_AGEMA_signal_16729 ;
    wire new_AGEMA_signal_16730 ;
    wire new_AGEMA_signal_16731 ;
    wire new_AGEMA_signal_16732 ;
    wire new_AGEMA_signal_16733 ;
    wire new_AGEMA_signal_16734 ;
    wire new_AGEMA_signal_16735 ;
    wire new_AGEMA_signal_16736 ;
    wire new_AGEMA_signal_16737 ;
    wire new_AGEMA_signal_16738 ;
    wire new_AGEMA_signal_16739 ;
    wire new_AGEMA_signal_16740 ;
    wire new_AGEMA_signal_16741 ;
    wire new_AGEMA_signal_16742 ;
    wire new_AGEMA_signal_16743 ;
    wire new_AGEMA_signal_16744 ;
    wire new_AGEMA_signal_16745 ;
    wire new_AGEMA_signal_16746 ;
    wire new_AGEMA_signal_16747 ;
    wire new_AGEMA_signal_16748 ;
    wire new_AGEMA_signal_16749 ;
    wire new_AGEMA_signal_16750 ;
    wire new_AGEMA_signal_16751 ;
    wire new_AGEMA_signal_16752 ;
    wire new_AGEMA_signal_16753 ;
    wire new_AGEMA_signal_16754 ;
    wire new_AGEMA_signal_16755 ;
    wire new_AGEMA_signal_16756 ;
    wire new_AGEMA_signal_16757 ;
    wire new_AGEMA_signal_16758 ;
    wire new_AGEMA_signal_16759 ;
    wire new_AGEMA_signal_16760 ;
    wire new_AGEMA_signal_16761 ;
    wire new_AGEMA_signal_16762 ;
    wire new_AGEMA_signal_16763 ;
    wire new_AGEMA_signal_16764 ;
    wire new_AGEMA_signal_16765 ;
    wire new_AGEMA_signal_16766 ;
    wire new_AGEMA_signal_16767 ;
    wire new_AGEMA_signal_16768 ;
    wire new_AGEMA_signal_16769 ;
    wire new_AGEMA_signal_16770 ;
    wire new_AGEMA_signal_16771 ;
    wire new_AGEMA_signal_16772 ;
    wire new_AGEMA_signal_16773 ;
    wire new_AGEMA_signal_16774 ;
    wire new_AGEMA_signal_16775 ;
    wire new_AGEMA_signal_16776 ;
    wire new_AGEMA_signal_16777 ;
    wire new_AGEMA_signal_16778 ;
    wire new_AGEMA_signal_16779 ;
    wire new_AGEMA_signal_16780 ;
    wire new_AGEMA_signal_16781 ;
    wire new_AGEMA_signal_16782 ;
    wire new_AGEMA_signal_16783 ;
    wire new_AGEMA_signal_16784 ;
    wire new_AGEMA_signal_16785 ;
    wire new_AGEMA_signal_16786 ;
    wire new_AGEMA_signal_16787 ;
    wire new_AGEMA_signal_16788 ;
    wire new_AGEMA_signal_16789 ;
    wire new_AGEMA_signal_16790 ;
    wire new_AGEMA_signal_16791 ;
    wire new_AGEMA_signal_16792 ;
    wire new_AGEMA_signal_16793 ;
    wire new_AGEMA_signal_16794 ;
    wire new_AGEMA_signal_16795 ;
    wire new_AGEMA_signal_16796 ;
    wire new_AGEMA_signal_16797 ;
    wire new_AGEMA_signal_16798 ;
    wire new_AGEMA_signal_16799 ;
    wire new_AGEMA_signal_16800 ;
    wire new_AGEMA_signal_16801 ;
    wire new_AGEMA_signal_16802 ;
    wire new_AGEMA_signal_16803 ;
    wire new_AGEMA_signal_16804 ;
    wire new_AGEMA_signal_16805 ;
    wire new_AGEMA_signal_16806 ;
    wire new_AGEMA_signal_16807 ;
    wire new_AGEMA_signal_16808 ;
    wire new_AGEMA_signal_16809 ;
    wire new_AGEMA_signal_16810 ;
    wire new_AGEMA_signal_16811 ;
    wire new_AGEMA_signal_16812 ;
    wire new_AGEMA_signal_16813 ;
    wire new_AGEMA_signal_16814 ;
    wire new_AGEMA_signal_16815 ;
    wire new_AGEMA_signal_16816 ;
    wire new_AGEMA_signal_16817 ;
    wire new_AGEMA_signal_16818 ;
    wire new_AGEMA_signal_16819 ;
    wire new_AGEMA_signal_16820 ;
    wire new_AGEMA_signal_16821 ;
    wire new_AGEMA_signal_16822 ;
    wire new_AGEMA_signal_16823 ;
    wire new_AGEMA_signal_16824 ;
    wire new_AGEMA_signal_16825 ;
    wire new_AGEMA_signal_16826 ;
    wire new_AGEMA_signal_16827 ;
    wire new_AGEMA_signal_16828 ;
    wire new_AGEMA_signal_16829 ;
    wire new_AGEMA_signal_16830 ;
    wire new_AGEMA_signal_16831 ;
    wire new_AGEMA_signal_16832 ;
    wire new_AGEMA_signal_16833 ;
    wire new_AGEMA_signal_16834 ;
    wire new_AGEMA_signal_16835 ;
    wire new_AGEMA_signal_16836 ;
    wire new_AGEMA_signal_16837 ;
    wire new_AGEMA_signal_16838 ;
    wire new_AGEMA_signal_16839 ;
    wire new_AGEMA_signal_16840 ;
    wire new_AGEMA_signal_16841 ;
    wire new_AGEMA_signal_16842 ;
    wire new_AGEMA_signal_16843 ;
    wire new_AGEMA_signal_16844 ;
    wire new_AGEMA_signal_16845 ;
    wire new_AGEMA_signal_16846 ;
    wire new_AGEMA_signal_16847 ;
    wire new_AGEMA_signal_16848 ;
    wire new_AGEMA_signal_16849 ;
    wire new_AGEMA_signal_16850 ;
    wire new_AGEMA_signal_16851 ;
    wire new_AGEMA_signal_16852 ;
    wire new_AGEMA_signal_16853 ;
    wire new_AGEMA_signal_16854 ;
    wire new_AGEMA_signal_16855 ;
    wire new_AGEMA_signal_16856 ;
    wire new_AGEMA_signal_16857 ;
    wire new_AGEMA_signal_16858 ;
    wire new_AGEMA_signal_16859 ;
    wire new_AGEMA_signal_16860 ;
    wire new_AGEMA_signal_16861 ;
    wire new_AGEMA_signal_16862 ;
    wire new_AGEMA_signal_16863 ;
    wire new_AGEMA_signal_16864 ;
    wire new_AGEMA_signal_16865 ;
    wire new_AGEMA_signal_16866 ;
    wire new_AGEMA_signal_16867 ;
    wire new_AGEMA_signal_16868 ;
    wire new_AGEMA_signal_16869 ;
    wire new_AGEMA_signal_16870 ;
    wire new_AGEMA_signal_16871 ;
    wire new_AGEMA_signal_16872 ;
    wire new_AGEMA_signal_16873 ;
    wire new_AGEMA_signal_16874 ;
    wire new_AGEMA_signal_16875 ;
    wire new_AGEMA_signal_16876 ;
    wire new_AGEMA_signal_16877 ;
    wire new_AGEMA_signal_16878 ;
    wire new_AGEMA_signal_16879 ;
    wire new_AGEMA_signal_16880 ;
    wire new_AGEMA_signal_16881 ;
    wire new_AGEMA_signal_16882 ;
    wire new_AGEMA_signal_16883 ;
    wire new_AGEMA_signal_16884 ;
    wire new_AGEMA_signal_16885 ;
    wire new_AGEMA_signal_16886 ;
    wire new_AGEMA_signal_16887 ;
    wire new_AGEMA_signal_16888 ;
    wire new_AGEMA_signal_16889 ;
    wire new_AGEMA_signal_16890 ;
    wire new_AGEMA_signal_16891 ;
    wire new_AGEMA_signal_16892 ;
    wire new_AGEMA_signal_16893 ;
    wire new_AGEMA_signal_16894 ;
    wire new_AGEMA_signal_16895 ;
    wire new_AGEMA_signal_16896 ;
    wire new_AGEMA_signal_16897 ;
    wire new_AGEMA_signal_16898 ;
    wire new_AGEMA_signal_16899 ;
    wire new_AGEMA_signal_16900 ;
    wire new_AGEMA_signal_16901 ;
    wire new_AGEMA_signal_16902 ;
    wire new_AGEMA_signal_16903 ;
    wire new_AGEMA_signal_16904 ;
    wire new_AGEMA_signal_16905 ;
    wire new_AGEMA_signal_16906 ;
    wire new_AGEMA_signal_16907 ;
    wire new_AGEMA_signal_16908 ;
    wire new_AGEMA_signal_16909 ;
    wire new_AGEMA_signal_16910 ;
    wire new_AGEMA_signal_16911 ;
    wire new_AGEMA_signal_16912 ;
    wire new_AGEMA_signal_16913 ;
    wire new_AGEMA_signal_16914 ;
    wire new_AGEMA_signal_16915 ;
    wire new_AGEMA_signal_16916 ;
    wire new_AGEMA_signal_16917 ;
    wire new_AGEMA_signal_16918 ;
    wire new_AGEMA_signal_16919 ;
    wire new_AGEMA_signal_16920 ;
    wire new_AGEMA_signal_16921 ;
    wire new_AGEMA_signal_16922 ;
    wire new_AGEMA_signal_16923 ;
    wire new_AGEMA_signal_16924 ;
    wire new_AGEMA_signal_16925 ;
    wire new_AGEMA_signal_16926 ;
    wire new_AGEMA_signal_16927 ;
    wire new_AGEMA_signal_16928 ;
    wire new_AGEMA_signal_16929 ;
    wire new_AGEMA_signal_16930 ;
    wire new_AGEMA_signal_16931 ;
    wire new_AGEMA_signal_16932 ;
    wire new_AGEMA_signal_16933 ;
    wire new_AGEMA_signal_16934 ;
    wire new_AGEMA_signal_16935 ;
    wire new_AGEMA_signal_16936 ;
    wire new_AGEMA_signal_16937 ;
    wire new_AGEMA_signal_16938 ;
    wire new_AGEMA_signal_16939 ;
    wire new_AGEMA_signal_16940 ;
    wire new_AGEMA_signal_16941 ;
    wire new_AGEMA_signal_16942 ;
    wire new_AGEMA_signal_16943 ;
    wire new_AGEMA_signal_16944 ;
    wire new_AGEMA_signal_16945 ;
    wire new_AGEMA_signal_16946 ;
    wire new_AGEMA_signal_16947 ;
    wire new_AGEMA_signal_16948 ;
    wire new_AGEMA_signal_16949 ;
    wire new_AGEMA_signal_16950 ;
    wire new_AGEMA_signal_16951 ;
    wire new_AGEMA_signal_16952 ;
    wire new_AGEMA_signal_16953 ;
    wire new_AGEMA_signal_16954 ;
    wire new_AGEMA_signal_16955 ;
    wire new_AGEMA_signal_16956 ;
    wire new_AGEMA_signal_16957 ;
    wire new_AGEMA_signal_16958 ;
    wire new_AGEMA_signal_16959 ;
    wire new_AGEMA_signal_16960 ;
    wire new_AGEMA_signal_16961 ;
    wire new_AGEMA_signal_16962 ;
    wire new_AGEMA_signal_16963 ;
    wire new_AGEMA_signal_16964 ;
    wire new_AGEMA_signal_16965 ;
    wire new_AGEMA_signal_16966 ;
    wire new_AGEMA_signal_16967 ;
    wire new_AGEMA_signal_16968 ;
    wire new_AGEMA_signal_16969 ;
    wire new_AGEMA_signal_16970 ;
    wire new_AGEMA_signal_16971 ;
    wire new_AGEMA_signal_16972 ;
    wire new_AGEMA_signal_16973 ;
    wire new_AGEMA_signal_16974 ;
    wire new_AGEMA_signal_16975 ;
    wire new_AGEMA_signal_16976 ;
    wire new_AGEMA_signal_16977 ;
    wire new_AGEMA_signal_16978 ;
    wire new_AGEMA_signal_16979 ;
    wire new_AGEMA_signal_16980 ;
    wire new_AGEMA_signal_16981 ;
    wire new_AGEMA_signal_16982 ;
    wire new_AGEMA_signal_16983 ;
    wire new_AGEMA_signal_16984 ;
    wire new_AGEMA_signal_16985 ;
    wire new_AGEMA_signal_16986 ;
    wire new_AGEMA_signal_16987 ;
    wire new_AGEMA_signal_16988 ;
    wire new_AGEMA_signal_16989 ;
    wire new_AGEMA_signal_16990 ;
    wire new_AGEMA_signal_16991 ;
    wire new_AGEMA_signal_16992 ;
    wire new_AGEMA_signal_16993 ;
    wire new_AGEMA_signal_16994 ;
    wire new_AGEMA_signal_16995 ;
    wire new_AGEMA_signal_16996 ;
    wire new_AGEMA_signal_16997 ;
    wire new_AGEMA_signal_16998 ;
    wire new_AGEMA_signal_16999 ;
    wire new_AGEMA_signal_17000 ;
    wire new_AGEMA_signal_17001 ;
    wire new_AGEMA_signal_17002 ;
    wire new_AGEMA_signal_17003 ;
    wire new_AGEMA_signal_17004 ;
    wire new_AGEMA_signal_17005 ;
    wire new_AGEMA_signal_17006 ;
    wire new_AGEMA_signal_17007 ;
    wire new_AGEMA_signal_17008 ;
    wire new_AGEMA_signal_17009 ;
    wire new_AGEMA_signal_17010 ;
    wire new_AGEMA_signal_17011 ;
    wire new_AGEMA_signal_17012 ;
    wire new_AGEMA_signal_17013 ;
    wire new_AGEMA_signal_17014 ;
    wire new_AGEMA_signal_17015 ;
    wire new_AGEMA_signal_17016 ;
    wire new_AGEMA_signal_17017 ;
    wire new_AGEMA_signal_17018 ;
    wire new_AGEMA_signal_17019 ;
    wire new_AGEMA_signal_17020 ;
    wire new_AGEMA_signal_17021 ;
    wire new_AGEMA_signal_17022 ;
    wire new_AGEMA_signal_17023 ;
    wire new_AGEMA_signal_17024 ;
    wire new_AGEMA_signal_17025 ;
    wire new_AGEMA_signal_17026 ;
    wire new_AGEMA_signal_17027 ;
    wire new_AGEMA_signal_17028 ;
    wire new_AGEMA_signal_17029 ;
    wire new_AGEMA_signal_17030 ;
    wire new_AGEMA_signal_17031 ;
    wire new_AGEMA_signal_17032 ;
    wire new_AGEMA_signal_17033 ;
    wire new_AGEMA_signal_17034 ;
    wire new_AGEMA_signal_17035 ;
    wire new_AGEMA_signal_17036 ;
    wire new_AGEMA_signal_17037 ;
    wire new_AGEMA_signal_17038 ;
    wire new_AGEMA_signal_17039 ;
    wire new_AGEMA_signal_17040 ;
    wire new_AGEMA_signal_17041 ;
    wire new_AGEMA_signal_17042 ;
    wire new_AGEMA_signal_17043 ;
    wire new_AGEMA_signal_17044 ;
    wire new_AGEMA_signal_17045 ;
    wire new_AGEMA_signal_17046 ;
    wire new_AGEMA_signal_17047 ;
    wire new_AGEMA_signal_17048 ;
    wire new_AGEMA_signal_17049 ;
    wire new_AGEMA_signal_17050 ;
    wire new_AGEMA_signal_17051 ;
    wire new_AGEMA_signal_17052 ;
    wire new_AGEMA_signal_17053 ;
    wire new_AGEMA_signal_17054 ;
    wire new_AGEMA_signal_17055 ;
    wire new_AGEMA_signal_17056 ;
    wire new_AGEMA_signal_17057 ;
    wire new_AGEMA_signal_17058 ;
    wire new_AGEMA_signal_17059 ;
    wire new_AGEMA_signal_17060 ;
    wire new_AGEMA_signal_17061 ;
    wire new_AGEMA_signal_17062 ;
    wire new_AGEMA_signal_17063 ;
    wire new_AGEMA_signal_17064 ;
    wire new_AGEMA_signal_17065 ;
    wire new_AGEMA_signal_17066 ;
    wire new_AGEMA_signal_17067 ;
    wire new_AGEMA_signal_17068 ;
    wire new_AGEMA_signal_17069 ;
    wire new_AGEMA_signal_17070 ;
    wire new_AGEMA_signal_17071 ;
    wire new_AGEMA_signal_17072 ;
    wire new_AGEMA_signal_17073 ;
    wire new_AGEMA_signal_17074 ;
    wire new_AGEMA_signal_17075 ;
    wire new_AGEMA_signal_17076 ;
    wire new_AGEMA_signal_17077 ;
    wire new_AGEMA_signal_17078 ;
    wire new_AGEMA_signal_17079 ;
    wire new_AGEMA_signal_17080 ;
    wire new_AGEMA_signal_17081 ;
    wire new_AGEMA_signal_17082 ;
    wire new_AGEMA_signal_17083 ;
    wire new_AGEMA_signal_17084 ;
    wire new_AGEMA_signal_17085 ;
    wire new_AGEMA_signal_17086 ;
    wire new_AGEMA_signal_17087 ;
    wire new_AGEMA_signal_17088 ;
    wire new_AGEMA_signal_17089 ;
    wire new_AGEMA_signal_17090 ;
    wire new_AGEMA_signal_17091 ;
    wire new_AGEMA_signal_17092 ;
    wire new_AGEMA_signal_17093 ;
    wire new_AGEMA_signal_17094 ;
    wire new_AGEMA_signal_17095 ;
    wire new_AGEMA_signal_17096 ;
    wire new_AGEMA_signal_17097 ;
    wire new_AGEMA_signal_17098 ;
    wire new_AGEMA_signal_17099 ;
    wire new_AGEMA_signal_17100 ;
    wire new_AGEMA_signal_17101 ;
    wire new_AGEMA_signal_17102 ;
    wire new_AGEMA_signal_17103 ;
    wire new_AGEMA_signal_17104 ;
    wire new_AGEMA_signal_17105 ;
    wire new_AGEMA_signal_17106 ;
    wire new_AGEMA_signal_17107 ;
    wire new_AGEMA_signal_17108 ;
    wire new_AGEMA_signal_17109 ;
    wire new_AGEMA_signal_17110 ;
    wire new_AGEMA_signal_17111 ;
    wire new_AGEMA_signal_17112 ;
    wire new_AGEMA_signal_17113 ;
    wire new_AGEMA_signal_17114 ;
    wire new_AGEMA_signal_17115 ;
    wire new_AGEMA_signal_17116 ;
    wire new_AGEMA_signal_17117 ;
    wire new_AGEMA_signal_17118 ;
    wire new_AGEMA_signal_17119 ;
    wire new_AGEMA_signal_17120 ;
    wire new_AGEMA_signal_17121 ;
    wire new_AGEMA_signal_17122 ;
    wire new_AGEMA_signal_17123 ;
    wire new_AGEMA_signal_17124 ;
    wire new_AGEMA_signal_17125 ;
    wire new_AGEMA_signal_17126 ;
    wire new_AGEMA_signal_17127 ;
    wire new_AGEMA_signal_17128 ;
    wire new_AGEMA_signal_17129 ;
    wire new_AGEMA_signal_17130 ;
    wire new_AGEMA_signal_17131 ;
    wire new_AGEMA_signal_17132 ;
    wire new_AGEMA_signal_17133 ;
    wire new_AGEMA_signal_17134 ;
    wire new_AGEMA_signal_17135 ;
    wire new_AGEMA_signal_17136 ;
    wire new_AGEMA_signal_17137 ;
    wire new_AGEMA_signal_17138 ;
    wire new_AGEMA_signal_17139 ;
    wire new_AGEMA_signal_17140 ;
    wire new_AGEMA_signal_17141 ;
    wire new_AGEMA_signal_17142 ;
    wire new_AGEMA_signal_17143 ;
    wire new_AGEMA_signal_17144 ;
    wire new_AGEMA_signal_17145 ;
    wire new_AGEMA_signal_17146 ;
    wire new_AGEMA_signal_17147 ;
    wire new_AGEMA_signal_17148 ;
    wire new_AGEMA_signal_17149 ;
    wire new_AGEMA_signal_17150 ;
    wire new_AGEMA_signal_17151 ;
    wire new_AGEMA_signal_17152 ;
    wire new_AGEMA_signal_17153 ;
    wire new_AGEMA_signal_17154 ;
    wire new_AGEMA_signal_17155 ;
    wire new_AGEMA_signal_17156 ;
    wire new_AGEMA_signal_17157 ;
    wire new_AGEMA_signal_17158 ;
    wire new_AGEMA_signal_17159 ;
    wire new_AGEMA_signal_17160 ;
    wire new_AGEMA_signal_17161 ;
    wire new_AGEMA_signal_17162 ;
    wire new_AGEMA_signal_17163 ;
    wire new_AGEMA_signal_17164 ;
    wire new_AGEMA_signal_17165 ;
    wire new_AGEMA_signal_17166 ;
    wire new_AGEMA_signal_17167 ;
    wire new_AGEMA_signal_17168 ;
    wire new_AGEMA_signal_17169 ;
    wire new_AGEMA_signal_17170 ;
    wire new_AGEMA_signal_17171 ;
    wire new_AGEMA_signal_17172 ;
    wire new_AGEMA_signal_17173 ;
    wire new_AGEMA_signal_17174 ;
    wire new_AGEMA_signal_17175 ;
    wire new_AGEMA_signal_17176 ;
    wire new_AGEMA_signal_17177 ;
    wire new_AGEMA_signal_17178 ;
    wire new_AGEMA_signal_17179 ;
    wire new_AGEMA_signal_17180 ;
    wire new_AGEMA_signal_17181 ;
    wire new_AGEMA_signal_17182 ;
    wire new_AGEMA_signal_17183 ;
    wire new_AGEMA_signal_17184 ;
    wire new_AGEMA_signal_17185 ;
    wire new_AGEMA_signal_17186 ;
    wire new_AGEMA_signal_17187 ;
    wire new_AGEMA_signal_17188 ;
    wire new_AGEMA_signal_17189 ;
    wire new_AGEMA_signal_17190 ;
    wire new_AGEMA_signal_17191 ;
    wire new_AGEMA_signal_17192 ;
    wire new_AGEMA_signal_17193 ;
    wire new_AGEMA_signal_17194 ;
    wire new_AGEMA_signal_17195 ;
    wire new_AGEMA_signal_17196 ;
    wire new_AGEMA_signal_17197 ;
    wire new_AGEMA_signal_17198 ;
    wire new_AGEMA_signal_17199 ;
    wire new_AGEMA_signal_17200 ;
    wire new_AGEMA_signal_17201 ;
    wire new_AGEMA_signal_17202 ;
    wire new_AGEMA_signal_17203 ;
    wire new_AGEMA_signal_17204 ;
    wire new_AGEMA_signal_17205 ;
    wire new_AGEMA_signal_17206 ;
    wire new_AGEMA_signal_17207 ;
    wire new_AGEMA_signal_17208 ;
    wire new_AGEMA_signal_17209 ;
    wire new_AGEMA_signal_17210 ;
    wire new_AGEMA_signal_17211 ;
    wire new_AGEMA_signal_17212 ;
    wire new_AGEMA_signal_17213 ;
    wire new_AGEMA_signal_17214 ;
    wire new_AGEMA_signal_17215 ;
    wire new_AGEMA_signal_17216 ;
    wire new_AGEMA_signal_17217 ;
    wire new_AGEMA_signal_17218 ;
    wire new_AGEMA_signal_17219 ;
    wire new_AGEMA_signal_17220 ;
    wire new_AGEMA_signal_17221 ;
    wire new_AGEMA_signal_17222 ;
    wire new_AGEMA_signal_17223 ;
    wire new_AGEMA_signal_17224 ;
    wire new_AGEMA_signal_17225 ;
    wire new_AGEMA_signal_17226 ;
    wire new_AGEMA_signal_17227 ;
    wire new_AGEMA_signal_17228 ;
    wire new_AGEMA_signal_17229 ;
    wire new_AGEMA_signal_17230 ;
    wire new_AGEMA_signal_17231 ;
    wire new_AGEMA_signal_17232 ;
    wire new_AGEMA_signal_17233 ;
    wire new_AGEMA_signal_17234 ;
    wire new_AGEMA_signal_17235 ;
    wire new_AGEMA_signal_17236 ;
    wire new_AGEMA_signal_17237 ;
    wire new_AGEMA_signal_17238 ;
    wire new_AGEMA_signal_17239 ;
    wire new_AGEMA_signal_17240 ;
    wire new_AGEMA_signal_17241 ;
    wire new_AGEMA_signal_17242 ;
    wire new_AGEMA_signal_17243 ;
    wire new_AGEMA_signal_17244 ;
    wire new_AGEMA_signal_17245 ;
    wire new_AGEMA_signal_17246 ;
    wire new_AGEMA_signal_17247 ;
    wire new_AGEMA_signal_17248 ;
    wire new_AGEMA_signal_17249 ;
    wire new_AGEMA_signal_17250 ;
    wire new_AGEMA_signal_17251 ;
    wire new_AGEMA_signal_17252 ;
    wire new_AGEMA_signal_17253 ;
    wire new_AGEMA_signal_17254 ;
    wire new_AGEMA_signal_17255 ;
    wire new_AGEMA_signal_17256 ;
    wire new_AGEMA_signal_17257 ;
    wire new_AGEMA_signal_17258 ;
    wire new_AGEMA_signal_17259 ;
    wire new_AGEMA_signal_17260 ;
    wire new_AGEMA_signal_17261 ;
    wire new_AGEMA_signal_17262 ;
    wire new_AGEMA_signal_17263 ;
    wire new_AGEMA_signal_17264 ;
    wire new_AGEMA_signal_17265 ;
    wire new_AGEMA_signal_17266 ;
    wire new_AGEMA_signal_17267 ;
    wire new_AGEMA_signal_17268 ;
    wire new_AGEMA_signal_17269 ;
    wire new_AGEMA_signal_17270 ;
    wire new_AGEMA_signal_17271 ;
    wire new_AGEMA_signal_17272 ;
    wire new_AGEMA_signal_17273 ;
    wire new_AGEMA_signal_17274 ;
    wire new_AGEMA_signal_17275 ;
    wire new_AGEMA_signal_17276 ;
    wire new_AGEMA_signal_17277 ;
    wire new_AGEMA_signal_17278 ;
    wire new_AGEMA_signal_17279 ;
    wire new_AGEMA_signal_17280 ;
    wire new_AGEMA_signal_17281 ;
    wire new_AGEMA_signal_17282 ;
    wire new_AGEMA_signal_17283 ;
    wire new_AGEMA_signal_17284 ;
    wire new_AGEMA_signal_17285 ;
    wire new_AGEMA_signal_17286 ;
    wire new_AGEMA_signal_17287 ;
    wire new_AGEMA_signal_17288 ;
    wire new_AGEMA_signal_17289 ;
    wire new_AGEMA_signal_17290 ;
    wire new_AGEMA_signal_17291 ;
    wire new_AGEMA_signal_17292 ;
    wire new_AGEMA_signal_17293 ;
    wire new_AGEMA_signal_17294 ;
    wire new_AGEMA_signal_17295 ;
    wire new_AGEMA_signal_17296 ;
    wire new_AGEMA_signal_17297 ;
    wire new_AGEMA_signal_17298 ;
    wire new_AGEMA_signal_17299 ;
    wire new_AGEMA_signal_17300 ;
    wire new_AGEMA_signal_17301 ;
    wire new_AGEMA_signal_17302 ;
    wire new_AGEMA_signal_17303 ;
    wire new_AGEMA_signal_17304 ;
    wire new_AGEMA_signal_17305 ;
    wire new_AGEMA_signal_17306 ;
    wire new_AGEMA_signal_17307 ;
    wire new_AGEMA_signal_17308 ;
    wire new_AGEMA_signal_17309 ;
    wire new_AGEMA_signal_17310 ;
    wire new_AGEMA_signal_17311 ;
    wire new_AGEMA_signal_17312 ;
    wire new_AGEMA_signal_17313 ;
    wire new_AGEMA_signal_17314 ;
    wire new_AGEMA_signal_17315 ;
    wire new_AGEMA_signal_17316 ;
    wire new_AGEMA_signal_17317 ;
    wire new_AGEMA_signal_17318 ;
    wire new_AGEMA_signal_17319 ;
    wire new_AGEMA_signal_17320 ;
    wire new_AGEMA_signal_17321 ;
    wire new_AGEMA_signal_17322 ;
    wire new_AGEMA_signal_17323 ;
    wire new_AGEMA_signal_17324 ;
    wire new_AGEMA_signal_17325 ;
    wire new_AGEMA_signal_17326 ;
    wire new_AGEMA_signal_17327 ;
    wire new_AGEMA_signal_17328 ;
    wire new_AGEMA_signal_17329 ;
    wire new_AGEMA_signal_17330 ;
    wire new_AGEMA_signal_17331 ;
    wire new_AGEMA_signal_17332 ;
    wire new_AGEMA_signal_17333 ;
    wire new_AGEMA_signal_17334 ;
    wire new_AGEMA_signal_17335 ;
    wire new_AGEMA_signal_17336 ;
    wire new_AGEMA_signal_17337 ;
    wire new_AGEMA_signal_17338 ;
    wire new_AGEMA_signal_17339 ;
    wire new_AGEMA_signal_17340 ;
    wire new_AGEMA_signal_17341 ;
    wire new_AGEMA_signal_17342 ;
    wire new_AGEMA_signal_17343 ;
    wire new_AGEMA_signal_17344 ;
    wire new_AGEMA_signal_17345 ;
    wire new_AGEMA_signal_17346 ;
    wire new_AGEMA_signal_17347 ;
    wire new_AGEMA_signal_17348 ;
    wire new_AGEMA_signal_17349 ;
    wire new_AGEMA_signal_17350 ;
    wire new_AGEMA_signal_17351 ;
    wire new_AGEMA_signal_17352 ;
    wire new_AGEMA_signal_17353 ;
    wire new_AGEMA_signal_17354 ;
    wire new_AGEMA_signal_17355 ;
    wire new_AGEMA_signal_17356 ;
    wire new_AGEMA_signal_17357 ;
    wire new_AGEMA_signal_17358 ;
    wire new_AGEMA_signal_17359 ;
    wire new_AGEMA_signal_17360 ;
    wire new_AGEMA_signal_17361 ;
    wire new_AGEMA_signal_17362 ;
    wire new_AGEMA_signal_17363 ;
    wire new_AGEMA_signal_17364 ;
    wire new_AGEMA_signal_17365 ;
    wire new_AGEMA_signal_17366 ;
    wire new_AGEMA_signal_17367 ;
    wire new_AGEMA_signal_17368 ;
    wire new_AGEMA_signal_17369 ;
    wire new_AGEMA_signal_17370 ;
    wire new_AGEMA_signal_17371 ;
    wire new_AGEMA_signal_17372 ;
    wire new_AGEMA_signal_17373 ;
    wire new_AGEMA_signal_17374 ;
    wire new_AGEMA_signal_17375 ;
    wire new_AGEMA_signal_17376 ;
    wire new_AGEMA_signal_17377 ;
    wire new_AGEMA_signal_17378 ;
    wire new_AGEMA_signal_17379 ;
    wire new_AGEMA_signal_17380 ;
    wire new_AGEMA_signal_17381 ;
    wire new_AGEMA_signal_17382 ;
    wire new_AGEMA_signal_17383 ;
    wire new_AGEMA_signal_17384 ;
    wire new_AGEMA_signal_17385 ;
    wire new_AGEMA_signal_17386 ;
    wire new_AGEMA_signal_17387 ;
    wire new_AGEMA_signal_17388 ;
    wire new_AGEMA_signal_17389 ;
    wire new_AGEMA_signal_17390 ;
    wire new_AGEMA_signal_17391 ;
    wire new_AGEMA_signal_17392 ;
    wire new_AGEMA_signal_17393 ;
    wire new_AGEMA_signal_17394 ;
    wire new_AGEMA_signal_17395 ;
    wire new_AGEMA_signal_17396 ;
    wire new_AGEMA_signal_17397 ;
    wire new_AGEMA_signal_17398 ;
    wire new_AGEMA_signal_17399 ;
    wire new_AGEMA_signal_17400 ;
    wire new_AGEMA_signal_17401 ;
    wire new_AGEMA_signal_17402 ;
    wire new_AGEMA_signal_17403 ;
    wire new_AGEMA_signal_17404 ;
    wire new_AGEMA_signal_17405 ;
    wire new_AGEMA_signal_17406 ;
    wire new_AGEMA_signal_17407 ;
    wire new_AGEMA_signal_17408 ;
    wire new_AGEMA_signal_17409 ;
    wire new_AGEMA_signal_17410 ;
    wire new_AGEMA_signal_17411 ;
    wire new_AGEMA_signal_17412 ;
    wire new_AGEMA_signal_17413 ;
    wire new_AGEMA_signal_17414 ;
    wire new_AGEMA_signal_17415 ;
    wire new_AGEMA_signal_17416 ;
    wire new_AGEMA_signal_17417 ;
    wire new_AGEMA_signal_17418 ;
    wire new_AGEMA_signal_17419 ;
    wire new_AGEMA_signal_17420 ;
    wire new_AGEMA_signal_17421 ;
    wire new_AGEMA_signal_17422 ;
    wire new_AGEMA_signal_17423 ;
    wire new_AGEMA_signal_17424 ;
    wire new_AGEMA_signal_17425 ;
    wire new_AGEMA_signal_17426 ;
    wire new_AGEMA_signal_17427 ;
    wire new_AGEMA_signal_17428 ;
    wire new_AGEMA_signal_17429 ;
    wire new_AGEMA_signal_17430 ;
    wire new_AGEMA_signal_17431 ;
    wire new_AGEMA_signal_17432 ;
    wire new_AGEMA_signal_17433 ;
    wire new_AGEMA_signal_17434 ;
    wire new_AGEMA_signal_17435 ;
    wire new_AGEMA_signal_17436 ;
    wire new_AGEMA_signal_17437 ;
    wire new_AGEMA_signal_17438 ;
    wire new_AGEMA_signal_17439 ;
    wire new_AGEMA_signal_17440 ;
    wire new_AGEMA_signal_17441 ;
    wire new_AGEMA_signal_17442 ;
    wire new_AGEMA_signal_17443 ;
    wire new_AGEMA_signal_17444 ;
    wire new_AGEMA_signal_17445 ;
    wire new_AGEMA_signal_17446 ;
    wire new_AGEMA_signal_17447 ;
    wire new_AGEMA_signal_17448 ;
    wire new_AGEMA_signal_17449 ;
    wire new_AGEMA_signal_17450 ;
    wire new_AGEMA_signal_17451 ;
    wire new_AGEMA_signal_17452 ;
    wire new_AGEMA_signal_17453 ;
    wire new_AGEMA_signal_17454 ;
    wire new_AGEMA_signal_17455 ;
    wire new_AGEMA_signal_17456 ;
    wire new_AGEMA_signal_17457 ;
    wire new_AGEMA_signal_17458 ;
    wire new_AGEMA_signal_17459 ;
    wire new_AGEMA_signal_17460 ;
    wire new_AGEMA_signal_17461 ;
    wire new_AGEMA_signal_17462 ;
    wire new_AGEMA_signal_17463 ;
    wire new_AGEMA_signal_17464 ;
    wire new_AGEMA_signal_17465 ;
    wire new_AGEMA_signal_17466 ;
    wire new_AGEMA_signal_17467 ;
    wire new_AGEMA_signal_17468 ;
    wire new_AGEMA_signal_17469 ;
    wire new_AGEMA_signal_17470 ;
    wire new_AGEMA_signal_17471 ;
    wire new_AGEMA_signal_17472 ;
    wire new_AGEMA_signal_17473 ;
    wire new_AGEMA_signal_17474 ;
    wire new_AGEMA_signal_17475 ;
    wire new_AGEMA_signal_17476 ;
    wire new_AGEMA_signal_17477 ;
    wire new_AGEMA_signal_17478 ;
    wire new_AGEMA_signal_17479 ;
    wire new_AGEMA_signal_17480 ;
    wire new_AGEMA_signal_17481 ;
    wire new_AGEMA_signal_17482 ;
    wire new_AGEMA_signal_17483 ;
    wire new_AGEMA_signal_17484 ;
    wire new_AGEMA_signal_17485 ;
    wire new_AGEMA_signal_17486 ;
    wire new_AGEMA_signal_17487 ;
    wire new_AGEMA_signal_17488 ;
    wire new_AGEMA_signal_17489 ;
    wire new_AGEMA_signal_17490 ;
    wire new_AGEMA_signal_17491 ;
    wire new_AGEMA_signal_17492 ;
    wire new_AGEMA_signal_17493 ;
    wire new_AGEMA_signal_17494 ;
    wire new_AGEMA_signal_17495 ;
    wire new_AGEMA_signal_17496 ;
    wire new_AGEMA_signal_17497 ;
    wire new_AGEMA_signal_17498 ;
    wire new_AGEMA_signal_17499 ;
    wire new_AGEMA_signal_17500 ;
    wire new_AGEMA_signal_17501 ;
    wire new_AGEMA_signal_17502 ;
    wire new_AGEMA_signal_17503 ;
    wire new_AGEMA_signal_17504 ;
    wire new_AGEMA_signal_17505 ;
    wire new_AGEMA_signal_17506 ;
    wire new_AGEMA_signal_17507 ;
    wire new_AGEMA_signal_17508 ;
    wire new_AGEMA_signal_17509 ;
    wire new_AGEMA_signal_17510 ;
    wire new_AGEMA_signal_17511 ;
    wire new_AGEMA_signal_17512 ;
    wire new_AGEMA_signal_17513 ;
    wire new_AGEMA_signal_17514 ;
    wire new_AGEMA_signal_17515 ;
    wire new_AGEMA_signal_17516 ;
    wire new_AGEMA_signal_17517 ;
    wire new_AGEMA_signal_17518 ;
    wire new_AGEMA_signal_17519 ;
    wire new_AGEMA_signal_17520 ;
    wire new_AGEMA_signal_17521 ;
    wire new_AGEMA_signal_17522 ;
    wire new_AGEMA_signal_17523 ;
    wire new_AGEMA_signal_17524 ;
    wire new_AGEMA_signal_17525 ;
    wire new_AGEMA_signal_17526 ;
    wire new_AGEMA_signal_17527 ;
    wire new_AGEMA_signal_17528 ;
    wire new_AGEMA_signal_17529 ;
    wire new_AGEMA_signal_17530 ;
    wire new_AGEMA_signal_17531 ;
    wire new_AGEMA_signal_17532 ;
    wire new_AGEMA_signal_17533 ;
    wire new_AGEMA_signal_17534 ;
    wire new_AGEMA_signal_17535 ;
    wire new_AGEMA_signal_17536 ;
    wire new_AGEMA_signal_17537 ;
    wire new_AGEMA_signal_17538 ;
    wire new_AGEMA_signal_17539 ;
    wire new_AGEMA_signal_17540 ;
    wire new_AGEMA_signal_17541 ;
    wire new_AGEMA_signal_17542 ;
    wire new_AGEMA_signal_17543 ;
    wire new_AGEMA_signal_17544 ;
    wire new_AGEMA_signal_17545 ;
    wire new_AGEMA_signal_17546 ;
    wire new_AGEMA_signal_17547 ;
    wire new_AGEMA_signal_17548 ;
    wire new_AGEMA_signal_17549 ;
    wire new_AGEMA_signal_17550 ;
    wire new_AGEMA_signal_17551 ;
    wire new_AGEMA_signal_17552 ;
    wire new_AGEMA_signal_17553 ;
    wire new_AGEMA_signal_17554 ;
    wire new_AGEMA_signal_17555 ;
    wire new_AGEMA_signal_17556 ;
    wire new_AGEMA_signal_17557 ;
    wire new_AGEMA_signal_17558 ;
    wire new_AGEMA_signal_17559 ;
    wire new_AGEMA_signal_17560 ;
    wire new_AGEMA_signal_17561 ;
    wire new_AGEMA_signal_17562 ;
    wire new_AGEMA_signal_17563 ;
    wire new_AGEMA_signal_17564 ;
    wire new_AGEMA_signal_17565 ;
    wire new_AGEMA_signal_17566 ;
    wire new_AGEMA_signal_17567 ;
    wire new_AGEMA_signal_17568 ;
    wire new_AGEMA_signal_17569 ;
    wire new_AGEMA_signal_17570 ;
    wire new_AGEMA_signal_17571 ;
    wire new_AGEMA_signal_17572 ;
    wire new_AGEMA_signal_17573 ;
    wire new_AGEMA_signal_17574 ;
    wire new_AGEMA_signal_17575 ;
    wire new_AGEMA_signal_17576 ;
    wire new_AGEMA_signal_17577 ;
    wire new_AGEMA_signal_17578 ;
    wire new_AGEMA_signal_17579 ;
    wire new_AGEMA_signal_17580 ;
    wire new_AGEMA_signal_17581 ;
    wire new_AGEMA_signal_17582 ;
    wire new_AGEMA_signal_17583 ;
    wire new_AGEMA_signal_17584 ;
    wire new_AGEMA_signal_17585 ;
    wire new_AGEMA_signal_17586 ;
    wire new_AGEMA_signal_17587 ;
    wire new_AGEMA_signal_17588 ;
    wire new_AGEMA_signal_17589 ;
    wire new_AGEMA_signal_17590 ;
    wire new_AGEMA_signal_17591 ;
    wire new_AGEMA_signal_17592 ;
    wire new_AGEMA_signal_17593 ;
    wire new_AGEMA_signal_17594 ;
    wire new_AGEMA_signal_17595 ;
    wire new_AGEMA_signal_17596 ;
    wire new_AGEMA_signal_17597 ;
    wire new_AGEMA_signal_17598 ;
    wire new_AGEMA_signal_17599 ;
    wire new_AGEMA_signal_17600 ;
    wire new_AGEMA_signal_17601 ;
    wire new_AGEMA_signal_17602 ;
    wire new_AGEMA_signal_17603 ;
    wire new_AGEMA_signal_17604 ;
    wire new_AGEMA_signal_17605 ;
    wire new_AGEMA_signal_17606 ;
    wire new_AGEMA_signal_17607 ;
    wire new_AGEMA_signal_17608 ;
    wire new_AGEMA_signal_17609 ;
    wire new_AGEMA_signal_17610 ;
    wire new_AGEMA_signal_17611 ;
    wire new_AGEMA_signal_17612 ;
    wire new_AGEMA_signal_17613 ;
    wire new_AGEMA_signal_17614 ;
    wire new_AGEMA_signal_17615 ;
    wire new_AGEMA_signal_17616 ;
    wire new_AGEMA_signal_17617 ;
    wire new_AGEMA_signal_17618 ;
    wire new_AGEMA_signal_17619 ;
    wire new_AGEMA_signal_17620 ;
    wire new_AGEMA_signal_17621 ;
    wire new_AGEMA_signal_17622 ;
    wire new_AGEMA_signal_17623 ;
    wire new_AGEMA_signal_17624 ;
    wire new_AGEMA_signal_17625 ;
    wire new_AGEMA_signal_17626 ;
    wire new_AGEMA_signal_17627 ;
    wire new_AGEMA_signal_17628 ;
    wire new_AGEMA_signal_17629 ;
    wire new_AGEMA_signal_17630 ;
    wire new_AGEMA_signal_17631 ;
    wire new_AGEMA_signal_17632 ;
    wire new_AGEMA_signal_17633 ;
    wire new_AGEMA_signal_17634 ;
    wire new_AGEMA_signal_17635 ;
    wire new_AGEMA_signal_17636 ;
    wire new_AGEMA_signal_17637 ;
    wire new_AGEMA_signal_17638 ;
    wire new_AGEMA_signal_17639 ;
    wire new_AGEMA_signal_17640 ;
    wire new_AGEMA_signal_17641 ;
    wire new_AGEMA_signal_17642 ;
    wire new_AGEMA_signal_17643 ;
    wire new_AGEMA_signal_17644 ;
    wire new_AGEMA_signal_17645 ;
    wire new_AGEMA_signal_17646 ;
    wire new_AGEMA_signal_17647 ;
    wire new_AGEMA_signal_17648 ;
    wire new_AGEMA_signal_17649 ;
    wire new_AGEMA_signal_17650 ;
    wire new_AGEMA_signal_17651 ;
    wire new_AGEMA_signal_17652 ;
    wire new_AGEMA_signal_17653 ;
    wire new_AGEMA_signal_17654 ;
    wire new_AGEMA_signal_17655 ;
    wire new_AGEMA_signal_17656 ;
    wire new_AGEMA_signal_17657 ;
    wire new_AGEMA_signal_17658 ;
    wire new_AGEMA_signal_17659 ;
    wire new_AGEMA_signal_17660 ;
    wire new_AGEMA_signal_17661 ;
    wire new_AGEMA_signal_17662 ;
    wire new_AGEMA_signal_17663 ;
    wire new_AGEMA_signal_17664 ;
    wire new_AGEMA_signal_17665 ;
    wire new_AGEMA_signal_17666 ;
    wire new_AGEMA_signal_17667 ;
    wire new_AGEMA_signal_17668 ;
    wire new_AGEMA_signal_17669 ;
    wire new_AGEMA_signal_17670 ;
    wire new_AGEMA_signal_17671 ;
    wire new_AGEMA_signal_17672 ;
    wire new_AGEMA_signal_17673 ;
    wire new_AGEMA_signal_17674 ;
    wire new_AGEMA_signal_17675 ;
    wire new_AGEMA_signal_17676 ;
    wire new_AGEMA_signal_17677 ;
    wire new_AGEMA_signal_17678 ;
    wire new_AGEMA_signal_17679 ;
    wire new_AGEMA_signal_17680 ;
    wire new_AGEMA_signal_17681 ;
    wire new_AGEMA_signal_17682 ;
    wire new_AGEMA_signal_17683 ;
    wire new_AGEMA_signal_17684 ;
    wire new_AGEMA_signal_17685 ;
    wire new_AGEMA_signal_17686 ;
    wire new_AGEMA_signal_17687 ;
    wire new_AGEMA_signal_17688 ;
    wire new_AGEMA_signal_17689 ;
    wire new_AGEMA_signal_17690 ;
    wire new_AGEMA_signal_17691 ;
    wire new_AGEMA_signal_17692 ;
    wire new_AGEMA_signal_17693 ;
    wire new_AGEMA_signal_17694 ;
    wire new_AGEMA_signal_17695 ;
    wire new_AGEMA_signal_17696 ;
    wire new_AGEMA_signal_17697 ;
    wire new_AGEMA_signal_17698 ;
    wire new_AGEMA_signal_17699 ;
    wire new_AGEMA_signal_17700 ;
    wire new_AGEMA_signal_17701 ;
    wire new_AGEMA_signal_17702 ;
    wire new_AGEMA_signal_17703 ;
    wire new_AGEMA_signal_17704 ;
    wire new_AGEMA_signal_17705 ;
    wire new_AGEMA_signal_17706 ;
    wire new_AGEMA_signal_17707 ;
    wire new_AGEMA_signal_17708 ;
    wire new_AGEMA_signal_17709 ;
    wire new_AGEMA_signal_17710 ;
    wire new_AGEMA_signal_17711 ;
    wire new_AGEMA_signal_17712 ;
    wire new_AGEMA_signal_17713 ;
    wire new_AGEMA_signal_17714 ;
    wire new_AGEMA_signal_17715 ;
    wire new_AGEMA_signal_17716 ;
    wire new_AGEMA_signal_17717 ;
    wire new_AGEMA_signal_17718 ;
    wire new_AGEMA_signal_17719 ;
    wire new_AGEMA_signal_17720 ;
    wire new_AGEMA_signal_17721 ;
    wire new_AGEMA_signal_17722 ;
    wire new_AGEMA_signal_17723 ;
    wire new_AGEMA_signal_17724 ;
    wire new_AGEMA_signal_17725 ;
    wire new_AGEMA_signal_17726 ;
    wire new_AGEMA_signal_17727 ;
    wire new_AGEMA_signal_17728 ;
    wire new_AGEMA_signal_17729 ;
    wire new_AGEMA_signal_17730 ;
    wire new_AGEMA_signal_17731 ;
    wire new_AGEMA_signal_17732 ;
    wire new_AGEMA_signal_17733 ;
    wire new_AGEMA_signal_17734 ;
    wire new_AGEMA_signal_17735 ;
    wire new_AGEMA_signal_17736 ;
    wire new_AGEMA_signal_17737 ;
    wire new_AGEMA_signal_17738 ;
    wire new_AGEMA_signal_17739 ;
    wire new_AGEMA_signal_17740 ;
    wire new_AGEMA_signal_17741 ;
    wire new_AGEMA_signal_17742 ;
    wire new_AGEMA_signal_17743 ;
    wire new_AGEMA_signal_17744 ;
    wire new_AGEMA_signal_17745 ;
    wire new_AGEMA_signal_17746 ;
    wire new_AGEMA_signal_17747 ;
    wire new_AGEMA_signal_17748 ;
    wire new_AGEMA_signal_17749 ;
    wire new_AGEMA_signal_17750 ;
    wire new_AGEMA_signal_17751 ;
    wire new_AGEMA_signal_17752 ;
    wire new_AGEMA_signal_17753 ;
    wire new_AGEMA_signal_17754 ;
    wire new_AGEMA_signal_17755 ;
    wire new_AGEMA_signal_17756 ;
    wire new_AGEMA_signal_17757 ;
    wire new_AGEMA_signal_17758 ;
    wire new_AGEMA_signal_17759 ;
    wire new_AGEMA_signal_17760 ;
    wire new_AGEMA_signal_17761 ;
    wire new_AGEMA_signal_17762 ;
    wire new_AGEMA_signal_17763 ;
    wire new_AGEMA_signal_17764 ;
    wire new_AGEMA_signal_17765 ;
    wire new_AGEMA_signal_17766 ;
    wire new_AGEMA_signal_17767 ;
    wire new_AGEMA_signal_17768 ;
    wire new_AGEMA_signal_17769 ;
    wire new_AGEMA_signal_17770 ;
    wire new_AGEMA_signal_17771 ;
    wire new_AGEMA_signal_17772 ;
    wire new_AGEMA_signal_17773 ;
    wire new_AGEMA_signal_17774 ;
    wire new_AGEMA_signal_17775 ;
    wire new_AGEMA_signal_17776 ;
    wire new_AGEMA_signal_17777 ;
    wire new_AGEMA_signal_17778 ;
    wire new_AGEMA_signal_17779 ;
    wire new_AGEMA_signal_17780 ;
    wire new_AGEMA_signal_17781 ;
    wire new_AGEMA_signal_17782 ;
    wire new_AGEMA_signal_17783 ;
    wire new_AGEMA_signal_17784 ;
    wire new_AGEMA_signal_17785 ;
    wire new_AGEMA_signal_17786 ;
    wire new_AGEMA_signal_17787 ;
    wire new_AGEMA_signal_17788 ;
    wire new_AGEMA_signal_17789 ;
    wire new_AGEMA_signal_17790 ;
    wire new_AGEMA_signal_17791 ;
    wire new_AGEMA_signal_17792 ;
    wire new_AGEMA_signal_17793 ;
    wire new_AGEMA_signal_17794 ;
    wire new_AGEMA_signal_17795 ;
    wire new_AGEMA_signal_17796 ;
    wire new_AGEMA_signal_17797 ;
    wire new_AGEMA_signal_17798 ;
    wire new_AGEMA_signal_17799 ;
    wire new_AGEMA_signal_17800 ;
    wire new_AGEMA_signal_17801 ;
    wire new_AGEMA_signal_17802 ;
    wire new_AGEMA_signal_17803 ;
    wire new_AGEMA_signal_17804 ;
    wire new_AGEMA_signal_17805 ;
    wire new_AGEMA_signal_17806 ;
    wire new_AGEMA_signal_17807 ;
    wire new_AGEMA_signal_17808 ;
    wire new_AGEMA_signal_17809 ;
    wire new_AGEMA_signal_17810 ;
    wire new_AGEMA_signal_17811 ;
    wire new_AGEMA_signal_17812 ;
    wire new_AGEMA_signal_17813 ;
    wire new_AGEMA_signal_17814 ;
    wire new_AGEMA_signal_17815 ;
    wire new_AGEMA_signal_17816 ;
    wire new_AGEMA_signal_17817 ;
    wire new_AGEMA_signal_17818 ;
    wire new_AGEMA_signal_17819 ;
    wire new_AGEMA_signal_17820 ;
    wire new_AGEMA_signal_17821 ;
    wire new_AGEMA_signal_17822 ;
    wire new_AGEMA_signal_17823 ;
    wire new_AGEMA_signal_17824 ;
    wire new_AGEMA_signal_17825 ;
    wire new_AGEMA_signal_17826 ;
    wire new_AGEMA_signal_17827 ;
    wire new_AGEMA_signal_17828 ;
    wire new_AGEMA_signal_17829 ;
    wire new_AGEMA_signal_17830 ;
    wire new_AGEMA_signal_17831 ;
    wire new_AGEMA_signal_17832 ;
    wire new_AGEMA_signal_17833 ;
    wire new_AGEMA_signal_17834 ;
    wire new_AGEMA_signal_17835 ;
    wire new_AGEMA_signal_17836 ;
    wire new_AGEMA_signal_17837 ;
    wire new_AGEMA_signal_17838 ;
    wire new_AGEMA_signal_17839 ;
    wire new_AGEMA_signal_17840 ;
    wire new_AGEMA_signal_17841 ;
    wire new_AGEMA_signal_17842 ;
    wire new_AGEMA_signal_17843 ;
    wire new_AGEMA_signal_17844 ;
    wire new_AGEMA_signal_17845 ;
    wire new_AGEMA_signal_17846 ;
    wire new_AGEMA_signal_17847 ;
    wire new_AGEMA_signal_17848 ;
    wire new_AGEMA_signal_17849 ;
    wire new_AGEMA_signal_17850 ;
    wire new_AGEMA_signal_17851 ;
    wire new_AGEMA_signal_17852 ;
    wire new_AGEMA_signal_17853 ;
    wire new_AGEMA_signal_17854 ;
    wire new_AGEMA_signal_17855 ;
    wire new_AGEMA_signal_17856 ;
    wire new_AGEMA_signal_17857 ;
    wire new_AGEMA_signal_17858 ;
    wire new_AGEMA_signal_17859 ;
    wire new_AGEMA_signal_17860 ;
    wire new_AGEMA_signal_17861 ;
    wire new_AGEMA_signal_17862 ;
    wire new_AGEMA_signal_17863 ;
    wire new_AGEMA_signal_17864 ;
    wire new_AGEMA_signal_17865 ;
    wire new_AGEMA_signal_17866 ;
    wire new_AGEMA_signal_17867 ;
    wire new_AGEMA_signal_17868 ;
    wire new_AGEMA_signal_17869 ;
    wire new_AGEMA_signal_17870 ;
    wire new_AGEMA_signal_17871 ;
    wire new_AGEMA_signal_17872 ;
    wire new_AGEMA_signal_17873 ;
    wire new_AGEMA_signal_17874 ;
    wire new_AGEMA_signal_17875 ;
    wire new_AGEMA_signal_17876 ;
    wire new_AGEMA_signal_17877 ;
    wire new_AGEMA_signal_17878 ;
    wire new_AGEMA_signal_17879 ;
    wire new_AGEMA_signal_17880 ;
    wire new_AGEMA_signal_17881 ;
    wire new_AGEMA_signal_17882 ;
    wire new_AGEMA_signal_17883 ;
    wire new_AGEMA_signal_17884 ;
    wire new_AGEMA_signal_17885 ;
    wire new_AGEMA_signal_17886 ;
    wire new_AGEMA_signal_17887 ;
    wire new_AGEMA_signal_17888 ;
    wire new_AGEMA_signal_17889 ;
    wire new_AGEMA_signal_17890 ;
    wire new_AGEMA_signal_17891 ;
    wire new_AGEMA_signal_17892 ;
    wire new_AGEMA_signal_17893 ;
    wire new_AGEMA_signal_17894 ;
    wire new_AGEMA_signal_17895 ;
    wire new_AGEMA_signal_17896 ;
    wire new_AGEMA_signal_17897 ;
    wire new_AGEMA_signal_17898 ;
    wire new_AGEMA_signal_17899 ;
    wire new_AGEMA_signal_17900 ;
    wire new_AGEMA_signal_17901 ;
    wire new_AGEMA_signal_17902 ;
    wire new_AGEMA_signal_17903 ;
    wire new_AGEMA_signal_17904 ;
    wire new_AGEMA_signal_17905 ;
    wire new_AGEMA_signal_17906 ;
    wire new_AGEMA_signal_17907 ;
    wire new_AGEMA_signal_17908 ;
    wire new_AGEMA_signal_17909 ;
    wire new_AGEMA_signal_17910 ;
    wire new_AGEMA_signal_17911 ;
    wire new_AGEMA_signal_17912 ;
    wire new_AGEMA_signal_17913 ;
    wire new_AGEMA_signal_17914 ;
    wire new_AGEMA_signal_17915 ;
    wire new_AGEMA_signal_17916 ;
    wire new_AGEMA_signal_17917 ;
    wire new_AGEMA_signal_17918 ;
    wire new_AGEMA_signal_17919 ;
    wire new_AGEMA_signal_17920 ;
    wire new_AGEMA_signal_17921 ;
    wire new_AGEMA_signal_17922 ;
    wire new_AGEMA_signal_17923 ;
    wire new_AGEMA_signal_17924 ;
    wire new_AGEMA_signal_17925 ;
    wire new_AGEMA_signal_17926 ;
    wire new_AGEMA_signal_17927 ;
    wire new_AGEMA_signal_17928 ;
    wire new_AGEMA_signal_17929 ;
    wire new_AGEMA_signal_17930 ;
    wire new_AGEMA_signal_17931 ;
    wire new_AGEMA_signal_17932 ;
    wire new_AGEMA_signal_17933 ;
    wire new_AGEMA_signal_17934 ;
    wire new_AGEMA_signal_17935 ;
    wire new_AGEMA_signal_17936 ;
    wire new_AGEMA_signal_17937 ;
    wire new_AGEMA_signal_17938 ;
    wire new_AGEMA_signal_17939 ;
    wire new_AGEMA_signal_17940 ;
    wire new_AGEMA_signal_17941 ;
    wire new_AGEMA_signal_17942 ;
    wire new_AGEMA_signal_17943 ;
    wire new_AGEMA_signal_17944 ;
    wire new_AGEMA_signal_17945 ;
    wire new_AGEMA_signal_17946 ;
    wire new_AGEMA_signal_17947 ;
    wire new_AGEMA_signal_17948 ;
    wire new_AGEMA_signal_17949 ;
    wire new_AGEMA_signal_17950 ;
    wire new_AGEMA_signal_17951 ;
    wire new_AGEMA_signal_17952 ;
    wire new_AGEMA_signal_17953 ;
    wire new_AGEMA_signal_17954 ;
    wire new_AGEMA_signal_17955 ;
    wire new_AGEMA_signal_17956 ;
    wire new_AGEMA_signal_17957 ;
    wire new_AGEMA_signal_17958 ;
    wire new_AGEMA_signal_17959 ;
    wire new_AGEMA_signal_17960 ;
    wire new_AGEMA_signal_17961 ;
    wire new_AGEMA_signal_17962 ;
    wire new_AGEMA_signal_17963 ;
    wire new_AGEMA_signal_17964 ;
    wire new_AGEMA_signal_17965 ;
    wire new_AGEMA_signal_17966 ;
    wire new_AGEMA_signal_17967 ;
    wire new_AGEMA_signal_17968 ;
    wire new_AGEMA_signal_17969 ;
    wire new_AGEMA_signal_17970 ;
    wire new_AGEMA_signal_17971 ;
    wire new_AGEMA_signal_17972 ;
    wire new_AGEMA_signal_17973 ;
    wire new_AGEMA_signal_17974 ;
    wire new_AGEMA_signal_17975 ;
    wire new_AGEMA_signal_17976 ;
    wire new_AGEMA_signal_17977 ;
    wire new_AGEMA_signal_17978 ;
    wire new_AGEMA_signal_17979 ;
    wire new_AGEMA_signal_17980 ;
    wire new_AGEMA_signal_17981 ;
    wire new_AGEMA_signal_17982 ;
    wire new_AGEMA_signal_17983 ;
    wire new_AGEMA_signal_17984 ;
    wire new_AGEMA_signal_17985 ;
    wire new_AGEMA_signal_17986 ;
    wire new_AGEMA_signal_17987 ;
    wire new_AGEMA_signal_17988 ;
    wire new_AGEMA_signal_17989 ;
    wire new_AGEMA_signal_17990 ;
    wire new_AGEMA_signal_17991 ;
    wire new_AGEMA_signal_17992 ;
    wire new_AGEMA_signal_17993 ;
    wire new_AGEMA_signal_17994 ;
    wire new_AGEMA_signal_17995 ;
    wire new_AGEMA_signal_17996 ;
    wire new_AGEMA_signal_17997 ;
    wire new_AGEMA_signal_17998 ;
    wire new_AGEMA_signal_17999 ;
    wire new_AGEMA_signal_18000 ;
    wire new_AGEMA_signal_18001 ;
    wire new_AGEMA_signal_18002 ;
    wire new_AGEMA_signal_18003 ;
    wire new_AGEMA_signal_18004 ;
    wire new_AGEMA_signal_18005 ;
    wire new_AGEMA_signal_18006 ;
    wire new_AGEMA_signal_18007 ;
    wire new_AGEMA_signal_18008 ;
    wire new_AGEMA_signal_18009 ;
    wire new_AGEMA_signal_18010 ;
    wire new_AGEMA_signal_18011 ;
    wire new_AGEMA_signal_18012 ;
    wire new_AGEMA_signal_18013 ;
    wire new_AGEMA_signal_18014 ;
    wire new_AGEMA_signal_18015 ;
    wire new_AGEMA_signal_18016 ;
    wire new_AGEMA_signal_18017 ;
    wire new_AGEMA_signal_18018 ;
    wire new_AGEMA_signal_18019 ;
    wire new_AGEMA_signal_18020 ;
    wire new_AGEMA_signal_18021 ;
    wire new_AGEMA_signal_18022 ;
    wire new_AGEMA_signal_18023 ;
    wire new_AGEMA_signal_18024 ;
    wire new_AGEMA_signal_18025 ;
    wire new_AGEMA_signal_18026 ;
    wire new_AGEMA_signal_18027 ;
    wire new_AGEMA_signal_18028 ;
    wire new_AGEMA_signal_18029 ;
    wire new_AGEMA_signal_18030 ;
    wire new_AGEMA_signal_18031 ;
    wire new_AGEMA_signal_18032 ;
    wire new_AGEMA_signal_18033 ;
    wire new_AGEMA_signal_18034 ;
    wire new_AGEMA_signal_18035 ;
    wire new_AGEMA_signal_18036 ;
    wire new_AGEMA_signal_18037 ;
    wire new_AGEMA_signal_18038 ;
    wire new_AGEMA_signal_18039 ;
    wire new_AGEMA_signal_18040 ;
    wire new_AGEMA_signal_18041 ;
    wire new_AGEMA_signal_18042 ;
    wire new_AGEMA_signal_18043 ;
    wire new_AGEMA_signal_18044 ;
    wire new_AGEMA_signal_18045 ;
    wire new_AGEMA_signal_18046 ;
    wire new_AGEMA_signal_18047 ;
    wire new_AGEMA_signal_18048 ;
    wire new_AGEMA_signal_18049 ;
    wire new_AGEMA_signal_18050 ;
    wire new_AGEMA_signal_18051 ;
    wire new_AGEMA_signal_18052 ;
    wire new_AGEMA_signal_18053 ;
    wire new_AGEMA_signal_18054 ;
    wire new_AGEMA_signal_18055 ;
    wire new_AGEMA_signal_18056 ;
    wire new_AGEMA_signal_18057 ;
    wire new_AGEMA_signal_18058 ;
    wire new_AGEMA_signal_18059 ;
    wire new_AGEMA_signal_18060 ;
    wire new_AGEMA_signal_18061 ;
    wire new_AGEMA_signal_18062 ;
    wire new_AGEMA_signal_18063 ;
    wire new_AGEMA_signal_18064 ;
    wire new_AGEMA_signal_18065 ;
    wire new_AGEMA_signal_18066 ;
    wire new_AGEMA_signal_18067 ;
    wire new_AGEMA_signal_18068 ;
    wire new_AGEMA_signal_18069 ;
    wire new_AGEMA_signal_18070 ;
    wire new_AGEMA_signal_18071 ;
    wire new_AGEMA_signal_18072 ;
    wire new_AGEMA_signal_18073 ;
    wire new_AGEMA_signal_18074 ;
    wire new_AGEMA_signal_18075 ;
    wire new_AGEMA_signal_18076 ;
    wire new_AGEMA_signal_18077 ;
    wire new_AGEMA_signal_18078 ;
    wire new_AGEMA_signal_18079 ;
    wire new_AGEMA_signal_18080 ;
    wire new_AGEMA_signal_18081 ;
    wire new_AGEMA_signal_18082 ;
    wire new_AGEMA_signal_18083 ;
    wire new_AGEMA_signal_18084 ;
    wire new_AGEMA_signal_18085 ;
    wire new_AGEMA_signal_18086 ;
    wire new_AGEMA_signal_18087 ;
    wire new_AGEMA_signal_18088 ;
    wire new_AGEMA_signal_18089 ;
    wire new_AGEMA_signal_18090 ;
    wire new_AGEMA_signal_18091 ;
    wire new_AGEMA_signal_18092 ;
    wire new_AGEMA_signal_18093 ;
    wire new_AGEMA_signal_18094 ;
    wire new_AGEMA_signal_18095 ;
    wire new_AGEMA_signal_18096 ;
    wire new_AGEMA_signal_18097 ;
    wire new_AGEMA_signal_18098 ;
    wire new_AGEMA_signal_18099 ;
    wire new_AGEMA_signal_18100 ;
    wire new_AGEMA_signal_18101 ;
    wire new_AGEMA_signal_18102 ;
    wire new_AGEMA_signal_18103 ;
    wire new_AGEMA_signal_18104 ;
    wire new_AGEMA_signal_18105 ;
    wire new_AGEMA_signal_18106 ;
    wire new_AGEMA_signal_18107 ;
    wire new_AGEMA_signal_18108 ;
    wire new_AGEMA_signal_18109 ;
    wire new_AGEMA_signal_18110 ;
    wire new_AGEMA_signal_18111 ;
    wire new_AGEMA_signal_18112 ;
    wire new_AGEMA_signal_18113 ;
    wire new_AGEMA_signal_18114 ;
    wire new_AGEMA_signal_18115 ;
    wire new_AGEMA_signal_18116 ;
    wire new_AGEMA_signal_18117 ;
    wire new_AGEMA_signal_18118 ;
    wire new_AGEMA_signal_18119 ;
    wire new_AGEMA_signal_18120 ;
    wire new_AGEMA_signal_18121 ;
    wire new_AGEMA_signal_18122 ;
    wire new_AGEMA_signal_18123 ;
    wire new_AGEMA_signal_18124 ;
    wire new_AGEMA_signal_18125 ;
    wire new_AGEMA_signal_18126 ;
    wire new_AGEMA_signal_18127 ;
    wire new_AGEMA_signal_18128 ;
    wire new_AGEMA_signal_18129 ;
    wire new_AGEMA_signal_18130 ;
    wire new_AGEMA_signal_18131 ;
    wire new_AGEMA_signal_18132 ;
    wire new_AGEMA_signal_18133 ;
    wire new_AGEMA_signal_18134 ;
    wire new_AGEMA_signal_18135 ;
    wire new_AGEMA_signal_18136 ;
    wire new_AGEMA_signal_18137 ;
    wire new_AGEMA_signal_18138 ;
    wire new_AGEMA_signal_18139 ;
    wire new_AGEMA_signal_18140 ;
    wire new_AGEMA_signal_18141 ;
    wire new_AGEMA_signal_18142 ;
    wire new_AGEMA_signal_18143 ;
    wire new_AGEMA_signal_18144 ;
    wire new_AGEMA_signal_18145 ;
    wire new_AGEMA_signal_18146 ;
    wire new_AGEMA_signal_18147 ;
    wire new_AGEMA_signal_18148 ;
    wire new_AGEMA_signal_18149 ;
    wire new_AGEMA_signal_18150 ;
    wire new_AGEMA_signal_18151 ;
    wire new_AGEMA_signal_18152 ;
    wire new_AGEMA_signal_18153 ;
    wire new_AGEMA_signal_18154 ;
    wire new_AGEMA_signal_18155 ;
    wire new_AGEMA_signal_18156 ;
    wire new_AGEMA_signal_18157 ;
    wire new_AGEMA_signal_18158 ;
    wire new_AGEMA_signal_18159 ;
    wire new_AGEMA_signal_18160 ;
    wire new_AGEMA_signal_18161 ;
    wire new_AGEMA_signal_18162 ;
    wire new_AGEMA_signal_18163 ;
    wire new_AGEMA_signal_18164 ;
    wire new_AGEMA_signal_18165 ;
    wire new_AGEMA_signal_18166 ;
    wire new_AGEMA_signal_18167 ;
    wire new_AGEMA_signal_18168 ;
    wire new_AGEMA_signal_18169 ;
    wire new_AGEMA_signal_18170 ;
    wire new_AGEMA_signal_18171 ;
    wire new_AGEMA_signal_18172 ;
    wire new_AGEMA_signal_18173 ;
    wire new_AGEMA_signal_18174 ;
    wire new_AGEMA_signal_18175 ;
    wire new_AGEMA_signal_18176 ;
    wire new_AGEMA_signal_18177 ;
    wire new_AGEMA_signal_18178 ;
    wire new_AGEMA_signal_18179 ;
    wire new_AGEMA_signal_18180 ;
    wire new_AGEMA_signal_18181 ;
    wire new_AGEMA_signal_18182 ;
    wire new_AGEMA_signal_18183 ;
    wire new_AGEMA_signal_18184 ;
    wire new_AGEMA_signal_18185 ;
    wire new_AGEMA_signal_18186 ;
    wire new_AGEMA_signal_18187 ;
    wire new_AGEMA_signal_18188 ;
    wire new_AGEMA_signal_18189 ;
    wire new_AGEMA_signal_18190 ;
    wire new_AGEMA_signal_18191 ;
    wire new_AGEMA_signal_18192 ;
    wire new_AGEMA_signal_18193 ;
    wire new_AGEMA_signal_18194 ;
    wire new_AGEMA_signal_18195 ;
    wire new_AGEMA_signal_18196 ;
    wire new_AGEMA_signal_18197 ;
    wire new_AGEMA_signal_18198 ;
    wire new_AGEMA_signal_18199 ;
    wire new_AGEMA_signal_18200 ;
    wire new_AGEMA_signal_18201 ;
    wire new_AGEMA_signal_18202 ;
    wire new_AGEMA_signal_18203 ;
    wire new_AGEMA_signal_18204 ;
    wire new_AGEMA_signal_18205 ;
    wire new_AGEMA_signal_18206 ;
    wire new_AGEMA_signal_18207 ;
    wire new_AGEMA_signal_18208 ;
    wire new_AGEMA_signal_18209 ;
    wire new_AGEMA_signal_18210 ;
    wire new_AGEMA_signal_18211 ;
    wire new_AGEMA_signal_18212 ;
    wire new_AGEMA_signal_18213 ;
    wire new_AGEMA_signal_18214 ;
    wire new_AGEMA_signal_18215 ;
    wire new_AGEMA_signal_18216 ;
    wire new_AGEMA_signal_18217 ;
    wire new_AGEMA_signal_18218 ;
    wire new_AGEMA_signal_18219 ;
    wire new_AGEMA_signal_18220 ;
    wire new_AGEMA_signal_18221 ;
    wire new_AGEMA_signal_18222 ;
    wire new_AGEMA_signal_18223 ;
    wire new_AGEMA_signal_18224 ;
    wire new_AGEMA_signal_18225 ;
    wire new_AGEMA_signal_18226 ;
    wire new_AGEMA_signal_18227 ;
    wire new_AGEMA_signal_18228 ;
    wire new_AGEMA_signal_18229 ;
    wire new_AGEMA_signal_18230 ;
    wire new_AGEMA_signal_18231 ;
    wire new_AGEMA_signal_18232 ;
    wire new_AGEMA_signal_18233 ;
    wire new_AGEMA_signal_18234 ;
    wire new_AGEMA_signal_18235 ;
    wire new_AGEMA_signal_18236 ;
    wire new_AGEMA_signal_18237 ;
    wire new_AGEMA_signal_18238 ;
    wire new_AGEMA_signal_18239 ;
    wire new_AGEMA_signal_18240 ;
    wire new_AGEMA_signal_18241 ;
    wire new_AGEMA_signal_18242 ;
    wire new_AGEMA_signal_18243 ;
    wire new_AGEMA_signal_18244 ;
    wire new_AGEMA_signal_18245 ;
    wire new_AGEMA_signal_18246 ;
    wire new_AGEMA_signal_18247 ;
    wire new_AGEMA_signal_18248 ;
    wire new_AGEMA_signal_18249 ;
    wire new_AGEMA_signal_18250 ;
    wire new_AGEMA_signal_18251 ;
    wire new_AGEMA_signal_18252 ;
    wire new_AGEMA_signal_18253 ;
    wire new_AGEMA_signal_18254 ;
    wire new_AGEMA_signal_18255 ;
    wire new_AGEMA_signal_18256 ;
    wire new_AGEMA_signal_18257 ;
    wire new_AGEMA_signal_18258 ;
    wire new_AGEMA_signal_18259 ;
    wire new_AGEMA_signal_18260 ;
    wire new_AGEMA_signal_18261 ;
    wire new_AGEMA_signal_18262 ;
    wire new_AGEMA_signal_18263 ;
    wire new_AGEMA_signal_18264 ;
    wire new_AGEMA_signal_18265 ;
    wire new_AGEMA_signal_18266 ;
    wire new_AGEMA_signal_18267 ;
    wire new_AGEMA_signal_18268 ;
    wire new_AGEMA_signal_18269 ;
    wire new_AGEMA_signal_18270 ;
    wire new_AGEMA_signal_18271 ;
    wire new_AGEMA_signal_18272 ;
    wire new_AGEMA_signal_18273 ;
    wire new_AGEMA_signal_18274 ;
    wire new_AGEMA_signal_18275 ;
    wire new_AGEMA_signal_18276 ;
    wire new_AGEMA_signal_18277 ;
    wire new_AGEMA_signal_18278 ;
    wire new_AGEMA_signal_18279 ;
    wire new_AGEMA_signal_18280 ;
    wire new_AGEMA_signal_18281 ;
    wire new_AGEMA_signal_18282 ;
    wire new_AGEMA_signal_18283 ;
    wire new_AGEMA_signal_18284 ;
    wire new_AGEMA_signal_18285 ;
    wire new_AGEMA_signal_18286 ;
    wire new_AGEMA_signal_18287 ;
    wire new_AGEMA_signal_18288 ;
    wire new_AGEMA_signal_18289 ;
    wire new_AGEMA_signal_18290 ;
    wire new_AGEMA_signal_18291 ;
    wire new_AGEMA_signal_18292 ;
    wire new_AGEMA_signal_18293 ;
    wire new_AGEMA_signal_18294 ;
    wire new_AGEMA_signal_18295 ;
    wire new_AGEMA_signal_18296 ;
    wire new_AGEMA_signal_18297 ;
    wire new_AGEMA_signal_18298 ;
    wire new_AGEMA_signal_18299 ;
    wire new_AGEMA_signal_18300 ;
    wire new_AGEMA_signal_18301 ;
    wire new_AGEMA_signal_18302 ;
    wire new_AGEMA_signal_18303 ;
    wire new_AGEMA_signal_18304 ;
    wire new_AGEMA_signal_18305 ;
    wire new_AGEMA_signal_18306 ;
    wire new_AGEMA_signal_18307 ;
    wire new_AGEMA_signal_18308 ;
    wire new_AGEMA_signal_18309 ;
    wire new_AGEMA_signal_18310 ;
    wire new_AGEMA_signal_18311 ;
    wire new_AGEMA_signal_18312 ;
    wire new_AGEMA_signal_18313 ;
    wire new_AGEMA_signal_18314 ;
    wire new_AGEMA_signal_18315 ;
    wire new_AGEMA_signal_18316 ;
    wire new_AGEMA_signal_18317 ;
    wire new_AGEMA_signal_18318 ;
    wire new_AGEMA_signal_18319 ;
    wire new_AGEMA_signal_18320 ;
    wire new_AGEMA_signal_18321 ;
    wire new_AGEMA_signal_18322 ;
    wire new_AGEMA_signal_18323 ;
    wire new_AGEMA_signal_18324 ;
    wire new_AGEMA_signal_18325 ;
    wire new_AGEMA_signal_18326 ;
    wire new_AGEMA_signal_18327 ;
    wire new_AGEMA_signal_18328 ;
    wire new_AGEMA_signal_18329 ;
    wire new_AGEMA_signal_18330 ;
    wire new_AGEMA_signal_18331 ;
    wire new_AGEMA_signal_18332 ;
    wire new_AGEMA_signal_18333 ;
    wire new_AGEMA_signal_18334 ;
    wire new_AGEMA_signal_18335 ;
    wire new_AGEMA_signal_18336 ;
    wire new_AGEMA_signal_18337 ;
    wire new_AGEMA_signal_18338 ;
    wire new_AGEMA_signal_18339 ;
    wire new_AGEMA_signal_18340 ;
    wire new_AGEMA_signal_18341 ;
    wire new_AGEMA_signal_18342 ;
    wire new_AGEMA_signal_18343 ;
    wire new_AGEMA_signal_18344 ;
    wire new_AGEMA_signal_18345 ;
    wire new_AGEMA_signal_18346 ;
    wire new_AGEMA_signal_18347 ;
    wire new_AGEMA_signal_18348 ;
    wire new_AGEMA_signal_18349 ;
    wire new_AGEMA_signal_18350 ;
    wire new_AGEMA_signal_18351 ;
    wire new_AGEMA_signal_18352 ;
    wire new_AGEMA_signal_18353 ;
    wire new_AGEMA_signal_18354 ;
    wire new_AGEMA_signal_18355 ;
    wire new_AGEMA_signal_18356 ;
    wire new_AGEMA_signal_18357 ;
    wire new_AGEMA_signal_18358 ;
    wire new_AGEMA_signal_18359 ;
    wire new_AGEMA_signal_18360 ;
    wire new_AGEMA_signal_18361 ;
    wire new_AGEMA_signal_18362 ;
    wire new_AGEMA_signal_18363 ;
    wire new_AGEMA_signal_18364 ;
    wire new_AGEMA_signal_18365 ;
    wire new_AGEMA_signal_18366 ;
    wire new_AGEMA_signal_18367 ;
    wire new_AGEMA_signal_18368 ;
    wire new_AGEMA_signal_18369 ;
    wire new_AGEMA_signal_18370 ;
    wire new_AGEMA_signal_18371 ;
    wire new_AGEMA_signal_18372 ;
    wire new_AGEMA_signal_18373 ;
    wire new_AGEMA_signal_18374 ;
    wire new_AGEMA_signal_18375 ;
    wire new_AGEMA_signal_18376 ;
    wire new_AGEMA_signal_18377 ;
    wire new_AGEMA_signal_18378 ;
    wire new_AGEMA_signal_18379 ;
    wire new_AGEMA_signal_18380 ;
    wire new_AGEMA_signal_18381 ;
    wire new_AGEMA_signal_18382 ;
    wire new_AGEMA_signal_18383 ;
    wire new_AGEMA_signal_18384 ;
    wire new_AGEMA_signal_18385 ;
    wire new_AGEMA_signal_18386 ;
    wire new_AGEMA_signal_18387 ;
    wire new_AGEMA_signal_18388 ;
    wire new_AGEMA_signal_18389 ;
    wire new_AGEMA_signal_18390 ;
    wire new_AGEMA_signal_18391 ;
    wire new_AGEMA_signal_18392 ;
    wire new_AGEMA_signal_18393 ;
    wire new_AGEMA_signal_18394 ;
    wire new_AGEMA_signal_18395 ;
    wire new_AGEMA_signal_18396 ;
    wire new_AGEMA_signal_18397 ;
    wire new_AGEMA_signal_18398 ;
    wire new_AGEMA_signal_18399 ;
    wire new_AGEMA_signal_18400 ;
    wire new_AGEMA_signal_18401 ;
    wire new_AGEMA_signal_18402 ;
    wire new_AGEMA_signal_18403 ;
    wire new_AGEMA_signal_18404 ;
    wire new_AGEMA_signal_18405 ;
    wire new_AGEMA_signal_18406 ;
    wire new_AGEMA_signal_18407 ;
    wire new_AGEMA_signal_18408 ;
    wire new_AGEMA_signal_18409 ;
    wire new_AGEMA_signal_18410 ;
    wire new_AGEMA_signal_18411 ;
    wire new_AGEMA_signal_18412 ;
    wire new_AGEMA_signal_18413 ;
    wire new_AGEMA_signal_18414 ;
    wire new_AGEMA_signal_18415 ;
    wire new_AGEMA_signal_18416 ;
    wire new_AGEMA_signal_18417 ;
    wire new_AGEMA_signal_18418 ;
    wire new_AGEMA_signal_18419 ;
    wire new_AGEMA_signal_18420 ;
    wire new_AGEMA_signal_18421 ;
    wire new_AGEMA_signal_18422 ;
    wire new_AGEMA_signal_18423 ;
    wire new_AGEMA_signal_18424 ;
    wire new_AGEMA_signal_18425 ;
    wire new_AGEMA_signal_18426 ;
    wire new_AGEMA_signal_18427 ;
    wire new_AGEMA_signal_18428 ;
    wire new_AGEMA_signal_18429 ;
    wire new_AGEMA_signal_18430 ;
    wire new_AGEMA_signal_18431 ;
    wire new_AGEMA_signal_18432 ;
    wire new_AGEMA_signal_18433 ;
    wire new_AGEMA_signal_18434 ;
    wire new_AGEMA_signal_18435 ;
    wire new_AGEMA_signal_18436 ;
    wire new_AGEMA_signal_18437 ;
    wire new_AGEMA_signal_18438 ;
    wire new_AGEMA_signal_18439 ;
    wire new_AGEMA_signal_18440 ;
    wire new_AGEMA_signal_18441 ;
    wire new_AGEMA_signal_18442 ;
    wire new_AGEMA_signal_18443 ;
    wire new_AGEMA_signal_18444 ;
    wire new_AGEMA_signal_18445 ;
    wire new_AGEMA_signal_18446 ;
    wire new_AGEMA_signal_18447 ;
    wire new_AGEMA_signal_18448 ;
    wire new_AGEMA_signal_18449 ;
    wire new_AGEMA_signal_18450 ;
    wire new_AGEMA_signal_18451 ;
    wire new_AGEMA_signal_18452 ;
    wire new_AGEMA_signal_18453 ;
    wire new_AGEMA_signal_18454 ;
    wire new_AGEMA_signal_18455 ;
    wire new_AGEMA_signal_18456 ;
    wire new_AGEMA_signal_18457 ;
    wire new_AGEMA_signal_18458 ;
    wire new_AGEMA_signal_18459 ;
    wire new_AGEMA_signal_18460 ;
    wire new_AGEMA_signal_18461 ;
    wire new_AGEMA_signal_18462 ;
    wire new_AGEMA_signal_18463 ;
    wire new_AGEMA_signal_18464 ;
    wire new_AGEMA_signal_18465 ;
    wire new_AGEMA_signal_18466 ;
    wire new_AGEMA_signal_18467 ;
    wire new_AGEMA_signal_18468 ;
    wire new_AGEMA_signal_18469 ;
    wire new_AGEMA_signal_18470 ;
    wire new_AGEMA_signal_18471 ;
    wire new_AGEMA_signal_18472 ;
    wire new_AGEMA_signal_18473 ;
    wire new_AGEMA_signal_18474 ;
    wire new_AGEMA_signal_18475 ;
    wire new_AGEMA_signal_18476 ;
    wire new_AGEMA_signal_18477 ;
    wire new_AGEMA_signal_18478 ;
    wire new_AGEMA_signal_18479 ;
    wire new_AGEMA_signal_18480 ;
    wire new_AGEMA_signal_18481 ;
    wire new_AGEMA_signal_18482 ;
    wire new_AGEMA_signal_18483 ;
    wire new_AGEMA_signal_18484 ;
    wire new_AGEMA_signal_18485 ;
    wire new_AGEMA_signal_18486 ;
    wire new_AGEMA_signal_18487 ;
    wire new_AGEMA_signal_18488 ;
    wire new_AGEMA_signal_18489 ;
    wire new_AGEMA_signal_18490 ;
    wire new_AGEMA_signal_18491 ;
    wire new_AGEMA_signal_18492 ;
    wire new_AGEMA_signal_18493 ;
    wire new_AGEMA_signal_18494 ;
    wire new_AGEMA_signal_18495 ;
    wire new_AGEMA_signal_18496 ;
    wire new_AGEMA_signal_18497 ;
    wire new_AGEMA_signal_18498 ;
    wire new_AGEMA_signal_18499 ;
    wire new_AGEMA_signal_18500 ;
    wire new_AGEMA_signal_18501 ;
    wire new_AGEMA_signal_18502 ;
    wire new_AGEMA_signal_18503 ;
    wire new_AGEMA_signal_18504 ;
    wire new_AGEMA_signal_18505 ;
    wire new_AGEMA_signal_18506 ;
    wire new_AGEMA_signal_18507 ;
    wire new_AGEMA_signal_18508 ;
    wire new_AGEMA_signal_18509 ;
    wire new_AGEMA_signal_18510 ;
    wire new_AGEMA_signal_18511 ;
    wire new_AGEMA_signal_18512 ;
    wire new_AGEMA_signal_18513 ;
    wire new_AGEMA_signal_18514 ;
    wire new_AGEMA_signal_18515 ;
    wire new_AGEMA_signal_18516 ;
    wire new_AGEMA_signal_18517 ;
    wire new_AGEMA_signal_18518 ;
    wire new_AGEMA_signal_18519 ;
    wire new_AGEMA_signal_18520 ;
    wire new_AGEMA_signal_18521 ;
    wire new_AGEMA_signal_18522 ;
    wire new_AGEMA_signal_18523 ;
    wire new_AGEMA_signal_18524 ;
    wire new_AGEMA_signal_18525 ;
    wire new_AGEMA_signal_18526 ;
    wire new_AGEMA_signal_18527 ;
    wire new_AGEMA_signal_18528 ;
    wire new_AGEMA_signal_18529 ;
    wire new_AGEMA_signal_18530 ;
    wire new_AGEMA_signal_18531 ;
    wire new_AGEMA_signal_18532 ;
    wire new_AGEMA_signal_18533 ;
    wire new_AGEMA_signal_18534 ;
    wire new_AGEMA_signal_18535 ;
    wire new_AGEMA_signal_18536 ;
    wire new_AGEMA_signal_18537 ;
    wire new_AGEMA_signal_18538 ;
    wire new_AGEMA_signal_18539 ;
    wire new_AGEMA_signal_18540 ;
    wire new_AGEMA_signal_18541 ;
    wire new_AGEMA_signal_18542 ;
    wire new_AGEMA_signal_18543 ;
    wire new_AGEMA_signal_18544 ;
    wire new_AGEMA_signal_18545 ;
    wire new_AGEMA_signal_18546 ;
    wire new_AGEMA_signal_18547 ;
    wire new_AGEMA_signal_18548 ;
    wire new_AGEMA_signal_18549 ;
    wire new_AGEMA_signal_18550 ;
    wire new_AGEMA_signal_18551 ;
    wire new_AGEMA_signal_18552 ;
    wire new_AGEMA_signal_18553 ;
    wire new_AGEMA_signal_18554 ;
    wire new_AGEMA_signal_18555 ;
    wire new_AGEMA_signal_18556 ;
    wire new_AGEMA_signal_18557 ;
    wire new_AGEMA_signal_18558 ;
    wire new_AGEMA_signal_18559 ;
    wire new_AGEMA_signal_18560 ;
    wire new_AGEMA_signal_18561 ;
    wire new_AGEMA_signal_18562 ;
    wire new_AGEMA_signal_18563 ;
    wire new_AGEMA_signal_18564 ;
    wire new_AGEMA_signal_18565 ;
    wire new_AGEMA_signal_18566 ;
    wire new_AGEMA_signal_18567 ;
    wire new_AGEMA_signal_18568 ;
    wire new_AGEMA_signal_18569 ;
    wire new_AGEMA_signal_18570 ;
    wire new_AGEMA_signal_18571 ;
    wire new_AGEMA_signal_18572 ;
    wire new_AGEMA_signal_18573 ;
    wire new_AGEMA_signal_18574 ;
    wire new_AGEMA_signal_18575 ;
    wire new_AGEMA_signal_18576 ;
    wire new_AGEMA_signal_18577 ;
    wire new_AGEMA_signal_18578 ;
    wire new_AGEMA_signal_18579 ;
    wire new_AGEMA_signal_18580 ;
    wire new_AGEMA_signal_18581 ;
    wire new_AGEMA_signal_18582 ;
    wire new_AGEMA_signal_18583 ;
    wire new_AGEMA_signal_18584 ;
    wire new_AGEMA_signal_18585 ;
    wire new_AGEMA_signal_18586 ;
    wire new_AGEMA_signal_18587 ;
    wire new_AGEMA_signal_18588 ;
    wire new_AGEMA_signal_18589 ;
    wire new_AGEMA_signal_18590 ;
    wire new_AGEMA_signal_18591 ;
    wire new_AGEMA_signal_18592 ;
    wire new_AGEMA_signal_18593 ;
    wire new_AGEMA_signal_18594 ;
    wire new_AGEMA_signal_18595 ;
    wire new_AGEMA_signal_18596 ;
    wire new_AGEMA_signal_18597 ;
    wire new_AGEMA_signal_18598 ;
    wire new_AGEMA_signal_18599 ;
    wire new_AGEMA_signal_18600 ;
    wire new_AGEMA_signal_18601 ;
    wire new_AGEMA_signal_18602 ;
    wire new_AGEMA_signal_18603 ;
    wire new_AGEMA_signal_18604 ;
    wire new_AGEMA_signal_18605 ;
    wire new_AGEMA_signal_18606 ;
    wire new_AGEMA_signal_18607 ;
    wire new_AGEMA_signal_18608 ;
    wire new_AGEMA_signal_18609 ;
    wire new_AGEMA_signal_18610 ;
    wire new_AGEMA_signal_18611 ;
    wire new_AGEMA_signal_18612 ;
    wire new_AGEMA_signal_18613 ;
    wire new_AGEMA_signal_18614 ;
    wire new_AGEMA_signal_18615 ;
    wire new_AGEMA_signal_18616 ;
    wire new_AGEMA_signal_18617 ;
    wire new_AGEMA_signal_18618 ;
    wire new_AGEMA_signal_18619 ;
    wire new_AGEMA_signal_18620 ;
    wire new_AGEMA_signal_18621 ;
    wire new_AGEMA_signal_18622 ;
    wire new_AGEMA_signal_18623 ;
    wire new_AGEMA_signal_18624 ;
    wire new_AGEMA_signal_18625 ;
    wire new_AGEMA_signal_18626 ;
    wire new_AGEMA_signal_18627 ;
    wire new_AGEMA_signal_18628 ;
    wire new_AGEMA_signal_18629 ;
    wire new_AGEMA_signal_18630 ;
    wire new_AGEMA_signal_18631 ;
    wire new_AGEMA_signal_18632 ;
    wire new_AGEMA_signal_18633 ;
    wire new_AGEMA_signal_18634 ;
    wire new_AGEMA_signal_18635 ;
    wire new_AGEMA_signal_18636 ;
    wire new_AGEMA_signal_18637 ;
    wire new_AGEMA_signal_18638 ;
    wire new_AGEMA_signal_18639 ;
    wire new_AGEMA_signal_18640 ;
    wire new_AGEMA_signal_18641 ;
    wire new_AGEMA_signal_18642 ;
    wire new_AGEMA_signal_18643 ;
    wire new_AGEMA_signal_18644 ;
    wire new_AGEMA_signal_18645 ;
    wire new_AGEMA_signal_18646 ;
    wire new_AGEMA_signal_18647 ;
    wire new_AGEMA_signal_18648 ;
    wire new_AGEMA_signal_18649 ;
    wire new_AGEMA_signal_18650 ;
    wire new_AGEMA_signal_18651 ;
    wire new_AGEMA_signal_18652 ;
    wire new_AGEMA_signal_18653 ;
    wire new_AGEMA_signal_18654 ;
    wire new_AGEMA_signal_18655 ;
    wire new_AGEMA_signal_18656 ;
    wire new_AGEMA_signal_18657 ;
    wire new_AGEMA_signal_18658 ;
    wire new_AGEMA_signal_18659 ;
    wire new_AGEMA_signal_18660 ;
    wire new_AGEMA_signal_18661 ;
    wire new_AGEMA_signal_18662 ;
    wire new_AGEMA_signal_18663 ;
    wire new_AGEMA_signal_18664 ;
    wire new_AGEMA_signal_18665 ;
    wire new_AGEMA_signal_18666 ;
    wire new_AGEMA_signal_18667 ;
    wire new_AGEMA_signal_18668 ;
    wire new_AGEMA_signal_18669 ;
    wire new_AGEMA_signal_18670 ;
    wire new_AGEMA_signal_18671 ;
    wire new_AGEMA_signal_18672 ;
    wire new_AGEMA_signal_18673 ;
    wire new_AGEMA_signal_18674 ;
    wire new_AGEMA_signal_18675 ;
    wire new_AGEMA_signal_18676 ;
    wire new_AGEMA_signal_18677 ;
    wire new_AGEMA_signal_18678 ;
    wire new_AGEMA_signal_18679 ;
    wire new_AGEMA_signal_18680 ;
    wire new_AGEMA_signal_18681 ;
    wire new_AGEMA_signal_18682 ;
    wire new_AGEMA_signal_18683 ;
    wire new_AGEMA_signal_18684 ;
    wire new_AGEMA_signal_18685 ;
    wire new_AGEMA_signal_18686 ;
    wire new_AGEMA_signal_18687 ;
    wire new_AGEMA_signal_18688 ;
    wire new_AGEMA_signal_18689 ;
    wire new_AGEMA_signal_18690 ;
    wire new_AGEMA_signal_18691 ;
    wire new_AGEMA_signal_18692 ;
    wire new_AGEMA_signal_18693 ;
    wire new_AGEMA_signal_18694 ;
    wire new_AGEMA_signal_18695 ;
    wire new_AGEMA_signal_18696 ;
    wire new_AGEMA_signal_18697 ;
    wire new_AGEMA_signal_18698 ;
    wire new_AGEMA_signal_18699 ;
    wire new_AGEMA_signal_18700 ;
    wire new_AGEMA_signal_18701 ;
    wire new_AGEMA_signal_18702 ;
    wire new_AGEMA_signal_18703 ;
    wire new_AGEMA_signal_18704 ;
    wire new_AGEMA_signal_18705 ;
    wire new_AGEMA_signal_18706 ;
    wire new_AGEMA_signal_18707 ;
    wire new_AGEMA_signal_18708 ;
    wire new_AGEMA_signal_18709 ;
    wire new_AGEMA_signal_18710 ;
    wire new_AGEMA_signal_18711 ;
    wire new_AGEMA_signal_18712 ;
    wire new_AGEMA_signal_18713 ;
    wire new_AGEMA_signal_18714 ;
    wire new_AGEMA_signal_18715 ;
    wire new_AGEMA_signal_18716 ;
    wire new_AGEMA_signal_18717 ;
    wire new_AGEMA_signal_18718 ;
    wire new_AGEMA_signal_18719 ;
    wire new_AGEMA_signal_18720 ;
    wire new_AGEMA_signal_18721 ;
    wire new_AGEMA_signal_18722 ;
    wire new_AGEMA_signal_18723 ;
    wire new_AGEMA_signal_18724 ;
    wire new_AGEMA_signal_18725 ;
    wire new_AGEMA_signal_18726 ;
    wire new_AGEMA_signal_18727 ;
    wire new_AGEMA_signal_18728 ;
    wire new_AGEMA_signal_18729 ;
    wire new_AGEMA_signal_18730 ;
    wire new_AGEMA_signal_18731 ;
    wire new_AGEMA_signal_18732 ;
    wire new_AGEMA_signal_18733 ;
    wire new_AGEMA_signal_18734 ;
    wire new_AGEMA_signal_18735 ;
    wire new_AGEMA_signal_18736 ;
    wire new_AGEMA_signal_18737 ;
    wire new_AGEMA_signal_18738 ;
    wire new_AGEMA_signal_18739 ;
    wire new_AGEMA_signal_18740 ;
    wire new_AGEMA_signal_18741 ;
    wire new_AGEMA_signal_18742 ;
    wire new_AGEMA_signal_18743 ;
    wire new_AGEMA_signal_18744 ;
    wire new_AGEMA_signal_18745 ;
    wire new_AGEMA_signal_18746 ;
    wire new_AGEMA_signal_18747 ;
    wire new_AGEMA_signal_18748 ;
    wire new_AGEMA_signal_18749 ;
    wire new_AGEMA_signal_18750 ;
    wire new_AGEMA_signal_18751 ;
    wire new_AGEMA_signal_18752 ;
    wire new_AGEMA_signal_18753 ;
    wire new_AGEMA_signal_18754 ;
    wire new_AGEMA_signal_18755 ;
    wire new_AGEMA_signal_18756 ;
    wire new_AGEMA_signal_18757 ;
    wire new_AGEMA_signal_18758 ;
    wire new_AGEMA_signal_18759 ;
    wire new_AGEMA_signal_18760 ;
    wire new_AGEMA_signal_18761 ;
    wire new_AGEMA_signal_18762 ;
    wire new_AGEMA_signal_18763 ;
    wire new_AGEMA_signal_18764 ;
    wire new_AGEMA_signal_18765 ;
    wire new_AGEMA_signal_18766 ;
    wire new_AGEMA_signal_18767 ;
    wire new_AGEMA_signal_18768 ;
    wire new_AGEMA_signal_18769 ;
    wire new_AGEMA_signal_18770 ;
    wire new_AGEMA_signal_18771 ;
    wire new_AGEMA_signal_18772 ;
    wire new_AGEMA_signal_18773 ;
    wire new_AGEMA_signal_18774 ;
    wire new_AGEMA_signal_18775 ;
    wire new_AGEMA_signal_18776 ;
    wire new_AGEMA_signal_18777 ;
    wire new_AGEMA_signal_18778 ;
    wire new_AGEMA_signal_18779 ;
    wire new_AGEMA_signal_18780 ;
    wire new_AGEMA_signal_18781 ;
    wire new_AGEMA_signal_18782 ;
    wire new_AGEMA_signal_18783 ;
    wire new_AGEMA_signal_18784 ;
    wire new_AGEMA_signal_18785 ;
    wire new_AGEMA_signal_18786 ;
    wire new_AGEMA_signal_18787 ;
    wire new_AGEMA_signal_18788 ;
    wire new_AGEMA_signal_18789 ;
    wire new_AGEMA_signal_18790 ;
    wire new_AGEMA_signal_18791 ;
    wire new_AGEMA_signal_18792 ;
    wire new_AGEMA_signal_18793 ;
    wire new_AGEMA_signal_18794 ;
    wire new_AGEMA_signal_18795 ;
    wire new_AGEMA_signal_18796 ;
    wire new_AGEMA_signal_18797 ;
    wire new_AGEMA_signal_18798 ;
    wire new_AGEMA_signal_18799 ;
    wire new_AGEMA_signal_18800 ;
    wire new_AGEMA_signal_18801 ;
    wire new_AGEMA_signal_18802 ;
    wire new_AGEMA_signal_18803 ;
    wire new_AGEMA_signal_18804 ;
    wire new_AGEMA_signal_18805 ;
    wire new_AGEMA_signal_18806 ;
    wire new_AGEMA_signal_18807 ;
    wire new_AGEMA_signal_18808 ;
    wire new_AGEMA_signal_18809 ;
    wire new_AGEMA_signal_18810 ;
    wire new_AGEMA_signal_18811 ;
    wire new_AGEMA_signal_18812 ;
    wire new_AGEMA_signal_18813 ;
    wire new_AGEMA_signal_18814 ;
    wire new_AGEMA_signal_18815 ;
    wire new_AGEMA_signal_18816 ;
    wire new_AGEMA_signal_18817 ;
    wire new_AGEMA_signal_18818 ;
    wire new_AGEMA_signal_18819 ;
    wire new_AGEMA_signal_18820 ;
    wire new_AGEMA_signal_18821 ;
    wire new_AGEMA_signal_18822 ;
    wire new_AGEMA_signal_18823 ;
    wire new_AGEMA_signal_18824 ;
    wire new_AGEMA_signal_18825 ;
    wire new_AGEMA_signal_18826 ;
    wire new_AGEMA_signal_18827 ;
    wire new_AGEMA_signal_18828 ;
    wire new_AGEMA_signal_18829 ;
    wire new_AGEMA_signal_18830 ;
    wire new_AGEMA_signal_18831 ;
    wire new_AGEMA_signal_18832 ;
    wire new_AGEMA_signal_18833 ;
    wire new_AGEMA_signal_18834 ;
    wire new_AGEMA_signal_18835 ;
    wire new_AGEMA_signal_18836 ;
    wire new_AGEMA_signal_18837 ;
    wire new_AGEMA_signal_18838 ;
    wire new_AGEMA_signal_18839 ;
    wire new_AGEMA_signal_18840 ;
    wire new_AGEMA_signal_18841 ;
    wire new_AGEMA_signal_18842 ;
    wire new_AGEMA_signal_18843 ;
    wire new_AGEMA_signal_18844 ;
    wire new_AGEMA_signal_18845 ;
    wire new_AGEMA_signal_18846 ;
    wire new_AGEMA_signal_18847 ;
    wire new_AGEMA_signal_18848 ;
    wire new_AGEMA_signal_18849 ;
    wire new_AGEMA_signal_18850 ;
    wire new_AGEMA_signal_18851 ;
    wire new_AGEMA_signal_18852 ;
    wire new_AGEMA_signal_18853 ;
    wire new_AGEMA_signal_18854 ;
    wire new_AGEMA_signal_18855 ;
    wire new_AGEMA_signal_18856 ;
    wire new_AGEMA_signal_18857 ;
    wire new_AGEMA_signal_18858 ;
    wire new_AGEMA_signal_18859 ;
    wire new_AGEMA_signal_18860 ;
    wire new_AGEMA_signal_18861 ;
    wire new_AGEMA_signal_18862 ;
    wire new_AGEMA_signal_18863 ;
    wire new_AGEMA_signal_18864 ;
    wire new_AGEMA_signal_18865 ;
    wire new_AGEMA_signal_18866 ;
    wire new_AGEMA_signal_18867 ;
    wire new_AGEMA_signal_18868 ;
    wire new_AGEMA_signal_18869 ;
    wire new_AGEMA_signal_18870 ;
    wire new_AGEMA_signal_18871 ;
    wire new_AGEMA_signal_18872 ;
    wire new_AGEMA_signal_18873 ;
    wire new_AGEMA_signal_18874 ;
    wire new_AGEMA_signal_18875 ;
    wire new_AGEMA_signal_18876 ;
    wire new_AGEMA_signal_18877 ;
    wire new_AGEMA_signal_18878 ;
    wire new_AGEMA_signal_18879 ;
    wire new_AGEMA_signal_18880 ;
    wire new_AGEMA_signal_18881 ;
    wire new_AGEMA_signal_18882 ;
    wire new_AGEMA_signal_18883 ;
    wire new_AGEMA_signal_18884 ;
    wire new_AGEMA_signal_18885 ;
    wire new_AGEMA_signal_18886 ;
    wire new_AGEMA_signal_18887 ;
    wire new_AGEMA_signal_18888 ;
    wire new_AGEMA_signal_18889 ;
    wire new_AGEMA_signal_18890 ;
    wire new_AGEMA_signal_18891 ;
    wire new_AGEMA_signal_18892 ;
    wire new_AGEMA_signal_18893 ;
    wire new_AGEMA_signal_18894 ;
    wire new_AGEMA_signal_18895 ;
    wire new_AGEMA_signal_18896 ;
    wire new_AGEMA_signal_18897 ;
    wire new_AGEMA_signal_18898 ;
    wire new_AGEMA_signal_18899 ;
    wire new_AGEMA_signal_18900 ;
    wire new_AGEMA_signal_18901 ;
    wire new_AGEMA_signal_18902 ;
    wire new_AGEMA_signal_18903 ;
    wire new_AGEMA_signal_18904 ;
    wire new_AGEMA_signal_18905 ;
    wire new_AGEMA_signal_18906 ;
    wire new_AGEMA_signal_18907 ;
    wire new_AGEMA_signal_18908 ;
    wire new_AGEMA_signal_18909 ;
    wire new_AGEMA_signal_18910 ;
    wire new_AGEMA_signal_18911 ;
    wire new_AGEMA_signal_18912 ;
    wire new_AGEMA_signal_18913 ;
    wire new_AGEMA_signal_18914 ;
    wire new_AGEMA_signal_18915 ;
    wire new_AGEMA_signal_18916 ;
    wire new_AGEMA_signal_18917 ;
    wire new_AGEMA_signal_18918 ;
    wire new_AGEMA_signal_18919 ;
    wire new_AGEMA_signal_18920 ;
    wire new_AGEMA_signal_18921 ;
    wire new_AGEMA_signal_18922 ;
    wire new_AGEMA_signal_18923 ;
    wire new_AGEMA_signal_18924 ;
    wire new_AGEMA_signal_18925 ;
    wire new_AGEMA_signal_18926 ;
    wire new_AGEMA_signal_18927 ;
    wire new_AGEMA_signal_18928 ;
    wire new_AGEMA_signal_18929 ;
    wire new_AGEMA_signal_18930 ;
    wire new_AGEMA_signal_18931 ;
    wire new_AGEMA_signal_18932 ;
    wire new_AGEMA_signal_18933 ;
    wire new_AGEMA_signal_18934 ;
    wire new_AGEMA_signal_18935 ;
    wire new_AGEMA_signal_18936 ;
    wire new_AGEMA_signal_18937 ;
    wire new_AGEMA_signal_18938 ;
    wire new_AGEMA_signal_18939 ;
    wire new_AGEMA_signal_18940 ;
    wire new_AGEMA_signal_18941 ;
    wire new_AGEMA_signal_18942 ;
    wire new_AGEMA_signal_18943 ;
    wire new_AGEMA_signal_18944 ;
    wire new_AGEMA_signal_18945 ;
    wire new_AGEMA_signal_18946 ;
    wire new_AGEMA_signal_18947 ;
    wire new_AGEMA_signal_18948 ;
    wire new_AGEMA_signal_18949 ;
    wire new_AGEMA_signal_18950 ;
    wire new_AGEMA_signal_18951 ;
    wire new_AGEMA_signal_18952 ;
    wire new_AGEMA_signal_18953 ;
    wire new_AGEMA_signal_18954 ;
    wire new_AGEMA_signal_18955 ;
    wire new_AGEMA_signal_18956 ;
    wire new_AGEMA_signal_18957 ;
    wire new_AGEMA_signal_18958 ;
    wire new_AGEMA_signal_18959 ;
    wire new_AGEMA_signal_18960 ;
    wire new_AGEMA_signal_18961 ;
    wire new_AGEMA_signal_18962 ;
    wire new_AGEMA_signal_18963 ;
    wire new_AGEMA_signal_18964 ;
    wire new_AGEMA_signal_18965 ;
    wire new_AGEMA_signal_18966 ;
    wire new_AGEMA_signal_18967 ;
    wire new_AGEMA_signal_18968 ;
    wire new_AGEMA_signal_18969 ;
    wire new_AGEMA_signal_18970 ;
    wire new_AGEMA_signal_18971 ;
    wire new_AGEMA_signal_18972 ;
    wire new_AGEMA_signal_18973 ;
    wire new_AGEMA_signal_18974 ;
    wire new_AGEMA_signal_18975 ;
    wire new_AGEMA_signal_18976 ;
    wire new_AGEMA_signal_18977 ;
    wire new_AGEMA_signal_18978 ;
    wire new_AGEMA_signal_18979 ;
    wire new_AGEMA_signal_18980 ;
    wire new_AGEMA_signal_18981 ;
    wire new_AGEMA_signal_18982 ;
    wire new_AGEMA_signal_18983 ;
    wire new_AGEMA_signal_18984 ;
    wire new_AGEMA_signal_18985 ;
    wire new_AGEMA_signal_18986 ;
    wire new_AGEMA_signal_18987 ;
    wire new_AGEMA_signal_18988 ;
    wire new_AGEMA_signal_18989 ;
    wire new_AGEMA_signal_18990 ;
    wire new_AGEMA_signal_18991 ;
    wire new_AGEMA_signal_18992 ;
    wire new_AGEMA_signal_18993 ;
    wire new_AGEMA_signal_18994 ;
    wire new_AGEMA_signal_18995 ;
    wire new_AGEMA_signal_18996 ;
    wire new_AGEMA_signal_18997 ;
    wire new_AGEMA_signal_18998 ;
    wire new_AGEMA_signal_18999 ;
    wire new_AGEMA_signal_19000 ;
    wire new_AGEMA_signal_19001 ;
    wire new_AGEMA_signal_19002 ;
    wire new_AGEMA_signal_19003 ;
    wire new_AGEMA_signal_19004 ;
    wire new_AGEMA_signal_19005 ;
    wire new_AGEMA_signal_19006 ;
    wire new_AGEMA_signal_19007 ;
    wire new_AGEMA_signal_19008 ;
    wire new_AGEMA_signal_19009 ;
    wire new_AGEMA_signal_19010 ;
    wire new_AGEMA_signal_19011 ;
    wire new_AGEMA_signal_19012 ;
    wire new_AGEMA_signal_19013 ;
    wire new_AGEMA_signal_19014 ;
    wire new_AGEMA_signal_19015 ;
    wire new_AGEMA_signal_19016 ;
    wire new_AGEMA_signal_19017 ;
    wire new_AGEMA_signal_19018 ;
    wire new_AGEMA_signal_19019 ;
    wire new_AGEMA_signal_19020 ;
    wire new_AGEMA_signal_19021 ;
    wire new_AGEMA_signal_19022 ;
    wire new_AGEMA_signal_19023 ;
    wire new_AGEMA_signal_19024 ;
    wire new_AGEMA_signal_19025 ;
    wire new_AGEMA_signal_19026 ;
    wire new_AGEMA_signal_19027 ;
    wire new_AGEMA_signal_19028 ;
    wire new_AGEMA_signal_19029 ;
    wire new_AGEMA_signal_19030 ;
    wire new_AGEMA_signal_19031 ;
    wire new_AGEMA_signal_19032 ;
    wire new_AGEMA_signal_19033 ;
    wire new_AGEMA_signal_19034 ;
    wire new_AGEMA_signal_19035 ;
    wire new_AGEMA_signal_19036 ;
    wire new_AGEMA_signal_19037 ;
    wire new_AGEMA_signal_19038 ;
    wire new_AGEMA_signal_19039 ;
    wire new_AGEMA_signal_19040 ;
    wire new_AGEMA_signal_19041 ;
    wire new_AGEMA_signal_19042 ;
    wire new_AGEMA_signal_19043 ;
    wire new_AGEMA_signal_19044 ;
    wire new_AGEMA_signal_19045 ;
    wire new_AGEMA_signal_19046 ;
    wire new_AGEMA_signal_19047 ;
    wire new_AGEMA_signal_19048 ;
    wire new_AGEMA_signal_19049 ;
    wire new_AGEMA_signal_19050 ;
    wire new_AGEMA_signal_19051 ;
    wire new_AGEMA_signal_19052 ;
    wire new_AGEMA_signal_19053 ;
    wire new_AGEMA_signal_19054 ;
    wire new_AGEMA_signal_19055 ;
    wire new_AGEMA_signal_19056 ;
    wire new_AGEMA_signal_19057 ;
    wire new_AGEMA_signal_19058 ;
    wire new_AGEMA_signal_19059 ;
    wire new_AGEMA_signal_19060 ;
    wire new_AGEMA_signal_19061 ;
    wire new_AGEMA_signal_19062 ;
    wire new_AGEMA_signal_19063 ;
    wire new_AGEMA_signal_19064 ;
    wire new_AGEMA_signal_19065 ;
    wire new_AGEMA_signal_19066 ;
    wire new_AGEMA_signal_19067 ;
    wire new_AGEMA_signal_19068 ;
    wire new_AGEMA_signal_19069 ;
    wire new_AGEMA_signal_19070 ;
    wire new_AGEMA_signal_19071 ;
    wire new_AGEMA_signal_19072 ;
    wire new_AGEMA_signal_19073 ;
    wire new_AGEMA_signal_19074 ;
    wire new_AGEMA_signal_19075 ;
    wire new_AGEMA_signal_19076 ;
    wire new_AGEMA_signal_19077 ;
    wire new_AGEMA_signal_19078 ;
    wire new_AGEMA_signal_19079 ;
    wire new_AGEMA_signal_19080 ;
    wire new_AGEMA_signal_19081 ;
    wire new_AGEMA_signal_19082 ;
    wire new_AGEMA_signal_19083 ;
    wire new_AGEMA_signal_19084 ;
    wire new_AGEMA_signal_19085 ;
    wire new_AGEMA_signal_19086 ;
    wire new_AGEMA_signal_19087 ;
    wire new_AGEMA_signal_19088 ;
    wire new_AGEMA_signal_19089 ;
    wire new_AGEMA_signal_19090 ;
    wire new_AGEMA_signal_19091 ;
    wire new_AGEMA_signal_19092 ;
    wire new_AGEMA_signal_19093 ;
    wire new_AGEMA_signal_19094 ;
    wire new_AGEMA_signal_19095 ;
    wire new_AGEMA_signal_19096 ;
    wire new_AGEMA_signal_19097 ;
    wire new_AGEMA_signal_19098 ;
    wire new_AGEMA_signal_19099 ;
    wire new_AGEMA_signal_19100 ;
    wire new_AGEMA_signal_19101 ;
    wire new_AGEMA_signal_19102 ;
    wire new_AGEMA_signal_19103 ;
    wire new_AGEMA_signal_19104 ;
    wire new_AGEMA_signal_19105 ;
    wire new_AGEMA_signal_19106 ;
    wire new_AGEMA_signal_19107 ;
    wire new_AGEMA_signal_19108 ;
    wire new_AGEMA_signal_19109 ;
    wire new_AGEMA_signal_19110 ;
    wire new_AGEMA_signal_19111 ;
    wire new_AGEMA_signal_19112 ;
    wire new_AGEMA_signal_19113 ;
    wire new_AGEMA_signal_19114 ;
    wire new_AGEMA_signal_19115 ;
    wire new_AGEMA_signal_19116 ;
    wire new_AGEMA_signal_19117 ;
    wire new_AGEMA_signal_19118 ;
    wire new_AGEMA_signal_19119 ;
    wire new_AGEMA_signal_19120 ;
    wire new_AGEMA_signal_19121 ;
    wire new_AGEMA_signal_19122 ;
    wire new_AGEMA_signal_19123 ;
    wire new_AGEMA_signal_19124 ;
    wire new_AGEMA_signal_19125 ;
    wire new_AGEMA_signal_19126 ;
    wire new_AGEMA_signal_19127 ;
    wire new_AGEMA_signal_19128 ;
    wire new_AGEMA_signal_19129 ;
    wire new_AGEMA_signal_19130 ;
    wire new_AGEMA_signal_19131 ;
    wire new_AGEMA_signal_19132 ;
    wire new_AGEMA_signal_19133 ;
    wire new_AGEMA_signal_19134 ;
    wire new_AGEMA_signal_19135 ;
    wire new_AGEMA_signal_19136 ;
    wire new_AGEMA_signal_19137 ;
    wire new_AGEMA_signal_19138 ;
    wire new_AGEMA_signal_19139 ;
    wire new_AGEMA_signal_19140 ;
    wire new_AGEMA_signal_19141 ;
    wire new_AGEMA_signal_19142 ;
    wire new_AGEMA_signal_19143 ;
    wire new_AGEMA_signal_19144 ;
    wire new_AGEMA_signal_19145 ;
    wire new_AGEMA_signal_19146 ;
    wire new_AGEMA_signal_19147 ;
    wire new_AGEMA_signal_19148 ;
    wire new_AGEMA_signal_19149 ;
    wire new_AGEMA_signal_19150 ;
    wire new_AGEMA_signal_19151 ;
    wire new_AGEMA_signal_19152 ;
    wire new_AGEMA_signal_19153 ;
    wire new_AGEMA_signal_19154 ;
    wire new_AGEMA_signal_19155 ;
    wire new_AGEMA_signal_19156 ;
    wire new_AGEMA_signal_19157 ;
    wire new_AGEMA_signal_19158 ;
    wire new_AGEMA_signal_19159 ;
    wire new_AGEMA_signal_19160 ;
    wire new_AGEMA_signal_19161 ;
    wire new_AGEMA_signal_19162 ;

    /* cells in depth 0 */
    not_masked #(.security_order(3), .pipeline(1)) U1938 ( .a ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({new_AGEMA_signal_947, new_AGEMA_signal_946, new_AGEMA_signal_945, n2796}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1939 ( .a ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({new_AGEMA_signal_953, new_AGEMA_signal_952, new_AGEMA_signal_951, n2810}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1940 ( .a ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({new_AGEMA_signal_959, new_AGEMA_signal_958, new_AGEMA_signal_957, n2462}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1941 ( .a ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, n2760}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1942 ( .a ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({new_AGEMA_signal_971, new_AGEMA_signal_970, new_AGEMA_signal_969, n2791}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1944 ( .a ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1945 ( .a ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({new_AGEMA_signal_983, new_AGEMA_signal_982, new_AGEMA_signal_981, n2630}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1946 ( .a ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}) ) ;

    /* cells in depth 1 */
    buf_clk new_AGEMA_reg_buffer_927 ( .C ( clk ), .D ( SI_s0[4] ), .Q ( new_AGEMA_signal_12427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_929 ( .C ( clk ), .D ( SI_s1[4] ), .Q ( new_AGEMA_signal_12429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_931 ( .C ( clk ), .D ( SI_s2[4] ), .Q ( new_AGEMA_signal_12431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_933 ( .C ( clk ), .D ( SI_s3[4] ), .Q ( new_AGEMA_signal_12433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_935 ( .C ( clk ), .D ( SI_s0[6] ), .Q ( new_AGEMA_signal_12435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_937 ( .C ( clk ), .D ( SI_s1[6] ), .Q ( new_AGEMA_signal_12437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_939 ( .C ( clk ), .D ( SI_s2[6] ), .Q ( new_AGEMA_signal_12439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_941 ( .C ( clk ), .D ( SI_s3[6] ), .Q ( new_AGEMA_signal_12441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_943 ( .C ( clk ), .D ( SI_s0[7] ), .Q ( new_AGEMA_signal_12443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_945 ( .C ( clk ), .D ( SI_s1[7] ), .Q ( new_AGEMA_signal_12445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_947 ( .C ( clk ), .D ( SI_s2[7] ), .Q ( new_AGEMA_signal_12447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_949 ( .C ( clk ), .D ( SI_s3[7] ), .Q ( new_AGEMA_signal_12449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_951 ( .C ( clk ), .D ( SI_s0[0] ), .Q ( new_AGEMA_signal_12451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_953 ( .C ( clk ), .D ( SI_s1[0] ), .Q ( new_AGEMA_signal_12453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_955 ( .C ( clk ), .D ( SI_s2[0] ), .Q ( new_AGEMA_signal_12455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_957 ( .C ( clk ), .D ( SI_s3[0] ), .Q ( new_AGEMA_signal_12457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_959 ( .C ( clk ), .D ( SI_s0[1] ), .Q ( new_AGEMA_signal_12459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_961 ( .C ( clk ), .D ( SI_s1[1] ), .Q ( new_AGEMA_signal_12461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_963 ( .C ( clk ), .D ( SI_s2[1] ), .Q ( new_AGEMA_signal_12463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_965 ( .C ( clk ), .D ( SI_s3[1] ), .Q ( new_AGEMA_signal_12465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_967 ( .C ( clk ), .D ( n2630 ), .Q ( new_AGEMA_signal_12467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_969 ( .C ( clk ), .D ( new_AGEMA_signal_981 ), .Q ( new_AGEMA_signal_12469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_971 ( .C ( clk ), .D ( new_AGEMA_signal_982 ), .Q ( new_AGEMA_signal_12471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_973 ( .C ( clk ), .D ( new_AGEMA_signal_983 ), .Q ( new_AGEMA_signal_12473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_975 ( .C ( clk ), .D ( SI_s0[5] ), .Q ( new_AGEMA_signal_12475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_977 ( .C ( clk ), .D ( SI_s1[5] ), .Q ( new_AGEMA_signal_12477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_979 ( .C ( clk ), .D ( SI_s2[5] ), .Q ( new_AGEMA_signal_12479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_981 ( .C ( clk ), .D ( SI_s3[5] ), .Q ( new_AGEMA_signal_12481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_983 ( .C ( clk ), .D ( n2462 ), .Q ( new_AGEMA_signal_12483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_985 ( .C ( clk ), .D ( new_AGEMA_signal_957 ), .Q ( new_AGEMA_signal_12485 ) ) ;
    buf_clk new_AGEMA_reg_buffer_987 ( .C ( clk ), .D ( new_AGEMA_signal_958 ), .Q ( new_AGEMA_signal_12487 ) ) ;
    buf_clk new_AGEMA_reg_buffer_989 ( .C ( clk ), .D ( new_AGEMA_signal_959 ), .Q ( new_AGEMA_signal_12489 ) ) ;
    buf_clk new_AGEMA_reg_buffer_991 ( .C ( clk ), .D ( n2760 ), .Q ( new_AGEMA_signal_12491 ) ) ;
    buf_clk new_AGEMA_reg_buffer_993 ( .C ( clk ), .D ( new_AGEMA_signal_963 ), .Q ( new_AGEMA_signal_12493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_995 ( .C ( clk ), .D ( new_AGEMA_signal_964 ), .Q ( new_AGEMA_signal_12495 ) ) ;
    buf_clk new_AGEMA_reg_buffer_997 ( .C ( clk ), .D ( new_AGEMA_signal_965 ), .Q ( new_AGEMA_signal_12497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_999 ( .C ( clk ), .D ( n2796 ), .Q ( new_AGEMA_signal_12499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1001 ( .C ( clk ), .D ( new_AGEMA_signal_945 ), .Q ( new_AGEMA_signal_12501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1003 ( .C ( clk ), .D ( new_AGEMA_signal_946 ), .Q ( new_AGEMA_signal_12503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1005 ( .C ( clk ), .D ( new_AGEMA_signal_947 ), .Q ( new_AGEMA_signal_12505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1007 ( .C ( clk ), .D ( n2765 ), .Q ( new_AGEMA_signal_12507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1009 ( .C ( clk ), .D ( new_AGEMA_signal_987 ), .Q ( new_AGEMA_signal_12509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1011 ( .C ( clk ), .D ( new_AGEMA_signal_988 ), .Q ( new_AGEMA_signal_12511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1013 ( .C ( clk ), .D ( new_AGEMA_signal_989 ), .Q ( new_AGEMA_signal_12513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1015 ( .C ( clk ), .D ( n2791 ), .Q ( new_AGEMA_signal_12515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1017 ( .C ( clk ), .D ( new_AGEMA_signal_969 ), .Q ( new_AGEMA_signal_12517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1019 ( .C ( clk ), .D ( new_AGEMA_signal_970 ), .Q ( new_AGEMA_signal_12519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1021 ( .C ( clk ), .D ( new_AGEMA_signal_971 ), .Q ( new_AGEMA_signal_12521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1023 ( .C ( clk ), .D ( SI_s0[3] ), .Q ( new_AGEMA_signal_12523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1025 ( .C ( clk ), .D ( SI_s1[3] ), .Q ( new_AGEMA_signal_12525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1027 ( .C ( clk ), .D ( SI_s2[3] ), .Q ( new_AGEMA_signal_12527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1029 ( .C ( clk ), .D ( SI_s3[3] ), .Q ( new_AGEMA_signal_12529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1031 ( .C ( clk ), .D ( n2813 ), .Q ( new_AGEMA_signal_12531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1033 ( .C ( clk ), .D ( new_AGEMA_signal_975 ), .Q ( new_AGEMA_signal_12533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1035 ( .C ( clk ), .D ( new_AGEMA_signal_976 ), .Q ( new_AGEMA_signal_12535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1037 ( .C ( clk ), .D ( new_AGEMA_signal_977 ), .Q ( new_AGEMA_signal_12537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1039 ( .C ( clk ), .D ( n2810 ), .Q ( new_AGEMA_signal_12539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1041 ( .C ( clk ), .D ( new_AGEMA_signal_951 ), .Q ( new_AGEMA_signal_12541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1043 ( .C ( clk ), .D ( new_AGEMA_signal_952 ), .Q ( new_AGEMA_signal_12543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1045 ( .C ( clk ), .D ( new_AGEMA_signal_953 ), .Q ( new_AGEMA_signal_12545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2071 ( .C ( clk ), .D ( SI_s0[2] ), .Q ( new_AGEMA_signal_13571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2077 ( .C ( clk ), .D ( SI_s1[2] ), .Q ( new_AGEMA_signal_13577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2083 ( .C ( clk ), .D ( SI_s2[2] ), .Q ( new_AGEMA_signal_13583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2089 ( .C ( clk ), .D ( SI_s3[2] ), .Q ( new_AGEMA_signal_13589 ) ) ;

    /* cells in depth 2 */
    nor_HPC1 #(.security_order(3), .pipeline(1)) U1937 ( .ina ({new_AGEMA_signal_947, new_AGEMA_signal_946, new_AGEMA_signal_945, n2796}), .inb ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .clk ( clk ), .rnd ({Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .outt ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2719}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1943 ( .a ({new_AGEMA_signal_1127, new_AGEMA_signal_1126, new_AGEMA_signal_1125, n2624}), .b ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U1947 ( .ina ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .inb ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .rnd ({Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10]}), .outt ({new_AGEMA_signal_992, new_AGEMA_signal_991, new_AGEMA_signal_990, n2635}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U1948 ( .ina ({new_AGEMA_signal_959, new_AGEMA_signal_958, new_AGEMA_signal_957, n2462}), .inb ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .clk ( clk ), .rnd ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20]}), .outt ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, new_AGEMA_signal_1029, n2641}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U1949 ( .ina ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .inb ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .outt ({new_AGEMA_signal_995, new_AGEMA_signal_994, new_AGEMA_signal_993, n2790}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U1950 ( .ina ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .inb ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .clk ( clk ), .rnd ({Fresh[49], Fresh[48], Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40]}), .outt ({new_AGEMA_signal_998, new_AGEMA_signal_997, new_AGEMA_signal_996, n2519}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1951 ( .a ({new_AGEMA_signal_998, new_AGEMA_signal_997, new_AGEMA_signal_996, n2519}), .b ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, new_AGEMA_signal_1032, n2750}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U1952 ( .ina ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, n2760}), .inb ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50]}), .outt ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, new_AGEMA_signal_1035, n2615}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1953 ( .a ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, new_AGEMA_signal_1035, n2615}), .b ({new_AGEMA_signal_1190, new_AGEMA_signal_1189, new_AGEMA_signal_1188, n2640}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U1955 ( .ina ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .inb ({new_AGEMA_signal_983, new_AGEMA_signal_982, new_AGEMA_signal_981, n2630}), .clk ( clk ), .rnd ({Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .outt ({new_AGEMA_signal_1040, new_AGEMA_signal_1039, new_AGEMA_signal_1038, n2699}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1956 ( .a ({new_AGEMA_signal_1040, new_AGEMA_signal_1039, new_AGEMA_signal_1038, n2699}), .b ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, new_AGEMA_signal_1191, n2737}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U1957 ( .ina ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .inb ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}), .clk ( clk ), .rnd ({Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72], Fresh[71], Fresh[70]}), .outt ({new_AGEMA_signal_1043, new_AGEMA_signal_1042, new_AGEMA_signal_1041, n2816}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1958 ( .a ({new_AGEMA_signal_1043, new_AGEMA_signal_1042, new_AGEMA_signal_1041, n2816}), .b ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2767}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U1961 ( .ina ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .inb ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .rnd ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84], Fresh[83], Fresh[82], Fresh[81], Fresh[80]}), .outt ({new_AGEMA_signal_1046, new_AGEMA_signal_1045, new_AGEMA_signal_1044, n2780}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1962 ( .a ({new_AGEMA_signal_1046, new_AGEMA_signal_1045, new_AGEMA_signal_1044, n2780}), .b ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, new_AGEMA_signal_1197, n2789}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U1963 ( .ina ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .inb ({new_AGEMA_signal_953, new_AGEMA_signal_952, new_AGEMA_signal_951, n2810}), .clk ( clk ), .rnd ({Fresh[99], Fresh[98], Fresh[97], Fresh[96], Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .outt ({new_AGEMA_signal_1049, new_AGEMA_signal_1048, new_AGEMA_signal_1047, n2317}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U1965 ( .ina ({new_AGEMA_signal_971, new_AGEMA_signal_970, new_AGEMA_signal_969, n2791}), .inb ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, n2760}), .clk ( clk ), .rnd ({Fresh[109], Fresh[108], Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100]}), .outt ({new_AGEMA_signal_1052, new_AGEMA_signal_1051, new_AGEMA_signal_1050, n2694}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1966 ( .a ({new_AGEMA_signal_1052, new_AGEMA_signal_1051, new_AGEMA_signal_1050, n2694}), .b ({new_AGEMA_signal_1202, new_AGEMA_signal_1201, new_AGEMA_signal_1200, n2769}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U1969 ( .ina ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, n2760}), .inb ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .clk ( clk ), .rnd ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114], Fresh[113], Fresh[112], Fresh[111], Fresh[110]}), .outt ({new_AGEMA_signal_1055, new_AGEMA_signal_1054, new_AGEMA_signal_1053, n2073}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1970 ( .a ({new_AGEMA_signal_1055, new_AGEMA_signal_1054, new_AGEMA_signal_1053, n2073}), .b ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U1971 ( .ina ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .inb ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[129], Fresh[128], Fresh[127], Fresh[126], Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .outt ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, new_AGEMA_signal_999, n2315}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U1972 ( .ina ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .inb ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .rnd ({Fresh[139], Fresh[138], Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132], Fresh[131], Fresh[130]}), .outt ({new_AGEMA_signal_1004, new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2682}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1973 ( .a ({new_AGEMA_signal_1004, new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2682}), .b ({new_AGEMA_signal_1058, new_AGEMA_signal_1057, new_AGEMA_signal_1056, n2713}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U1975 ( .ina ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}), .inb ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .rnd ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144], Fresh[143], Fresh[142], Fresh[141], Fresh[140]}), .outt ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, new_AGEMA_signal_1059, n2723}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1976 ( .a ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, new_AGEMA_signal_1059, n2723}), .b ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, new_AGEMA_signal_1209, n2688}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U1978 ( .ina ({new_AGEMA_signal_953, new_AGEMA_signal_952, new_AGEMA_signal_951, n2810}), .inb ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .clk ( clk ), .rnd ({Fresh[159], Fresh[158], Fresh[157], Fresh[156], Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .outt ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2725}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1979 ( .a ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2725}), .b ({new_AGEMA_signal_1214, new_AGEMA_signal_1213, new_AGEMA_signal_1212, n2541}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U1984 ( .ina ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, n2760}), .inb ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .clk ( clk ), .rnd ({Fresh[169], Fresh[168], Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162], Fresh[161], Fresh[160]}), .outt ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, new_AGEMA_signal_1065, n2815}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1985 ( .a ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, new_AGEMA_signal_1065, n2815}), .b ({new_AGEMA_signal_1217, new_AGEMA_signal_1216, new_AGEMA_signal_1215, n2086}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U1987 ( .ina ({new_AGEMA_signal_953, new_AGEMA_signal_952, new_AGEMA_signal_951, n2810}), .inb ({new_AGEMA_signal_971, new_AGEMA_signal_970, new_AGEMA_signal_969, n2791}), .clk ( clk ), .rnd ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174], Fresh[173], Fresh[172], Fresh[171], Fresh[170]}), .outt ({new_AGEMA_signal_1070, new_AGEMA_signal_1069, new_AGEMA_signal_1068, n2600}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U1990 ( .ina ({new_AGEMA_signal_959, new_AGEMA_signal_958, new_AGEMA_signal_957, n2462}), .inb ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[189], Fresh[188], Fresh[187], Fresh[186], Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .outt ({new_AGEMA_signal_1073, new_AGEMA_signal_1072, new_AGEMA_signal_1071, n2538}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1991 ( .a ({new_AGEMA_signal_1073, new_AGEMA_signal_1072, new_AGEMA_signal_1071, n2538}), .b ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, n2786}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U1995 ( .ina ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .inb ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .rnd ({Fresh[199], Fresh[198], Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192], Fresh[191], Fresh[190]}), .outt ({new_AGEMA_signal_1007, new_AGEMA_signal_1006, new_AGEMA_signal_1005, n2595}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1996 ( .a ({new_AGEMA_signal_1007, new_AGEMA_signal_1006, new_AGEMA_signal_1005, n2595}), .b ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2742}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U1999 ( .ina ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .inb ({new_AGEMA_signal_983, new_AGEMA_signal_982, new_AGEMA_signal_981, n2630}), .clk ( clk ), .rnd ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204], Fresh[203], Fresh[202], Fresh[201], Fresh[200]}), .outt ({new_AGEMA_signal_1079, new_AGEMA_signal_1078, new_AGEMA_signal_1077, n2753}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2000 ( .a ({new_AGEMA_signal_1079, new_AGEMA_signal_1078, new_AGEMA_signal_1077, n2753}), .b ({new_AGEMA_signal_1229, new_AGEMA_signal_1228, new_AGEMA_signal_1227, n2577}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2004 ( .ina ({new_AGEMA_signal_953, new_AGEMA_signal_952, new_AGEMA_signal_951, n2810}), .inb ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .clk ( clk ), .rnd ({Fresh[219], Fresh[218], Fresh[217], Fresh[216], Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .outt ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, new_AGEMA_signal_1080, n2400}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2008 ( .ina ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .inb ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .rnd ({Fresh[229], Fresh[228], Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222], Fresh[221], Fresh[220]}), .outt ({new_AGEMA_signal_1085, new_AGEMA_signal_1084, new_AGEMA_signal_1083, n2785}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2009 ( .a ({new_AGEMA_signal_1085, new_AGEMA_signal_1084, new_AGEMA_signal_1083, n2785}), .b ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, n2792}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2013 ( .ina ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}), .inb ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .rnd ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234], Fresh[233], Fresh[232], Fresh[231], Fresh[230]}), .outt ({new_AGEMA_signal_1088, new_AGEMA_signal_1087, new_AGEMA_signal_1086, n2609}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2014 ( .a ({new_AGEMA_signal_1088, new_AGEMA_signal_1087, new_AGEMA_signal_1086, n2609}), .b ({new_AGEMA_signal_1238, new_AGEMA_signal_1237, new_AGEMA_signal_1236, n2724}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2017 ( .ina ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, n2760}), .inb ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}), .clk ( clk ), .rnd ({Fresh[249], Fresh[248], Fresh[247], Fresh[246], Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .outt ({new_AGEMA_signal_1091, new_AGEMA_signal_1090, new_AGEMA_signal_1089, n2661}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2018 ( .a ({new_AGEMA_signal_1091, new_AGEMA_signal_1090, new_AGEMA_signal_1089, n2661}), .b ({new_AGEMA_signal_1241, new_AGEMA_signal_1240, new_AGEMA_signal_1239, n2174}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2020 ( .ina ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .inb ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .rnd ({Fresh[259], Fresh[258], Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252], Fresh[251], Fresh[250]}), .outt ({new_AGEMA_signal_1010, new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2708}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2021 ( .a ({new_AGEMA_signal_1010, new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2708}), .b ({new_AGEMA_signal_1094, new_AGEMA_signal_1093, new_AGEMA_signal_1092, n2493}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2025 ( .ina ({new_AGEMA_signal_947, new_AGEMA_signal_946, new_AGEMA_signal_945, n2796}), .inb ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264], Fresh[263], Fresh[262], Fresh[261], Fresh[260]}), .outt ({new_AGEMA_signal_1097, new_AGEMA_signal_1096, new_AGEMA_signal_1095, n2587}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2028 ( .a ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2719}), .b ({new_AGEMA_signal_1250, new_AGEMA_signal_1249, new_AGEMA_signal_1248, n2570}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2029 ( .ina ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .inb ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .rnd ({Fresh[279], Fresh[278], Fresh[277], Fresh[276], Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .outt ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, new_AGEMA_signal_1011, n2559}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2035 ( .ina ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .inb ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .rnd ({Fresh[289], Fresh[288], Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282], Fresh[281], Fresh[280]}), .outt ({new_AGEMA_signal_1100, new_AGEMA_signal_1099, new_AGEMA_signal_1098, n2643}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2036 ( .a ({new_AGEMA_signal_1100, new_AGEMA_signal_1099, new_AGEMA_signal_1098, n2643}), .b ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, n2442}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2038 ( .a ({new_AGEMA_signal_995, new_AGEMA_signal_994, new_AGEMA_signal_993, n2790}), .b ({new_AGEMA_signal_1103, new_AGEMA_signal_1102, new_AGEMA_signal_1101, n2739}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2044 ( .ina ({new_AGEMA_signal_959, new_AGEMA_signal_958, new_AGEMA_signal_957, n2462}), .inb ({new_AGEMA_signal_947, new_AGEMA_signal_946, new_AGEMA_signal_945, n2796}), .clk ( clk ), .rnd ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294], Fresh[293], Fresh[292], Fresh[291], Fresh[290]}), .outt ({new_AGEMA_signal_1106, new_AGEMA_signal_1105, new_AGEMA_signal_1104, n2437}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2045 ( .ina ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .inb ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .clk ( clk ), .rnd ({Fresh[309], Fresh[308], Fresh[307], Fresh[306], Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .outt ({new_AGEMA_signal_1016, new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2261}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2046 ( .a ({new_AGEMA_signal_1016, new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2261}), .b ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, new_AGEMA_signal_1107, n2778}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2052 ( .ina ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .inb ({new_AGEMA_signal_971, new_AGEMA_signal_970, new_AGEMA_signal_969, n2791}), .clk ( clk ), .rnd ({Fresh[319], Fresh[318], Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312], Fresh[311], Fresh[310]}), .outt ({new_AGEMA_signal_1112, new_AGEMA_signal_1111, new_AGEMA_signal_1110, n2452}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2055 ( .a ({new_AGEMA_signal_1106, new_AGEMA_signal_1105, new_AGEMA_signal_1104, n2437}), .b ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2766}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2068 ( .ina ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .inb ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .rnd ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324], Fresh[323], Fresh[322], Fresh[321], Fresh[320]}), .outt ({new_AGEMA_signal_1118, new_AGEMA_signal_1117, new_AGEMA_signal_1116, n2772}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2070 ( .ina ({new_AGEMA_signal_971, new_AGEMA_signal_970, new_AGEMA_signal_969, n2791}), .inb ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[339], Fresh[338], Fresh[337], Fresh[336], Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .outt ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, new_AGEMA_signal_1119, n2824}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2071 ( .a ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, new_AGEMA_signal_1119, n2824}), .b ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, n2612}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2074 ( .a ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, new_AGEMA_signal_1080, n2400}), .b ({new_AGEMA_signal_1280, new_AGEMA_signal_1279, new_AGEMA_signal_1278, n2313}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2089 ( .ina ({new_AGEMA_signal_953, new_AGEMA_signal_952, new_AGEMA_signal_951, n2810}), .inb ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, n2760}), .clk ( clk ), .rnd ({Fresh[349], Fresh[348], Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342], Fresh[341], Fresh[340]}), .outt ({new_AGEMA_signal_1124, new_AGEMA_signal_1123, new_AGEMA_signal_1122, n2395}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2090 ( .a ({new_AGEMA_signal_1124, new_AGEMA_signal_1123, new_AGEMA_signal_1122, n2395}), .b ({new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2818}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2094 ( .ina ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .inb ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354], Fresh[353], Fresh[352], Fresh[351], Fresh[350]}), .outt ({new_AGEMA_signal_1019, new_AGEMA_signal_1018, new_AGEMA_signal_1017, n2779}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2096 ( .ina ({new_AGEMA_signal_983, new_AGEMA_signal_982, new_AGEMA_signal_981, n2630}), .inb ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}), .clk ( clk ), .rnd ({Fresh[369], Fresh[368], Fresh[367], Fresh[366], Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .outt ({new_AGEMA_signal_1127, new_AGEMA_signal_1126, new_AGEMA_signal_1125, n2624}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2097 ( .ina ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .inb ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .rnd ({Fresh[379], Fresh[378], Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372], Fresh[371], Fresh[370]}), .outt ({new_AGEMA_signal_1022, new_AGEMA_signal_1021, new_AGEMA_signal_1020, n2242}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2100 ( .ina ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .inb ({new_AGEMA_signal_971, new_AGEMA_signal_970, new_AGEMA_signal_969, n2791}), .clk ( clk ), .rnd ({Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384], Fresh[383], Fresh[382], Fresh[381], Fresh[380]}), .outt ({new_AGEMA_signal_1130, new_AGEMA_signal_1129, new_AGEMA_signal_1128, n2356}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2119 ( .a ({new_AGEMA_signal_1118, new_AGEMA_signal_1117, new_AGEMA_signal_1116, n2772}), .b ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, new_AGEMA_signal_1305, n2823}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2122 ( .ina ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, n2760}), .inb ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[399], Fresh[398], Fresh[397], Fresh[396], Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390]}), .outt ({new_AGEMA_signal_1133, new_AGEMA_signal_1132, new_AGEMA_signal_1131, n2611}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2131 ( .a ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, new_AGEMA_signal_1029, n2641}), .b ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, new_AGEMA_signal_1311, n2828}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2133 ( .ina ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .inb ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .rnd ({Fresh[409], Fresh[408], Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402], Fresh[401], Fresh[400]}), .outt ({new_AGEMA_signal_1136, new_AGEMA_signal_1135, new_AGEMA_signal_1134, n2616}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2134 ( .a ({new_AGEMA_signal_1136, new_AGEMA_signal_1135, new_AGEMA_signal_1134, n2616}), .b ({new_AGEMA_signal_1316, new_AGEMA_signal_1315, new_AGEMA_signal_1314, n2679}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2138 ( .ina ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .inb ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, n2760}), .clk ( clk ), .rnd ({Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414], Fresh[413], Fresh[412], Fresh[411], Fresh[410]}), .outt ({new_AGEMA_signal_1139, new_AGEMA_signal_1138, new_AGEMA_signal_1137, n2563}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2139 ( .a ({new_AGEMA_signal_1139, new_AGEMA_signal_1138, new_AGEMA_signal_1137, n2563}), .b ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, new_AGEMA_signal_1317, n2809}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2150 ( .a ({new_AGEMA_signal_1133, new_AGEMA_signal_1132, new_AGEMA_signal_1131, n2611}), .b ({new_AGEMA_signal_1322, new_AGEMA_signal_1321, new_AGEMA_signal_1320, n2709}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2163 ( .ina ({new_AGEMA_signal_947, new_AGEMA_signal_946, new_AGEMA_signal_945, n2796}), .inb ({new_AGEMA_signal_953, new_AGEMA_signal_952, new_AGEMA_signal_951, n2810}), .clk ( clk ), .rnd ({Fresh[429], Fresh[428], Fresh[427], Fresh[426], Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420]}), .outt ({new_AGEMA_signal_1142, new_AGEMA_signal_1141, new_AGEMA_signal_1140, n2401}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2211 ( .ina ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .inb ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[439], Fresh[438], Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432], Fresh[431], Fresh[430]}), .outt ({new_AGEMA_signal_1148, new_AGEMA_signal_1147, new_AGEMA_signal_1146, n2061}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2232 ( .ina ({new_AGEMA_signal_947, new_AGEMA_signal_946, new_AGEMA_signal_945, n2796}), .inb ({new_AGEMA_signal_971, new_AGEMA_signal_970, new_AGEMA_signal_969, n2791}), .clk ( clk ), .rnd ({Fresh[449], Fresh[448], Fresh[447], Fresh[446], Fresh[445], Fresh[444], Fresh[443], Fresh[442], Fresh[441], Fresh[440]}), .outt ({new_AGEMA_signal_1151, new_AGEMA_signal_1150, new_AGEMA_signal_1149, n2721}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2276 ( .ina ({new_AGEMA_signal_971, new_AGEMA_signal_970, new_AGEMA_signal_969, n2791}), .inb ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .clk ( clk ), .rnd ({Fresh[459], Fresh[458], Fresh[457], Fresh[456], Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450]}), .outt ({new_AGEMA_signal_1154, new_AGEMA_signal_1153, new_AGEMA_signal_1152, n2298}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2278 ( .a ({new_AGEMA_signal_1142, new_AGEMA_signal_1141, new_AGEMA_signal_1140, n2401}), .b ({new_AGEMA_signal_1358, new_AGEMA_signal_1357, new_AGEMA_signal_1356, n2118}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2307 ( .ina ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .inb ({new_AGEMA_signal_983, new_AGEMA_signal_982, new_AGEMA_signal_981, n2630}), .clk ( clk ), .rnd ({Fresh[469], Fresh[468], Fresh[467], Fresh[466], Fresh[465], Fresh[464], Fresh[463], Fresh[462], Fresh[461], Fresh[460]}), .outt ({new_AGEMA_signal_1157, new_AGEMA_signal_1156, new_AGEMA_signal_1155, n2346}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2341 ( .ina ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .inb ({new_AGEMA_signal_971, new_AGEMA_signal_970, new_AGEMA_signal_969, n2791}), .clk ( clk ), .rnd ({Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474], Fresh[473], Fresh[472], Fresh[471], Fresh[470]}), .outt ({new_AGEMA_signal_1163, new_AGEMA_signal_1162, new_AGEMA_signal_1161, n2430}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2383 ( .ina ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .inb ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .rnd ({Fresh[489], Fresh[488], Fresh[487], Fresh[486], Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .outt ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, new_AGEMA_signal_1023, n2712}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2402 ( .ina ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .inb ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}), .clk ( clk ), .rnd ({Fresh[499], Fresh[498], Fresh[497], Fresh[496], Fresh[495], Fresh[494], Fresh[493], Fresh[492], Fresh[491], Fresh[490]}), .outt ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, new_AGEMA_signal_1167, n2777}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2615 ( .ina ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .inb ({new_AGEMA_signal_959, new_AGEMA_signal_958, new_AGEMA_signal_957, n2462}), .clk ( clk ), .rnd ({Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504], Fresh[503], Fresh[502], Fresh[501], Fresh[500]}), .outt ({new_AGEMA_signal_1175, new_AGEMA_signal_1174, new_AGEMA_signal_1173, n2463}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2627 ( .ina ({new_AGEMA_signal_953, new_AGEMA_signal_952, new_AGEMA_signal_951, n2810}), .inb ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .rnd ({Fresh[519], Fresh[518], Fresh[517], Fresh[516], Fresh[515], Fresh[514], Fresh[513], Fresh[512], Fresh[511], Fresh[510]}), .outt ({new_AGEMA_signal_1178, new_AGEMA_signal_1177, new_AGEMA_signal_1176, n2474}) ) ;
    buf_clk new_AGEMA_reg_buffer_928 ( .C ( clk ), .D ( new_AGEMA_signal_12427 ), .Q ( new_AGEMA_signal_12428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_930 ( .C ( clk ), .D ( new_AGEMA_signal_12429 ), .Q ( new_AGEMA_signal_12430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_932 ( .C ( clk ), .D ( new_AGEMA_signal_12431 ), .Q ( new_AGEMA_signal_12432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_934 ( .C ( clk ), .D ( new_AGEMA_signal_12433 ), .Q ( new_AGEMA_signal_12434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_936 ( .C ( clk ), .D ( new_AGEMA_signal_12435 ), .Q ( new_AGEMA_signal_12436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_938 ( .C ( clk ), .D ( new_AGEMA_signal_12437 ), .Q ( new_AGEMA_signal_12438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_940 ( .C ( clk ), .D ( new_AGEMA_signal_12439 ), .Q ( new_AGEMA_signal_12440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_942 ( .C ( clk ), .D ( new_AGEMA_signal_12441 ), .Q ( new_AGEMA_signal_12442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_944 ( .C ( clk ), .D ( new_AGEMA_signal_12443 ), .Q ( new_AGEMA_signal_12444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_946 ( .C ( clk ), .D ( new_AGEMA_signal_12445 ), .Q ( new_AGEMA_signal_12446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_948 ( .C ( clk ), .D ( new_AGEMA_signal_12447 ), .Q ( new_AGEMA_signal_12448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_950 ( .C ( clk ), .D ( new_AGEMA_signal_12449 ), .Q ( new_AGEMA_signal_12450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_952 ( .C ( clk ), .D ( new_AGEMA_signal_12451 ), .Q ( new_AGEMA_signal_12452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_954 ( .C ( clk ), .D ( new_AGEMA_signal_12453 ), .Q ( new_AGEMA_signal_12454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_956 ( .C ( clk ), .D ( new_AGEMA_signal_12455 ), .Q ( new_AGEMA_signal_12456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_958 ( .C ( clk ), .D ( new_AGEMA_signal_12457 ), .Q ( new_AGEMA_signal_12458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_960 ( .C ( clk ), .D ( new_AGEMA_signal_12459 ), .Q ( new_AGEMA_signal_12460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_962 ( .C ( clk ), .D ( new_AGEMA_signal_12461 ), .Q ( new_AGEMA_signal_12462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_964 ( .C ( clk ), .D ( new_AGEMA_signal_12463 ), .Q ( new_AGEMA_signal_12464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_966 ( .C ( clk ), .D ( new_AGEMA_signal_12465 ), .Q ( new_AGEMA_signal_12466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_968 ( .C ( clk ), .D ( new_AGEMA_signal_12467 ), .Q ( new_AGEMA_signal_12468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_970 ( .C ( clk ), .D ( new_AGEMA_signal_12469 ), .Q ( new_AGEMA_signal_12470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_972 ( .C ( clk ), .D ( new_AGEMA_signal_12471 ), .Q ( new_AGEMA_signal_12472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_974 ( .C ( clk ), .D ( new_AGEMA_signal_12473 ), .Q ( new_AGEMA_signal_12474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_976 ( .C ( clk ), .D ( new_AGEMA_signal_12475 ), .Q ( new_AGEMA_signal_12476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_978 ( .C ( clk ), .D ( new_AGEMA_signal_12477 ), .Q ( new_AGEMA_signal_12478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_980 ( .C ( clk ), .D ( new_AGEMA_signal_12479 ), .Q ( new_AGEMA_signal_12480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_982 ( .C ( clk ), .D ( new_AGEMA_signal_12481 ), .Q ( new_AGEMA_signal_12482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_984 ( .C ( clk ), .D ( new_AGEMA_signal_12483 ), .Q ( new_AGEMA_signal_12484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_986 ( .C ( clk ), .D ( new_AGEMA_signal_12485 ), .Q ( new_AGEMA_signal_12486 ) ) ;
    buf_clk new_AGEMA_reg_buffer_988 ( .C ( clk ), .D ( new_AGEMA_signal_12487 ), .Q ( new_AGEMA_signal_12488 ) ) ;
    buf_clk new_AGEMA_reg_buffer_990 ( .C ( clk ), .D ( new_AGEMA_signal_12489 ), .Q ( new_AGEMA_signal_12490 ) ) ;
    buf_clk new_AGEMA_reg_buffer_992 ( .C ( clk ), .D ( new_AGEMA_signal_12491 ), .Q ( new_AGEMA_signal_12492 ) ) ;
    buf_clk new_AGEMA_reg_buffer_994 ( .C ( clk ), .D ( new_AGEMA_signal_12493 ), .Q ( new_AGEMA_signal_12494 ) ) ;
    buf_clk new_AGEMA_reg_buffer_996 ( .C ( clk ), .D ( new_AGEMA_signal_12495 ), .Q ( new_AGEMA_signal_12496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_998 ( .C ( clk ), .D ( new_AGEMA_signal_12497 ), .Q ( new_AGEMA_signal_12498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1000 ( .C ( clk ), .D ( new_AGEMA_signal_12499 ), .Q ( new_AGEMA_signal_12500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1002 ( .C ( clk ), .D ( new_AGEMA_signal_12501 ), .Q ( new_AGEMA_signal_12502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1004 ( .C ( clk ), .D ( new_AGEMA_signal_12503 ), .Q ( new_AGEMA_signal_12504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1006 ( .C ( clk ), .D ( new_AGEMA_signal_12505 ), .Q ( new_AGEMA_signal_12506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1008 ( .C ( clk ), .D ( new_AGEMA_signal_12507 ), .Q ( new_AGEMA_signal_12508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1010 ( .C ( clk ), .D ( new_AGEMA_signal_12509 ), .Q ( new_AGEMA_signal_12510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1012 ( .C ( clk ), .D ( new_AGEMA_signal_12511 ), .Q ( new_AGEMA_signal_12512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1014 ( .C ( clk ), .D ( new_AGEMA_signal_12513 ), .Q ( new_AGEMA_signal_12514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1016 ( .C ( clk ), .D ( new_AGEMA_signal_12515 ), .Q ( new_AGEMA_signal_12516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1018 ( .C ( clk ), .D ( new_AGEMA_signal_12517 ), .Q ( new_AGEMA_signal_12518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1020 ( .C ( clk ), .D ( new_AGEMA_signal_12519 ), .Q ( new_AGEMA_signal_12520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1022 ( .C ( clk ), .D ( new_AGEMA_signal_12521 ), .Q ( new_AGEMA_signal_12522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1024 ( .C ( clk ), .D ( new_AGEMA_signal_12523 ), .Q ( new_AGEMA_signal_12524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1026 ( .C ( clk ), .D ( new_AGEMA_signal_12525 ), .Q ( new_AGEMA_signal_12526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1028 ( .C ( clk ), .D ( new_AGEMA_signal_12527 ), .Q ( new_AGEMA_signal_12528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1030 ( .C ( clk ), .D ( new_AGEMA_signal_12529 ), .Q ( new_AGEMA_signal_12530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1032 ( .C ( clk ), .D ( new_AGEMA_signal_12531 ), .Q ( new_AGEMA_signal_12532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1034 ( .C ( clk ), .D ( new_AGEMA_signal_12533 ), .Q ( new_AGEMA_signal_12534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1036 ( .C ( clk ), .D ( new_AGEMA_signal_12535 ), .Q ( new_AGEMA_signal_12536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1038 ( .C ( clk ), .D ( new_AGEMA_signal_12537 ), .Q ( new_AGEMA_signal_12538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1040 ( .C ( clk ), .D ( new_AGEMA_signal_12539 ), .Q ( new_AGEMA_signal_12540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1042 ( .C ( clk ), .D ( new_AGEMA_signal_12541 ), .Q ( new_AGEMA_signal_12542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1044 ( .C ( clk ), .D ( new_AGEMA_signal_12543 ), .Q ( new_AGEMA_signal_12544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1046 ( .C ( clk ), .D ( new_AGEMA_signal_12545 ), .Q ( new_AGEMA_signal_12546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2072 ( .C ( clk ), .D ( new_AGEMA_signal_13571 ), .Q ( new_AGEMA_signal_13572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2078 ( .C ( clk ), .D ( new_AGEMA_signal_13577 ), .Q ( new_AGEMA_signal_13578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2084 ( .C ( clk ), .D ( new_AGEMA_signal_13583 ), .Q ( new_AGEMA_signal_13584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2090 ( .C ( clk ), .D ( new_AGEMA_signal_13589 ), .Q ( new_AGEMA_signal_13590 ) ) ;

    /* cells in depth 3 */
    buf_clk new_AGEMA_reg_buffer_1047 ( .C ( clk ), .D ( n2769 ), .Q ( new_AGEMA_signal_12547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1049 ( .C ( clk ), .D ( new_AGEMA_signal_1200 ), .Q ( new_AGEMA_signal_12549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1051 ( .C ( clk ), .D ( new_AGEMA_signal_1201 ), .Q ( new_AGEMA_signal_12551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1053 ( .C ( clk ), .D ( new_AGEMA_signal_1202 ), .Q ( new_AGEMA_signal_12553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1055 ( .C ( clk ), .D ( new_AGEMA_signal_12524 ), .Q ( new_AGEMA_signal_12555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1057 ( .C ( clk ), .D ( new_AGEMA_signal_12526 ), .Q ( new_AGEMA_signal_12557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1059 ( .C ( clk ), .D ( new_AGEMA_signal_12528 ), .Q ( new_AGEMA_signal_12559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1061 ( .C ( clk ), .D ( new_AGEMA_signal_12530 ), .Q ( new_AGEMA_signal_12561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1063 ( .C ( clk ), .D ( new_AGEMA_signal_12436 ), .Q ( new_AGEMA_signal_12563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1065 ( .C ( clk ), .D ( new_AGEMA_signal_12438 ), .Q ( new_AGEMA_signal_12565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1067 ( .C ( clk ), .D ( new_AGEMA_signal_12440 ), .Q ( new_AGEMA_signal_12567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1069 ( .C ( clk ), .D ( new_AGEMA_signal_12442 ), .Q ( new_AGEMA_signal_12569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1071 ( .C ( clk ), .D ( n2174 ), .Q ( new_AGEMA_signal_12571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1073 ( .C ( clk ), .D ( new_AGEMA_signal_1239 ), .Q ( new_AGEMA_signal_12573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1075 ( .C ( clk ), .D ( new_AGEMA_signal_1240 ), .Q ( new_AGEMA_signal_12575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1077 ( .C ( clk ), .D ( new_AGEMA_signal_1241 ), .Q ( new_AGEMA_signal_12577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1079 ( .C ( clk ), .D ( new_AGEMA_signal_12428 ), .Q ( new_AGEMA_signal_12579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1081 ( .C ( clk ), .D ( new_AGEMA_signal_12430 ), .Q ( new_AGEMA_signal_12581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1083 ( .C ( clk ), .D ( new_AGEMA_signal_12432 ), .Q ( new_AGEMA_signal_12583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1085 ( .C ( clk ), .D ( new_AGEMA_signal_12434 ), .Q ( new_AGEMA_signal_12585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1087 ( .C ( clk ), .D ( new_AGEMA_signal_12452 ), .Q ( new_AGEMA_signal_12587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1089 ( .C ( clk ), .D ( new_AGEMA_signal_12454 ), .Q ( new_AGEMA_signal_12589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1091 ( .C ( clk ), .D ( new_AGEMA_signal_12456 ), .Q ( new_AGEMA_signal_12591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1093 ( .C ( clk ), .D ( new_AGEMA_signal_12458 ), .Q ( new_AGEMA_signal_12593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1095 ( .C ( clk ), .D ( n2570 ), .Q ( new_AGEMA_signal_12595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1097 ( .C ( clk ), .D ( new_AGEMA_signal_1248 ), .Q ( new_AGEMA_signal_12597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1099 ( .C ( clk ), .D ( new_AGEMA_signal_1249 ), .Q ( new_AGEMA_signal_12599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1101 ( .C ( clk ), .D ( new_AGEMA_signal_1250 ), .Q ( new_AGEMA_signal_12601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1103 ( .C ( clk ), .D ( n2792 ), .Q ( new_AGEMA_signal_12603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1105 ( .C ( clk ), .D ( new_AGEMA_signal_1233 ), .Q ( new_AGEMA_signal_12605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1107 ( .C ( clk ), .D ( new_AGEMA_signal_1234 ), .Q ( new_AGEMA_signal_12607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1109 ( .C ( clk ), .D ( new_AGEMA_signal_1235 ), .Q ( new_AGEMA_signal_12609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1111 ( .C ( clk ), .D ( n2635 ), .Q ( new_AGEMA_signal_12611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1113 ( .C ( clk ), .D ( new_AGEMA_signal_990 ), .Q ( new_AGEMA_signal_12613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1115 ( .C ( clk ), .D ( new_AGEMA_signal_991 ), .Q ( new_AGEMA_signal_12615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1117 ( .C ( clk ), .D ( new_AGEMA_signal_992 ), .Q ( new_AGEMA_signal_12617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1119 ( .C ( clk ), .D ( n2587 ), .Q ( new_AGEMA_signal_12619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1121 ( .C ( clk ), .D ( new_AGEMA_signal_1095 ), .Q ( new_AGEMA_signal_12621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1123 ( .C ( clk ), .D ( new_AGEMA_signal_1096 ), .Q ( new_AGEMA_signal_12623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1125 ( .C ( clk ), .D ( new_AGEMA_signal_1097 ), .Q ( new_AGEMA_signal_12625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1127 ( .C ( clk ), .D ( n2725 ), .Q ( new_AGEMA_signal_12627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1129 ( .C ( clk ), .D ( new_AGEMA_signal_1062 ), .Q ( new_AGEMA_signal_12629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1131 ( .C ( clk ), .D ( new_AGEMA_signal_1063 ), .Q ( new_AGEMA_signal_12631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1133 ( .C ( clk ), .D ( new_AGEMA_signal_1064 ), .Q ( new_AGEMA_signal_12633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1135 ( .C ( clk ), .D ( n2708 ), .Q ( new_AGEMA_signal_12635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1137 ( .C ( clk ), .D ( new_AGEMA_signal_1008 ), .Q ( new_AGEMA_signal_12637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1139 ( .C ( clk ), .D ( new_AGEMA_signal_1009 ), .Q ( new_AGEMA_signal_12639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1141 ( .C ( clk ), .D ( new_AGEMA_signal_1010 ), .Q ( new_AGEMA_signal_12641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1143 ( .C ( clk ), .D ( n2818 ), .Q ( new_AGEMA_signal_12643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1145 ( .C ( clk ), .D ( new_AGEMA_signal_1290 ), .Q ( new_AGEMA_signal_12645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1147 ( .C ( clk ), .D ( new_AGEMA_signal_1291 ), .Q ( new_AGEMA_signal_12647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1149 ( .C ( clk ), .D ( new_AGEMA_signal_1292 ), .Q ( new_AGEMA_signal_12649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1151 ( .C ( clk ), .D ( n2790 ), .Q ( new_AGEMA_signal_12651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1153 ( .C ( clk ), .D ( new_AGEMA_signal_993 ), .Q ( new_AGEMA_signal_12653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1155 ( .C ( clk ), .D ( new_AGEMA_signal_994 ), .Q ( new_AGEMA_signal_12655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1157 ( .C ( clk ), .D ( new_AGEMA_signal_995 ), .Q ( new_AGEMA_signal_12657 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1159 ( .C ( clk ), .D ( n2786 ), .Q ( new_AGEMA_signal_12659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1161 ( .C ( clk ), .D ( new_AGEMA_signal_1221 ), .Q ( new_AGEMA_signal_12661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1163 ( .C ( clk ), .D ( new_AGEMA_signal_1222 ), .Q ( new_AGEMA_signal_12663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1165 ( .C ( clk ), .D ( new_AGEMA_signal_1223 ), .Q ( new_AGEMA_signal_12665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1167 ( .C ( clk ), .D ( n2400 ), .Q ( new_AGEMA_signal_12667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1169 ( .C ( clk ), .D ( new_AGEMA_signal_1080 ), .Q ( new_AGEMA_signal_12669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1171 ( .C ( clk ), .D ( new_AGEMA_signal_1081 ), .Q ( new_AGEMA_signal_12671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1173 ( .C ( clk ), .D ( new_AGEMA_signal_1082 ), .Q ( new_AGEMA_signal_12673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1175 ( .C ( clk ), .D ( new_AGEMA_signal_12460 ), .Q ( new_AGEMA_signal_12675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1177 ( .C ( clk ), .D ( new_AGEMA_signal_12462 ), .Q ( new_AGEMA_signal_12677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1179 ( .C ( clk ), .D ( new_AGEMA_signal_12464 ), .Q ( new_AGEMA_signal_12679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1181 ( .C ( clk ), .D ( new_AGEMA_signal_12466 ), .Q ( new_AGEMA_signal_12681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1183 ( .C ( clk ), .D ( n2815 ), .Q ( new_AGEMA_signal_12683 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1185 ( .C ( clk ), .D ( new_AGEMA_signal_1065 ), .Q ( new_AGEMA_signal_12685 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1187 ( .C ( clk ), .D ( new_AGEMA_signal_1066 ), .Q ( new_AGEMA_signal_12687 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1189 ( .C ( clk ), .D ( new_AGEMA_signal_1067 ), .Q ( new_AGEMA_signal_12689 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1191 ( .C ( clk ), .D ( n2723 ), .Q ( new_AGEMA_signal_12691 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1193 ( .C ( clk ), .D ( new_AGEMA_signal_1059 ), .Q ( new_AGEMA_signal_12693 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1195 ( .C ( clk ), .D ( new_AGEMA_signal_1060 ), .Q ( new_AGEMA_signal_12695 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1197 ( .C ( clk ), .D ( new_AGEMA_signal_1061 ), .Q ( new_AGEMA_signal_12697 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1199 ( .C ( clk ), .D ( n2709 ), .Q ( new_AGEMA_signal_12699 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1201 ( .C ( clk ), .D ( new_AGEMA_signal_1320 ), .Q ( new_AGEMA_signal_12701 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1203 ( .C ( clk ), .D ( new_AGEMA_signal_1321 ), .Q ( new_AGEMA_signal_12703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1205 ( .C ( clk ), .D ( new_AGEMA_signal_1322 ), .Q ( new_AGEMA_signal_12705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1207 ( .C ( clk ), .D ( n2753 ), .Q ( new_AGEMA_signal_12707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1209 ( .C ( clk ), .D ( new_AGEMA_signal_1077 ), .Q ( new_AGEMA_signal_12709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1211 ( .C ( clk ), .D ( new_AGEMA_signal_1078 ), .Q ( new_AGEMA_signal_12711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1213 ( .C ( clk ), .D ( new_AGEMA_signal_1079 ), .Q ( new_AGEMA_signal_12713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1215 ( .C ( clk ), .D ( n2401 ), .Q ( new_AGEMA_signal_12715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1217 ( .C ( clk ), .D ( new_AGEMA_signal_1140 ), .Q ( new_AGEMA_signal_12717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1219 ( .C ( clk ), .D ( new_AGEMA_signal_1141 ), .Q ( new_AGEMA_signal_12719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1221 ( .C ( clk ), .D ( new_AGEMA_signal_1142 ), .Q ( new_AGEMA_signal_12721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1223 ( .C ( clk ), .D ( new_AGEMA_signal_12508 ), .Q ( new_AGEMA_signal_12723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1225 ( .C ( clk ), .D ( new_AGEMA_signal_12510 ), .Q ( new_AGEMA_signal_12725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1227 ( .C ( clk ), .D ( new_AGEMA_signal_12512 ), .Q ( new_AGEMA_signal_12727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1229 ( .C ( clk ), .D ( new_AGEMA_signal_12514 ), .Q ( new_AGEMA_signal_12729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1231 ( .C ( clk ), .D ( new_AGEMA_signal_12468 ), .Q ( new_AGEMA_signal_12731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1233 ( .C ( clk ), .D ( new_AGEMA_signal_12470 ), .Q ( new_AGEMA_signal_12733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1235 ( .C ( clk ), .D ( new_AGEMA_signal_12472 ), .Q ( new_AGEMA_signal_12735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1237 ( .C ( clk ), .D ( new_AGEMA_signal_12474 ), .Q ( new_AGEMA_signal_12737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1239 ( .C ( clk ), .D ( n2615 ), .Q ( new_AGEMA_signal_12739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1241 ( .C ( clk ), .D ( new_AGEMA_signal_1035 ), .Q ( new_AGEMA_signal_12741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1243 ( .C ( clk ), .D ( new_AGEMA_signal_1036 ), .Q ( new_AGEMA_signal_12743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1245 ( .C ( clk ), .D ( new_AGEMA_signal_1037 ), .Q ( new_AGEMA_signal_12745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1247 ( .C ( clk ), .D ( n2643 ), .Q ( new_AGEMA_signal_12747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1249 ( .C ( clk ), .D ( new_AGEMA_signal_1098 ), .Q ( new_AGEMA_signal_12749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1251 ( .C ( clk ), .D ( new_AGEMA_signal_1099 ), .Q ( new_AGEMA_signal_12751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1253 ( .C ( clk ), .D ( new_AGEMA_signal_1100 ), .Q ( new_AGEMA_signal_12753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1255 ( .C ( clk ), .D ( n2563 ), .Q ( new_AGEMA_signal_12755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1257 ( .C ( clk ), .D ( new_AGEMA_signal_1137 ), .Q ( new_AGEMA_signal_12757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1259 ( .C ( clk ), .D ( new_AGEMA_signal_1138 ), .Q ( new_AGEMA_signal_12759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1261 ( .C ( clk ), .D ( new_AGEMA_signal_1139 ), .Q ( new_AGEMA_signal_12761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1263 ( .C ( clk ), .D ( n2612 ), .Q ( new_AGEMA_signal_12763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1265 ( .C ( clk ), .D ( new_AGEMA_signal_1275 ), .Q ( new_AGEMA_signal_12765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1267 ( .C ( clk ), .D ( new_AGEMA_signal_1276 ), .Q ( new_AGEMA_signal_12767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1269 ( .C ( clk ), .D ( new_AGEMA_signal_1277 ), .Q ( new_AGEMA_signal_12769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1271 ( .C ( clk ), .D ( n2824 ), .Q ( new_AGEMA_signal_12771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1273 ( .C ( clk ), .D ( new_AGEMA_signal_1119 ), .Q ( new_AGEMA_signal_12773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1275 ( .C ( clk ), .D ( new_AGEMA_signal_1120 ), .Q ( new_AGEMA_signal_12775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1277 ( .C ( clk ), .D ( new_AGEMA_signal_1121 ), .Q ( new_AGEMA_signal_12777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1279 ( .C ( clk ), .D ( n2816 ), .Q ( new_AGEMA_signal_12779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1281 ( .C ( clk ), .D ( new_AGEMA_signal_1041 ), .Q ( new_AGEMA_signal_12781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1283 ( .C ( clk ), .D ( new_AGEMA_signal_1042 ), .Q ( new_AGEMA_signal_12783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1285 ( .C ( clk ), .D ( new_AGEMA_signal_1043 ), .Q ( new_AGEMA_signal_12785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1287 ( .C ( clk ), .D ( n2073 ), .Q ( new_AGEMA_signal_12787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1289 ( .C ( clk ), .D ( new_AGEMA_signal_1053 ), .Q ( new_AGEMA_signal_12789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1291 ( .C ( clk ), .D ( new_AGEMA_signal_1054 ), .Q ( new_AGEMA_signal_12791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1293 ( .C ( clk ), .D ( new_AGEMA_signal_1055 ), .Q ( new_AGEMA_signal_12793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1295 ( .C ( clk ), .D ( n2519 ), .Q ( new_AGEMA_signal_12795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1297 ( .C ( clk ), .D ( new_AGEMA_signal_996 ), .Q ( new_AGEMA_signal_12797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1299 ( .C ( clk ), .D ( new_AGEMA_signal_997 ), .Q ( new_AGEMA_signal_12799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1301 ( .C ( clk ), .D ( new_AGEMA_signal_998 ), .Q ( new_AGEMA_signal_12801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1303 ( .C ( clk ), .D ( n2616 ), .Q ( new_AGEMA_signal_12803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1305 ( .C ( clk ), .D ( new_AGEMA_signal_1134 ), .Q ( new_AGEMA_signal_12805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1307 ( .C ( clk ), .D ( new_AGEMA_signal_1135 ), .Q ( new_AGEMA_signal_12807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1309 ( .C ( clk ), .D ( new_AGEMA_signal_1136 ), .Q ( new_AGEMA_signal_12809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1311 ( .C ( clk ), .D ( new_AGEMA_signal_12516 ), .Q ( new_AGEMA_signal_12811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1313 ( .C ( clk ), .D ( new_AGEMA_signal_12518 ), .Q ( new_AGEMA_signal_12813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1315 ( .C ( clk ), .D ( new_AGEMA_signal_12520 ), .Q ( new_AGEMA_signal_12815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1317 ( .C ( clk ), .D ( new_AGEMA_signal_12522 ), .Q ( new_AGEMA_signal_12817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1319 ( .C ( clk ), .D ( n2780 ), .Q ( new_AGEMA_signal_12819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1321 ( .C ( clk ), .D ( new_AGEMA_signal_1044 ), .Q ( new_AGEMA_signal_12821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1323 ( .C ( clk ), .D ( new_AGEMA_signal_1045 ), .Q ( new_AGEMA_signal_12823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1325 ( .C ( clk ), .D ( new_AGEMA_signal_1046 ), .Q ( new_AGEMA_signal_12825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1327 ( .C ( clk ), .D ( new_AGEMA_signal_12532 ), .Q ( new_AGEMA_signal_12827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1329 ( .C ( clk ), .D ( new_AGEMA_signal_12534 ), .Q ( new_AGEMA_signal_12829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1331 ( .C ( clk ), .D ( new_AGEMA_signal_12536 ), .Q ( new_AGEMA_signal_12831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1333 ( .C ( clk ), .D ( new_AGEMA_signal_12538 ), .Q ( new_AGEMA_signal_12833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1335 ( .C ( clk ), .D ( n2742 ), .Q ( new_AGEMA_signal_12835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1337 ( .C ( clk ), .D ( new_AGEMA_signal_1074 ), .Q ( new_AGEMA_signal_12837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1339 ( .C ( clk ), .D ( new_AGEMA_signal_1075 ), .Q ( new_AGEMA_signal_12839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1341 ( .C ( clk ), .D ( new_AGEMA_signal_1076 ), .Q ( new_AGEMA_signal_12841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1343 ( .C ( clk ), .D ( n2724 ), .Q ( new_AGEMA_signal_12843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1345 ( .C ( clk ), .D ( new_AGEMA_signal_1236 ), .Q ( new_AGEMA_signal_12845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1347 ( .C ( clk ), .D ( new_AGEMA_signal_1237 ), .Q ( new_AGEMA_signal_12847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1349 ( .C ( clk ), .D ( new_AGEMA_signal_1238 ), .Q ( new_AGEMA_signal_12849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1351 ( .C ( clk ), .D ( n2317 ), .Q ( new_AGEMA_signal_12851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1353 ( .C ( clk ), .D ( new_AGEMA_signal_1047 ), .Q ( new_AGEMA_signal_12853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1355 ( .C ( clk ), .D ( new_AGEMA_signal_1048 ), .Q ( new_AGEMA_signal_12855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1357 ( .C ( clk ), .D ( new_AGEMA_signal_1049 ), .Q ( new_AGEMA_signal_12857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1359 ( .C ( clk ), .D ( n2688 ), .Q ( new_AGEMA_signal_12859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1361 ( .C ( clk ), .D ( new_AGEMA_signal_1209 ), .Q ( new_AGEMA_signal_12861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1363 ( .C ( clk ), .D ( new_AGEMA_signal_1210 ), .Q ( new_AGEMA_signal_12863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1365 ( .C ( clk ), .D ( new_AGEMA_signal_1211 ), .Q ( new_AGEMA_signal_12865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1367 ( .C ( clk ), .D ( n2609 ), .Q ( new_AGEMA_signal_12867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1369 ( .C ( clk ), .D ( new_AGEMA_signal_1086 ), .Q ( new_AGEMA_signal_12869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1371 ( .C ( clk ), .D ( new_AGEMA_signal_1087 ), .Q ( new_AGEMA_signal_12871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1373 ( .C ( clk ), .D ( new_AGEMA_signal_1088 ), .Q ( new_AGEMA_signal_12873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1375 ( .C ( clk ), .D ( n2672 ), .Q ( new_AGEMA_signal_12875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1377 ( .C ( clk ), .D ( new_AGEMA_signal_1185 ), .Q ( new_AGEMA_signal_12877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1379 ( .C ( clk ), .D ( new_AGEMA_signal_1186 ), .Q ( new_AGEMA_signal_12879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1381 ( .C ( clk ), .D ( new_AGEMA_signal_1187 ), .Q ( new_AGEMA_signal_12881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1383 ( .C ( clk ), .D ( n2640 ), .Q ( new_AGEMA_signal_12883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1385 ( .C ( clk ), .D ( new_AGEMA_signal_1188 ), .Q ( new_AGEMA_signal_12885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1387 ( .C ( clk ), .D ( new_AGEMA_signal_1189 ), .Q ( new_AGEMA_signal_12887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1389 ( .C ( clk ), .D ( new_AGEMA_signal_1190 ), .Q ( new_AGEMA_signal_12889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1391 ( .C ( clk ), .D ( n2713 ), .Q ( new_AGEMA_signal_12891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1393 ( .C ( clk ), .D ( new_AGEMA_signal_1056 ), .Q ( new_AGEMA_signal_12893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1395 ( .C ( clk ), .D ( new_AGEMA_signal_1057 ), .Q ( new_AGEMA_signal_12895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1397 ( .C ( clk ), .D ( new_AGEMA_signal_1058 ), .Q ( new_AGEMA_signal_12897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1399 ( .C ( clk ), .D ( n2777 ), .Q ( new_AGEMA_signal_12899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1401 ( .C ( clk ), .D ( new_AGEMA_signal_1167 ), .Q ( new_AGEMA_signal_12901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1403 ( .C ( clk ), .D ( new_AGEMA_signal_1168 ), .Q ( new_AGEMA_signal_12903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1405 ( .C ( clk ), .D ( new_AGEMA_signal_1169 ), .Q ( new_AGEMA_signal_12905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1407 ( .C ( clk ), .D ( n2789 ), .Q ( new_AGEMA_signal_12907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1409 ( .C ( clk ), .D ( new_AGEMA_signal_1197 ), .Q ( new_AGEMA_signal_12909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1411 ( .C ( clk ), .D ( new_AGEMA_signal_1198 ), .Q ( new_AGEMA_signal_12911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1413 ( .C ( clk ), .D ( new_AGEMA_signal_1199 ), .Q ( new_AGEMA_signal_12913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1415 ( .C ( clk ), .D ( n2661 ), .Q ( new_AGEMA_signal_12915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1417 ( .C ( clk ), .D ( new_AGEMA_signal_1089 ), .Q ( new_AGEMA_signal_12917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1419 ( .C ( clk ), .D ( new_AGEMA_signal_1090 ), .Q ( new_AGEMA_signal_12919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1421 ( .C ( clk ), .D ( new_AGEMA_signal_1091 ), .Q ( new_AGEMA_signal_12921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1423 ( .C ( clk ), .D ( new_AGEMA_signal_12484 ), .Q ( new_AGEMA_signal_12923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1425 ( .C ( clk ), .D ( new_AGEMA_signal_12486 ), .Q ( new_AGEMA_signal_12925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1427 ( .C ( clk ), .D ( new_AGEMA_signal_12488 ), .Q ( new_AGEMA_signal_12927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1429 ( .C ( clk ), .D ( new_AGEMA_signal_12490 ), .Q ( new_AGEMA_signal_12929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1431 ( .C ( clk ), .D ( n2694 ), .Q ( new_AGEMA_signal_12931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1433 ( .C ( clk ), .D ( new_AGEMA_signal_1050 ), .Q ( new_AGEMA_signal_12933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1435 ( .C ( clk ), .D ( new_AGEMA_signal_1051 ), .Q ( new_AGEMA_signal_12935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1437 ( .C ( clk ), .D ( new_AGEMA_signal_1052 ), .Q ( new_AGEMA_signal_12937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1439 ( .C ( clk ), .D ( new_AGEMA_signal_12492 ), .Q ( new_AGEMA_signal_12939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1441 ( .C ( clk ), .D ( new_AGEMA_signal_12494 ), .Q ( new_AGEMA_signal_12941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1443 ( .C ( clk ), .D ( new_AGEMA_signal_12496 ), .Q ( new_AGEMA_signal_12943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1445 ( .C ( clk ), .D ( new_AGEMA_signal_12498 ), .Q ( new_AGEMA_signal_12945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1447 ( .C ( clk ), .D ( n2682 ), .Q ( new_AGEMA_signal_12947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1449 ( .C ( clk ), .D ( new_AGEMA_signal_1002 ), .Q ( new_AGEMA_signal_12949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1451 ( .C ( clk ), .D ( new_AGEMA_signal_1003 ), .Q ( new_AGEMA_signal_12951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1453 ( .C ( clk ), .D ( new_AGEMA_signal_1004 ), .Q ( new_AGEMA_signal_12953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1455 ( .C ( clk ), .D ( new_AGEMA_signal_12540 ), .Q ( new_AGEMA_signal_12955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1457 ( .C ( clk ), .D ( new_AGEMA_signal_12542 ), .Q ( new_AGEMA_signal_12957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1459 ( .C ( clk ), .D ( new_AGEMA_signal_12544 ), .Q ( new_AGEMA_signal_12959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1461 ( .C ( clk ), .D ( new_AGEMA_signal_12546 ), .Q ( new_AGEMA_signal_12961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1463 ( .C ( clk ), .D ( n2624 ), .Q ( new_AGEMA_signal_12963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1465 ( .C ( clk ), .D ( new_AGEMA_signal_1125 ), .Q ( new_AGEMA_signal_12965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1467 ( .C ( clk ), .D ( new_AGEMA_signal_1126 ), .Q ( new_AGEMA_signal_12967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1469 ( .C ( clk ), .D ( new_AGEMA_signal_1127 ), .Q ( new_AGEMA_signal_12969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1471 ( .C ( clk ), .D ( n2356 ), .Q ( new_AGEMA_signal_12971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1473 ( .C ( clk ), .D ( new_AGEMA_signal_1128 ), .Q ( new_AGEMA_signal_12973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1475 ( .C ( clk ), .D ( new_AGEMA_signal_1129 ), .Q ( new_AGEMA_signal_12975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1477 ( .C ( clk ), .D ( new_AGEMA_signal_1130 ), .Q ( new_AGEMA_signal_12977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1479 ( .C ( clk ), .D ( n2778 ), .Q ( new_AGEMA_signal_12979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1481 ( .C ( clk ), .D ( new_AGEMA_signal_1107 ), .Q ( new_AGEMA_signal_12981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1483 ( .C ( clk ), .D ( new_AGEMA_signal_1108 ), .Q ( new_AGEMA_signal_12983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1485 ( .C ( clk ), .D ( new_AGEMA_signal_1109 ), .Q ( new_AGEMA_signal_12985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1487 ( .C ( clk ), .D ( n2766 ), .Q ( new_AGEMA_signal_12987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1489 ( .C ( clk ), .D ( new_AGEMA_signal_1266 ), .Q ( new_AGEMA_signal_12989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1491 ( .C ( clk ), .D ( new_AGEMA_signal_1267 ), .Q ( new_AGEMA_signal_12991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1493 ( .C ( clk ), .D ( new_AGEMA_signal_1268 ), .Q ( new_AGEMA_signal_12993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1495 ( .C ( clk ), .D ( n2767 ), .Q ( new_AGEMA_signal_12995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1497 ( .C ( clk ), .D ( new_AGEMA_signal_1194 ), .Q ( new_AGEMA_signal_12997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1499 ( .C ( clk ), .D ( new_AGEMA_signal_1195 ), .Q ( new_AGEMA_signal_12999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1501 ( .C ( clk ), .D ( new_AGEMA_signal_1196 ), .Q ( new_AGEMA_signal_13001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1503 ( .C ( clk ), .D ( n2641 ), .Q ( new_AGEMA_signal_13003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1505 ( .C ( clk ), .D ( new_AGEMA_signal_1029 ), .Q ( new_AGEMA_signal_13005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1507 ( .C ( clk ), .D ( new_AGEMA_signal_1030 ), .Q ( new_AGEMA_signal_13007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1509 ( .C ( clk ), .D ( new_AGEMA_signal_1031 ), .Q ( new_AGEMA_signal_13009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1511 ( .C ( clk ), .D ( n2719 ), .Q ( new_AGEMA_signal_13011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1513 ( .C ( clk ), .D ( new_AGEMA_signal_1026 ), .Q ( new_AGEMA_signal_13013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1515 ( .C ( clk ), .D ( new_AGEMA_signal_1027 ), .Q ( new_AGEMA_signal_13015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1517 ( .C ( clk ), .D ( new_AGEMA_signal_1028 ), .Q ( new_AGEMA_signal_13017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1519 ( .C ( clk ), .D ( n2707 ), .Q ( new_AGEMA_signal_13019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1521 ( .C ( clk ), .D ( new_AGEMA_signal_1203 ), .Q ( new_AGEMA_signal_13021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1523 ( .C ( clk ), .D ( new_AGEMA_signal_1204 ), .Q ( new_AGEMA_signal_13023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1525 ( .C ( clk ), .D ( new_AGEMA_signal_1205 ), .Q ( new_AGEMA_signal_13025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1527 ( .C ( clk ), .D ( n2493 ), .Q ( new_AGEMA_signal_13027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1529 ( .C ( clk ), .D ( new_AGEMA_signal_1092 ), .Q ( new_AGEMA_signal_13029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1531 ( .C ( clk ), .D ( new_AGEMA_signal_1093 ), .Q ( new_AGEMA_signal_13031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1533 ( .C ( clk ), .D ( new_AGEMA_signal_1094 ), .Q ( new_AGEMA_signal_13033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1535 ( .C ( clk ), .D ( n2577 ), .Q ( new_AGEMA_signal_13035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1537 ( .C ( clk ), .D ( new_AGEMA_signal_1227 ), .Q ( new_AGEMA_signal_13037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1539 ( .C ( clk ), .D ( new_AGEMA_signal_1228 ), .Q ( new_AGEMA_signal_13039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1541 ( .C ( clk ), .D ( new_AGEMA_signal_1229 ), .Q ( new_AGEMA_signal_13041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1543 ( .C ( clk ), .D ( n2541 ), .Q ( new_AGEMA_signal_13043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1545 ( .C ( clk ), .D ( new_AGEMA_signal_1212 ), .Q ( new_AGEMA_signal_13045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1547 ( .C ( clk ), .D ( new_AGEMA_signal_1213 ), .Q ( new_AGEMA_signal_13047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1549 ( .C ( clk ), .D ( new_AGEMA_signal_1214 ), .Q ( new_AGEMA_signal_13049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1551 ( .C ( clk ), .D ( n2679 ), .Q ( new_AGEMA_signal_13051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1553 ( .C ( clk ), .D ( new_AGEMA_signal_1314 ), .Q ( new_AGEMA_signal_13053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1555 ( .C ( clk ), .D ( new_AGEMA_signal_1315 ), .Q ( new_AGEMA_signal_13055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1557 ( .C ( clk ), .D ( new_AGEMA_signal_1316 ), .Q ( new_AGEMA_signal_13057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1559 ( .C ( clk ), .D ( n2699 ), .Q ( new_AGEMA_signal_13059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1561 ( .C ( clk ), .D ( new_AGEMA_signal_1038 ), .Q ( new_AGEMA_signal_13061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1563 ( .C ( clk ), .D ( new_AGEMA_signal_1039 ), .Q ( new_AGEMA_signal_13063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1565 ( .C ( clk ), .D ( new_AGEMA_signal_1040 ), .Q ( new_AGEMA_signal_13065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1567 ( .C ( clk ), .D ( n2611 ), .Q ( new_AGEMA_signal_13067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1569 ( .C ( clk ), .D ( new_AGEMA_signal_1131 ), .Q ( new_AGEMA_signal_13069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1571 ( .C ( clk ), .D ( new_AGEMA_signal_1132 ), .Q ( new_AGEMA_signal_13071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1573 ( .C ( clk ), .D ( new_AGEMA_signal_1133 ), .Q ( new_AGEMA_signal_13073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1575 ( .C ( clk ), .D ( n2739 ), .Q ( new_AGEMA_signal_13075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1577 ( .C ( clk ), .D ( new_AGEMA_signal_1101 ), .Q ( new_AGEMA_signal_13077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1579 ( .C ( clk ), .D ( new_AGEMA_signal_1102 ), .Q ( new_AGEMA_signal_13079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1581 ( .C ( clk ), .D ( new_AGEMA_signal_1103 ), .Q ( new_AGEMA_signal_13081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1583 ( .C ( clk ), .D ( n2772 ), .Q ( new_AGEMA_signal_13083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1585 ( .C ( clk ), .D ( new_AGEMA_signal_1116 ), .Q ( new_AGEMA_signal_13085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1587 ( .C ( clk ), .D ( new_AGEMA_signal_1117 ), .Q ( new_AGEMA_signal_13087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1589 ( .C ( clk ), .D ( new_AGEMA_signal_1118 ), .Q ( new_AGEMA_signal_13089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1607 ( .C ( clk ), .D ( n2442 ), .Q ( new_AGEMA_signal_13107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1611 ( .C ( clk ), .D ( new_AGEMA_signal_1251 ), .Q ( new_AGEMA_signal_13111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1615 ( .C ( clk ), .D ( new_AGEMA_signal_1252 ), .Q ( new_AGEMA_signal_13115 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1619 ( .C ( clk ), .D ( new_AGEMA_signal_1253 ), .Q ( new_AGEMA_signal_13119 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1711 ( .C ( clk ), .D ( n2779 ), .Q ( new_AGEMA_signal_13211 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1715 ( .C ( clk ), .D ( new_AGEMA_signal_1017 ), .Q ( new_AGEMA_signal_13215 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1719 ( .C ( clk ), .D ( new_AGEMA_signal_1018 ), .Q ( new_AGEMA_signal_13219 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1723 ( .C ( clk ), .D ( new_AGEMA_signal_1019 ), .Q ( new_AGEMA_signal_13223 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1783 ( .C ( clk ), .D ( n2721 ), .Q ( new_AGEMA_signal_13283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1787 ( .C ( clk ), .D ( new_AGEMA_signal_1149 ), .Q ( new_AGEMA_signal_13287 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1791 ( .C ( clk ), .D ( new_AGEMA_signal_1150 ), .Q ( new_AGEMA_signal_13291 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1795 ( .C ( clk ), .D ( new_AGEMA_signal_1151 ), .Q ( new_AGEMA_signal_13295 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1839 ( .C ( clk ), .D ( n2823 ), .Q ( new_AGEMA_signal_13339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1843 ( .C ( clk ), .D ( new_AGEMA_signal_1305 ), .Q ( new_AGEMA_signal_13343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1847 ( .C ( clk ), .D ( new_AGEMA_signal_1306 ), .Q ( new_AGEMA_signal_13347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1851 ( .C ( clk ), .D ( new_AGEMA_signal_1307 ), .Q ( new_AGEMA_signal_13351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1879 ( .C ( clk ), .D ( n2346 ), .Q ( new_AGEMA_signal_13379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1883 ( .C ( clk ), .D ( new_AGEMA_signal_1155 ), .Q ( new_AGEMA_signal_13383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1887 ( .C ( clk ), .D ( new_AGEMA_signal_1156 ), .Q ( new_AGEMA_signal_13387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1891 ( .C ( clk ), .D ( new_AGEMA_signal_1157 ), .Q ( new_AGEMA_signal_13391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1919 ( .C ( clk ), .D ( n2315 ), .Q ( new_AGEMA_signal_13419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1923 ( .C ( clk ), .D ( new_AGEMA_signal_999 ), .Q ( new_AGEMA_signal_13423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1927 ( .C ( clk ), .D ( new_AGEMA_signal_1000 ), .Q ( new_AGEMA_signal_13427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1931 ( .C ( clk ), .D ( new_AGEMA_signal_1001 ), .Q ( new_AGEMA_signal_13431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2073 ( .C ( clk ), .D ( new_AGEMA_signal_13572 ), .Q ( new_AGEMA_signal_13573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2079 ( .C ( clk ), .D ( new_AGEMA_signal_13578 ), .Q ( new_AGEMA_signal_13579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2085 ( .C ( clk ), .D ( new_AGEMA_signal_13584 ), .Q ( new_AGEMA_signal_13585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2091 ( .C ( clk ), .D ( new_AGEMA_signal_13590 ), .Q ( new_AGEMA_signal_13591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2119 ( .C ( clk ), .D ( new_AGEMA_signal_12444 ), .Q ( new_AGEMA_signal_13619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2123 ( .C ( clk ), .D ( new_AGEMA_signal_12446 ), .Q ( new_AGEMA_signal_13623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2127 ( .C ( clk ), .D ( new_AGEMA_signal_12448 ), .Q ( new_AGEMA_signal_13627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2131 ( .C ( clk ), .D ( new_AGEMA_signal_12450 ), .Q ( new_AGEMA_signal_13631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2159 ( .C ( clk ), .D ( n2600 ), .Q ( new_AGEMA_signal_13659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2163 ( .C ( clk ), .D ( new_AGEMA_signal_1068 ), .Q ( new_AGEMA_signal_13663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2167 ( .C ( clk ), .D ( new_AGEMA_signal_1069 ), .Q ( new_AGEMA_signal_13667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2171 ( .C ( clk ), .D ( new_AGEMA_signal_1070 ), .Q ( new_AGEMA_signal_13671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2231 ( .C ( clk ), .D ( n2750 ), .Q ( new_AGEMA_signal_13731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2235 ( .C ( clk ), .D ( new_AGEMA_signal_1032 ), .Q ( new_AGEMA_signal_13735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2239 ( .C ( clk ), .D ( new_AGEMA_signal_1033 ), .Q ( new_AGEMA_signal_13739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2243 ( .C ( clk ), .D ( new_AGEMA_signal_1034 ), .Q ( new_AGEMA_signal_13743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2263 ( .C ( clk ), .D ( new_AGEMA_signal_12500 ), .Q ( new_AGEMA_signal_13763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2267 ( .C ( clk ), .D ( new_AGEMA_signal_12502 ), .Q ( new_AGEMA_signal_13767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2271 ( .C ( clk ), .D ( new_AGEMA_signal_12504 ), .Q ( new_AGEMA_signal_13771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2275 ( .C ( clk ), .D ( new_AGEMA_signal_12506 ), .Q ( new_AGEMA_signal_13775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2559 ( .C ( clk ), .D ( n2737 ), .Q ( new_AGEMA_signal_14059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2565 ( .C ( clk ), .D ( new_AGEMA_signal_1191 ), .Q ( new_AGEMA_signal_14065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2571 ( .C ( clk ), .D ( new_AGEMA_signal_1192 ), .Q ( new_AGEMA_signal_14071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2577 ( .C ( clk ), .D ( new_AGEMA_signal_1193 ), .Q ( new_AGEMA_signal_14077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2663 ( .C ( clk ), .D ( n2785 ), .Q ( new_AGEMA_signal_14163 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2669 ( .C ( clk ), .D ( new_AGEMA_signal_1083 ), .Q ( new_AGEMA_signal_14169 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2675 ( .C ( clk ), .D ( new_AGEMA_signal_1084 ), .Q ( new_AGEMA_signal_14175 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2681 ( .C ( clk ), .D ( new_AGEMA_signal_1085 ), .Q ( new_AGEMA_signal_14181 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3127 ( .C ( clk ), .D ( n2595 ), .Q ( new_AGEMA_signal_14627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3135 ( .C ( clk ), .D ( new_AGEMA_signal_1005 ), .Q ( new_AGEMA_signal_14635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3143 ( .C ( clk ), .D ( new_AGEMA_signal_1006 ), .Q ( new_AGEMA_signal_14643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3151 ( .C ( clk ), .D ( new_AGEMA_signal_1007 ), .Q ( new_AGEMA_signal_14651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3167 ( .C ( clk ), .D ( n2437 ), .Q ( new_AGEMA_signal_14667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3175 ( .C ( clk ), .D ( new_AGEMA_signal_1104 ), .Q ( new_AGEMA_signal_14675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3183 ( .C ( clk ), .D ( new_AGEMA_signal_1105 ), .Q ( new_AGEMA_signal_14683 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3191 ( .C ( clk ), .D ( new_AGEMA_signal_1106 ), .Q ( new_AGEMA_signal_14691 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3471 ( .C ( clk ), .D ( n2828 ), .Q ( new_AGEMA_signal_14971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3479 ( .C ( clk ), .D ( new_AGEMA_signal_1311 ), .Q ( new_AGEMA_signal_14979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3487 ( .C ( clk ), .D ( new_AGEMA_signal_1312 ), .Q ( new_AGEMA_signal_14987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3495 ( .C ( clk ), .D ( new_AGEMA_signal_1313 ), .Q ( new_AGEMA_signal_14995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3815 ( .C ( clk ), .D ( n2538 ), .Q ( new_AGEMA_signal_15315 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3823 ( .C ( clk ), .D ( new_AGEMA_signal_1071 ), .Q ( new_AGEMA_signal_15323 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3831 ( .C ( clk ), .D ( new_AGEMA_signal_1072 ), .Q ( new_AGEMA_signal_15331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3839 ( .C ( clk ), .D ( new_AGEMA_signal_1073 ), .Q ( new_AGEMA_signal_15339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3935 ( .C ( clk ), .D ( n2809 ), .Q ( new_AGEMA_signal_15435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3943 ( .C ( clk ), .D ( new_AGEMA_signal_1317 ), .Q ( new_AGEMA_signal_15443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3951 ( .C ( clk ), .D ( new_AGEMA_signal_1318 ), .Q ( new_AGEMA_signal_15451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3959 ( .C ( clk ), .D ( new_AGEMA_signal_1319 ), .Q ( new_AGEMA_signal_15459 ) ) ;

    /* cells in depth 4 */
    nand_HPC1 #(.security_order(3), .pipeline(1)) U1954 ( .ina ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, new_AGEMA_signal_1032, n2750}), .inb ({new_AGEMA_signal_1190, new_AGEMA_signal_1189, new_AGEMA_signal_1188, n2640}), .clk ( clk ), .rnd ({Fresh[529], Fresh[528], Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522], Fresh[521], Fresh[520]}), .outt ({new_AGEMA_signal_1499, new_AGEMA_signal_1498, new_AGEMA_signal_1497, n2575}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U1959 ( .ina ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, new_AGEMA_signal_1191, n2737}), .inb ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2767}), .clk ( clk ), .rnd ({Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534], Fresh[533], Fresh[532], Fresh[531], Fresh[530]}), .outt ({new_AGEMA_signal_1502, new_AGEMA_signal_1501, new_AGEMA_signal_1500, n1962}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U1964 ( .ina ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, new_AGEMA_signal_1197, n2789}), .inb ({new_AGEMA_signal_1049, new_AGEMA_signal_1048, new_AGEMA_signal_1047, n2317}), .clk ( clk ), .rnd ({Fresh[549], Fresh[548], Fresh[547], Fresh[546], Fresh[545], Fresh[544], Fresh[543], Fresh[542], Fresh[541], Fresh[540]}), .outt ({new_AGEMA_signal_1505, new_AGEMA_signal_1504, new_AGEMA_signal_1503, n1922}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U1974 ( .ina ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, new_AGEMA_signal_999, n2315}), .inb ({new_AGEMA_signal_1058, new_AGEMA_signal_1057, new_AGEMA_signal_1056, n2713}), .clk ( clk ), .rnd ({Fresh[559], Fresh[558], Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552], Fresh[551], Fresh[550]}), .outt ({new_AGEMA_signal_1208, new_AGEMA_signal_1207, new_AGEMA_signal_1206, n2755}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U1977 ( .ina ({new_AGEMA_signal_1049, new_AGEMA_signal_1048, new_AGEMA_signal_1047, n2317}), .inb ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, new_AGEMA_signal_1209, n2688}), .clk ( clk ), .rnd ({Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564], Fresh[563], Fresh[562], Fresh[561], Fresh[560]}), .outt ({new_AGEMA_signal_1508, new_AGEMA_signal_1507, new_AGEMA_signal_1506, n1926}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U1980 ( .ina ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2767}), .inb ({new_AGEMA_signal_1214, new_AGEMA_signal_1213, new_AGEMA_signal_1212, n2541}), .clk ( clk ), .rnd ({Fresh[579], Fresh[578], Fresh[577], Fresh[576], Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570]}), .outt ({new_AGEMA_signal_1511, new_AGEMA_signal_1510, new_AGEMA_signal_1509, n1925}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U1986 ( .ina ({new_AGEMA_signal_1217, new_AGEMA_signal_1216, new_AGEMA_signal_1215, n2086}), .inb ({new_AGEMA_signal_1049, new_AGEMA_signal_1048, new_AGEMA_signal_1047, n2317}), .clk ( clk ), .rnd ({Fresh[589], Fresh[588], Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582], Fresh[581], Fresh[580]}), .outt ({new_AGEMA_signal_1514, new_AGEMA_signal_1513, new_AGEMA_signal_1512, n2151}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U1988 ( .ina ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, new_AGEMA_signal_1029, n2641}), .inb ({new_AGEMA_signal_1070, new_AGEMA_signal_1069, new_AGEMA_signal_1068, n2600}), .clk ( clk ), .rnd ({Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594], Fresh[593], Fresh[592], Fresh[591], Fresh[590]}), .outt ({new_AGEMA_signal_1220, new_AGEMA_signal_1219, new_AGEMA_signal_1218, n2631}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1989 ( .a ({new_AGEMA_signal_1220, new_AGEMA_signal_1219, new_AGEMA_signal_1218, n2631}), .b ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, new_AGEMA_signal_1515, n2734}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U1992 ( .ina ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .inb ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, n2786}), .clk ( clk ), .rnd ({Fresh[609], Fresh[608], Fresh[607], Fresh[606], Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600]}), .outt ({new_AGEMA_signal_1520, new_AGEMA_signal_1519, new_AGEMA_signal_1518, n2763}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U1997 ( .ina ({new_AGEMA_signal_998, new_AGEMA_signal_997, new_AGEMA_signal_996, n2519}), .inb ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2742}), .clk ( clk ), .rnd ({Fresh[619], Fresh[618], Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612], Fresh[611], Fresh[610]}), .outt ({new_AGEMA_signal_1226, new_AGEMA_signal_1225, new_AGEMA_signal_1224, n1930}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2005 ( .ina ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, new_AGEMA_signal_1080, n2400}), .inb ({new_AGEMA_signal_998, new_AGEMA_signal_997, new_AGEMA_signal_996, n2519}), .clk ( clk ), .rnd ({Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624], Fresh[623], Fresh[622], Fresh[621], Fresh[620]}), .outt ({new_AGEMA_signal_1232, new_AGEMA_signal_1231, new_AGEMA_signal_1230, n2492}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2006 ( .a ({new_AGEMA_signal_1232, new_AGEMA_signal_1231, new_AGEMA_signal_1230, n2492}), .b ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, new_AGEMA_signal_1521, n2732}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2010 ( .ina ({new_AGEMA_signal_12434, new_AGEMA_signal_12432, new_AGEMA_signal_12430, new_AGEMA_signal_12428}), .inb ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, n2792}), .clk ( clk ), .rnd ({Fresh[639], Fresh[638], Fresh[637], Fresh[636], Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630]}), .outt ({new_AGEMA_signal_1526, new_AGEMA_signal_1525, new_AGEMA_signal_1524, n1937}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2022 ( .ina ({new_AGEMA_signal_12442, new_AGEMA_signal_12440, new_AGEMA_signal_12438, new_AGEMA_signal_12436}), .inb ({new_AGEMA_signal_1094, new_AGEMA_signal_1093, new_AGEMA_signal_1092, n2493}), .clk ( clk ), .rnd ({Fresh[649], Fresh[648], Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642], Fresh[641], Fresh[640]}), .outt ({new_AGEMA_signal_1244, new_AGEMA_signal_1243, new_AGEMA_signal_1242, n1942}) ) ;
    or_HPC1 #(.security_order(3), .pipeline(1)) U2026 ( .ina ({new_AGEMA_signal_1097, new_AGEMA_signal_1096, new_AGEMA_signal_1095, n2587}), .inb ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, new_AGEMA_signal_1065, n2815}), .clk ( clk ), .rnd ({Fresh[659], Fresh[658], Fresh[657], Fresh[656], Fresh[655], Fresh[654], Fresh[653], Fresh[652], Fresh[651], Fresh[650]}), .outt ({new_AGEMA_signal_1247, new_AGEMA_signal_1246, new_AGEMA_signal_1245, n2676}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2030 ( .ina ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, new_AGEMA_signal_1197, n2789}), .inb ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, new_AGEMA_signal_1011, n2559}), .clk ( clk ), .rnd ({Fresh[669], Fresh[668], Fresh[667], Fresh[666], Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660]}), .outt ({new_AGEMA_signal_1535, new_AGEMA_signal_1534, new_AGEMA_signal_1533, n1944}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2037 ( .ina ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2725}), .inb ({new_AGEMA_signal_1202, new_AGEMA_signal_1201, new_AGEMA_signal_1200, n2769}), .clk ( clk ), .rnd ({Fresh[679], Fresh[678], Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672], Fresh[671], Fresh[670]}), .outt ({new_AGEMA_signal_1538, new_AGEMA_signal_1537, new_AGEMA_signal_1536, n1950}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2039 ( .ina ({new_AGEMA_signal_12450, new_AGEMA_signal_12448, new_AGEMA_signal_12446, new_AGEMA_signal_12444}), .inb ({new_AGEMA_signal_1103, new_AGEMA_signal_1102, new_AGEMA_signal_1101, n2739}), .clk ( clk ), .rnd ({Fresh[689], Fresh[688], Fresh[687], Fresh[686], Fresh[685], Fresh[684], Fresh[683], Fresh[682], Fresh[681], Fresh[680]}), .outt ({new_AGEMA_signal_1256, new_AGEMA_signal_1255, new_AGEMA_signal_1254, n1949}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2042 ( .ina ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, new_AGEMA_signal_1032, n2750}), .inb ({new_AGEMA_signal_1070, new_AGEMA_signal_1069, new_AGEMA_signal_1068, n2600}), .clk ( clk ), .rnd ({Fresh[699], Fresh[698], Fresh[697], Fresh[696], Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690]}), .outt ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, new_AGEMA_signal_1257, n2677}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2043 ( .a ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, new_AGEMA_signal_1257, n2677}), .b ({new_AGEMA_signal_1541, new_AGEMA_signal_1540, new_AGEMA_signal_1539, n2662}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2047 ( .ina ({new_AGEMA_signal_1106, new_AGEMA_signal_1105, new_AGEMA_signal_1104, n2437}), .inb ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, new_AGEMA_signal_1107, n2778}), .clk ( clk ), .rnd ({Fresh[709], Fresh[708], Fresh[707], Fresh[706], Fresh[705], Fresh[704], Fresh[703], Fresh[702], Fresh[701], Fresh[700]}), .outt ({new_AGEMA_signal_1262, new_AGEMA_signal_1261, new_AGEMA_signal_1260, n2627}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2053 ( .ina ({new_AGEMA_signal_1043, new_AGEMA_signal_1042, new_AGEMA_signal_1041, n2816}), .inb ({new_AGEMA_signal_1112, new_AGEMA_signal_1111, new_AGEMA_signal_1110, n2452}), .clk ( clk ), .rnd ({Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714], Fresh[713], Fresh[712], Fresh[711], Fresh[710]}), .outt ({new_AGEMA_signal_1265, new_AGEMA_signal_1264, new_AGEMA_signal_1263, n1957}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2056 ( .ina ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2766}), .inb ({new_AGEMA_signal_1070, new_AGEMA_signal_1069, new_AGEMA_signal_1068, n2600}), .clk ( clk ), .rnd ({Fresh[729], Fresh[728], Fresh[727], Fresh[726], Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720]}), .outt ({new_AGEMA_signal_1544, new_AGEMA_signal_1543, new_AGEMA_signal_1542, n2088}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2062 ( .ina ({new_AGEMA_signal_998, new_AGEMA_signal_997, new_AGEMA_signal_996, n2519}), .inb ({new_AGEMA_signal_1010, new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2708}), .clk ( clk ), .rnd ({Fresh[739], Fresh[738], Fresh[737], Fresh[736], Fresh[735], Fresh[734], Fresh[733], Fresh[732], Fresh[731], Fresh[730]}), .outt ({new_AGEMA_signal_1115, new_AGEMA_signal_1114, new_AGEMA_signal_1113, n1964}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2063 ( .ina ({new_AGEMA_signal_12458, new_AGEMA_signal_12456, new_AGEMA_signal_12454, new_AGEMA_signal_12452}), .inb ({new_AGEMA_signal_1100, new_AGEMA_signal_1099, new_AGEMA_signal_1098, n2643}), .clk ( clk ), .rnd ({Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744], Fresh[743], Fresh[742], Fresh[741], Fresh[740]}), .outt ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, new_AGEMA_signal_1269, n2736}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2069 ( .ina ({new_AGEMA_signal_1118, new_AGEMA_signal_1117, new_AGEMA_signal_1116, n2772}), .inb ({new_AGEMA_signal_12466, new_AGEMA_signal_12464, new_AGEMA_signal_12462, new_AGEMA_signal_12460}), .clk ( clk ), .rnd ({Fresh[759], Fresh[758], Fresh[757], Fresh[756], Fresh[755], Fresh[754], Fresh[753], Fresh[752], Fresh[751], Fresh[750]}), .outt ({new_AGEMA_signal_1274, new_AGEMA_signal_1273, new_AGEMA_signal_1272, n2673}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2072 ( .ina ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2766}), .inb ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, n2612}), .clk ( clk ), .rnd ({Fresh[769], Fresh[768], Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762], Fresh[761], Fresh[760]}), .outt ({new_AGEMA_signal_1550, new_AGEMA_signal_1549, new_AGEMA_signal_1548, n2761}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2073 ( .a ({new_AGEMA_signal_1550, new_AGEMA_signal_1549, new_AGEMA_signal_1548, n2761}), .b ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, new_AGEMA_signal_2085, n2720}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2075 ( .ina ({new_AGEMA_signal_1280, new_AGEMA_signal_1279, new_AGEMA_signal_1278, n2313}), .inb ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2719}), .clk ( clk ), .rnd ({Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774], Fresh[773], Fresh[772], Fresh[771], Fresh[770]}), .outt ({new_AGEMA_signal_1553, new_AGEMA_signal_1552, new_AGEMA_signal_1551, n2412}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2076 ( .a ({new_AGEMA_signal_1553, new_AGEMA_signal_1552, new_AGEMA_signal_1551, n2412}), .b ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, new_AGEMA_signal_2088, n2417}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2079 ( .ina ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, new_AGEMA_signal_1029, n2641}), .inb ({new_AGEMA_signal_1016, new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2261}), .clk ( clk ), .rnd ({Fresh[789], Fresh[788], Fresh[787], Fresh[786], Fresh[785], Fresh[784], Fresh[783], Fresh[782], Fresh[781], Fresh[780]}), .outt ({new_AGEMA_signal_1283, new_AGEMA_signal_1282, new_AGEMA_signal_1281, n2571}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2080 ( .a ({new_AGEMA_signal_1283, new_AGEMA_signal_1282, new_AGEMA_signal_1281, n2571}), .b ({new_AGEMA_signal_1556, new_AGEMA_signal_1555, new_AGEMA_signal_1554, n2505}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2081 ( .ina ({new_AGEMA_signal_998, new_AGEMA_signal_997, new_AGEMA_signal_996, n2519}), .inb ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, new_AGEMA_signal_1119, n2824}), .clk ( clk ), .rnd ({Fresh[799], Fresh[798], Fresh[797], Fresh[796], Fresh[795], Fresh[794], Fresh[793], Fresh[792], Fresh[791], Fresh[790]}), .outt ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2083 ( .ina ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, n2792}), .inb ({new_AGEMA_signal_12466, new_AGEMA_signal_12464, new_AGEMA_signal_12462, new_AGEMA_signal_12460}), .clk ( clk ), .rnd ({Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804], Fresh[803], Fresh[802], Fresh[801], Fresh[800]}), .outt ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, new_AGEMA_signal_1557, n2359}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2086 ( .ina ({new_AGEMA_signal_998, new_AGEMA_signal_997, new_AGEMA_signal_996, n2519}), .inb ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, new_AGEMA_signal_1107, n2778}), .clk ( clk ), .rnd ({Fresh[819], Fresh[818], Fresh[817], Fresh[816], Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810]}), .outt ({new_AGEMA_signal_1289, new_AGEMA_signal_1288, new_AGEMA_signal_1287, n2101}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2087 ( .a ({new_AGEMA_signal_1289, new_AGEMA_signal_1288, new_AGEMA_signal_1287, n2101}), .b ({new_AGEMA_signal_1562, new_AGEMA_signal_1561, new_AGEMA_signal_1560, n2625}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2091 ( .ina ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2719}), .inb ({new_AGEMA_signal_1088, new_AGEMA_signal_1087, new_AGEMA_signal_1086, n2609}), .clk ( clk ), .rnd ({Fresh[829], Fresh[828], Fresh[827], Fresh[826], Fresh[825], Fresh[824], Fresh[823], Fresh[822], Fresh[821], Fresh[820]}), .outt ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, new_AGEMA_signal_1293, n2190}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2095 ( .ina ({new_AGEMA_signal_1103, new_AGEMA_signal_1102, new_AGEMA_signal_1101, n2739}), .inb ({new_AGEMA_signal_1019, new_AGEMA_signal_1018, new_AGEMA_signal_1017, n2779}), .clk ( clk ), .rnd ({Fresh[839], Fresh[838], Fresh[837], Fresh[836], Fresh[835], Fresh[834], Fresh[833], Fresh[832], Fresh[831], Fresh[830]}), .outt ({new_AGEMA_signal_1298, new_AGEMA_signal_1297, new_AGEMA_signal_1296, n1976}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2098 ( .ina ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}), .inb ({new_AGEMA_signal_1022, new_AGEMA_signal_1021, new_AGEMA_signal_1020, n2242}), .clk ( clk ), .rnd ({Fresh[849], Fresh[848], Fresh[847], Fresh[846], Fresh[845], Fresh[844], Fresh[843], Fresh[842], Fresh[841], Fresh[840]}), .outt ({new_AGEMA_signal_1568, new_AGEMA_signal_1567, new_AGEMA_signal_1566, n2535}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2101 ( .ina ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, new_AGEMA_signal_1209, n2688}), .inb ({new_AGEMA_signal_1130, new_AGEMA_signal_1129, new_AGEMA_signal_1128, n2356}), .clk ( clk ), .rnd ({Fresh[859], Fresh[858], Fresh[857], Fresh[856], Fresh[855], Fresh[854], Fresh[853], Fresh[852], Fresh[851], Fresh[850]}), .outt ({new_AGEMA_signal_1571, new_AGEMA_signal_1570, new_AGEMA_signal_1569, n1973}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2105 ( .ina ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, new_AGEMA_signal_1065, n2815}), .inb ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, new_AGEMA_signal_999, n2315}), .clk ( clk ), .rnd ({Fresh[869], Fresh[868], Fresh[867], Fresh[866], Fresh[865], Fresh[864], Fresh[863], Fresh[862], Fresh[861], Fresh[860]}), .outt ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, new_AGEMA_signal_1299, n2690}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2111 ( .ina ({new_AGEMA_signal_1094, new_AGEMA_signal_1093, new_AGEMA_signal_1092, n2493}), .inb ({new_AGEMA_signal_12474, new_AGEMA_signal_12472, new_AGEMA_signal_12470, new_AGEMA_signal_12468}), .clk ( clk ), .rnd ({Fresh[879], Fresh[878], Fresh[877], Fresh[876], Fresh[875], Fresh[874], Fresh[873], Fresh[872], Fresh[871], Fresh[870]}), .outt ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, new_AGEMA_signal_1302, n2817}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2113 ( .ina ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, n2442}), .inb ({new_AGEMA_signal_1019, new_AGEMA_signal_1018, new_AGEMA_signal_1017, n2779}), .clk ( clk ), .rnd ({Fresh[889], Fresh[888], Fresh[887], Fresh[886], Fresh[885], Fresh[884], Fresh[883], Fresh[882], Fresh[881], Fresh[880]}), .outt ({new_AGEMA_signal_1577, new_AGEMA_signal_1576, new_AGEMA_signal_1575, n2741}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2118 ( .ina ({new_AGEMA_signal_1046, new_AGEMA_signal_1045, new_AGEMA_signal_1044, n2780}), .inb ({new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2818}), .clk ( clk ), .rnd ({Fresh[899], Fresh[898], Fresh[897], Fresh[896], Fresh[895], Fresh[894], Fresh[893], Fresh[892], Fresh[891], Fresh[890]}), .outt ({new_AGEMA_signal_1580, new_AGEMA_signal_1579, new_AGEMA_signal_1578, n1992}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2120 ( .ina ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, new_AGEMA_signal_1305, n2823}), .inb ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}), .clk ( clk ), .rnd ({Fresh[909], Fresh[908], Fresh[907], Fresh[906], Fresh[905], Fresh[904], Fresh[903], Fresh[902], Fresh[901], Fresh[900]}), .outt ({new_AGEMA_signal_1583, new_AGEMA_signal_1582, new_AGEMA_signal_1581, n1991}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2123 ( .ina ({new_AGEMA_signal_1100, new_AGEMA_signal_1099, new_AGEMA_signal_1098, n2643}), .inb ({new_AGEMA_signal_1133, new_AGEMA_signal_1132, new_AGEMA_signal_1131, n2611}), .clk ( clk ), .rnd ({Fresh[919], Fresh[918], Fresh[917], Fresh[916], Fresh[915], Fresh[914], Fresh[913], Fresh[912], Fresh[911], Fresh[910]}), .outt ({new_AGEMA_signal_1310, new_AGEMA_signal_1309, new_AGEMA_signal_1308, n1993}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2125 ( .ina ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, new_AGEMA_signal_1191, n2737}), .inb ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, n2792}), .clk ( clk ), .rnd ({Fresh[929], Fresh[928], Fresh[927], Fresh[926], Fresh[925], Fresh[924], Fresh[923], Fresh[922], Fresh[921], Fresh[920]}), .outt ({new_AGEMA_signal_1586, new_AGEMA_signal_1585, new_AGEMA_signal_1584, n1995}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2132 ( .ina ({new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2818}), .inb ({new_AGEMA_signal_1010, new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2708}), .clk ( clk ), .rnd ({Fresh[939], Fresh[938], Fresh[937], Fresh[936], Fresh[935], Fresh[934], Fresh[933], Fresh[932], Fresh[931], Fresh[930]}), .outt ({new_AGEMA_signal_1589, new_AGEMA_signal_1588, new_AGEMA_signal_1587, n2241}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2135 ( .ina ({new_AGEMA_signal_12482, new_AGEMA_signal_12480, new_AGEMA_signal_12478, new_AGEMA_signal_12476}), .inb ({new_AGEMA_signal_1316, new_AGEMA_signal_1315, new_AGEMA_signal_1314, n2679}), .clk ( clk ), .rnd ({Fresh[949], Fresh[948], Fresh[947], Fresh[946], Fresh[945], Fresh[944], Fresh[943], Fresh[942], Fresh[941], Fresh[940]}), .outt ({new_AGEMA_signal_1592, new_AGEMA_signal_1591, new_AGEMA_signal_1590, n2003}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2140 ( .ina ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, n2612}), .inb ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, new_AGEMA_signal_1317, n2809}), .clk ( clk ), .rnd ({Fresh[959], Fresh[958], Fresh[957], Fresh[956], Fresh[955], Fresh[954], Fresh[953], Fresh[952], Fresh[951], Fresh[950]}), .outt ({new_AGEMA_signal_1595, new_AGEMA_signal_1594, new_AGEMA_signal_1593, n2008}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2141 ( .ina ({new_AGEMA_signal_1316, new_AGEMA_signal_1315, new_AGEMA_signal_1314, n2679}), .inb ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, new_AGEMA_signal_1209, n2688}), .clk ( clk ), .rnd ({Fresh[969], Fresh[968], Fresh[967], Fresh[966], Fresh[965], Fresh[964], Fresh[963], Fresh[962], Fresh[961], Fresh[960]}), .outt ({new_AGEMA_signal_1598, new_AGEMA_signal_1597, new_AGEMA_signal_1596, n2572}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2143 ( .ina ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, new_AGEMA_signal_1317, n2809}), .inb ({new_AGEMA_signal_1130, new_AGEMA_signal_1129, new_AGEMA_signal_1128, n2356}), .clk ( clk ), .rnd ({Fresh[979], Fresh[978], Fresh[977], Fresh[976], Fresh[975], Fresh[974], Fresh[973], Fresh[972], Fresh[971], Fresh[970]}), .outt ({new_AGEMA_signal_1601, new_AGEMA_signal_1600, new_AGEMA_signal_1599, n2004}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2147 ( .ina ({new_AGEMA_signal_992, new_AGEMA_signal_991, new_AGEMA_signal_990, n2635}), .inb ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}), .clk ( clk ), .rnd ({Fresh[989], Fresh[988], Fresh[987], Fresh[986], Fresh[985], Fresh[984], Fresh[983], Fresh[982], Fresh[981], Fresh[980]}), .outt ({new_AGEMA_signal_1604, new_AGEMA_signal_1603, new_AGEMA_signal_1602, n2009}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2151 ( .ina ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, new_AGEMA_signal_1197, n2789}), .inb ({new_AGEMA_signal_12474, new_AGEMA_signal_12472, new_AGEMA_signal_12470, new_AGEMA_signal_12468}), .clk ( clk ), .rnd ({Fresh[999], Fresh[998], Fresh[997], Fresh[996], Fresh[995], Fresh[994], Fresh[993], Fresh[992], Fresh[991], Fresh[990]}), .outt ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, new_AGEMA_signal_1605, n2533}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2157 ( .ina ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2719}), .inb ({new_AGEMA_signal_1004, new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2682}), .clk ( clk ), .rnd ({Fresh[1009], Fresh[1008], Fresh[1007], Fresh[1006], Fresh[1005], Fresh[1004], Fresh[1003], Fresh[1002], Fresh[1001], Fresh[1000]}), .outt ({new_AGEMA_signal_1325, new_AGEMA_signal_1324, new_AGEMA_signal_1323, n2026}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2158 ( .ina ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2766}), .inb ({new_AGEMA_signal_1094, new_AGEMA_signal_1093, new_AGEMA_signal_1092, n2493}), .clk ( clk ), .rnd ({Fresh[1019], Fresh[1018], Fresh[1017], Fresh[1016], Fresh[1015], Fresh[1014], Fresh[1013], Fresh[1012], Fresh[1011], Fresh[1010]}), .outt ({new_AGEMA_signal_1610, new_AGEMA_signal_1609, new_AGEMA_signal_1608, n2022}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2159 ( .ina ({new_AGEMA_signal_12490, new_AGEMA_signal_12488, new_AGEMA_signal_12486, new_AGEMA_signal_12484}), .inb ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2725}), .clk ( clk ), .rnd ({Fresh[1029], Fresh[1028], Fresh[1027], Fresh[1026], Fresh[1025], Fresh[1024], Fresh[1023], Fresh[1022], Fresh[1021], Fresh[1020]}), .outt ({new_AGEMA_signal_1328, new_AGEMA_signal_1327, new_AGEMA_signal_1326, n2227}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2167 ( .ina ({new_AGEMA_signal_995, new_AGEMA_signal_994, new_AGEMA_signal_993, n2790}), .inb ({new_AGEMA_signal_12474, new_AGEMA_signal_12472, new_AGEMA_signal_12470, new_AGEMA_signal_12468}), .clk ( clk ), .rnd ({Fresh[1039], Fresh[1038], Fresh[1037], Fresh[1036], Fresh[1035], Fresh[1034], Fresh[1033], Fresh[1032], Fresh[1031], Fresh[1030]}), .outt ({new_AGEMA_signal_1145, new_AGEMA_signal_1144, new_AGEMA_signal_1143, n2027}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2171 ( .ina ({new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2818}), .inb ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, n2442}), .clk ( clk ), .rnd ({Fresh[1049], Fresh[1048], Fresh[1047], Fresh[1046], Fresh[1045], Fresh[1044], Fresh[1043], Fresh[1042], Fresh[1041], Fresh[1040]}), .outt ({new_AGEMA_signal_1619, new_AGEMA_signal_1618, new_AGEMA_signal_1617, n2214}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2173 ( .ina ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, n2442}), .inb ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .clk ( clk ), .rnd ({Fresh[1059], Fresh[1058], Fresh[1057], Fresh[1056], Fresh[1055], Fresh[1054], Fresh[1053], Fresh[1052], Fresh[1051], Fresh[1050]}), .outt ({new_AGEMA_signal_1622, new_AGEMA_signal_1621, new_AGEMA_signal_1620, n2290}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2174 ( .ina ({new_AGEMA_signal_12458, new_AGEMA_signal_12456, new_AGEMA_signal_12454, new_AGEMA_signal_12452}), .inb ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2767}), .clk ( clk ), .rnd ({Fresh[1069], Fresh[1068], Fresh[1067], Fresh[1066], Fresh[1065], Fresh[1064], Fresh[1063], Fresh[1062], Fresh[1061], Fresh[1060]}), .outt ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, new_AGEMA_signal_1623, n2376}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2178 ( .ina ({new_AGEMA_signal_1010, new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2708}), .inb ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, new_AGEMA_signal_1080, n2400}), .clk ( clk ), .rnd ({Fresh[1079], Fresh[1078], Fresh[1077], Fresh[1076], Fresh[1075], Fresh[1074], Fresh[1073], Fresh[1072], Fresh[1071], Fresh[1070]}), .outt ({new_AGEMA_signal_1334, new_AGEMA_signal_1333, new_AGEMA_signal_1332, n2034}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2182 ( .ina ({new_AGEMA_signal_1133, new_AGEMA_signal_1132, new_AGEMA_signal_1131, n2611}), .inb ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2719}), .clk ( clk ), .rnd ({Fresh[1089], Fresh[1088], Fresh[1087], Fresh[1086], Fresh[1085], Fresh[1084], Fresh[1083], Fresh[1082], Fresh[1081], Fresh[1080]}), .outt ({new_AGEMA_signal_1337, new_AGEMA_signal_1336, new_AGEMA_signal_1335, n2171}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2183 ( .ina ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, new_AGEMA_signal_1311, n2828}), .inb ({new_AGEMA_signal_1202, new_AGEMA_signal_1201, new_AGEMA_signal_1200, n2769}), .clk ( clk ), .rnd ({Fresh[1099], Fresh[1098], Fresh[1097], Fresh[1096], Fresh[1095], Fresh[1094], Fresh[1093], Fresh[1092], Fresh[1091], Fresh[1090]}), .outt ({new_AGEMA_signal_1628, new_AGEMA_signal_1627, new_AGEMA_signal_1626, n2039}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2188 ( .ina ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2725}), .inb ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .clk ( clk ), .rnd ({Fresh[1109], Fresh[1108], Fresh[1107], Fresh[1106], Fresh[1105], Fresh[1104], Fresh[1103], Fresh[1102], Fresh[1101], Fresh[1100]}), .outt ({new_AGEMA_signal_1634, new_AGEMA_signal_1633, new_AGEMA_signal_1632, n2042}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2191 ( .ina ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .inb ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, new_AGEMA_signal_999, n2315}), .clk ( clk ), .rnd ({Fresh[1119], Fresh[1118], Fresh[1117], Fresh[1116], Fresh[1115], Fresh[1114], Fresh[1113], Fresh[1112], Fresh[1111], Fresh[1110]}), .outt ({new_AGEMA_signal_1637, new_AGEMA_signal_1636, new_AGEMA_signal_1635, n2754}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2192 ( .ina ({new_AGEMA_signal_1280, new_AGEMA_signal_1279, new_AGEMA_signal_1278, n2313}), .inb ({new_AGEMA_signal_995, new_AGEMA_signal_994, new_AGEMA_signal_993, n2790}), .clk ( clk ), .rnd ({Fresh[1129], Fresh[1128], Fresh[1127], Fresh[1126], Fresh[1125], Fresh[1124], Fresh[1123], Fresh[1122], Fresh[1121], Fresh[1120]}), .outt ({new_AGEMA_signal_1640, new_AGEMA_signal_1639, new_AGEMA_signal_1638, n2044}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2198 ( .ina ({new_AGEMA_signal_1280, new_AGEMA_signal_1279, new_AGEMA_signal_1278, n2313}), .inb ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, new_AGEMA_signal_1029, n2641}), .clk ( clk ), .rnd ({Fresh[1139], Fresh[1138], Fresh[1137], Fresh[1136], Fresh[1135], Fresh[1134], Fresh[1133], Fresh[1132], Fresh[1131], Fresh[1130]}), .outt ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, new_AGEMA_signal_1641, n2654}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2202 ( .ina ({new_AGEMA_signal_992, new_AGEMA_signal_991, new_AGEMA_signal_990, n2635}), .inb ({new_AGEMA_signal_1229, new_AGEMA_signal_1228, new_AGEMA_signal_1227, n2577}), .clk ( clk ), .rnd ({Fresh[1149], Fresh[1148], Fresh[1147], Fresh[1146], Fresh[1145], Fresh[1144], Fresh[1143], Fresh[1142], Fresh[1141], Fresh[1140]}), .outt ({new_AGEMA_signal_1646, new_AGEMA_signal_1645, new_AGEMA_signal_1644, n2055}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2205 ( .ina ({new_AGEMA_signal_1124, new_AGEMA_signal_1123, new_AGEMA_signal_1122, n2395}), .inb ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2767}), .clk ( clk ), .rnd ({Fresh[1159], Fresh[1158], Fresh[1157], Fresh[1156], Fresh[1155], Fresh[1154], Fresh[1153], Fresh[1152], Fresh[1151], Fresh[1150]}), .outt ({new_AGEMA_signal_1649, new_AGEMA_signal_1648, new_AGEMA_signal_1647, n2057}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2208 ( .ina ({new_AGEMA_signal_1316, new_AGEMA_signal_1315, new_AGEMA_signal_1314, n2679}), .inb ({new_AGEMA_signal_1004, new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2682}), .clk ( clk ), .rnd ({Fresh[1169], Fresh[1168], Fresh[1167], Fresh[1166], Fresh[1165], Fresh[1164], Fresh[1163], Fresh[1162], Fresh[1161], Fresh[1160]}), .outt ({new_AGEMA_signal_1652, new_AGEMA_signal_1651, new_AGEMA_signal_1650, n2407}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2212 ( .ina ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, new_AGEMA_signal_1209, n2688}), .inb ({new_AGEMA_signal_1148, new_AGEMA_signal_1147, new_AGEMA_signal_1146, n2061}), .clk ( clk ), .rnd ({Fresh[1179], Fresh[1178], Fresh[1177], Fresh[1176], Fresh[1175], Fresh[1174], Fresh[1173], Fresh[1172], Fresh[1171], Fresh[1170]}), .outt ({new_AGEMA_signal_1655, new_AGEMA_signal_1654, new_AGEMA_signal_1653, n2062}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2216 ( .ina ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2766}), .inb ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, new_AGEMA_signal_1011, n2559}), .clk ( clk ), .rnd ({Fresh[1189], Fresh[1188], Fresh[1187], Fresh[1186], Fresh[1185], Fresh[1184], Fresh[1183], Fresh[1182], Fresh[1181], Fresh[1180]}), .outt ({new_AGEMA_signal_1658, new_AGEMA_signal_1657, new_AGEMA_signal_1656, n2731}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2220 ( .a ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, new_AGEMA_signal_1299, n2690}), .b ({new_AGEMA_signal_1661, new_AGEMA_signal_1660, new_AGEMA_signal_1659, n2068}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2224 ( .ina ({new_AGEMA_signal_1133, new_AGEMA_signal_1132, new_AGEMA_signal_1131, n2611}), .inb ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, new_AGEMA_signal_1032, n2750}), .clk ( clk ), .rnd ({Fresh[1199], Fresh[1198], Fresh[1197], Fresh[1196], Fresh[1195], Fresh[1194], Fresh[1193], Fresh[1192], Fresh[1191], Fresh[1190]}), .outt ({new_AGEMA_signal_1340, new_AGEMA_signal_1339, new_AGEMA_signal_1338, n2642}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2225 ( .ina ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2725}), .inb ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, n2786}), .clk ( clk ), .rnd ({Fresh[1209], Fresh[1208], Fresh[1207], Fresh[1206], Fresh[1205], Fresh[1204], Fresh[1203], Fresh[1202], Fresh[1201], Fresh[1200]}), .outt ({new_AGEMA_signal_1664, new_AGEMA_signal_1663, new_AGEMA_signal_1662, n2252}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2228 ( .ina ({new_AGEMA_signal_1103, new_AGEMA_signal_1102, new_AGEMA_signal_1101, n2739}), .inb ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, new_AGEMA_signal_1065, n2815}), .clk ( clk ), .rnd ({Fresh[1219], Fresh[1218], Fresh[1217], Fresh[1216], Fresh[1215], Fresh[1214], Fresh[1213], Fresh[1212], Fresh[1211], Fresh[1210]}), .outt ({new_AGEMA_signal_1343, new_AGEMA_signal_1342, new_AGEMA_signal_1341, n2075}) ) ;
    or_HPC1 #(.security_order(3), .pipeline(1)) U2233 ( .ina ({new_AGEMA_signal_992, new_AGEMA_signal_991, new_AGEMA_signal_990, n2635}), .inb ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, new_AGEMA_signal_1059, n2723}), .clk ( clk ), .rnd ({Fresh[1229], Fresh[1228], Fresh[1227], Fresh[1226], Fresh[1225], Fresh[1224], Fresh[1223], Fresh[1222], Fresh[1221], Fresh[1220]}), .outt ({new_AGEMA_signal_1346, new_AGEMA_signal_1345, new_AGEMA_signal_1344, n2081}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2234 ( .ina ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, n2792}), .inb ({new_AGEMA_signal_1004, new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2682}), .clk ( clk ), .rnd ({Fresh[1239], Fresh[1238], Fresh[1237], Fresh[1236], Fresh[1235], Fresh[1234], Fresh[1233], Fresh[1232], Fresh[1231], Fresh[1230]}), .outt ({new_AGEMA_signal_1667, new_AGEMA_signal_1666, new_AGEMA_signal_1665, n2080}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2237 ( .ina ({new_AGEMA_signal_1070, new_AGEMA_signal_1069, new_AGEMA_signal_1068, n2600}), .inb ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2719}), .clk ( clk ), .rnd ({Fresh[1249], Fresh[1248], Fresh[1247], Fresh[1246], Fresh[1245], Fresh[1244], Fresh[1243], Fresh[1242], Fresh[1241], Fresh[1240]}), .outt ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, n2498}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2238 ( .a ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, n2498}), .b ({new_AGEMA_signal_1670, new_AGEMA_signal_1669, new_AGEMA_signal_1668, n2773}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2239 ( .ina ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2767}), .inb ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, n2792}), .clk ( clk ), .rnd ({Fresh[1259], Fresh[1258], Fresh[1257], Fresh[1256], Fresh[1255], Fresh[1254], Fresh[1253], Fresh[1252], Fresh[1251], Fresh[1250]}), .outt ({new_AGEMA_signal_1673, new_AGEMA_signal_1672, new_AGEMA_signal_1671, n2083}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2244 ( .ina ({new_AGEMA_signal_12482, new_AGEMA_signal_12480, new_AGEMA_signal_12478, new_AGEMA_signal_12476}), .inb ({new_AGEMA_signal_1217, new_AGEMA_signal_1216, new_AGEMA_signal_1215, n2086}), .clk ( clk ), .rnd ({Fresh[1269], Fresh[1268], Fresh[1267], Fresh[1266], Fresh[1265], Fresh[1264], Fresh[1263], Fresh[1262], Fresh[1261], Fresh[1260]}), .outt ({new_AGEMA_signal_1676, new_AGEMA_signal_1675, new_AGEMA_signal_1674, n2562}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2247 ( .ina ({new_AGEMA_signal_12458, new_AGEMA_signal_12456, new_AGEMA_signal_12454, new_AGEMA_signal_12452}), .inb ({new_AGEMA_signal_1091, new_AGEMA_signal_1090, new_AGEMA_signal_1089, n2661}), .clk ( clk ), .rnd ({Fresh[1279], Fresh[1278], Fresh[1277], Fresh[1276], Fresh[1275], Fresh[1274], Fresh[1273], Fresh[1272], Fresh[1271], Fresh[1270]}), .outt ({new_AGEMA_signal_1352, new_AGEMA_signal_1351, new_AGEMA_signal_1350, n2087}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2251 ( .ina ({new_AGEMA_signal_1139, new_AGEMA_signal_1138, new_AGEMA_signal_1137, n2563}), .inb ({new_AGEMA_signal_1241, new_AGEMA_signal_1240, new_AGEMA_signal_1239, n2174}), .clk ( clk ), .rnd ({Fresh[1289], Fresh[1288], Fresh[1287], Fresh[1286], Fresh[1285], Fresh[1284], Fresh[1283], Fresh[1282], Fresh[1281], Fresh[1280]}), .outt ({new_AGEMA_signal_1679, new_AGEMA_signal_1678, new_AGEMA_signal_1677, n2156}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2260 ( .ina ({new_AGEMA_signal_1202, new_AGEMA_signal_1201, new_AGEMA_signal_1200, n2769}), .inb ({new_AGEMA_signal_1142, new_AGEMA_signal_1141, new_AGEMA_signal_1140, n2401}), .clk ( clk ), .rnd ({Fresh[1299], Fresh[1298], Fresh[1297], Fresh[1296], Fresh[1295], Fresh[1294], Fresh[1293], Fresh[1292], Fresh[1291], Fresh[1290]}), .outt ({new_AGEMA_signal_1682, new_AGEMA_signal_1681, new_AGEMA_signal_1680, n2100}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2277 ( .ina ({new_AGEMA_signal_1103, new_AGEMA_signal_1102, new_AGEMA_signal_1101, n2739}), .inb ({new_AGEMA_signal_1154, new_AGEMA_signal_1153, new_AGEMA_signal_1152, n2298}), .clk ( clk ), .rnd ({Fresh[1309], Fresh[1308], Fresh[1307], Fresh[1306], Fresh[1305], Fresh[1304], Fresh[1303], Fresh[1302], Fresh[1301], Fresh[1300]}), .outt ({new_AGEMA_signal_1355, new_AGEMA_signal_1354, new_AGEMA_signal_1353, n2544}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2279 ( .ina ({new_AGEMA_signal_1130, new_AGEMA_signal_1129, new_AGEMA_signal_1128, n2356}), .inb ({new_AGEMA_signal_1358, new_AGEMA_signal_1357, new_AGEMA_signal_1356, n2118}), .clk ( clk ), .rnd ({Fresh[1319], Fresh[1318], Fresh[1317], Fresh[1316], Fresh[1315], Fresh[1314], Fresh[1313], Fresh[1312], Fresh[1311], Fresh[1310]}), .outt ({new_AGEMA_signal_1691, new_AGEMA_signal_1690, new_AGEMA_signal_1689, n2121}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2284 ( .ina ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .inb ({new_AGEMA_signal_1250, new_AGEMA_signal_1249, new_AGEMA_signal_1248, n2570}), .clk ( clk ), .rnd ({Fresh[1329], Fresh[1328], Fresh[1327], Fresh[1326], Fresh[1325], Fresh[1324], Fresh[1323], Fresh[1322], Fresh[1321], Fresh[1320]}), .outt ({new_AGEMA_signal_1697, new_AGEMA_signal_1696, new_AGEMA_signal_1695, n2122}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2286 ( .ina ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, n2792}), .inb ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, n2612}), .clk ( clk ), .rnd ({Fresh[1339], Fresh[1338], Fresh[1337], Fresh[1336], Fresh[1335], Fresh[1334], Fresh[1333], Fresh[1332], Fresh[1331], Fresh[1330]}), .outt ({new_AGEMA_signal_1700, new_AGEMA_signal_1699, new_AGEMA_signal_1698, n2811}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2294 ( .ina ({new_AGEMA_signal_1106, new_AGEMA_signal_1105, new_AGEMA_signal_1104, n2437}), .inb ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2742}), .clk ( clk ), .rnd ({Fresh[1349], Fresh[1348], Fresh[1347], Fresh[1346], Fresh[1345], Fresh[1344], Fresh[1343], Fresh[1342], Fresh[1341], Fresh[1340]}), .outt ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, new_AGEMA_signal_1359, n2647}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2297 ( .ina ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2742}), .inb ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, new_AGEMA_signal_999, n2315}), .clk ( clk ), .rnd ({Fresh[1359], Fresh[1358], Fresh[1357], Fresh[1356], Fresh[1355], Fresh[1354], Fresh[1353], Fresh[1352], Fresh[1351], Fresh[1350]}), .outt ({new_AGEMA_signal_1364, new_AGEMA_signal_1363, new_AGEMA_signal_1362, n2132}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2304 ( .ina ({new_AGEMA_signal_1136, new_AGEMA_signal_1135, new_AGEMA_signal_1134, n2616}), .inb ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .clk ( clk ), .rnd ({Fresh[1369], Fresh[1368], Fresh[1367], Fresh[1366], Fresh[1365], Fresh[1364], Fresh[1363], Fresh[1362], Fresh[1361], Fresh[1360]}), .outt ({new_AGEMA_signal_1715, new_AGEMA_signal_1714, new_AGEMA_signal_1713, n2220}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2305 ( .ina ({new_AGEMA_signal_12434, new_AGEMA_signal_12432, new_AGEMA_signal_12430, new_AGEMA_signal_12428}), .inb ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2767}), .clk ( clk ), .rnd ({Fresh[1379], Fresh[1378], Fresh[1377], Fresh[1376], Fresh[1375], Fresh[1374], Fresh[1373], Fresh[1372], Fresh[1371], Fresh[1370]}), .outt ({new_AGEMA_signal_1718, new_AGEMA_signal_1717, new_AGEMA_signal_1716, n2138}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2312 ( .ina ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, n2612}), .inb ({new_AGEMA_signal_12498, new_AGEMA_signal_12496, new_AGEMA_signal_12494, new_AGEMA_signal_12492}), .clk ( clk ), .rnd ({Fresh[1389], Fresh[1388], Fresh[1387], Fresh[1386], Fresh[1385], Fresh[1384], Fresh[1383], Fresh[1382], Fresh[1381], Fresh[1380]}), .outt ({new_AGEMA_signal_1721, new_AGEMA_signal_1720, new_AGEMA_signal_1719, n2555}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2322 ( .ina ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, n2612}), .inb ({new_AGEMA_signal_12506, new_AGEMA_signal_12504, new_AGEMA_signal_12502, new_AGEMA_signal_12500}), .clk ( clk ), .rnd ({Fresh[1399], Fresh[1398], Fresh[1397], Fresh[1396], Fresh[1395], Fresh[1394], Fresh[1393], Fresh[1392], Fresh[1391], Fresh[1390]}), .outt ({new_AGEMA_signal_1724, new_AGEMA_signal_1723, new_AGEMA_signal_1722, n2429}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2328 ( .ina ({new_AGEMA_signal_1106, new_AGEMA_signal_1105, new_AGEMA_signal_1104, n2437}), .inb ({new_AGEMA_signal_12474, new_AGEMA_signal_12472, new_AGEMA_signal_12470, new_AGEMA_signal_12468}), .clk ( clk ), .rnd ({Fresh[1409], Fresh[1408], Fresh[1407], Fresh[1406], Fresh[1405], Fresh[1404], Fresh[1403], Fresh[1402], Fresh[1401], Fresh[1400]}), .outt ({new_AGEMA_signal_1367, new_AGEMA_signal_1366, new_AGEMA_signal_1365, n2162}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2337 ( .ina ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, new_AGEMA_signal_999, n2315}), .inb ({new_AGEMA_signal_1022, new_AGEMA_signal_1021, new_AGEMA_signal_1020, n2242}), .clk ( clk ), .rnd ({Fresh[1419], Fresh[1418], Fresh[1417], Fresh[1416], Fresh[1415], Fresh[1414], Fresh[1413], Fresh[1412], Fresh[1411], Fresh[1410]}), .outt ({new_AGEMA_signal_1160, new_AGEMA_signal_1159, new_AGEMA_signal_1158, n2545}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2340 ( .ina ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, new_AGEMA_signal_1011, n2559}), .inb ({new_AGEMA_signal_1100, new_AGEMA_signal_1099, new_AGEMA_signal_1098, n2643}), .clk ( clk ), .rnd ({Fresh[1429], Fresh[1428], Fresh[1427], Fresh[1426], Fresh[1425], Fresh[1424], Fresh[1423], Fresh[1422], Fresh[1421], Fresh[1420]}), .outt ({new_AGEMA_signal_1373, new_AGEMA_signal_1372, new_AGEMA_signal_1371, n2178}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2342 ( .ina ({new_AGEMA_signal_1163, new_AGEMA_signal_1162, new_AGEMA_signal_1161, n2430}), .inb ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .clk ( clk ), .rnd ({Fresh[1439], Fresh[1438], Fresh[1437], Fresh[1436], Fresh[1435], Fresh[1434], Fresh[1433], Fresh[1432], Fresh[1431], Fresh[1430]}), .outt ({new_AGEMA_signal_1730, new_AGEMA_signal_1729, new_AGEMA_signal_1728, n2176}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2343 ( .ina ({new_AGEMA_signal_1241, new_AGEMA_signal_1240, new_AGEMA_signal_1239, n2174}), .inb ({new_AGEMA_signal_12482, new_AGEMA_signal_12480, new_AGEMA_signal_12478, new_AGEMA_signal_12476}), .clk ( clk ), .rnd ({Fresh[1449], Fresh[1448], Fresh[1447], Fresh[1446], Fresh[1445], Fresh[1444], Fresh[1443], Fresh[1442], Fresh[1441], Fresh[1440]}), .outt ({new_AGEMA_signal_1733, new_AGEMA_signal_1732, new_AGEMA_signal_1731, n2175}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2348 ( .ina ({new_AGEMA_signal_1016, new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2261}), .inb ({new_AGEMA_signal_12506, new_AGEMA_signal_12504, new_AGEMA_signal_12502, new_AGEMA_signal_12500}), .clk ( clk ), .rnd ({Fresh[1459], Fresh[1458], Fresh[1457], Fresh[1456], Fresh[1455], Fresh[1454], Fresh[1453], Fresh[1452], Fresh[1451], Fresh[1450]}), .outt ({new_AGEMA_signal_1166, new_AGEMA_signal_1165, new_AGEMA_signal_1164, n2182}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2353 ( .ina ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, n2786}), .inb ({new_AGEMA_signal_1163, new_AGEMA_signal_1162, new_AGEMA_signal_1161, n2430}), .clk ( clk ), .rnd ({Fresh[1469], Fresh[1468], Fresh[1467], Fresh[1466], Fresh[1465], Fresh[1464], Fresh[1463], Fresh[1462], Fresh[1461], Fresh[1460]}), .outt ({new_AGEMA_signal_1736, new_AGEMA_signal_1735, new_AGEMA_signal_1734, n2188}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2355 ( .ina ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, n2792}), .inb ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, n2612}), .clk ( clk ), .rnd ({Fresh[1479], Fresh[1478], Fresh[1477], Fresh[1476], Fresh[1475], Fresh[1474], Fresh[1473], Fresh[1472], Fresh[1471], Fresh[1470]}), .outt ({new_AGEMA_signal_1739, new_AGEMA_signal_1738, new_AGEMA_signal_1737, n2189}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2357 ( .ina ({new_AGEMA_signal_992, new_AGEMA_signal_991, new_AGEMA_signal_990, n2635}), .inb ({new_AGEMA_signal_1202, new_AGEMA_signal_1201, new_AGEMA_signal_1200, n2769}), .clk ( clk ), .rnd ({Fresh[1489], Fresh[1488], Fresh[1487], Fresh[1486], Fresh[1485], Fresh[1484], Fresh[1483], Fresh[1482], Fresh[1481], Fresh[1480]}), .outt ({new_AGEMA_signal_1742, new_AGEMA_signal_1741, new_AGEMA_signal_1740, n2446}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2362 ( .ina ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, new_AGEMA_signal_1032, n2750}), .inb ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, new_AGEMA_signal_1011, n2559}), .clk ( clk ), .rnd ({Fresh[1499], Fresh[1498], Fresh[1497], Fresh[1496], Fresh[1495], Fresh[1494], Fresh[1493], Fresh[1492], Fresh[1491], Fresh[1490]}), .outt ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, new_AGEMA_signal_1377, n2576}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2363 ( .ina ({new_AGEMA_signal_1088, new_AGEMA_signal_1087, new_AGEMA_signal_1086, n2609}), .inb ({new_AGEMA_signal_12514, new_AGEMA_signal_12512, new_AGEMA_signal_12510, new_AGEMA_signal_12508}), .clk ( clk ), .rnd ({Fresh[1509], Fresh[1508], Fresh[1507], Fresh[1506], Fresh[1505], Fresh[1504], Fresh[1503], Fresh[1502], Fresh[1501], Fresh[1500]}), .outt ({new_AGEMA_signal_1382, new_AGEMA_signal_1381, new_AGEMA_signal_1380, n2748}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2368 ( .a ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, new_AGEMA_signal_1641, n2654}), .b ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, new_AGEMA_signal_2241, n2674}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2378 ( .ina ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, new_AGEMA_signal_1065, n2815}), .inb ({new_AGEMA_signal_1010, new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2708}), .clk ( clk ), .rnd ({Fresh[1519], Fresh[1518], Fresh[1517], Fresh[1516], Fresh[1515], Fresh[1514], Fresh[1513], Fresh[1512], Fresh[1511], Fresh[1510]}), .outt ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, new_AGEMA_signal_1383, n2213}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2380 ( .ina ({new_AGEMA_signal_1043, new_AGEMA_signal_1042, new_AGEMA_signal_1041, n2816}), .inb ({new_AGEMA_signal_12458, new_AGEMA_signal_12456, new_AGEMA_signal_12454, new_AGEMA_signal_12452}), .clk ( clk ), .rnd ({Fresh[1529], Fresh[1528], Fresh[1527], Fresh[1526], Fresh[1525], Fresh[1524], Fresh[1523], Fresh[1522], Fresh[1521], Fresh[1520]}), .outt ({new_AGEMA_signal_1388, new_AGEMA_signal_1387, new_AGEMA_signal_1386, n2215}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2384 ( .ina ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, new_AGEMA_signal_1023, n2712}), .inb ({new_AGEMA_signal_1202, new_AGEMA_signal_1201, new_AGEMA_signal_1200, n2769}), .clk ( clk ), .rnd ({Fresh[1539], Fresh[1538], Fresh[1537], Fresh[1536], Fresh[1535], Fresh[1534], Fresh[1533], Fresh[1532], Fresh[1531], Fresh[1530]}), .outt ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, new_AGEMA_signal_1749, n2218}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2386 ( .ina ({new_AGEMA_signal_1154, new_AGEMA_signal_1153, new_AGEMA_signal_1152, n2298}), .inb ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}), .clk ( clk ), .rnd ({Fresh[1549], Fresh[1548], Fresh[1547], Fresh[1546], Fresh[1545], Fresh[1544], Fresh[1543], Fresh[1542], Fresh[1541], Fresh[1540]}), .outt ({new_AGEMA_signal_1754, new_AGEMA_signal_1753, new_AGEMA_signal_1752, n2219}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2405 ( .ina ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .inb ({new_AGEMA_signal_1058, new_AGEMA_signal_1057, new_AGEMA_signal_1056, n2713}), .clk ( clk ), .rnd ({Fresh[1559], Fresh[1558], Fresh[1557], Fresh[1556], Fresh[1555], Fresh[1554], Fresh[1553], Fresh[1552], Fresh[1551], Fresh[1550]}), .outt ({new_AGEMA_signal_1769, new_AGEMA_signal_1768, new_AGEMA_signal_1767, n2240}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2407 ( .ina ({new_AGEMA_signal_1322, new_AGEMA_signal_1321, new_AGEMA_signal_1320, n2709}), .inb ({new_AGEMA_signal_1022, new_AGEMA_signal_1021, new_AGEMA_signal_1020, n2242}), .clk ( clk ), .rnd ({Fresh[1569], Fresh[1568], Fresh[1567], Fresh[1566], Fresh[1565], Fresh[1564], Fresh[1563], Fresh[1562], Fresh[1561], Fresh[1560]}), .outt ({new_AGEMA_signal_1772, new_AGEMA_signal_1771, new_AGEMA_signal_1770, n2561}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2408 ( .ina ({new_AGEMA_signal_12482, new_AGEMA_signal_12480, new_AGEMA_signal_12478, new_AGEMA_signal_12476}), .inb ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, n2442}), .clk ( clk ), .rnd ({Fresh[1579], Fresh[1578], Fresh[1577], Fresh[1576], Fresh[1575], Fresh[1574], Fresh[1573], Fresh[1572], Fresh[1571], Fresh[1570]}), .outt ({new_AGEMA_signal_1775, new_AGEMA_signal_1774, new_AGEMA_signal_1773, n2243}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2411 ( .ina ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, new_AGEMA_signal_1035, n2615}), .inb ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, n2442}), .clk ( clk ), .rnd ({Fresh[1589], Fresh[1588], Fresh[1587], Fresh[1586], Fresh[1585], Fresh[1584], Fresh[1583], Fresh[1582], Fresh[1581], Fresh[1580]}), .outt ({new_AGEMA_signal_1778, new_AGEMA_signal_1777, new_AGEMA_signal_1776, n2245}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2422 ( .ina ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}), .inb ({new_AGEMA_signal_1163, new_AGEMA_signal_1162, new_AGEMA_signal_1161, n2430}), .clk ( clk ), .rnd ({Fresh[1599], Fresh[1598], Fresh[1597], Fresh[1596], Fresh[1595], Fresh[1594], Fresh[1593], Fresh[1592], Fresh[1591], Fresh[1590]}), .outt ({new_AGEMA_signal_1781, new_AGEMA_signal_1780, new_AGEMA_signal_1779, n2540}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2423 ( .ina ({new_AGEMA_signal_1016, new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2261}), .inb ({new_AGEMA_signal_1190, new_AGEMA_signal_1189, new_AGEMA_signal_1188, n2640}), .clk ( clk ), .rnd ({Fresh[1609], Fresh[1608], Fresh[1607], Fresh[1606], Fresh[1605], Fresh[1604], Fresh[1603], Fresh[1602], Fresh[1601], Fresh[1600]}), .outt ({new_AGEMA_signal_1784, new_AGEMA_signal_1783, new_AGEMA_signal_1782, n2259}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2426 ( .ina ({new_AGEMA_signal_1016, new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2261}), .inb ({new_AGEMA_signal_1091, new_AGEMA_signal_1090, new_AGEMA_signal_1089, n2661}), .clk ( clk ), .rnd ({Fresh[1619], Fresh[1618], Fresh[1617], Fresh[1616], Fresh[1615], Fresh[1614], Fresh[1613], Fresh[1612], Fresh[1611], Fresh[1610]}), .outt ({new_AGEMA_signal_1391, new_AGEMA_signal_1390, new_AGEMA_signal_1389, n2262}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2431 ( .ina ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, new_AGEMA_signal_999, n2315}), .inb ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, new_AGEMA_signal_1167, n2777}), .clk ( clk ), .rnd ({Fresh[1629], Fresh[1628], Fresh[1627], Fresh[1626], Fresh[1625], Fresh[1624], Fresh[1623], Fresh[1622], Fresh[1621], Fresh[1620]}), .outt ({new_AGEMA_signal_1394, new_AGEMA_signal_1393, new_AGEMA_signal_1392, n2266}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2432 ( .ina ({new_AGEMA_signal_1118, new_AGEMA_signal_1117, new_AGEMA_signal_1116, n2772}), .inb ({new_AGEMA_signal_12506, new_AGEMA_signal_12504, new_AGEMA_signal_12502, new_AGEMA_signal_12500}), .clk ( clk ), .rnd ({Fresh[1639], Fresh[1638], Fresh[1637], Fresh[1636], Fresh[1635], Fresh[1634], Fresh[1633], Fresh[1632], Fresh[1631], Fresh[1630]}), .outt ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, new_AGEMA_signal_1395, n2645}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2436 ( .ina ({new_AGEMA_signal_12434, new_AGEMA_signal_12432, new_AGEMA_signal_12430, new_AGEMA_signal_12428}), .inb ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2725}), .clk ( clk ), .rnd ({Fresh[1649], Fresh[1648], Fresh[1647], Fresh[1646], Fresh[1645], Fresh[1644], Fresh[1643], Fresh[1642], Fresh[1641], Fresh[1640]}), .outt ({new_AGEMA_signal_1400, new_AGEMA_signal_1399, new_AGEMA_signal_1398, n2268}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2443 ( .ina ({new_AGEMA_signal_1043, new_AGEMA_signal_1042, new_AGEMA_signal_1041, n2816}), .inb ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, n2786}), .clk ( clk ), .rnd ({Fresh[1659], Fresh[1658], Fresh[1657], Fresh[1656], Fresh[1655], Fresh[1654], Fresh[1653], Fresh[1652], Fresh[1651], Fresh[1650]}), .outt ({new_AGEMA_signal_1793, new_AGEMA_signal_1792, new_AGEMA_signal_1791, n2278}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2448 ( .ina ({new_AGEMA_signal_12522, new_AGEMA_signal_12520, new_AGEMA_signal_12518, new_AGEMA_signal_12516}), .inb ({new_AGEMA_signal_1058, new_AGEMA_signal_1057, new_AGEMA_signal_1056, n2713}), .clk ( clk ), .rnd ({Fresh[1669], Fresh[1668], Fresh[1667], Fresh[1666], Fresh[1665], Fresh[1664], Fresh[1663], Fresh[1662], Fresh[1661], Fresh[1660]}), .outt ({new_AGEMA_signal_1403, new_AGEMA_signal_1402, new_AGEMA_signal_1401, n2383}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2455 ( .ina ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, new_AGEMA_signal_1107, n2778}), .inb ({new_AGEMA_signal_1250, new_AGEMA_signal_1249, new_AGEMA_signal_1248, n2570}), .clk ( clk ), .rnd ({Fresh[1679], Fresh[1678], Fresh[1677], Fresh[1676], Fresh[1675], Fresh[1674], Fresh[1673], Fresh[1672], Fresh[1671], Fresh[1670]}), .outt ({new_AGEMA_signal_1802, new_AGEMA_signal_1801, new_AGEMA_signal_1800, n2774}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2458 ( .ina ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, new_AGEMA_signal_1305, n2823}), .inb ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, new_AGEMA_signal_1107, n2778}), .clk ( clk ), .rnd ({Fresh[1689], Fresh[1688], Fresh[1687], Fresh[1686], Fresh[1685], Fresh[1684], Fresh[1683], Fresh[1682], Fresh[1681], Fresh[1680]}), .outt ({new_AGEMA_signal_1805, new_AGEMA_signal_1804, new_AGEMA_signal_1803, n2287}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2470 ( .ina ({new_AGEMA_signal_998, new_AGEMA_signal_997, new_AGEMA_signal_996, n2519}), .inb ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .clk ( clk ), .rnd ({Fresh[1699], Fresh[1698], Fresh[1697], Fresh[1696], Fresh[1695], Fresh[1694], Fresh[1693], Fresh[1692], Fresh[1691], Fresh[1690]}), .outt ({new_AGEMA_signal_1811, new_AGEMA_signal_1810, new_AGEMA_signal_1809, n2438}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2471 ( .ina ({new_AGEMA_signal_1154, new_AGEMA_signal_1153, new_AGEMA_signal_1152, n2298}), .inb ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, new_AGEMA_signal_999, n2315}), .clk ( clk ), .rnd ({Fresh[1709], Fresh[1708], Fresh[1707], Fresh[1706], Fresh[1705], Fresh[1704], Fresh[1703], Fresh[1702], Fresh[1701], Fresh[1700]}), .outt ({new_AGEMA_signal_1406, new_AGEMA_signal_1405, new_AGEMA_signal_1404, n2299}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2481 ( .ina ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2766}), .inb ({new_AGEMA_signal_1280, new_AGEMA_signal_1279, new_AGEMA_signal_1278, n2313}), .clk ( clk ), .rnd ({Fresh[1719], Fresh[1718], Fresh[1717], Fresh[1716], Fresh[1715], Fresh[1714], Fresh[1713], Fresh[1712], Fresh[1711], Fresh[1710]}), .outt ({new_AGEMA_signal_1814, new_AGEMA_signal_1813, new_AGEMA_signal_1812, n2371}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2484 ( .ina ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, new_AGEMA_signal_999, n2315}), .inb ({new_AGEMA_signal_998, new_AGEMA_signal_997, new_AGEMA_signal_996, n2519}), .clk ( clk ), .rnd ({Fresh[1729], Fresh[1728], Fresh[1727], Fresh[1726], Fresh[1725], Fresh[1724], Fresh[1723], Fresh[1722], Fresh[1721], Fresh[1720]}), .outt ({new_AGEMA_signal_1172, new_AGEMA_signal_1171, new_AGEMA_signal_1170, n2316}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2486 ( .ina ({new_AGEMA_signal_1127, new_AGEMA_signal_1126, new_AGEMA_signal_1125, n2624}), .inb ({new_AGEMA_signal_1049, new_AGEMA_signal_1048, new_AGEMA_signal_1047, n2317}), .clk ( clk ), .rnd ({Fresh[1739], Fresh[1738], Fresh[1737], Fresh[1736], Fresh[1735], Fresh[1734], Fresh[1733], Fresh[1732], Fresh[1731], Fresh[1730]}), .outt ({new_AGEMA_signal_1412, new_AGEMA_signal_1411, new_AGEMA_signal_1410, n2318}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2492 ( .ina ({new_AGEMA_signal_1010, new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2708}), .inb ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}), .clk ( clk ), .rnd ({Fresh[1749], Fresh[1748], Fresh[1747], Fresh[1746], Fresh[1745], Fresh[1744], Fresh[1743], Fresh[1742], Fresh[1741], Fresh[1740]}), .outt ({new_AGEMA_signal_1823, new_AGEMA_signal_1822, new_AGEMA_signal_1821, n2325}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2494 ( .ina ({new_AGEMA_signal_1010, new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2708}), .inb ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .clk ( clk ), .rnd ({Fresh[1759], Fresh[1758], Fresh[1757], Fresh[1756], Fresh[1755], Fresh[1754], Fresh[1753], Fresh[1752], Fresh[1751], Fresh[1750]}), .outt ({new_AGEMA_signal_1826, new_AGEMA_signal_1825, new_AGEMA_signal_1824, n2328}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2495 ( .ina ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2742}), .inb ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, new_AGEMA_signal_1059, n2723}), .clk ( clk ), .rnd ({Fresh[1769], Fresh[1768], Fresh[1767], Fresh[1766], Fresh[1765], Fresh[1764], Fresh[1763], Fresh[1762], Fresh[1761], Fresh[1760]}), .outt ({new_AGEMA_signal_1415, new_AGEMA_signal_1414, new_AGEMA_signal_1413, n2327}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2505 ( .ina ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, new_AGEMA_signal_1191, n2737}), .inb ({new_AGEMA_signal_1052, new_AGEMA_signal_1051, new_AGEMA_signal_1050, n2694}), .clk ( clk ), .rnd ({Fresh[1779], Fresh[1778], Fresh[1777], Fresh[1776], Fresh[1775], Fresh[1774], Fresh[1773], Fresh[1772], Fresh[1771], Fresh[1770]}), .outt ({new_AGEMA_signal_1829, new_AGEMA_signal_1828, new_AGEMA_signal_1827, n2343}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2510 ( .ina ({new_AGEMA_signal_1139, new_AGEMA_signal_1138, new_AGEMA_signal_1137, n2563}), .inb ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}), .clk ( clk ), .rnd ({Fresh[1789], Fresh[1788], Fresh[1787], Fresh[1786], Fresh[1785], Fresh[1784], Fresh[1783], Fresh[1782], Fresh[1781], Fresh[1780]}), .outt ({new_AGEMA_signal_1835, new_AGEMA_signal_1834, new_AGEMA_signal_1833, n2344}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) U2512 ( .ina ({new_AGEMA_signal_1124, new_AGEMA_signal_1123, new_AGEMA_signal_1122, n2395}), .inb ({new_AGEMA_signal_1157, new_AGEMA_signal_1156, new_AGEMA_signal_1155, n2346}), .clk ( clk ), .rnd ({Fresh[1799], Fresh[1798], Fresh[1797], Fresh[1796], Fresh[1795], Fresh[1794], Fresh[1793], Fresh[1792], Fresh[1791], Fresh[1790]}), .outt ({new_AGEMA_signal_1418, new_AGEMA_signal_1417, new_AGEMA_signal_1416, n2348}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2513 ( .ina ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2742}), .inb ({new_AGEMA_signal_1046, new_AGEMA_signal_1045, new_AGEMA_signal_1044, n2780}), .clk ( clk ), .rnd ({Fresh[1809], Fresh[1808], Fresh[1807], Fresh[1806], Fresh[1805], Fresh[1804], Fresh[1803], Fresh[1802], Fresh[1801], Fresh[1800]}), .outt ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, new_AGEMA_signal_1419, n2347}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2520 ( .ina ({new_AGEMA_signal_1052, new_AGEMA_signal_1051, new_AGEMA_signal_1050, n2694}), .inb ({new_AGEMA_signal_1079, new_AGEMA_signal_1078, new_AGEMA_signal_1077, n2753}), .clk ( clk ), .rnd ({Fresh[1819], Fresh[1818], Fresh[1817], Fresh[1816], Fresh[1815], Fresh[1814], Fresh[1813], Fresh[1812], Fresh[1811], Fresh[1810]}), .outt ({new_AGEMA_signal_1424, new_AGEMA_signal_1423, new_AGEMA_signal_1422, n2363}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2521 ( .ina ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, new_AGEMA_signal_1317, n2809}), .inb ({new_AGEMA_signal_12466, new_AGEMA_signal_12464, new_AGEMA_signal_12462, new_AGEMA_signal_12460}), .clk ( clk ), .rnd ({Fresh[1829], Fresh[1828], Fresh[1827], Fresh[1826], Fresh[1825], Fresh[1824], Fresh[1823], Fresh[1822], Fresh[1821], Fresh[1820]}), .outt ({new_AGEMA_signal_1847, new_AGEMA_signal_1846, new_AGEMA_signal_1845, n2353}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2524 ( .ina ({new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2818}), .inb ({new_AGEMA_signal_1058, new_AGEMA_signal_1057, new_AGEMA_signal_1056, n2713}), .clk ( clk ), .rnd ({Fresh[1839], Fresh[1838], Fresh[1837], Fresh[1836], Fresh[1835], Fresh[1834], Fresh[1833], Fresh[1832], Fresh[1831], Fresh[1830]}), .outt ({new_AGEMA_signal_1850, new_AGEMA_signal_1849, new_AGEMA_signal_1848, n2355}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2530 ( .ina ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, new_AGEMA_signal_1023, n2712}), .inb ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}), .clk ( clk ), .rnd ({Fresh[1849], Fresh[1848], Fresh[1847], Fresh[1846], Fresh[1845], Fresh[1844], Fresh[1843], Fresh[1842], Fresh[1841], Fresh[1840]}), .outt ({new_AGEMA_signal_1853, new_AGEMA_signal_1852, new_AGEMA_signal_1851, n2364}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2543 ( .ina ({new_AGEMA_signal_12434, new_AGEMA_signal_12432, new_AGEMA_signal_12430, new_AGEMA_signal_12428}), .inb ({new_AGEMA_signal_1142, new_AGEMA_signal_1141, new_AGEMA_signal_1140, n2401}), .clk ( clk ), .rnd ({Fresh[1859], Fresh[1858], Fresh[1857], Fresh[1856], Fresh[1855], Fresh[1854], Fresh[1853], Fresh[1852], Fresh[1851], Fresh[1850]}), .outt ({new_AGEMA_signal_1427, new_AGEMA_signal_1426, new_AGEMA_signal_1425, n2415}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2558 ( .ina ({new_AGEMA_signal_1124, new_AGEMA_signal_1123, new_AGEMA_signal_1122, n2395}), .inb ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, new_AGEMA_signal_1032, n2750}), .clk ( clk ), .rnd ({Fresh[1869], Fresh[1868], Fresh[1867], Fresh[1866], Fresh[1865], Fresh[1864], Fresh[1863], Fresh[1862], Fresh[1861], Fresh[1860]}), .outt ({new_AGEMA_signal_1430, new_AGEMA_signal_1429, new_AGEMA_signal_1428, n2700}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2563 ( .ina ({new_AGEMA_signal_12530, new_AGEMA_signal_12528, new_AGEMA_signal_12526, new_AGEMA_signal_12524}), .inb ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, new_AGEMA_signal_1080, n2400}), .clk ( clk ), .rnd ({Fresh[1879], Fresh[1878], Fresh[1877], Fresh[1876], Fresh[1875], Fresh[1874], Fresh[1873], Fresh[1872], Fresh[1871], Fresh[1870]}), .outt ({new_AGEMA_signal_1433, new_AGEMA_signal_1432, new_AGEMA_signal_1431, n2594}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2564 ( .ina ({new_AGEMA_signal_1142, new_AGEMA_signal_1141, new_AGEMA_signal_1140, n2401}), .inb ({new_AGEMA_signal_12474, new_AGEMA_signal_12472, new_AGEMA_signal_12470, new_AGEMA_signal_12468}), .clk ( clk ), .rnd ({Fresh[1889], Fresh[1888], Fresh[1887], Fresh[1886], Fresh[1885], Fresh[1884], Fresh[1883], Fresh[1882], Fresh[1881], Fresh[1880]}), .outt ({new_AGEMA_signal_1436, new_AGEMA_signal_1435, new_AGEMA_signal_1434, n2402}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2585 ( .ina ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, new_AGEMA_signal_1023, n2712}), .inb ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, new_AGEMA_signal_1305, n2823}), .clk ( clk ), .rnd ({Fresh[1899], Fresh[1898], Fresh[1897], Fresh[1896], Fresh[1895], Fresh[1894], Fresh[1893], Fresh[1892], Fresh[1891], Fresh[1890]}), .outt ({new_AGEMA_signal_1883, new_AGEMA_signal_1882, new_AGEMA_signal_1881, n2428}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2588 ( .ina ({new_AGEMA_signal_1163, new_AGEMA_signal_1162, new_AGEMA_signal_1161, n2430}), .inb ({new_AGEMA_signal_1250, new_AGEMA_signal_1249, new_AGEMA_signal_1248, n2570}), .clk ( clk ), .rnd ({Fresh[1909], Fresh[1908], Fresh[1907], Fresh[1906], Fresh[1905], Fresh[1904], Fresh[1903], Fresh[1902], Fresh[1901], Fresh[1900]}), .outt ({new_AGEMA_signal_1886, new_AGEMA_signal_1885, new_AGEMA_signal_1884, n2431}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2594 ( .ina ({new_AGEMA_signal_1106, new_AGEMA_signal_1105, new_AGEMA_signal_1104, n2437}), .inb ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, new_AGEMA_signal_1035, n2615}), .clk ( clk ), .rnd ({Fresh[1919], Fresh[1918], Fresh[1917], Fresh[1916], Fresh[1915], Fresh[1914], Fresh[1913], Fresh[1912], Fresh[1911], Fresh[1910]}), .outt ({new_AGEMA_signal_1439, new_AGEMA_signal_1438, new_AGEMA_signal_1437, n2483}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2599 ( .ina ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, n2442}), .inb ({new_AGEMA_signal_1058, new_AGEMA_signal_1057, new_AGEMA_signal_1056, n2713}), .clk ( clk ), .rnd ({Fresh[1929], Fresh[1928], Fresh[1927], Fresh[1926], Fresh[1925], Fresh[1924], Fresh[1923], Fresh[1922], Fresh[1921], Fresh[1920]}), .outt ({new_AGEMA_signal_1892, new_AGEMA_signal_1891, new_AGEMA_signal_1890, n2443}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2606 ( .ina ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2766}), .inb ({new_AGEMA_signal_1088, new_AGEMA_signal_1087, new_AGEMA_signal_1086, n2609}), .clk ( clk ), .rnd ({Fresh[1939], Fresh[1938], Fresh[1937], Fresh[1936], Fresh[1935], Fresh[1934], Fresh[1933], Fresh[1932], Fresh[1931], Fresh[1930]}), .outt ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, new_AGEMA_signal_1893, n2693}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2608 ( .ina ({new_AGEMA_signal_1112, new_AGEMA_signal_1111, new_AGEMA_signal_1110, n2452}), .inb ({new_AGEMA_signal_12538, new_AGEMA_signal_12536, new_AGEMA_signal_12534, new_AGEMA_signal_12532}), .clk ( clk ), .rnd ({Fresh[1949], Fresh[1948], Fresh[1947], Fresh[1946], Fresh[1945], Fresh[1944], Fresh[1943], Fresh[1942], Fresh[1941], Fresh[1940]}), .outt ({new_AGEMA_signal_1442, new_AGEMA_signal_1441, new_AGEMA_signal_1440, n2453}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2616 ( .ina ({new_AGEMA_signal_995, new_AGEMA_signal_994, new_AGEMA_signal_993, n2790}), .inb ({new_AGEMA_signal_1175, new_AGEMA_signal_1174, new_AGEMA_signal_1173, n2463}), .clk ( clk ), .rnd ({Fresh[1959], Fresh[1958], Fresh[1957], Fresh[1956], Fresh[1955], Fresh[1954], Fresh[1953], Fresh[1952], Fresh[1951], Fresh[1950]}), .outt ({new_AGEMA_signal_1445, new_AGEMA_signal_1444, new_AGEMA_signal_1443, n2464}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2620 ( .ina ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2725}), .inb ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2742}), .clk ( clk ), .rnd ({Fresh[1969], Fresh[1968], Fresh[1967], Fresh[1966], Fresh[1965], Fresh[1964], Fresh[1963], Fresh[1962], Fresh[1961], Fresh[1960]}), .outt ({new_AGEMA_signal_1448, new_AGEMA_signal_1447, new_AGEMA_signal_1446, n2468}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2624 ( .ina ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, new_AGEMA_signal_1107, n2778}), .inb ({new_AGEMA_signal_12466, new_AGEMA_signal_12464, new_AGEMA_signal_12462, new_AGEMA_signal_12460}), .clk ( clk ), .rnd ({Fresh[1979], Fresh[1978], Fresh[1977], Fresh[1976], Fresh[1975], Fresh[1974], Fresh[1973], Fresh[1972], Fresh[1971], Fresh[1970]}), .outt ({new_AGEMA_signal_1451, new_AGEMA_signal_1450, new_AGEMA_signal_1449, n2473}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2625 ( .ina ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, new_AGEMA_signal_1065, n2815}), .inb ({new_AGEMA_signal_1046, new_AGEMA_signal_1045, new_AGEMA_signal_1044, n2780}), .clk ( clk ), .rnd ({Fresh[1989], Fresh[1988], Fresh[1987], Fresh[1986], Fresh[1985], Fresh[1984], Fresh[1983], Fresh[1982], Fresh[1981], Fresh[1980]}), .outt ({new_AGEMA_signal_1454, new_AGEMA_signal_1453, new_AGEMA_signal_1452, n2472}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2628 ( .ina ({new_AGEMA_signal_1091, new_AGEMA_signal_1090, new_AGEMA_signal_1089, n2661}), .inb ({new_AGEMA_signal_1178, new_AGEMA_signal_1177, new_AGEMA_signal_1176, n2474}), .clk ( clk ), .rnd ({Fresh[1999], Fresh[1998], Fresh[1997], Fresh[1996], Fresh[1995], Fresh[1994], Fresh[1993], Fresh[1992], Fresh[1991], Fresh[1990]}), .outt ({new_AGEMA_signal_1457, new_AGEMA_signal_1456, new_AGEMA_signal_1455, n2475}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2632 ( .ina ({new_AGEMA_signal_12546, new_AGEMA_signal_12544, new_AGEMA_signal_12542, new_AGEMA_signal_12540}), .inb ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, new_AGEMA_signal_1311, n2828}), .clk ( clk ), .rnd ({Fresh[2009], Fresh[2008], Fresh[2007], Fresh[2006], Fresh[2005], Fresh[2004], Fresh[2003], Fresh[2002], Fresh[2001], Fresh[2000]}), .outt ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, new_AGEMA_signal_1905, n2480}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2638 ( .ina ({new_AGEMA_signal_1229, new_AGEMA_signal_1228, new_AGEMA_signal_1227, n2577}), .inb ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, new_AGEMA_signal_1035, n2615}), .clk ( clk ), .rnd ({Fresh[2019], Fresh[2018], Fresh[2017], Fresh[2016], Fresh[2015], Fresh[2014], Fresh[2013], Fresh[2012], Fresh[2011], Fresh[2010]}), .outt ({new_AGEMA_signal_1910, new_AGEMA_signal_1909, new_AGEMA_signal_1908, n2487}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2641 ( .ina ({new_AGEMA_signal_1136, new_AGEMA_signal_1135, new_AGEMA_signal_1134, n2616}), .inb ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, new_AGEMA_signal_1119, n2824}), .clk ( clk ), .rnd ({Fresh[2029], Fresh[2028], Fresh[2027], Fresh[2026], Fresh[2025], Fresh[2024], Fresh[2023], Fresh[2022], Fresh[2021], Fresh[2020]}), .outt ({new_AGEMA_signal_1460, new_AGEMA_signal_1459, new_AGEMA_signal_1458, n2488}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2665 ( .ina ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, n2786}), .inb ({new_AGEMA_signal_998, new_AGEMA_signal_997, new_AGEMA_signal_996, n2519}), .clk ( clk ), .rnd ({Fresh[2039], Fresh[2038], Fresh[2037], Fresh[2036], Fresh[2035], Fresh[2034], Fresh[2033], Fresh[2032], Fresh[2031], Fresh[2030]}), .outt ({new_AGEMA_signal_1928, new_AGEMA_signal_1927, new_AGEMA_signal_1926, n2520}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2667 ( .ina ({new_AGEMA_signal_1058, new_AGEMA_signal_1057, new_AGEMA_signal_1056, n2713}), .inb ({new_AGEMA_signal_1097, new_AGEMA_signal_1096, new_AGEMA_signal_1095, n2587}), .clk ( clk ), .rnd ({Fresh[2049], Fresh[2048], Fresh[2047], Fresh[2046], Fresh[2045], Fresh[2044], Fresh[2043], Fresh[2042], Fresh[2041], Fresh[2040]}), .outt ({new_AGEMA_signal_1463, new_AGEMA_signal_1462, new_AGEMA_signal_1461, n2521}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2674 ( .ina ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, new_AGEMA_signal_1191, n2737}), .inb ({new_AGEMA_signal_1007, new_AGEMA_signal_1006, new_AGEMA_signal_1005, n2595}), .clk ( clk ), .rnd ({Fresh[2059], Fresh[2058], Fresh[2057], Fresh[2056], Fresh[2055], Fresh[2054], Fresh[2053], Fresh[2052], Fresh[2051], Fresh[2050]}), .outt ({new_AGEMA_signal_1931, new_AGEMA_signal_1930, new_AGEMA_signal_1929, n2531}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2689 ( .ina ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, new_AGEMA_signal_1119, n2824}), .inb ({new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2818}), .clk ( clk ), .rnd ({Fresh[2069], Fresh[2068], Fresh[2067], Fresh[2066], Fresh[2065], Fresh[2064], Fresh[2063], Fresh[2062], Fresh[2061], Fresh[2060]}), .outt ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, new_AGEMA_signal_1935, n2553}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2691 ( .ina ({new_AGEMA_signal_1052, new_AGEMA_signal_1051, new_AGEMA_signal_1050, n2694}), .inb ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, n2792}), .clk ( clk ), .rnd ({Fresh[2079], Fresh[2078], Fresh[2077], Fresh[2076], Fresh[2075], Fresh[2074], Fresh[2073], Fresh[2072], Fresh[2071], Fresh[2070]}), .outt ({new_AGEMA_signal_1940, new_AGEMA_signal_1939, new_AGEMA_signal_1938, n2554}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) U2695 ( .ina ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, new_AGEMA_signal_1011, n2559}), .inb ({new_AGEMA_signal_1100, new_AGEMA_signal_1099, new_AGEMA_signal_1098, n2643}), .clk ( clk ), .rnd ({Fresh[2089], Fresh[2088], Fresh[2087], Fresh[2086], Fresh[2085], Fresh[2084], Fresh[2083], Fresh[2082], Fresh[2081], Fresh[2080]}), .outt ({new_AGEMA_signal_1466, new_AGEMA_signal_1465, new_AGEMA_signal_1464, n2560}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2698 ( .ina ({new_AGEMA_signal_1238, new_AGEMA_signal_1237, new_AGEMA_signal_1236, n2724}), .inb ({new_AGEMA_signal_1139, new_AGEMA_signal_1138, new_AGEMA_signal_1137, n2563}), .clk ( clk ), .rnd ({Fresh[2099], Fresh[2098], Fresh[2097], Fresh[2096], Fresh[2095], Fresh[2094], Fresh[2093], Fresh[2092], Fresh[2091], Fresh[2090]}), .outt ({new_AGEMA_signal_1943, new_AGEMA_signal_1942, new_AGEMA_signal_1941, n2564}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2714 ( .ina ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, new_AGEMA_signal_1209, n2688}), .inb ({new_AGEMA_signal_1052, new_AGEMA_signal_1051, new_AGEMA_signal_1050, n2694}), .clk ( clk ), .rnd ({Fresh[2109], Fresh[2108], Fresh[2107], Fresh[2106], Fresh[2105], Fresh[2104], Fresh[2103], Fresh[2102], Fresh[2101], Fresh[2100]}), .outt ({new_AGEMA_signal_1952, new_AGEMA_signal_1951, new_AGEMA_signal_1950, n2586}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2720 ( .ina ({new_AGEMA_signal_1007, new_AGEMA_signal_1006, new_AGEMA_signal_1005, n2595}), .inb ({new_AGEMA_signal_1100, new_AGEMA_signal_1099, new_AGEMA_signal_1098, n2643}), .clk ( clk ), .rnd ({Fresh[2119], Fresh[2118], Fresh[2117], Fresh[2116], Fresh[2115], Fresh[2114], Fresh[2113], Fresh[2112], Fresh[2111], Fresh[2110]}), .outt ({new_AGEMA_signal_1469, new_AGEMA_signal_1468, new_AGEMA_signal_1467, n2597}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2721 ( .ina ({new_AGEMA_signal_1190, new_AGEMA_signal_1189, new_AGEMA_signal_1188, n2640}), .inb ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, new_AGEMA_signal_1197, n2789}), .clk ( clk ), .rnd ({Fresh[2129], Fresh[2128], Fresh[2127], Fresh[2126], Fresh[2125], Fresh[2124], Fresh[2123], Fresh[2122], Fresh[2121], Fresh[2120]}), .outt ({new_AGEMA_signal_1958, new_AGEMA_signal_1957, new_AGEMA_signal_1956, n2596}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2723 ( .ina ({new_AGEMA_signal_1238, new_AGEMA_signal_1237, new_AGEMA_signal_1236, n2724}), .inb ({new_AGEMA_signal_1046, new_AGEMA_signal_1045, new_AGEMA_signal_1044, n2780}), .clk ( clk ), .rnd ({Fresh[2139], Fresh[2138], Fresh[2137], Fresh[2136], Fresh[2135], Fresh[2134], Fresh[2133], Fresh[2132], Fresh[2131], Fresh[2130]}), .outt ({new_AGEMA_signal_1961, new_AGEMA_signal_1960, new_AGEMA_signal_1959, n2598}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2725 ( .ina ({new_AGEMA_signal_992, new_AGEMA_signal_991, new_AGEMA_signal_990, n2635}), .inb ({new_AGEMA_signal_12458, new_AGEMA_signal_12456, new_AGEMA_signal_12454, new_AGEMA_signal_12452}), .clk ( clk ), .rnd ({Fresh[2149], Fresh[2148], Fresh[2147], Fresh[2146], Fresh[2145], Fresh[2144], Fresh[2143], Fresh[2142], Fresh[2141], Fresh[2140]}), .outt ({new_AGEMA_signal_1181, new_AGEMA_signal_1180, new_AGEMA_signal_1179, n2599}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2732 ( .ina ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .inb ({new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2818}), .clk ( clk ), .rnd ({Fresh[2159], Fresh[2158], Fresh[2157], Fresh[2156], Fresh[2155], Fresh[2154], Fresh[2153], Fresh[2152], Fresh[2151], Fresh[2150]}), .outt ({new_AGEMA_signal_1967, new_AGEMA_signal_1966, new_AGEMA_signal_1965, n2610}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2734 ( .ina ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2767}), .inb ({new_AGEMA_signal_1133, new_AGEMA_signal_1132, new_AGEMA_signal_1131, n2611}), .clk ( clk ), .rnd ({Fresh[2169], Fresh[2168], Fresh[2167], Fresh[2166], Fresh[2165], Fresh[2164], Fresh[2163], Fresh[2162], Fresh[2161], Fresh[2160]}), .outt ({new_AGEMA_signal_1970, new_AGEMA_signal_1969, new_AGEMA_signal_1968, n2614}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2735 ( .ina ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, n2612}), .inb ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, new_AGEMA_signal_1197, n2789}), .clk ( clk ), .rnd ({Fresh[2179], Fresh[2178], Fresh[2177], Fresh[2176], Fresh[2175], Fresh[2174], Fresh[2173], Fresh[2172], Fresh[2171], Fresh[2170]}), .outt ({new_AGEMA_signal_1973, new_AGEMA_signal_1972, new_AGEMA_signal_1971, n2613}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2737 ( .ina ({new_AGEMA_signal_1136, new_AGEMA_signal_1135, new_AGEMA_signal_1134, n2616}), .inb ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, new_AGEMA_signal_1035, n2615}), .clk ( clk ), .rnd ({Fresh[2189], Fresh[2188], Fresh[2187], Fresh[2186], Fresh[2185], Fresh[2184], Fresh[2183], Fresh[2182], Fresh[2181], Fresh[2180]}), .outt ({new_AGEMA_signal_1475, new_AGEMA_signal_1474, new_AGEMA_signal_1473, n2617}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2742 ( .ina ({new_AGEMA_signal_1127, new_AGEMA_signal_1126, new_AGEMA_signal_1125, n2624}), .inb ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, new_AGEMA_signal_1032, n2750}), .clk ( clk ), .rnd ({Fresh[2199], Fresh[2198], Fresh[2197], Fresh[2196], Fresh[2195], Fresh[2194], Fresh[2193], Fresh[2192], Fresh[2191], Fresh[2190]}), .outt ({new_AGEMA_signal_1478, new_AGEMA_signal_1477, new_AGEMA_signal_1476, n2629}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2751 ( .ina ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, new_AGEMA_signal_1029, n2641}), .inb ({new_AGEMA_signal_1190, new_AGEMA_signal_1189, new_AGEMA_signal_1188, n2640}), .clk ( clk ), .rnd ({Fresh[2209], Fresh[2208], Fresh[2207], Fresh[2206], Fresh[2205], Fresh[2204], Fresh[2203], Fresh[2202], Fresh[2201], Fresh[2200]}), .outt ({new_AGEMA_signal_1979, new_AGEMA_signal_1978, new_AGEMA_signal_1977, n2784}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2757 ( .ina ({new_AGEMA_signal_1085, new_AGEMA_signal_1084, new_AGEMA_signal_1083, n2785}), .inb ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, new_AGEMA_signal_1167, n2777}), .clk ( clk ), .rnd ({Fresh[2219], Fresh[2218], Fresh[2217], Fresh[2216], Fresh[2215], Fresh[2214], Fresh[2213], Fresh[2212], Fresh[2211], Fresh[2210]}), .outt ({new_AGEMA_signal_1481, new_AGEMA_signal_1480, new_AGEMA_signal_1479, n2650}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2775 ( .ina ({new_AGEMA_signal_12498, new_AGEMA_signal_12496, new_AGEMA_signal_12494, new_AGEMA_signal_12492}), .inb ({new_AGEMA_signal_1004, new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2682}), .clk ( clk ), .rnd ({Fresh[2229], Fresh[2228], Fresh[2227], Fresh[2226], Fresh[2225], Fresh[2224], Fresh[2223], Fresh[2222], Fresh[2221], Fresh[2220]}), .outt ({new_AGEMA_signal_1184, new_AGEMA_signal_1183, new_AGEMA_signal_1182, n2683}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2789 ( .ina ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, new_AGEMA_signal_1059, n2723}), .inb ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .clk ( clk ), .rnd ({Fresh[2239], Fresh[2238], Fresh[2237], Fresh[2236], Fresh[2235], Fresh[2234], Fresh[2233], Fresh[2232], Fresh[2231], Fresh[2230]}), .outt ({new_AGEMA_signal_2000, new_AGEMA_signal_1999, new_AGEMA_signal_1998, n2711}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2790 ( .ina ({new_AGEMA_signal_1322, new_AGEMA_signal_1321, new_AGEMA_signal_1320, n2709}), .inb ({new_AGEMA_signal_1010, new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2708}), .clk ( clk ), .rnd ({Fresh[2249], Fresh[2248], Fresh[2247], Fresh[2246], Fresh[2245], Fresh[2244], Fresh[2243], Fresh[2242], Fresh[2241], Fresh[2240]}), .outt ({new_AGEMA_signal_2003, new_AGEMA_signal_2002, new_AGEMA_signal_2001, n2710}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2792 ( .ina ({new_AGEMA_signal_1058, new_AGEMA_signal_1057, new_AGEMA_signal_1056, n2713}), .inb ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, new_AGEMA_signal_1023, n2712}), .clk ( clk ), .rnd ({Fresh[2259], Fresh[2258], Fresh[2257], Fresh[2256], Fresh[2255], Fresh[2254], Fresh[2253], Fresh[2252], Fresh[2251], Fresh[2250]}), .outt ({new_AGEMA_signal_1484, new_AGEMA_signal_1483, new_AGEMA_signal_1482, n2714}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2797 ( .ina ({new_AGEMA_signal_995, new_AGEMA_signal_994, new_AGEMA_signal_993, n2790}), .inb ({new_AGEMA_signal_1151, new_AGEMA_signal_1150, new_AGEMA_signal_1149, n2721}), .clk ( clk ), .rnd ({Fresh[2269], Fresh[2268], Fresh[2267], Fresh[2266], Fresh[2265], Fresh[2264], Fresh[2263], Fresh[2262], Fresh[2261], Fresh[2260]}), .outt ({new_AGEMA_signal_1487, new_AGEMA_signal_1486, new_AGEMA_signal_1485, n2722}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2799 ( .ina ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2725}), .inb ({new_AGEMA_signal_1238, new_AGEMA_signal_1237, new_AGEMA_signal_1236, n2724}), .clk ( clk ), .rnd ({Fresh[2279], Fresh[2278], Fresh[2277], Fresh[2276], Fresh[2275], Fresh[2274], Fresh[2273], Fresh[2272], Fresh[2271], Fresh[2270]}), .outt ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, new_AGEMA_signal_2007, n2726}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2806 ( .ina ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, new_AGEMA_signal_1191, n2737}), .inb ({new_AGEMA_signal_1079, new_AGEMA_signal_1078, new_AGEMA_signal_1077, n2753}), .clk ( clk ), .rnd ({Fresh[2289], Fresh[2288], Fresh[2287], Fresh[2286], Fresh[2285], Fresh[2284], Fresh[2283], Fresh[2282], Fresh[2281], Fresh[2280]}), .outt ({new_AGEMA_signal_2012, new_AGEMA_signal_2011, new_AGEMA_signal_2010, n2738}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2822 ( .ina ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2767}), .inb ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2766}), .clk ( clk ), .rnd ({Fresh[2299], Fresh[2298], Fresh[2297], Fresh[2296], Fresh[2295], Fresh[2294], Fresh[2293], Fresh[2292], Fresh[2291], Fresh[2290]}), .outt ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, new_AGEMA_signal_2019, n2768}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2828 ( .ina ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, new_AGEMA_signal_1107, n2778}), .inb ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, new_AGEMA_signal_1167, n2777}), .clk ( clk ), .rnd ({Fresh[2309], Fresh[2308], Fresh[2307], Fresh[2306], Fresh[2305], Fresh[2304], Fresh[2303], Fresh[2302], Fresh[2301], Fresh[2300]}), .outt ({new_AGEMA_signal_1490, new_AGEMA_signal_1489, new_AGEMA_signal_1488, n2782}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2829 ( .ina ({new_AGEMA_signal_1046, new_AGEMA_signal_1045, new_AGEMA_signal_1044, n2780}), .inb ({new_AGEMA_signal_1019, new_AGEMA_signal_1018, new_AGEMA_signal_1017, n2779}), .clk ( clk ), .rnd ({Fresh[2319], Fresh[2318], Fresh[2317], Fresh[2316], Fresh[2315], Fresh[2314], Fresh[2313], Fresh[2312], Fresh[2311], Fresh[2310]}), .outt ({new_AGEMA_signal_1493, new_AGEMA_signal_1492, new_AGEMA_signal_1491, n2781}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2832 ( .ina ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, n2786}), .inb ({new_AGEMA_signal_1085, new_AGEMA_signal_1084, new_AGEMA_signal_1083, n2785}), .clk ( clk ), .rnd ({Fresh[2329], Fresh[2328], Fresh[2327], Fresh[2326], Fresh[2325], Fresh[2324], Fresh[2323], Fresh[2322], Fresh[2321], Fresh[2320]}), .outt ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, new_AGEMA_signal_2025, n2787}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2834 ( .ina ({new_AGEMA_signal_995, new_AGEMA_signal_994, new_AGEMA_signal_993, n2790}), .inb ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, new_AGEMA_signal_1197, n2789}), .clk ( clk ), .rnd ({Fresh[2339], Fresh[2338], Fresh[2337], Fresh[2336], Fresh[2335], Fresh[2334], Fresh[2333], Fresh[2332], Fresh[2331], Fresh[2330]}), .outt ({new_AGEMA_signal_2030, new_AGEMA_signal_2029, new_AGEMA_signal_2028, n2794}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2835 ( .ina ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, n2792}), .inb ({new_AGEMA_signal_12522, new_AGEMA_signal_12520, new_AGEMA_signal_12518, new_AGEMA_signal_12516}), .clk ( clk ), .rnd ({Fresh[2349], Fresh[2348], Fresh[2347], Fresh[2346], Fresh[2345], Fresh[2344], Fresh[2343], Fresh[2342], Fresh[2341], Fresh[2340]}), .outt ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, new_AGEMA_signal_2031, n2793}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2844 ( .ina ({new_AGEMA_signal_12546, new_AGEMA_signal_12544, new_AGEMA_signal_12542, new_AGEMA_signal_12540}), .inb ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, new_AGEMA_signal_1317, n2809}), .clk ( clk ), .rnd ({Fresh[2359], Fresh[2358], Fresh[2357], Fresh[2356], Fresh[2355], Fresh[2354], Fresh[2353], Fresh[2352], Fresh[2351], Fresh[2350]}), .outt ({new_AGEMA_signal_2036, new_AGEMA_signal_2035, new_AGEMA_signal_2034, n2812}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2847 ( .ina ({new_AGEMA_signal_1043, new_AGEMA_signal_1042, new_AGEMA_signal_1041, n2816}), .inb ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, new_AGEMA_signal_1065, n2815}), .clk ( clk ), .rnd ({Fresh[2369], Fresh[2368], Fresh[2367], Fresh[2366], Fresh[2365], Fresh[2364], Fresh[2363], Fresh[2362], Fresh[2361], Fresh[2360]}), .outt ({new_AGEMA_signal_1496, new_AGEMA_signal_1495, new_AGEMA_signal_1494, n2820}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2851 ( .ina ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, new_AGEMA_signal_1119, n2824}), .inb ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, new_AGEMA_signal_1305, n2823}), .clk ( clk ), .rnd ({Fresh[2379], Fresh[2378], Fresh[2377], Fresh[2376], Fresh[2375], Fresh[2374], Fresh[2373], Fresh[2372], Fresh[2371], Fresh[2370]}), .outt ({new_AGEMA_signal_2042, new_AGEMA_signal_2041, new_AGEMA_signal_2040, n2825}) ) ;
    buf_clk new_AGEMA_reg_buffer_1048 ( .C ( clk ), .D ( new_AGEMA_signal_12547 ), .Q ( new_AGEMA_signal_12548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1050 ( .C ( clk ), .D ( new_AGEMA_signal_12549 ), .Q ( new_AGEMA_signal_12550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1052 ( .C ( clk ), .D ( new_AGEMA_signal_12551 ), .Q ( new_AGEMA_signal_12552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1054 ( .C ( clk ), .D ( new_AGEMA_signal_12553 ), .Q ( new_AGEMA_signal_12554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1056 ( .C ( clk ), .D ( new_AGEMA_signal_12555 ), .Q ( new_AGEMA_signal_12556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1058 ( .C ( clk ), .D ( new_AGEMA_signal_12557 ), .Q ( new_AGEMA_signal_12558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1060 ( .C ( clk ), .D ( new_AGEMA_signal_12559 ), .Q ( new_AGEMA_signal_12560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1062 ( .C ( clk ), .D ( new_AGEMA_signal_12561 ), .Q ( new_AGEMA_signal_12562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1064 ( .C ( clk ), .D ( new_AGEMA_signal_12563 ), .Q ( new_AGEMA_signal_12564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1066 ( .C ( clk ), .D ( new_AGEMA_signal_12565 ), .Q ( new_AGEMA_signal_12566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1068 ( .C ( clk ), .D ( new_AGEMA_signal_12567 ), .Q ( new_AGEMA_signal_12568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1070 ( .C ( clk ), .D ( new_AGEMA_signal_12569 ), .Q ( new_AGEMA_signal_12570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1072 ( .C ( clk ), .D ( new_AGEMA_signal_12571 ), .Q ( new_AGEMA_signal_12572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1074 ( .C ( clk ), .D ( new_AGEMA_signal_12573 ), .Q ( new_AGEMA_signal_12574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1076 ( .C ( clk ), .D ( new_AGEMA_signal_12575 ), .Q ( new_AGEMA_signal_12576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1078 ( .C ( clk ), .D ( new_AGEMA_signal_12577 ), .Q ( new_AGEMA_signal_12578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1080 ( .C ( clk ), .D ( new_AGEMA_signal_12579 ), .Q ( new_AGEMA_signal_12580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1082 ( .C ( clk ), .D ( new_AGEMA_signal_12581 ), .Q ( new_AGEMA_signal_12582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1084 ( .C ( clk ), .D ( new_AGEMA_signal_12583 ), .Q ( new_AGEMA_signal_12584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1086 ( .C ( clk ), .D ( new_AGEMA_signal_12585 ), .Q ( new_AGEMA_signal_12586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1088 ( .C ( clk ), .D ( new_AGEMA_signal_12587 ), .Q ( new_AGEMA_signal_12588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1090 ( .C ( clk ), .D ( new_AGEMA_signal_12589 ), .Q ( new_AGEMA_signal_12590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1092 ( .C ( clk ), .D ( new_AGEMA_signal_12591 ), .Q ( new_AGEMA_signal_12592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1094 ( .C ( clk ), .D ( new_AGEMA_signal_12593 ), .Q ( new_AGEMA_signal_12594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1096 ( .C ( clk ), .D ( new_AGEMA_signal_12595 ), .Q ( new_AGEMA_signal_12596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1098 ( .C ( clk ), .D ( new_AGEMA_signal_12597 ), .Q ( new_AGEMA_signal_12598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1100 ( .C ( clk ), .D ( new_AGEMA_signal_12599 ), .Q ( new_AGEMA_signal_12600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1102 ( .C ( clk ), .D ( new_AGEMA_signal_12601 ), .Q ( new_AGEMA_signal_12602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1104 ( .C ( clk ), .D ( new_AGEMA_signal_12603 ), .Q ( new_AGEMA_signal_12604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1106 ( .C ( clk ), .D ( new_AGEMA_signal_12605 ), .Q ( new_AGEMA_signal_12606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1108 ( .C ( clk ), .D ( new_AGEMA_signal_12607 ), .Q ( new_AGEMA_signal_12608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1110 ( .C ( clk ), .D ( new_AGEMA_signal_12609 ), .Q ( new_AGEMA_signal_12610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1112 ( .C ( clk ), .D ( new_AGEMA_signal_12611 ), .Q ( new_AGEMA_signal_12612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1114 ( .C ( clk ), .D ( new_AGEMA_signal_12613 ), .Q ( new_AGEMA_signal_12614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1116 ( .C ( clk ), .D ( new_AGEMA_signal_12615 ), .Q ( new_AGEMA_signal_12616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1118 ( .C ( clk ), .D ( new_AGEMA_signal_12617 ), .Q ( new_AGEMA_signal_12618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1120 ( .C ( clk ), .D ( new_AGEMA_signal_12619 ), .Q ( new_AGEMA_signal_12620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1122 ( .C ( clk ), .D ( new_AGEMA_signal_12621 ), .Q ( new_AGEMA_signal_12622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1124 ( .C ( clk ), .D ( new_AGEMA_signal_12623 ), .Q ( new_AGEMA_signal_12624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1126 ( .C ( clk ), .D ( new_AGEMA_signal_12625 ), .Q ( new_AGEMA_signal_12626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1128 ( .C ( clk ), .D ( new_AGEMA_signal_12627 ), .Q ( new_AGEMA_signal_12628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1130 ( .C ( clk ), .D ( new_AGEMA_signal_12629 ), .Q ( new_AGEMA_signal_12630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1132 ( .C ( clk ), .D ( new_AGEMA_signal_12631 ), .Q ( new_AGEMA_signal_12632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1134 ( .C ( clk ), .D ( new_AGEMA_signal_12633 ), .Q ( new_AGEMA_signal_12634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1136 ( .C ( clk ), .D ( new_AGEMA_signal_12635 ), .Q ( new_AGEMA_signal_12636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1138 ( .C ( clk ), .D ( new_AGEMA_signal_12637 ), .Q ( new_AGEMA_signal_12638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1140 ( .C ( clk ), .D ( new_AGEMA_signal_12639 ), .Q ( new_AGEMA_signal_12640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1142 ( .C ( clk ), .D ( new_AGEMA_signal_12641 ), .Q ( new_AGEMA_signal_12642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1144 ( .C ( clk ), .D ( new_AGEMA_signal_12643 ), .Q ( new_AGEMA_signal_12644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1146 ( .C ( clk ), .D ( new_AGEMA_signal_12645 ), .Q ( new_AGEMA_signal_12646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1148 ( .C ( clk ), .D ( new_AGEMA_signal_12647 ), .Q ( new_AGEMA_signal_12648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1150 ( .C ( clk ), .D ( new_AGEMA_signal_12649 ), .Q ( new_AGEMA_signal_12650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1152 ( .C ( clk ), .D ( new_AGEMA_signal_12651 ), .Q ( new_AGEMA_signal_12652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1154 ( .C ( clk ), .D ( new_AGEMA_signal_12653 ), .Q ( new_AGEMA_signal_12654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1156 ( .C ( clk ), .D ( new_AGEMA_signal_12655 ), .Q ( new_AGEMA_signal_12656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1158 ( .C ( clk ), .D ( new_AGEMA_signal_12657 ), .Q ( new_AGEMA_signal_12658 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1160 ( .C ( clk ), .D ( new_AGEMA_signal_12659 ), .Q ( new_AGEMA_signal_12660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1162 ( .C ( clk ), .D ( new_AGEMA_signal_12661 ), .Q ( new_AGEMA_signal_12662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1164 ( .C ( clk ), .D ( new_AGEMA_signal_12663 ), .Q ( new_AGEMA_signal_12664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1166 ( .C ( clk ), .D ( new_AGEMA_signal_12665 ), .Q ( new_AGEMA_signal_12666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1168 ( .C ( clk ), .D ( new_AGEMA_signal_12667 ), .Q ( new_AGEMA_signal_12668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1170 ( .C ( clk ), .D ( new_AGEMA_signal_12669 ), .Q ( new_AGEMA_signal_12670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1172 ( .C ( clk ), .D ( new_AGEMA_signal_12671 ), .Q ( new_AGEMA_signal_12672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1174 ( .C ( clk ), .D ( new_AGEMA_signal_12673 ), .Q ( new_AGEMA_signal_12674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1176 ( .C ( clk ), .D ( new_AGEMA_signal_12675 ), .Q ( new_AGEMA_signal_12676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1178 ( .C ( clk ), .D ( new_AGEMA_signal_12677 ), .Q ( new_AGEMA_signal_12678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1180 ( .C ( clk ), .D ( new_AGEMA_signal_12679 ), .Q ( new_AGEMA_signal_12680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1182 ( .C ( clk ), .D ( new_AGEMA_signal_12681 ), .Q ( new_AGEMA_signal_12682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1184 ( .C ( clk ), .D ( new_AGEMA_signal_12683 ), .Q ( new_AGEMA_signal_12684 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1186 ( .C ( clk ), .D ( new_AGEMA_signal_12685 ), .Q ( new_AGEMA_signal_12686 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1188 ( .C ( clk ), .D ( new_AGEMA_signal_12687 ), .Q ( new_AGEMA_signal_12688 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1190 ( .C ( clk ), .D ( new_AGEMA_signal_12689 ), .Q ( new_AGEMA_signal_12690 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1192 ( .C ( clk ), .D ( new_AGEMA_signal_12691 ), .Q ( new_AGEMA_signal_12692 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1194 ( .C ( clk ), .D ( new_AGEMA_signal_12693 ), .Q ( new_AGEMA_signal_12694 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1196 ( .C ( clk ), .D ( new_AGEMA_signal_12695 ), .Q ( new_AGEMA_signal_12696 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1198 ( .C ( clk ), .D ( new_AGEMA_signal_12697 ), .Q ( new_AGEMA_signal_12698 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1200 ( .C ( clk ), .D ( new_AGEMA_signal_12699 ), .Q ( new_AGEMA_signal_12700 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1202 ( .C ( clk ), .D ( new_AGEMA_signal_12701 ), .Q ( new_AGEMA_signal_12702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1204 ( .C ( clk ), .D ( new_AGEMA_signal_12703 ), .Q ( new_AGEMA_signal_12704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1206 ( .C ( clk ), .D ( new_AGEMA_signal_12705 ), .Q ( new_AGEMA_signal_12706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1208 ( .C ( clk ), .D ( new_AGEMA_signal_12707 ), .Q ( new_AGEMA_signal_12708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1210 ( .C ( clk ), .D ( new_AGEMA_signal_12709 ), .Q ( new_AGEMA_signal_12710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1212 ( .C ( clk ), .D ( new_AGEMA_signal_12711 ), .Q ( new_AGEMA_signal_12712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1214 ( .C ( clk ), .D ( new_AGEMA_signal_12713 ), .Q ( new_AGEMA_signal_12714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1216 ( .C ( clk ), .D ( new_AGEMA_signal_12715 ), .Q ( new_AGEMA_signal_12716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1218 ( .C ( clk ), .D ( new_AGEMA_signal_12717 ), .Q ( new_AGEMA_signal_12718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1220 ( .C ( clk ), .D ( new_AGEMA_signal_12719 ), .Q ( new_AGEMA_signal_12720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1222 ( .C ( clk ), .D ( new_AGEMA_signal_12721 ), .Q ( new_AGEMA_signal_12722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1224 ( .C ( clk ), .D ( new_AGEMA_signal_12723 ), .Q ( new_AGEMA_signal_12724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1226 ( .C ( clk ), .D ( new_AGEMA_signal_12725 ), .Q ( new_AGEMA_signal_12726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1228 ( .C ( clk ), .D ( new_AGEMA_signal_12727 ), .Q ( new_AGEMA_signal_12728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1230 ( .C ( clk ), .D ( new_AGEMA_signal_12729 ), .Q ( new_AGEMA_signal_12730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1232 ( .C ( clk ), .D ( new_AGEMA_signal_12731 ), .Q ( new_AGEMA_signal_12732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1234 ( .C ( clk ), .D ( new_AGEMA_signal_12733 ), .Q ( new_AGEMA_signal_12734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1236 ( .C ( clk ), .D ( new_AGEMA_signal_12735 ), .Q ( new_AGEMA_signal_12736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1238 ( .C ( clk ), .D ( new_AGEMA_signal_12737 ), .Q ( new_AGEMA_signal_12738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1240 ( .C ( clk ), .D ( new_AGEMA_signal_12739 ), .Q ( new_AGEMA_signal_12740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1242 ( .C ( clk ), .D ( new_AGEMA_signal_12741 ), .Q ( new_AGEMA_signal_12742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1244 ( .C ( clk ), .D ( new_AGEMA_signal_12743 ), .Q ( new_AGEMA_signal_12744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1246 ( .C ( clk ), .D ( new_AGEMA_signal_12745 ), .Q ( new_AGEMA_signal_12746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1248 ( .C ( clk ), .D ( new_AGEMA_signal_12747 ), .Q ( new_AGEMA_signal_12748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1250 ( .C ( clk ), .D ( new_AGEMA_signal_12749 ), .Q ( new_AGEMA_signal_12750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1252 ( .C ( clk ), .D ( new_AGEMA_signal_12751 ), .Q ( new_AGEMA_signal_12752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1254 ( .C ( clk ), .D ( new_AGEMA_signal_12753 ), .Q ( new_AGEMA_signal_12754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1256 ( .C ( clk ), .D ( new_AGEMA_signal_12755 ), .Q ( new_AGEMA_signal_12756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1258 ( .C ( clk ), .D ( new_AGEMA_signal_12757 ), .Q ( new_AGEMA_signal_12758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1260 ( .C ( clk ), .D ( new_AGEMA_signal_12759 ), .Q ( new_AGEMA_signal_12760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1262 ( .C ( clk ), .D ( new_AGEMA_signal_12761 ), .Q ( new_AGEMA_signal_12762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1264 ( .C ( clk ), .D ( new_AGEMA_signal_12763 ), .Q ( new_AGEMA_signal_12764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1266 ( .C ( clk ), .D ( new_AGEMA_signal_12765 ), .Q ( new_AGEMA_signal_12766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1268 ( .C ( clk ), .D ( new_AGEMA_signal_12767 ), .Q ( new_AGEMA_signal_12768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1270 ( .C ( clk ), .D ( new_AGEMA_signal_12769 ), .Q ( new_AGEMA_signal_12770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1272 ( .C ( clk ), .D ( new_AGEMA_signal_12771 ), .Q ( new_AGEMA_signal_12772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1274 ( .C ( clk ), .D ( new_AGEMA_signal_12773 ), .Q ( new_AGEMA_signal_12774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1276 ( .C ( clk ), .D ( new_AGEMA_signal_12775 ), .Q ( new_AGEMA_signal_12776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1278 ( .C ( clk ), .D ( new_AGEMA_signal_12777 ), .Q ( new_AGEMA_signal_12778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1280 ( .C ( clk ), .D ( new_AGEMA_signal_12779 ), .Q ( new_AGEMA_signal_12780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1282 ( .C ( clk ), .D ( new_AGEMA_signal_12781 ), .Q ( new_AGEMA_signal_12782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1284 ( .C ( clk ), .D ( new_AGEMA_signal_12783 ), .Q ( new_AGEMA_signal_12784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1286 ( .C ( clk ), .D ( new_AGEMA_signal_12785 ), .Q ( new_AGEMA_signal_12786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1288 ( .C ( clk ), .D ( new_AGEMA_signal_12787 ), .Q ( new_AGEMA_signal_12788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1290 ( .C ( clk ), .D ( new_AGEMA_signal_12789 ), .Q ( new_AGEMA_signal_12790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1292 ( .C ( clk ), .D ( new_AGEMA_signal_12791 ), .Q ( new_AGEMA_signal_12792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1294 ( .C ( clk ), .D ( new_AGEMA_signal_12793 ), .Q ( new_AGEMA_signal_12794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1296 ( .C ( clk ), .D ( new_AGEMA_signal_12795 ), .Q ( new_AGEMA_signal_12796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1298 ( .C ( clk ), .D ( new_AGEMA_signal_12797 ), .Q ( new_AGEMA_signal_12798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1300 ( .C ( clk ), .D ( new_AGEMA_signal_12799 ), .Q ( new_AGEMA_signal_12800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1302 ( .C ( clk ), .D ( new_AGEMA_signal_12801 ), .Q ( new_AGEMA_signal_12802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1304 ( .C ( clk ), .D ( new_AGEMA_signal_12803 ), .Q ( new_AGEMA_signal_12804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1306 ( .C ( clk ), .D ( new_AGEMA_signal_12805 ), .Q ( new_AGEMA_signal_12806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1308 ( .C ( clk ), .D ( new_AGEMA_signal_12807 ), .Q ( new_AGEMA_signal_12808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1310 ( .C ( clk ), .D ( new_AGEMA_signal_12809 ), .Q ( new_AGEMA_signal_12810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1312 ( .C ( clk ), .D ( new_AGEMA_signal_12811 ), .Q ( new_AGEMA_signal_12812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1314 ( .C ( clk ), .D ( new_AGEMA_signal_12813 ), .Q ( new_AGEMA_signal_12814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1316 ( .C ( clk ), .D ( new_AGEMA_signal_12815 ), .Q ( new_AGEMA_signal_12816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1318 ( .C ( clk ), .D ( new_AGEMA_signal_12817 ), .Q ( new_AGEMA_signal_12818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1320 ( .C ( clk ), .D ( new_AGEMA_signal_12819 ), .Q ( new_AGEMA_signal_12820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1322 ( .C ( clk ), .D ( new_AGEMA_signal_12821 ), .Q ( new_AGEMA_signal_12822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1324 ( .C ( clk ), .D ( new_AGEMA_signal_12823 ), .Q ( new_AGEMA_signal_12824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1326 ( .C ( clk ), .D ( new_AGEMA_signal_12825 ), .Q ( new_AGEMA_signal_12826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1328 ( .C ( clk ), .D ( new_AGEMA_signal_12827 ), .Q ( new_AGEMA_signal_12828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1330 ( .C ( clk ), .D ( new_AGEMA_signal_12829 ), .Q ( new_AGEMA_signal_12830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1332 ( .C ( clk ), .D ( new_AGEMA_signal_12831 ), .Q ( new_AGEMA_signal_12832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1334 ( .C ( clk ), .D ( new_AGEMA_signal_12833 ), .Q ( new_AGEMA_signal_12834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1336 ( .C ( clk ), .D ( new_AGEMA_signal_12835 ), .Q ( new_AGEMA_signal_12836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1338 ( .C ( clk ), .D ( new_AGEMA_signal_12837 ), .Q ( new_AGEMA_signal_12838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1340 ( .C ( clk ), .D ( new_AGEMA_signal_12839 ), .Q ( new_AGEMA_signal_12840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1342 ( .C ( clk ), .D ( new_AGEMA_signal_12841 ), .Q ( new_AGEMA_signal_12842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1344 ( .C ( clk ), .D ( new_AGEMA_signal_12843 ), .Q ( new_AGEMA_signal_12844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1346 ( .C ( clk ), .D ( new_AGEMA_signal_12845 ), .Q ( new_AGEMA_signal_12846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1348 ( .C ( clk ), .D ( new_AGEMA_signal_12847 ), .Q ( new_AGEMA_signal_12848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1350 ( .C ( clk ), .D ( new_AGEMA_signal_12849 ), .Q ( new_AGEMA_signal_12850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1352 ( .C ( clk ), .D ( new_AGEMA_signal_12851 ), .Q ( new_AGEMA_signal_12852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1354 ( .C ( clk ), .D ( new_AGEMA_signal_12853 ), .Q ( new_AGEMA_signal_12854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1356 ( .C ( clk ), .D ( new_AGEMA_signal_12855 ), .Q ( new_AGEMA_signal_12856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1358 ( .C ( clk ), .D ( new_AGEMA_signal_12857 ), .Q ( new_AGEMA_signal_12858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1360 ( .C ( clk ), .D ( new_AGEMA_signal_12859 ), .Q ( new_AGEMA_signal_12860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1362 ( .C ( clk ), .D ( new_AGEMA_signal_12861 ), .Q ( new_AGEMA_signal_12862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1364 ( .C ( clk ), .D ( new_AGEMA_signal_12863 ), .Q ( new_AGEMA_signal_12864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1366 ( .C ( clk ), .D ( new_AGEMA_signal_12865 ), .Q ( new_AGEMA_signal_12866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1368 ( .C ( clk ), .D ( new_AGEMA_signal_12867 ), .Q ( new_AGEMA_signal_12868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1370 ( .C ( clk ), .D ( new_AGEMA_signal_12869 ), .Q ( new_AGEMA_signal_12870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1372 ( .C ( clk ), .D ( new_AGEMA_signal_12871 ), .Q ( new_AGEMA_signal_12872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1374 ( .C ( clk ), .D ( new_AGEMA_signal_12873 ), .Q ( new_AGEMA_signal_12874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1376 ( .C ( clk ), .D ( new_AGEMA_signal_12875 ), .Q ( new_AGEMA_signal_12876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1378 ( .C ( clk ), .D ( new_AGEMA_signal_12877 ), .Q ( new_AGEMA_signal_12878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1380 ( .C ( clk ), .D ( new_AGEMA_signal_12879 ), .Q ( new_AGEMA_signal_12880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1382 ( .C ( clk ), .D ( new_AGEMA_signal_12881 ), .Q ( new_AGEMA_signal_12882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1384 ( .C ( clk ), .D ( new_AGEMA_signal_12883 ), .Q ( new_AGEMA_signal_12884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1386 ( .C ( clk ), .D ( new_AGEMA_signal_12885 ), .Q ( new_AGEMA_signal_12886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1388 ( .C ( clk ), .D ( new_AGEMA_signal_12887 ), .Q ( new_AGEMA_signal_12888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1390 ( .C ( clk ), .D ( new_AGEMA_signal_12889 ), .Q ( new_AGEMA_signal_12890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1392 ( .C ( clk ), .D ( new_AGEMA_signal_12891 ), .Q ( new_AGEMA_signal_12892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1394 ( .C ( clk ), .D ( new_AGEMA_signal_12893 ), .Q ( new_AGEMA_signal_12894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1396 ( .C ( clk ), .D ( new_AGEMA_signal_12895 ), .Q ( new_AGEMA_signal_12896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1398 ( .C ( clk ), .D ( new_AGEMA_signal_12897 ), .Q ( new_AGEMA_signal_12898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1400 ( .C ( clk ), .D ( new_AGEMA_signal_12899 ), .Q ( new_AGEMA_signal_12900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1402 ( .C ( clk ), .D ( new_AGEMA_signal_12901 ), .Q ( new_AGEMA_signal_12902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1404 ( .C ( clk ), .D ( new_AGEMA_signal_12903 ), .Q ( new_AGEMA_signal_12904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1406 ( .C ( clk ), .D ( new_AGEMA_signal_12905 ), .Q ( new_AGEMA_signal_12906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1408 ( .C ( clk ), .D ( new_AGEMA_signal_12907 ), .Q ( new_AGEMA_signal_12908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1410 ( .C ( clk ), .D ( new_AGEMA_signal_12909 ), .Q ( new_AGEMA_signal_12910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1412 ( .C ( clk ), .D ( new_AGEMA_signal_12911 ), .Q ( new_AGEMA_signal_12912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1414 ( .C ( clk ), .D ( new_AGEMA_signal_12913 ), .Q ( new_AGEMA_signal_12914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1416 ( .C ( clk ), .D ( new_AGEMA_signal_12915 ), .Q ( new_AGEMA_signal_12916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1418 ( .C ( clk ), .D ( new_AGEMA_signal_12917 ), .Q ( new_AGEMA_signal_12918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1420 ( .C ( clk ), .D ( new_AGEMA_signal_12919 ), .Q ( new_AGEMA_signal_12920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1422 ( .C ( clk ), .D ( new_AGEMA_signal_12921 ), .Q ( new_AGEMA_signal_12922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1424 ( .C ( clk ), .D ( new_AGEMA_signal_12923 ), .Q ( new_AGEMA_signal_12924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1426 ( .C ( clk ), .D ( new_AGEMA_signal_12925 ), .Q ( new_AGEMA_signal_12926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1428 ( .C ( clk ), .D ( new_AGEMA_signal_12927 ), .Q ( new_AGEMA_signal_12928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1430 ( .C ( clk ), .D ( new_AGEMA_signal_12929 ), .Q ( new_AGEMA_signal_12930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1432 ( .C ( clk ), .D ( new_AGEMA_signal_12931 ), .Q ( new_AGEMA_signal_12932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1434 ( .C ( clk ), .D ( new_AGEMA_signal_12933 ), .Q ( new_AGEMA_signal_12934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1436 ( .C ( clk ), .D ( new_AGEMA_signal_12935 ), .Q ( new_AGEMA_signal_12936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1438 ( .C ( clk ), .D ( new_AGEMA_signal_12937 ), .Q ( new_AGEMA_signal_12938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1440 ( .C ( clk ), .D ( new_AGEMA_signal_12939 ), .Q ( new_AGEMA_signal_12940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1442 ( .C ( clk ), .D ( new_AGEMA_signal_12941 ), .Q ( new_AGEMA_signal_12942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1444 ( .C ( clk ), .D ( new_AGEMA_signal_12943 ), .Q ( new_AGEMA_signal_12944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1446 ( .C ( clk ), .D ( new_AGEMA_signal_12945 ), .Q ( new_AGEMA_signal_12946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1448 ( .C ( clk ), .D ( new_AGEMA_signal_12947 ), .Q ( new_AGEMA_signal_12948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1450 ( .C ( clk ), .D ( new_AGEMA_signal_12949 ), .Q ( new_AGEMA_signal_12950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1452 ( .C ( clk ), .D ( new_AGEMA_signal_12951 ), .Q ( new_AGEMA_signal_12952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1454 ( .C ( clk ), .D ( new_AGEMA_signal_12953 ), .Q ( new_AGEMA_signal_12954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1456 ( .C ( clk ), .D ( new_AGEMA_signal_12955 ), .Q ( new_AGEMA_signal_12956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1458 ( .C ( clk ), .D ( new_AGEMA_signal_12957 ), .Q ( new_AGEMA_signal_12958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1460 ( .C ( clk ), .D ( new_AGEMA_signal_12959 ), .Q ( new_AGEMA_signal_12960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1462 ( .C ( clk ), .D ( new_AGEMA_signal_12961 ), .Q ( new_AGEMA_signal_12962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1464 ( .C ( clk ), .D ( new_AGEMA_signal_12963 ), .Q ( new_AGEMA_signal_12964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1466 ( .C ( clk ), .D ( new_AGEMA_signal_12965 ), .Q ( new_AGEMA_signal_12966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1468 ( .C ( clk ), .D ( new_AGEMA_signal_12967 ), .Q ( new_AGEMA_signal_12968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1470 ( .C ( clk ), .D ( new_AGEMA_signal_12969 ), .Q ( new_AGEMA_signal_12970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1472 ( .C ( clk ), .D ( new_AGEMA_signal_12971 ), .Q ( new_AGEMA_signal_12972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1474 ( .C ( clk ), .D ( new_AGEMA_signal_12973 ), .Q ( new_AGEMA_signal_12974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1476 ( .C ( clk ), .D ( new_AGEMA_signal_12975 ), .Q ( new_AGEMA_signal_12976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1478 ( .C ( clk ), .D ( new_AGEMA_signal_12977 ), .Q ( new_AGEMA_signal_12978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1480 ( .C ( clk ), .D ( new_AGEMA_signal_12979 ), .Q ( new_AGEMA_signal_12980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1482 ( .C ( clk ), .D ( new_AGEMA_signal_12981 ), .Q ( new_AGEMA_signal_12982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1484 ( .C ( clk ), .D ( new_AGEMA_signal_12983 ), .Q ( new_AGEMA_signal_12984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1486 ( .C ( clk ), .D ( new_AGEMA_signal_12985 ), .Q ( new_AGEMA_signal_12986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1488 ( .C ( clk ), .D ( new_AGEMA_signal_12987 ), .Q ( new_AGEMA_signal_12988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1490 ( .C ( clk ), .D ( new_AGEMA_signal_12989 ), .Q ( new_AGEMA_signal_12990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1492 ( .C ( clk ), .D ( new_AGEMA_signal_12991 ), .Q ( new_AGEMA_signal_12992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1494 ( .C ( clk ), .D ( new_AGEMA_signal_12993 ), .Q ( new_AGEMA_signal_12994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1496 ( .C ( clk ), .D ( new_AGEMA_signal_12995 ), .Q ( new_AGEMA_signal_12996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1498 ( .C ( clk ), .D ( new_AGEMA_signal_12997 ), .Q ( new_AGEMA_signal_12998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1500 ( .C ( clk ), .D ( new_AGEMA_signal_12999 ), .Q ( new_AGEMA_signal_13000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1502 ( .C ( clk ), .D ( new_AGEMA_signal_13001 ), .Q ( new_AGEMA_signal_13002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1504 ( .C ( clk ), .D ( new_AGEMA_signal_13003 ), .Q ( new_AGEMA_signal_13004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1506 ( .C ( clk ), .D ( new_AGEMA_signal_13005 ), .Q ( new_AGEMA_signal_13006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1508 ( .C ( clk ), .D ( new_AGEMA_signal_13007 ), .Q ( new_AGEMA_signal_13008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1510 ( .C ( clk ), .D ( new_AGEMA_signal_13009 ), .Q ( new_AGEMA_signal_13010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1512 ( .C ( clk ), .D ( new_AGEMA_signal_13011 ), .Q ( new_AGEMA_signal_13012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1514 ( .C ( clk ), .D ( new_AGEMA_signal_13013 ), .Q ( new_AGEMA_signal_13014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1516 ( .C ( clk ), .D ( new_AGEMA_signal_13015 ), .Q ( new_AGEMA_signal_13016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1518 ( .C ( clk ), .D ( new_AGEMA_signal_13017 ), .Q ( new_AGEMA_signal_13018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1520 ( .C ( clk ), .D ( new_AGEMA_signal_13019 ), .Q ( new_AGEMA_signal_13020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1522 ( .C ( clk ), .D ( new_AGEMA_signal_13021 ), .Q ( new_AGEMA_signal_13022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1524 ( .C ( clk ), .D ( new_AGEMA_signal_13023 ), .Q ( new_AGEMA_signal_13024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1526 ( .C ( clk ), .D ( new_AGEMA_signal_13025 ), .Q ( new_AGEMA_signal_13026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1528 ( .C ( clk ), .D ( new_AGEMA_signal_13027 ), .Q ( new_AGEMA_signal_13028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1530 ( .C ( clk ), .D ( new_AGEMA_signal_13029 ), .Q ( new_AGEMA_signal_13030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1532 ( .C ( clk ), .D ( new_AGEMA_signal_13031 ), .Q ( new_AGEMA_signal_13032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1534 ( .C ( clk ), .D ( new_AGEMA_signal_13033 ), .Q ( new_AGEMA_signal_13034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1536 ( .C ( clk ), .D ( new_AGEMA_signal_13035 ), .Q ( new_AGEMA_signal_13036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1538 ( .C ( clk ), .D ( new_AGEMA_signal_13037 ), .Q ( new_AGEMA_signal_13038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1540 ( .C ( clk ), .D ( new_AGEMA_signal_13039 ), .Q ( new_AGEMA_signal_13040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1542 ( .C ( clk ), .D ( new_AGEMA_signal_13041 ), .Q ( new_AGEMA_signal_13042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1544 ( .C ( clk ), .D ( new_AGEMA_signal_13043 ), .Q ( new_AGEMA_signal_13044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1546 ( .C ( clk ), .D ( new_AGEMA_signal_13045 ), .Q ( new_AGEMA_signal_13046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1548 ( .C ( clk ), .D ( new_AGEMA_signal_13047 ), .Q ( new_AGEMA_signal_13048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1550 ( .C ( clk ), .D ( new_AGEMA_signal_13049 ), .Q ( new_AGEMA_signal_13050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1552 ( .C ( clk ), .D ( new_AGEMA_signal_13051 ), .Q ( new_AGEMA_signal_13052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1554 ( .C ( clk ), .D ( new_AGEMA_signal_13053 ), .Q ( new_AGEMA_signal_13054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1556 ( .C ( clk ), .D ( new_AGEMA_signal_13055 ), .Q ( new_AGEMA_signal_13056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1558 ( .C ( clk ), .D ( new_AGEMA_signal_13057 ), .Q ( new_AGEMA_signal_13058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1560 ( .C ( clk ), .D ( new_AGEMA_signal_13059 ), .Q ( new_AGEMA_signal_13060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1562 ( .C ( clk ), .D ( new_AGEMA_signal_13061 ), .Q ( new_AGEMA_signal_13062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1564 ( .C ( clk ), .D ( new_AGEMA_signal_13063 ), .Q ( new_AGEMA_signal_13064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1566 ( .C ( clk ), .D ( new_AGEMA_signal_13065 ), .Q ( new_AGEMA_signal_13066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1568 ( .C ( clk ), .D ( new_AGEMA_signal_13067 ), .Q ( new_AGEMA_signal_13068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1570 ( .C ( clk ), .D ( new_AGEMA_signal_13069 ), .Q ( new_AGEMA_signal_13070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1572 ( .C ( clk ), .D ( new_AGEMA_signal_13071 ), .Q ( new_AGEMA_signal_13072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1574 ( .C ( clk ), .D ( new_AGEMA_signal_13073 ), .Q ( new_AGEMA_signal_13074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1576 ( .C ( clk ), .D ( new_AGEMA_signal_13075 ), .Q ( new_AGEMA_signal_13076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1578 ( .C ( clk ), .D ( new_AGEMA_signal_13077 ), .Q ( new_AGEMA_signal_13078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1580 ( .C ( clk ), .D ( new_AGEMA_signal_13079 ), .Q ( new_AGEMA_signal_13080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1582 ( .C ( clk ), .D ( new_AGEMA_signal_13081 ), .Q ( new_AGEMA_signal_13082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1584 ( .C ( clk ), .D ( new_AGEMA_signal_13083 ), .Q ( new_AGEMA_signal_13084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1586 ( .C ( clk ), .D ( new_AGEMA_signal_13085 ), .Q ( new_AGEMA_signal_13086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1588 ( .C ( clk ), .D ( new_AGEMA_signal_13087 ), .Q ( new_AGEMA_signal_13088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1590 ( .C ( clk ), .D ( new_AGEMA_signal_13089 ), .Q ( new_AGEMA_signal_13090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1608 ( .C ( clk ), .D ( new_AGEMA_signal_13107 ), .Q ( new_AGEMA_signal_13108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1612 ( .C ( clk ), .D ( new_AGEMA_signal_13111 ), .Q ( new_AGEMA_signal_13112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1616 ( .C ( clk ), .D ( new_AGEMA_signal_13115 ), .Q ( new_AGEMA_signal_13116 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1620 ( .C ( clk ), .D ( new_AGEMA_signal_13119 ), .Q ( new_AGEMA_signal_13120 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1712 ( .C ( clk ), .D ( new_AGEMA_signal_13211 ), .Q ( new_AGEMA_signal_13212 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1716 ( .C ( clk ), .D ( new_AGEMA_signal_13215 ), .Q ( new_AGEMA_signal_13216 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1720 ( .C ( clk ), .D ( new_AGEMA_signal_13219 ), .Q ( new_AGEMA_signal_13220 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1724 ( .C ( clk ), .D ( new_AGEMA_signal_13223 ), .Q ( new_AGEMA_signal_13224 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1784 ( .C ( clk ), .D ( new_AGEMA_signal_13283 ), .Q ( new_AGEMA_signal_13284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1788 ( .C ( clk ), .D ( new_AGEMA_signal_13287 ), .Q ( new_AGEMA_signal_13288 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1792 ( .C ( clk ), .D ( new_AGEMA_signal_13291 ), .Q ( new_AGEMA_signal_13292 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1796 ( .C ( clk ), .D ( new_AGEMA_signal_13295 ), .Q ( new_AGEMA_signal_13296 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1840 ( .C ( clk ), .D ( new_AGEMA_signal_13339 ), .Q ( new_AGEMA_signal_13340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1844 ( .C ( clk ), .D ( new_AGEMA_signal_13343 ), .Q ( new_AGEMA_signal_13344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1848 ( .C ( clk ), .D ( new_AGEMA_signal_13347 ), .Q ( new_AGEMA_signal_13348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1852 ( .C ( clk ), .D ( new_AGEMA_signal_13351 ), .Q ( new_AGEMA_signal_13352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1880 ( .C ( clk ), .D ( new_AGEMA_signal_13379 ), .Q ( new_AGEMA_signal_13380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1884 ( .C ( clk ), .D ( new_AGEMA_signal_13383 ), .Q ( new_AGEMA_signal_13384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1888 ( .C ( clk ), .D ( new_AGEMA_signal_13387 ), .Q ( new_AGEMA_signal_13388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1892 ( .C ( clk ), .D ( new_AGEMA_signal_13391 ), .Q ( new_AGEMA_signal_13392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1920 ( .C ( clk ), .D ( new_AGEMA_signal_13419 ), .Q ( new_AGEMA_signal_13420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1924 ( .C ( clk ), .D ( new_AGEMA_signal_13423 ), .Q ( new_AGEMA_signal_13424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1928 ( .C ( clk ), .D ( new_AGEMA_signal_13427 ), .Q ( new_AGEMA_signal_13428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1932 ( .C ( clk ), .D ( new_AGEMA_signal_13431 ), .Q ( new_AGEMA_signal_13432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2074 ( .C ( clk ), .D ( new_AGEMA_signal_13573 ), .Q ( new_AGEMA_signal_13574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2080 ( .C ( clk ), .D ( new_AGEMA_signal_13579 ), .Q ( new_AGEMA_signal_13580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2086 ( .C ( clk ), .D ( new_AGEMA_signal_13585 ), .Q ( new_AGEMA_signal_13586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2092 ( .C ( clk ), .D ( new_AGEMA_signal_13591 ), .Q ( new_AGEMA_signal_13592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2120 ( .C ( clk ), .D ( new_AGEMA_signal_13619 ), .Q ( new_AGEMA_signal_13620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2124 ( .C ( clk ), .D ( new_AGEMA_signal_13623 ), .Q ( new_AGEMA_signal_13624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2128 ( .C ( clk ), .D ( new_AGEMA_signal_13627 ), .Q ( new_AGEMA_signal_13628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2132 ( .C ( clk ), .D ( new_AGEMA_signal_13631 ), .Q ( new_AGEMA_signal_13632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2160 ( .C ( clk ), .D ( new_AGEMA_signal_13659 ), .Q ( new_AGEMA_signal_13660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2164 ( .C ( clk ), .D ( new_AGEMA_signal_13663 ), .Q ( new_AGEMA_signal_13664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2168 ( .C ( clk ), .D ( new_AGEMA_signal_13667 ), .Q ( new_AGEMA_signal_13668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2172 ( .C ( clk ), .D ( new_AGEMA_signal_13671 ), .Q ( new_AGEMA_signal_13672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2232 ( .C ( clk ), .D ( new_AGEMA_signal_13731 ), .Q ( new_AGEMA_signal_13732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2236 ( .C ( clk ), .D ( new_AGEMA_signal_13735 ), .Q ( new_AGEMA_signal_13736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2240 ( .C ( clk ), .D ( new_AGEMA_signal_13739 ), .Q ( new_AGEMA_signal_13740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2244 ( .C ( clk ), .D ( new_AGEMA_signal_13743 ), .Q ( new_AGEMA_signal_13744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2264 ( .C ( clk ), .D ( new_AGEMA_signal_13763 ), .Q ( new_AGEMA_signal_13764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2268 ( .C ( clk ), .D ( new_AGEMA_signal_13767 ), .Q ( new_AGEMA_signal_13768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2272 ( .C ( clk ), .D ( new_AGEMA_signal_13771 ), .Q ( new_AGEMA_signal_13772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2276 ( .C ( clk ), .D ( new_AGEMA_signal_13775 ), .Q ( new_AGEMA_signal_13776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2560 ( .C ( clk ), .D ( new_AGEMA_signal_14059 ), .Q ( new_AGEMA_signal_14060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2566 ( .C ( clk ), .D ( new_AGEMA_signal_14065 ), .Q ( new_AGEMA_signal_14066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2572 ( .C ( clk ), .D ( new_AGEMA_signal_14071 ), .Q ( new_AGEMA_signal_14072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2578 ( .C ( clk ), .D ( new_AGEMA_signal_14077 ), .Q ( new_AGEMA_signal_14078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2664 ( .C ( clk ), .D ( new_AGEMA_signal_14163 ), .Q ( new_AGEMA_signal_14164 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2670 ( .C ( clk ), .D ( new_AGEMA_signal_14169 ), .Q ( new_AGEMA_signal_14170 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2676 ( .C ( clk ), .D ( new_AGEMA_signal_14175 ), .Q ( new_AGEMA_signal_14176 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2682 ( .C ( clk ), .D ( new_AGEMA_signal_14181 ), .Q ( new_AGEMA_signal_14182 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3128 ( .C ( clk ), .D ( new_AGEMA_signal_14627 ), .Q ( new_AGEMA_signal_14628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3136 ( .C ( clk ), .D ( new_AGEMA_signal_14635 ), .Q ( new_AGEMA_signal_14636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3144 ( .C ( clk ), .D ( new_AGEMA_signal_14643 ), .Q ( new_AGEMA_signal_14644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3152 ( .C ( clk ), .D ( new_AGEMA_signal_14651 ), .Q ( new_AGEMA_signal_14652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3168 ( .C ( clk ), .D ( new_AGEMA_signal_14667 ), .Q ( new_AGEMA_signal_14668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3176 ( .C ( clk ), .D ( new_AGEMA_signal_14675 ), .Q ( new_AGEMA_signal_14676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3184 ( .C ( clk ), .D ( new_AGEMA_signal_14683 ), .Q ( new_AGEMA_signal_14684 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3192 ( .C ( clk ), .D ( new_AGEMA_signal_14691 ), .Q ( new_AGEMA_signal_14692 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3472 ( .C ( clk ), .D ( new_AGEMA_signal_14971 ), .Q ( new_AGEMA_signal_14972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3480 ( .C ( clk ), .D ( new_AGEMA_signal_14979 ), .Q ( new_AGEMA_signal_14980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3488 ( .C ( clk ), .D ( new_AGEMA_signal_14987 ), .Q ( new_AGEMA_signal_14988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3496 ( .C ( clk ), .D ( new_AGEMA_signal_14995 ), .Q ( new_AGEMA_signal_14996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3816 ( .C ( clk ), .D ( new_AGEMA_signal_15315 ), .Q ( new_AGEMA_signal_15316 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3824 ( .C ( clk ), .D ( new_AGEMA_signal_15323 ), .Q ( new_AGEMA_signal_15324 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3832 ( .C ( clk ), .D ( new_AGEMA_signal_15331 ), .Q ( new_AGEMA_signal_15332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3840 ( .C ( clk ), .D ( new_AGEMA_signal_15339 ), .Q ( new_AGEMA_signal_15340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3936 ( .C ( clk ), .D ( new_AGEMA_signal_15435 ), .Q ( new_AGEMA_signal_15436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3944 ( .C ( clk ), .D ( new_AGEMA_signal_15443 ), .Q ( new_AGEMA_signal_15444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3952 ( .C ( clk ), .D ( new_AGEMA_signal_15451 ), .Q ( new_AGEMA_signal_15452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3960 ( .C ( clk ), .D ( new_AGEMA_signal_15459 ), .Q ( new_AGEMA_signal_15460 ) ) ;

    /* cells in depth 5 */
    buf_clk new_AGEMA_reg_buffer_1591 ( .C ( clk ), .D ( n2755 ), .Q ( new_AGEMA_signal_13091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1593 ( .C ( clk ), .D ( new_AGEMA_signal_1206 ), .Q ( new_AGEMA_signal_13093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1595 ( .C ( clk ), .D ( new_AGEMA_signal_1207 ), .Q ( new_AGEMA_signal_13095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1597 ( .C ( clk ), .D ( new_AGEMA_signal_1208 ), .Q ( new_AGEMA_signal_13097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1599 ( .C ( clk ), .D ( n2151 ), .Q ( new_AGEMA_signal_13099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1601 ( .C ( clk ), .D ( new_AGEMA_signal_1512 ), .Q ( new_AGEMA_signal_13101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1603 ( .C ( clk ), .D ( new_AGEMA_signal_1513 ), .Q ( new_AGEMA_signal_13103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1605 ( .C ( clk ), .D ( new_AGEMA_signal_1514 ), .Q ( new_AGEMA_signal_13105 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1609 ( .C ( clk ), .D ( new_AGEMA_signal_13108 ), .Q ( new_AGEMA_signal_13109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1613 ( .C ( clk ), .D ( new_AGEMA_signal_13112 ), .Q ( new_AGEMA_signal_13113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1617 ( .C ( clk ), .D ( new_AGEMA_signal_13116 ), .Q ( new_AGEMA_signal_13117 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1621 ( .C ( clk ), .D ( new_AGEMA_signal_13120 ), .Q ( new_AGEMA_signal_13121 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1623 ( .C ( clk ), .D ( new_AGEMA_signal_12612 ), .Q ( new_AGEMA_signal_13123 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1625 ( .C ( clk ), .D ( new_AGEMA_signal_12614 ), .Q ( new_AGEMA_signal_13125 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1627 ( .C ( clk ), .D ( new_AGEMA_signal_12616 ), .Q ( new_AGEMA_signal_13127 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1629 ( .C ( clk ), .D ( new_AGEMA_signal_12618 ), .Q ( new_AGEMA_signal_13129 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1631 ( .C ( clk ), .D ( new_AGEMA_signal_12588 ), .Q ( new_AGEMA_signal_13131 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1633 ( .C ( clk ), .D ( new_AGEMA_signal_12590 ), .Q ( new_AGEMA_signal_13133 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1635 ( .C ( clk ), .D ( new_AGEMA_signal_12592 ), .Q ( new_AGEMA_signal_13135 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1637 ( .C ( clk ), .D ( new_AGEMA_signal_12594 ), .Q ( new_AGEMA_signal_13137 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1639 ( .C ( clk ), .D ( n1964 ), .Q ( new_AGEMA_signal_13139 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1641 ( .C ( clk ), .D ( new_AGEMA_signal_1113 ), .Q ( new_AGEMA_signal_13141 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1643 ( .C ( clk ), .D ( new_AGEMA_signal_1114 ), .Q ( new_AGEMA_signal_13143 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1645 ( .C ( clk ), .D ( new_AGEMA_signal_1115 ), .Q ( new_AGEMA_signal_13145 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1647 ( .C ( clk ), .D ( n2673 ), .Q ( new_AGEMA_signal_13147 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1649 ( .C ( clk ), .D ( new_AGEMA_signal_1272 ), .Q ( new_AGEMA_signal_13149 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1651 ( .C ( clk ), .D ( new_AGEMA_signal_1273 ), .Q ( new_AGEMA_signal_13151 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1653 ( .C ( clk ), .D ( new_AGEMA_signal_1274 ), .Q ( new_AGEMA_signal_13153 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1655 ( .C ( clk ), .D ( n2359 ), .Q ( new_AGEMA_signal_13155 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1657 ( .C ( clk ), .D ( new_AGEMA_signal_1557 ), .Q ( new_AGEMA_signal_13157 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1659 ( .C ( clk ), .D ( new_AGEMA_signal_1558 ), .Q ( new_AGEMA_signal_13159 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1661 ( .C ( clk ), .D ( new_AGEMA_signal_1559 ), .Q ( new_AGEMA_signal_13161 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1663 ( .C ( clk ), .D ( n1973 ), .Q ( new_AGEMA_signal_13163 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1665 ( .C ( clk ), .D ( new_AGEMA_signal_1569 ), .Q ( new_AGEMA_signal_13165 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1667 ( .C ( clk ), .D ( new_AGEMA_signal_1570 ), .Q ( new_AGEMA_signal_13167 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1669 ( .C ( clk ), .D ( new_AGEMA_signal_1571 ), .Q ( new_AGEMA_signal_13169 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1671 ( .C ( clk ), .D ( n2690 ), .Q ( new_AGEMA_signal_13171 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1673 ( .C ( clk ), .D ( new_AGEMA_signal_1299 ), .Q ( new_AGEMA_signal_13173 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1675 ( .C ( clk ), .D ( new_AGEMA_signal_1300 ), .Q ( new_AGEMA_signal_13175 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1677 ( .C ( clk ), .D ( new_AGEMA_signal_1301 ), .Q ( new_AGEMA_signal_13177 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1679 ( .C ( clk ), .D ( n2741 ), .Q ( new_AGEMA_signal_13179 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1681 ( .C ( clk ), .D ( new_AGEMA_signal_1575 ), .Q ( new_AGEMA_signal_13181 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1683 ( .C ( clk ), .D ( new_AGEMA_signal_1576 ), .Q ( new_AGEMA_signal_13183 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1685 ( .C ( clk ), .D ( new_AGEMA_signal_1577 ), .Q ( new_AGEMA_signal_13185 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1687 ( .C ( clk ), .D ( n1993 ), .Q ( new_AGEMA_signal_13187 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1689 ( .C ( clk ), .D ( new_AGEMA_signal_1308 ), .Q ( new_AGEMA_signal_13189 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1691 ( .C ( clk ), .D ( new_AGEMA_signal_1309 ), .Q ( new_AGEMA_signal_13191 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1693 ( .C ( clk ), .D ( new_AGEMA_signal_1310 ), .Q ( new_AGEMA_signal_13193 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1695 ( .C ( clk ), .D ( n2241 ), .Q ( new_AGEMA_signal_13195 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1697 ( .C ( clk ), .D ( new_AGEMA_signal_1587 ), .Q ( new_AGEMA_signal_13197 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1699 ( .C ( clk ), .D ( new_AGEMA_signal_1588 ), .Q ( new_AGEMA_signal_13199 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1701 ( .C ( clk ), .D ( new_AGEMA_signal_1589 ), .Q ( new_AGEMA_signal_13201 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1703 ( .C ( clk ), .D ( new_AGEMA_signal_12828 ), .Q ( new_AGEMA_signal_13203 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1705 ( .C ( clk ), .D ( new_AGEMA_signal_12830 ), .Q ( new_AGEMA_signal_13205 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1707 ( .C ( clk ), .D ( new_AGEMA_signal_12832 ), .Q ( new_AGEMA_signal_13207 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1709 ( .C ( clk ), .D ( new_AGEMA_signal_12834 ), .Q ( new_AGEMA_signal_13209 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1713 ( .C ( clk ), .D ( new_AGEMA_signal_13212 ), .Q ( new_AGEMA_signal_13213 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1717 ( .C ( clk ), .D ( new_AGEMA_signal_13216 ), .Q ( new_AGEMA_signal_13217 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1721 ( .C ( clk ), .D ( new_AGEMA_signal_13220 ), .Q ( new_AGEMA_signal_13221 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1725 ( .C ( clk ), .D ( new_AGEMA_signal_13224 ), .Q ( new_AGEMA_signal_13225 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1727 ( .C ( clk ), .D ( n2290 ), .Q ( new_AGEMA_signal_13227 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1729 ( .C ( clk ), .D ( new_AGEMA_signal_1620 ), .Q ( new_AGEMA_signal_13229 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1731 ( .C ( clk ), .D ( new_AGEMA_signal_1621 ), .Q ( new_AGEMA_signal_13231 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1733 ( .C ( clk ), .D ( new_AGEMA_signal_1622 ), .Q ( new_AGEMA_signal_13233 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1735 ( .C ( clk ), .D ( n2171 ), .Q ( new_AGEMA_signal_13235 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1737 ( .C ( clk ), .D ( new_AGEMA_signal_1335 ), .Q ( new_AGEMA_signal_13237 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1739 ( .C ( clk ), .D ( new_AGEMA_signal_1336 ), .Q ( new_AGEMA_signal_13239 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1741 ( .C ( clk ), .D ( new_AGEMA_signal_1337 ), .Q ( new_AGEMA_signal_13241 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1743 ( .C ( clk ), .D ( n2042 ), .Q ( new_AGEMA_signal_13243 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1745 ( .C ( clk ), .D ( new_AGEMA_signal_1632 ), .Q ( new_AGEMA_signal_13245 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1747 ( .C ( clk ), .D ( new_AGEMA_signal_1633 ), .Q ( new_AGEMA_signal_13247 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1749 ( .C ( clk ), .D ( new_AGEMA_signal_1634 ), .Q ( new_AGEMA_signal_13249 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1751 ( .C ( clk ), .D ( n2754 ), .Q ( new_AGEMA_signal_13251 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1753 ( .C ( clk ), .D ( new_AGEMA_signal_1635 ), .Q ( new_AGEMA_signal_13253 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1755 ( .C ( clk ), .D ( new_AGEMA_signal_1636 ), .Q ( new_AGEMA_signal_13255 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1757 ( .C ( clk ), .D ( new_AGEMA_signal_1637 ), .Q ( new_AGEMA_signal_13257 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1759 ( .C ( clk ), .D ( new_AGEMA_signal_12548 ), .Q ( new_AGEMA_signal_13259 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1761 ( .C ( clk ), .D ( new_AGEMA_signal_12550 ), .Q ( new_AGEMA_signal_13261 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1763 ( .C ( clk ), .D ( new_AGEMA_signal_12552 ), .Q ( new_AGEMA_signal_13263 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1765 ( .C ( clk ), .D ( new_AGEMA_signal_12554 ), .Q ( new_AGEMA_signal_13265 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1767 ( .C ( clk ), .D ( n2535 ), .Q ( new_AGEMA_signal_13267 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1769 ( .C ( clk ), .D ( new_AGEMA_signal_1566 ), .Q ( new_AGEMA_signal_13269 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1771 ( .C ( clk ), .D ( new_AGEMA_signal_1567 ), .Q ( new_AGEMA_signal_13271 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1773 ( .C ( clk ), .D ( new_AGEMA_signal_1568 ), .Q ( new_AGEMA_signal_13273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1775 ( .C ( clk ), .D ( n2642 ), .Q ( new_AGEMA_signal_13275 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1777 ( .C ( clk ), .D ( new_AGEMA_signal_1338 ), .Q ( new_AGEMA_signal_13277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1779 ( .C ( clk ), .D ( new_AGEMA_signal_1339 ), .Q ( new_AGEMA_signal_13279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1781 ( .C ( clk ), .D ( new_AGEMA_signal_1340 ), .Q ( new_AGEMA_signal_13281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1785 ( .C ( clk ), .D ( new_AGEMA_signal_13284 ), .Q ( new_AGEMA_signal_13285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1789 ( .C ( clk ), .D ( new_AGEMA_signal_13288 ), .Q ( new_AGEMA_signal_13289 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1793 ( .C ( clk ), .D ( new_AGEMA_signal_13292 ), .Q ( new_AGEMA_signal_13293 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1797 ( .C ( clk ), .D ( new_AGEMA_signal_13296 ), .Q ( new_AGEMA_signal_13297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1799 ( .C ( clk ), .D ( n2773 ), .Q ( new_AGEMA_signal_13299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1801 ( .C ( clk ), .D ( new_AGEMA_signal_1668 ), .Q ( new_AGEMA_signal_13301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1803 ( .C ( clk ), .D ( new_AGEMA_signal_1669 ), .Q ( new_AGEMA_signal_13303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1805 ( .C ( clk ), .D ( new_AGEMA_signal_1670 ), .Q ( new_AGEMA_signal_13305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1807 ( .C ( clk ), .D ( n2627 ), .Q ( new_AGEMA_signal_13307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1809 ( .C ( clk ), .D ( new_AGEMA_signal_1260 ), .Q ( new_AGEMA_signal_13309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1811 ( .C ( clk ), .D ( new_AGEMA_signal_1261 ), .Q ( new_AGEMA_signal_13311 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1813 ( .C ( clk ), .D ( new_AGEMA_signal_1262 ), .Q ( new_AGEMA_signal_13313 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1815 ( .C ( clk ), .D ( new_AGEMA_signal_12708 ), .Q ( new_AGEMA_signal_13315 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1817 ( .C ( clk ), .D ( new_AGEMA_signal_12710 ), .Q ( new_AGEMA_signal_13317 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1819 ( .C ( clk ), .D ( new_AGEMA_signal_12712 ), .Q ( new_AGEMA_signal_13319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1821 ( .C ( clk ), .D ( new_AGEMA_signal_12714 ), .Q ( new_AGEMA_signal_13321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1823 ( .C ( clk ), .D ( n2631 ), .Q ( new_AGEMA_signal_13323 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1825 ( .C ( clk ), .D ( new_AGEMA_signal_1218 ), .Q ( new_AGEMA_signal_13325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1827 ( .C ( clk ), .D ( new_AGEMA_signal_1219 ), .Q ( new_AGEMA_signal_13327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1829 ( .C ( clk ), .D ( new_AGEMA_signal_1220 ), .Q ( new_AGEMA_signal_13329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1831 ( .C ( clk ), .D ( n2376 ), .Q ( new_AGEMA_signal_13331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1833 ( .C ( clk ), .D ( new_AGEMA_signal_1623 ), .Q ( new_AGEMA_signal_13333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1835 ( .C ( clk ), .D ( new_AGEMA_signal_1624 ), .Q ( new_AGEMA_signal_13335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1837 ( .C ( clk ), .D ( new_AGEMA_signal_1625 ), .Q ( new_AGEMA_signal_13337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1841 ( .C ( clk ), .D ( new_AGEMA_signal_13340 ), .Q ( new_AGEMA_signal_13341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1845 ( .C ( clk ), .D ( new_AGEMA_signal_13344 ), .Q ( new_AGEMA_signal_13345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1849 ( .C ( clk ), .D ( new_AGEMA_signal_13348 ), .Q ( new_AGEMA_signal_13349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1853 ( .C ( clk ), .D ( new_AGEMA_signal_13352 ), .Q ( new_AGEMA_signal_13353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1855 ( .C ( clk ), .D ( new_AGEMA_signal_12892 ), .Q ( new_AGEMA_signal_13355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1857 ( .C ( clk ), .D ( new_AGEMA_signal_12894 ), .Q ( new_AGEMA_signal_13357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1859 ( .C ( clk ), .D ( new_AGEMA_signal_12896 ), .Q ( new_AGEMA_signal_13359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1861 ( .C ( clk ), .D ( new_AGEMA_signal_12898 ), .Q ( new_AGEMA_signal_13361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1863 ( .C ( clk ), .D ( new_AGEMA_signal_12748 ), .Q ( new_AGEMA_signal_13363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1865 ( .C ( clk ), .D ( new_AGEMA_signal_12750 ), .Q ( new_AGEMA_signal_13365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1867 ( .C ( clk ), .D ( new_AGEMA_signal_12752 ), .Q ( new_AGEMA_signal_13367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1869 ( .C ( clk ), .D ( new_AGEMA_signal_12754 ), .Q ( new_AGEMA_signal_13369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1871 ( .C ( clk ), .D ( new_AGEMA_signal_12780 ), .Q ( new_AGEMA_signal_13371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1873 ( .C ( clk ), .D ( new_AGEMA_signal_12782 ), .Q ( new_AGEMA_signal_13373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1875 ( .C ( clk ), .D ( new_AGEMA_signal_12784 ), .Q ( new_AGEMA_signal_13375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1877 ( .C ( clk ), .D ( new_AGEMA_signal_12786 ), .Q ( new_AGEMA_signal_13377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1881 ( .C ( clk ), .D ( new_AGEMA_signal_13380 ), .Q ( new_AGEMA_signal_13381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1885 ( .C ( clk ), .D ( new_AGEMA_signal_13384 ), .Q ( new_AGEMA_signal_13385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1889 ( .C ( clk ), .D ( new_AGEMA_signal_13388 ), .Q ( new_AGEMA_signal_13389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1893 ( .C ( clk ), .D ( new_AGEMA_signal_13392 ), .Q ( new_AGEMA_signal_13393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1895 ( .C ( clk ), .D ( new_AGEMA_signal_13052 ), .Q ( new_AGEMA_signal_13395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1897 ( .C ( clk ), .D ( new_AGEMA_signal_13054 ), .Q ( new_AGEMA_signal_13397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1899 ( .C ( clk ), .D ( new_AGEMA_signal_13056 ), .Q ( new_AGEMA_signal_13399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1901 ( .C ( clk ), .D ( new_AGEMA_signal_13058 ), .Q ( new_AGEMA_signal_13401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1903 ( .C ( clk ), .D ( n2498 ), .Q ( new_AGEMA_signal_13403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1905 ( .C ( clk ), .D ( new_AGEMA_signal_1347 ), .Q ( new_AGEMA_signal_13405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1907 ( .C ( clk ), .D ( new_AGEMA_signal_1348 ), .Q ( new_AGEMA_signal_13407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1909 ( .C ( clk ), .D ( new_AGEMA_signal_1349 ), .Q ( new_AGEMA_signal_13409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1911 ( .C ( clk ), .D ( n2178 ), .Q ( new_AGEMA_signal_13411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1913 ( .C ( clk ), .D ( new_AGEMA_signal_1371 ), .Q ( new_AGEMA_signal_13413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1915 ( .C ( clk ), .D ( new_AGEMA_signal_1372 ), .Q ( new_AGEMA_signal_13415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1917 ( .C ( clk ), .D ( new_AGEMA_signal_1373 ), .Q ( new_AGEMA_signal_13417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1921 ( .C ( clk ), .D ( new_AGEMA_signal_13420 ), .Q ( new_AGEMA_signal_13421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1925 ( .C ( clk ), .D ( new_AGEMA_signal_13424 ), .Q ( new_AGEMA_signal_13425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1929 ( .C ( clk ), .D ( new_AGEMA_signal_13428 ), .Q ( new_AGEMA_signal_13429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1933 ( .C ( clk ), .D ( new_AGEMA_signal_13432 ), .Q ( new_AGEMA_signal_13433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1935 ( .C ( clk ), .D ( n2505 ), .Q ( new_AGEMA_signal_13435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1937 ( .C ( clk ), .D ( new_AGEMA_signal_1554 ), .Q ( new_AGEMA_signal_13437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1939 ( .C ( clk ), .D ( new_AGEMA_signal_1555 ), .Q ( new_AGEMA_signal_13439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1941 ( .C ( clk ), .D ( new_AGEMA_signal_1556 ), .Q ( new_AGEMA_signal_13441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1943 ( .C ( clk ), .D ( n2540 ), .Q ( new_AGEMA_signal_13443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1945 ( .C ( clk ), .D ( new_AGEMA_signal_1779 ), .Q ( new_AGEMA_signal_13445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1947 ( .C ( clk ), .D ( new_AGEMA_signal_1780 ), .Q ( new_AGEMA_signal_13447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1949 ( .C ( clk ), .D ( new_AGEMA_signal_1781 ), .Q ( new_AGEMA_signal_13449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1951 ( .C ( clk ), .D ( n2266 ), .Q ( new_AGEMA_signal_13451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1953 ( .C ( clk ), .D ( new_AGEMA_signal_1392 ), .Q ( new_AGEMA_signal_13453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1955 ( .C ( clk ), .D ( new_AGEMA_signal_1393 ), .Q ( new_AGEMA_signal_13455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1957 ( .C ( clk ), .D ( new_AGEMA_signal_1394 ), .Q ( new_AGEMA_signal_13457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1959 ( .C ( clk ), .D ( n2278 ), .Q ( new_AGEMA_signal_13459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1961 ( .C ( clk ), .D ( new_AGEMA_signal_1791 ), .Q ( new_AGEMA_signal_13461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1963 ( .C ( clk ), .D ( new_AGEMA_signal_1792 ), .Q ( new_AGEMA_signal_13463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1965 ( .C ( clk ), .D ( new_AGEMA_signal_1793 ), .Q ( new_AGEMA_signal_13465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1967 ( .C ( clk ), .D ( new_AGEMA_signal_12876 ), .Q ( new_AGEMA_signal_13467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1969 ( .C ( clk ), .D ( new_AGEMA_signal_12878 ), .Q ( new_AGEMA_signal_13469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1971 ( .C ( clk ), .D ( new_AGEMA_signal_12880 ), .Q ( new_AGEMA_signal_13471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1973 ( .C ( clk ), .D ( new_AGEMA_signal_12882 ), .Q ( new_AGEMA_signal_13473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1975 ( .C ( clk ), .D ( new_AGEMA_signal_12964 ), .Q ( new_AGEMA_signal_13475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1977 ( .C ( clk ), .D ( new_AGEMA_signal_12966 ), .Q ( new_AGEMA_signal_13477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1979 ( .C ( clk ), .D ( new_AGEMA_signal_12968 ), .Q ( new_AGEMA_signal_13479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1981 ( .C ( clk ), .D ( new_AGEMA_signal_12970 ), .Q ( new_AGEMA_signal_13481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1983 ( .C ( clk ), .D ( new_AGEMA_signal_12692 ), .Q ( new_AGEMA_signal_13483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1985 ( .C ( clk ), .D ( new_AGEMA_signal_12694 ), .Q ( new_AGEMA_signal_13485 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1987 ( .C ( clk ), .D ( new_AGEMA_signal_12696 ), .Q ( new_AGEMA_signal_13487 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1989 ( .C ( clk ), .D ( new_AGEMA_signal_12698 ), .Q ( new_AGEMA_signal_13489 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1991 ( .C ( clk ), .D ( new_AGEMA_signal_12676 ), .Q ( new_AGEMA_signal_13491 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1993 ( .C ( clk ), .D ( new_AGEMA_signal_12678 ), .Q ( new_AGEMA_signal_13493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1995 ( .C ( clk ), .D ( new_AGEMA_signal_12680 ), .Q ( new_AGEMA_signal_13495 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1997 ( .C ( clk ), .D ( new_AGEMA_signal_12682 ), .Q ( new_AGEMA_signal_13497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1999 ( .C ( clk ), .D ( n2318 ), .Q ( new_AGEMA_signal_13499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2001 ( .C ( clk ), .D ( new_AGEMA_signal_1410 ), .Q ( new_AGEMA_signal_13501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2003 ( .C ( clk ), .D ( new_AGEMA_signal_1411 ), .Q ( new_AGEMA_signal_13503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2005 ( .C ( clk ), .D ( new_AGEMA_signal_1412 ), .Q ( new_AGEMA_signal_13505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2007 ( .C ( clk ), .D ( n2325 ), .Q ( new_AGEMA_signal_13507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2009 ( .C ( clk ), .D ( new_AGEMA_signal_1821 ), .Q ( new_AGEMA_signal_13509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2011 ( .C ( clk ), .D ( new_AGEMA_signal_1822 ), .Q ( new_AGEMA_signal_13511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2013 ( .C ( clk ), .D ( new_AGEMA_signal_1823 ), .Q ( new_AGEMA_signal_13513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2015 ( .C ( clk ), .D ( n2677 ), .Q ( new_AGEMA_signal_13515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2017 ( .C ( clk ), .D ( new_AGEMA_signal_1257 ), .Q ( new_AGEMA_signal_13517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2019 ( .C ( clk ), .D ( new_AGEMA_signal_1258 ), .Q ( new_AGEMA_signal_13519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2021 ( .C ( clk ), .D ( new_AGEMA_signal_1259 ), .Q ( new_AGEMA_signal_13521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2023 ( .C ( clk ), .D ( new_AGEMA_signal_13036 ), .Q ( new_AGEMA_signal_13523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2025 ( .C ( clk ), .D ( new_AGEMA_signal_13038 ), .Q ( new_AGEMA_signal_13525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2027 ( .C ( clk ), .D ( new_AGEMA_signal_13040 ), .Q ( new_AGEMA_signal_13527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2029 ( .C ( clk ), .D ( new_AGEMA_signal_13042 ), .Q ( new_AGEMA_signal_13529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2031 ( .C ( clk ), .D ( new_AGEMA_signal_13068 ), .Q ( new_AGEMA_signal_13531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2033 ( .C ( clk ), .D ( new_AGEMA_signal_13070 ), .Q ( new_AGEMA_signal_13533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2035 ( .C ( clk ), .D ( new_AGEMA_signal_13072 ), .Q ( new_AGEMA_signal_13535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2037 ( .C ( clk ), .D ( new_AGEMA_signal_13074 ), .Q ( new_AGEMA_signal_13537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2039 ( .C ( clk ), .D ( new_AGEMA_signal_12764 ), .Q ( new_AGEMA_signal_13539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2041 ( .C ( clk ), .D ( new_AGEMA_signal_12766 ), .Q ( new_AGEMA_signal_13541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2043 ( .C ( clk ), .D ( new_AGEMA_signal_12768 ), .Q ( new_AGEMA_signal_13543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2045 ( .C ( clk ), .D ( new_AGEMA_signal_12770 ), .Q ( new_AGEMA_signal_13545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2047 ( .C ( clk ), .D ( new_AGEMA_signal_12564 ), .Q ( new_AGEMA_signal_13547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2049 ( .C ( clk ), .D ( new_AGEMA_signal_12566 ), .Q ( new_AGEMA_signal_13549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2051 ( .C ( clk ), .D ( new_AGEMA_signal_12568 ), .Q ( new_AGEMA_signal_13551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2053 ( .C ( clk ), .D ( new_AGEMA_signal_12570 ), .Q ( new_AGEMA_signal_13553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2055 ( .C ( clk ), .D ( n2625 ), .Q ( new_AGEMA_signal_13555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2057 ( .C ( clk ), .D ( new_AGEMA_signal_1560 ), .Q ( new_AGEMA_signal_13557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2059 ( .C ( clk ), .D ( new_AGEMA_signal_1561 ), .Q ( new_AGEMA_signal_13559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2061 ( .C ( clk ), .D ( new_AGEMA_signal_1562 ), .Q ( new_AGEMA_signal_13561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2063 ( .C ( clk ), .D ( n2431 ), .Q ( new_AGEMA_signal_13563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2065 ( .C ( clk ), .D ( new_AGEMA_signal_1884 ), .Q ( new_AGEMA_signal_13565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2067 ( .C ( clk ), .D ( new_AGEMA_signal_1885 ), .Q ( new_AGEMA_signal_13567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2069 ( .C ( clk ), .D ( new_AGEMA_signal_1886 ), .Q ( new_AGEMA_signal_13569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2075 ( .C ( clk ), .D ( new_AGEMA_signal_13574 ), .Q ( new_AGEMA_signal_13575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2081 ( .C ( clk ), .D ( new_AGEMA_signal_13580 ), .Q ( new_AGEMA_signal_13581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2087 ( .C ( clk ), .D ( new_AGEMA_signal_13586 ), .Q ( new_AGEMA_signal_13587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2093 ( .C ( clk ), .D ( new_AGEMA_signal_13592 ), .Q ( new_AGEMA_signal_13593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2095 ( .C ( clk ), .D ( n2453 ), .Q ( new_AGEMA_signal_13595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2097 ( .C ( clk ), .D ( new_AGEMA_signal_1440 ), .Q ( new_AGEMA_signal_13597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2099 ( .C ( clk ), .D ( new_AGEMA_signal_1441 ), .Q ( new_AGEMA_signal_13599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2101 ( .C ( clk ), .D ( new_AGEMA_signal_1442 ), .Q ( new_AGEMA_signal_13601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2103 ( .C ( clk ), .D ( n2475 ), .Q ( new_AGEMA_signal_13603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2105 ( .C ( clk ), .D ( new_AGEMA_signal_1455 ), .Q ( new_AGEMA_signal_13605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2107 ( .C ( clk ), .D ( new_AGEMA_signal_1456 ), .Q ( new_AGEMA_signal_13607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2109 ( .C ( clk ), .D ( new_AGEMA_signal_1457 ), .Q ( new_AGEMA_signal_13609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2111 ( .C ( clk ), .D ( n2487 ), .Q ( new_AGEMA_signal_13611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2113 ( .C ( clk ), .D ( new_AGEMA_signal_1908 ), .Q ( new_AGEMA_signal_13613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2115 ( .C ( clk ), .D ( new_AGEMA_signal_1909 ), .Q ( new_AGEMA_signal_13615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2117 ( .C ( clk ), .D ( new_AGEMA_signal_1910 ), .Q ( new_AGEMA_signal_13617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2121 ( .C ( clk ), .D ( new_AGEMA_signal_13620 ), .Q ( new_AGEMA_signal_13621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2125 ( .C ( clk ), .D ( new_AGEMA_signal_13624 ), .Q ( new_AGEMA_signal_13625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2129 ( .C ( clk ), .D ( new_AGEMA_signal_13628 ), .Q ( new_AGEMA_signal_13629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2133 ( .C ( clk ), .D ( new_AGEMA_signal_13632 ), .Q ( new_AGEMA_signal_13633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2135 ( .C ( clk ), .D ( new_AGEMA_signal_12844 ), .Q ( new_AGEMA_signal_13635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2137 ( .C ( clk ), .D ( new_AGEMA_signal_12846 ), .Q ( new_AGEMA_signal_13637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2139 ( .C ( clk ), .D ( new_AGEMA_signal_12848 ), .Q ( new_AGEMA_signal_13639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2141 ( .C ( clk ), .D ( new_AGEMA_signal_12850 ), .Q ( new_AGEMA_signal_13641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2143 ( .C ( clk ), .D ( new_AGEMA_signal_12860 ), .Q ( new_AGEMA_signal_13643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2145 ( .C ( clk ), .D ( new_AGEMA_signal_12862 ), .Q ( new_AGEMA_signal_13645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2147 ( .C ( clk ), .D ( new_AGEMA_signal_12864 ), .Q ( new_AGEMA_signal_13647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2149 ( .C ( clk ), .D ( new_AGEMA_signal_12866 ), .Q ( new_AGEMA_signal_13649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2151 ( .C ( clk ), .D ( n2564 ), .Q ( new_AGEMA_signal_13651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2153 ( .C ( clk ), .D ( new_AGEMA_signal_1941 ), .Q ( new_AGEMA_signal_13653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2155 ( .C ( clk ), .D ( new_AGEMA_signal_1942 ), .Q ( new_AGEMA_signal_13655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2157 ( .C ( clk ), .D ( new_AGEMA_signal_1943 ), .Q ( new_AGEMA_signal_13657 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2161 ( .C ( clk ), .D ( new_AGEMA_signal_13660 ), .Q ( new_AGEMA_signal_13661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2165 ( .C ( clk ), .D ( new_AGEMA_signal_13664 ), .Q ( new_AGEMA_signal_13665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2169 ( .C ( clk ), .D ( new_AGEMA_signal_13668 ), .Q ( new_AGEMA_signal_13669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2173 ( .C ( clk ), .D ( new_AGEMA_signal_13672 ), .Q ( new_AGEMA_signal_13673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2175 ( .C ( clk ), .D ( n2617 ), .Q ( new_AGEMA_signal_13675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2177 ( .C ( clk ), .D ( new_AGEMA_signal_1473 ), .Q ( new_AGEMA_signal_13677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2179 ( .C ( clk ), .D ( new_AGEMA_signal_1474 ), .Q ( new_AGEMA_signal_13679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2181 ( .C ( clk ), .D ( new_AGEMA_signal_1475 ), .Q ( new_AGEMA_signal_13681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2183 ( .C ( clk ), .D ( n2647 ), .Q ( new_AGEMA_signal_13683 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2185 ( .C ( clk ), .D ( new_AGEMA_signal_1359 ), .Q ( new_AGEMA_signal_13685 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2187 ( .C ( clk ), .D ( new_AGEMA_signal_1360 ), .Q ( new_AGEMA_signal_13687 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2189 ( .C ( clk ), .D ( new_AGEMA_signal_1361 ), .Q ( new_AGEMA_signal_13689 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2191 ( .C ( clk ), .D ( n2674 ), .Q ( new_AGEMA_signal_13691 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2193 ( .C ( clk ), .D ( new_AGEMA_signal_2241 ), .Q ( new_AGEMA_signal_13693 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2195 ( .C ( clk ), .D ( new_AGEMA_signal_2242 ), .Q ( new_AGEMA_signal_13695 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2197 ( .C ( clk ), .D ( new_AGEMA_signal_2243 ), .Q ( new_AGEMA_signal_13697 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2199 ( .C ( clk ), .D ( n2683 ), .Q ( new_AGEMA_signal_13699 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2201 ( .C ( clk ), .D ( new_AGEMA_signal_1182 ), .Q ( new_AGEMA_signal_13701 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2203 ( .C ( clk ), .D ( new_AGEMA_signal_1183 ), .Q ( new_AGEMA_signal_13703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2205 ( .C ( clk ), .D ( new_AGEMA_signal_1184 ), .Q ( new_AGEMA_signal_13705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2207 ( .C ( clk ), .D ( n2714 ), .Q ( new_AGEMA_signal_13707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2209 ( .C ( clk ), .D ( new_AGEMA_signal_1482 ), .Q ( new_AGEMA_signal_13709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2211 ( .C ( clk ), .D ( new_AGEMA_signal_1483 ), .Q ( new_AGEMA_signal_13711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2213 ( .C ( clk ), .D ( new_AGEMA_signal_1484 ), .Q ( new_AGEMA_signal_13713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2215 ( .C ( clk ), .D ( n2726 ), .Q ( new_AGEMA_signal_13715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2217 ( .C ( clk ), .D ( new_AGEMA_signal_2007 ), .Q ( new_AGEMA_signal_13717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2219 ( .C ( clk ), .D ( new_AGEMA_signal_2008 ), .Q ( new_AGEMA_signal_13719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2221 ( .C ( clk ), .D ( new_AGEMA_signal_2009 ), .Q ( new_AGEMA_signal_13721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2223 ( .C ( clk ), .D ( n2734 ), .Q ( new_AGEMA_signal_13723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2225 ( .C ( clk ), .D ( new_AGEMA_signal_1515 ), .Q ( new_AGEMA_signal_13725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2227 ( .C ( clk ), .D ( new_AGEMA_signal_1516 ), .Q ( new_AGEMA_signal_13727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2229 ( .C ( clk ), .D ( new_AGEMA_signal_1517 ), .Q ( new_AGEMA_signal_13729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2233 ( .C ( clk ), .D ( new_AGEMA_signal_13732 ), .Q ( new_AGEMA_signal_13733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2237 ( .C ( clk ), .D ( new_AGEMA_signal_13736 ), .Q ( new_AGEMA_signal_13737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2241 ( .C ( clk ), .D ( new_AGEMA_signal_13740 ), .Q ( new_AGEMA_signal_13741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2245 ( .C ( clk ), .D ( new_AGEMA_signal_13744 ), .Q ( new_AGEMA_signal_13745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2247 ( .C ( clk ), .D ( n2763 ), .Q ( new_AGEMA_signal_13747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2249 ( .C ( clk ), .D ( new_AGEMA_signal_1518 ), .Q ( new_AGEMA_signal_13749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2251 ( .C ( clk ), .D ( new_AGEMA_signal_1519 ), .Q ( new_AGEMA_signal_13751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2253 ( .C ( clk ), .D ( new_AGEMA_signal_1520 ), .Q ( new_AGEMA_signal_13753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2255 ( .C ( clk ), .D ( n2784 ), .Q ( new_AGEMA_signal_13755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2257 ( .C ( clk ), .D ( new_AGEMA_signal_1977 ), .Q ( new_AGEMA_signal_13757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2259 ( .C ( clk ), .D ( new_AGEMA_signal_1978 ), .Q ( new_AGEMA_signal_13759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2261 ( .C ( clk ), .D ( new_AGEMA_signal_1979 ), .Q ( new_AGEMA_signal_13761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2265 ( .C ( clk ), .D ( new_AGEMA_signal_13764 ), .Q ( new_AGEMA_signal_13765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2269 ( .C ( clk ), .D ( new_AGEMA_signal_13768 ), .Q ( new_AGEMA_signal_13769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2273 ( .C ( clk ), .D ( new_AGEMA_signal_13772 ), .Q ( new_AGEMA_signal_13773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2277 ( .C ( clk ), .D ( new_AGEMA_signal_13776 ), .Q ( new_AGEMA_signal_13777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2279 ( .C ( clk ), .D ( n2820 ), .Q ( new_AGEMA_signal_13779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2281 ( .C ( clk ), .D ( new_AGEMA_signal_1494 ), .Q ( new_AGEMA_signal_13781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2283 ( .C ( clk ), .D ( new_AGEMA_signal_1495 ), .Q ( new_AGEMA_signal_13783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2285 ( .C ( clk ), .D ( new_AGEMA_signal_1496 ), .Q ( new_AGEMA_signal_13785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2287 ( .C ( clk ), .D ( new_AGEMA_signal_13020 ), .Q ( new_AGEMA_signal_13787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2291 ( .C ( clk ), .D ( new_AGEMA_signal_13022 ), .Q ( new_AGEMA_signal_13791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2295 ( .C ( clk ), .D ( new_AGEMA_signal_13024 ), .Q ( new_AGEMA_signal_13795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2299 ( .C ( clk ), .D ( new_AGEMA_signal_13026 ), .Q ( new_AGEMA_signal_13799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2303 ( .C ( clk ), .D ( n1930 ), .Q ( new_AGEMA_signal_13803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2307 ( .C ( clk ), .D ( new_AGEMA_signal_1224 ), .Q ( new_AGEMA_signal_13807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2311 ( .C ( clk ), .D ( new_AGEMA_signal_1225 ), .Q ( new_AGEMA_signal_13811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2315 ( .C ( clk ), .D ( new_AGEMA_signal_1226 ), .Q ( new_AGEMA_signal_13815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2335 ( .C ( clk ), .D ( n1976 ), .Q ( new_AGEMA_signal_13835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2339 ( .C ( clk ), .D ( new_AGEMA_signal_1296 ), .Q ( new_AGEMA_signal_13839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2343 ( .C ( clk ), .D ( new_AGEMA_signal_1297 ), .Q ( new_AGEMA_signal_13843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2347 ( .C ( clk ), .D ( new_AGEMA_signal_1298 ), .Q ( new_AGEMA_signal_13847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2359 ( .C ( clk ), .D ( new_AGEMA_signal_12684 ), .Q ( new_AGEMA_signal_13859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2363 ( .C ( clk ), .D ( new_AGEMA_signal_12686 ), .Q ( new_AGEMA_signal_13863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2367 ( .C ( clk ), .D ( new_AGEMA_signal_12688 ), .Q ( new_AGEMA_signal_13867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2371 ( .C ( clk ), .D ( new_AGEMA_signal_12690 ), .Q ( new_AGEMA_signal_13871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2383 ( .C ( clk ), .D ( n2008 ), .Q ( new_AGEMA_signal_13883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2387 ( .C ( clk ), .D ( new_AGEMA_signal_1593 ), .Q ( new_AGEMA_signal_13887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2391 ( .C ( clk ), .D ( new_AGEMA_signal_1594 ), .Q ( new_AGEMA_signal_13891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2395 ( .C ( clk ), .D ( new_AGEMA_signal_1595 ), .Q ( new_AGEMA_signal_13895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2399 ( .C ( clk ), .D ( n2022 ), .Q ( new_AGEMA_signal_13899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2403 ( .C ( clk ), .D ( new_AGEMA_signal_1608 ), .Q ( new_AGEMA_signal_13903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2407 ( .C ( clk ), .D ( new_AGEMA_signal_1609 ), .Q ( new_AGEMA_signal_13907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2411 ( .C ( clk ), .D ( new_AGEMA_signal_1610 ), .Q ( new_AGEMA_signal_13911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2447 ( .C ( clk ), .D ( n2057 ), .Q ( new_AGEMA_signal_13947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2451 ( .C ( clk ), .D ( new_AGEMA_signal_1647 ), .Q ( new_AGEMA_signal_13951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2455 ( .C ( clk ), .D ( new_AGEMA_signal_1648 ), .Q ( new_AGEMA_signal_13955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2459 ( .C ( clk ), .D ( new_AGEMA_signal_1649 ), .Q ( new_AGEMA_signal_13959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2463 ( .C ( clk ), .D ( n2062 ), .Q ( new_AGEMA_signal_13963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2467 ( .C ( clk ), .D ( new_AGEMA_signal_1653 ), .Q ( new_AGEMA_signal_13967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2471 ( .C ( clk ), .D ( new_AGEMA_signal_1654 ), .Q ( new_AGEMA_signal_13971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2475 ( .C ( clk ), .D ( new_AGEMA_signal_1655 ), .Q ( new_AGEMA_signal_13975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2479 ( .C ( clk ), .D ( n2075 ), .Q ( new_AGEMA_signal_13979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2483 ( .C ( clk ), .D ( new_AGEMA_signal_1341 ), .Q ( new_AGEMA_signal_13983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2487 ( .C ( clk ), .D ( new_AGEMA_signal_1342 ), .Q ( new_AGEMA_signal_13987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2491 ( .C ( clk ), .D ( new_AGEMA_signal_1343 ), .Q ( new_AGEMA_signal_13991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2519 ( .C ( clk ), .D ( n2121 ), .Q ( new_AGEMA_signal_14019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2523 ( .C ( clk ), .D ( new_AGEMA_signal_1689 ), .Q ( new_AGEMA_signal_14023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2527 ( .C ( clk ), .D ( new_AGEMA_signal_1690 ), .Q ( new_AGEMA_signal_14027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2531 ( .C ( clk ), .D ( new_AGEMA_signal_1691 ), .Q ( new_AGEMA_signal_14031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2543 ( .C ( clk ), .D ( new_AGEMA_signal_12644 ), .Q ( new_AGEMA_signal_14043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2547 ( .C ( clk ), .D ( new_AGEMA_signal_12646 ), .Q ( new_AGEMA_signal_14047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2551 ( .C ( clk ), .D ( new_AGEMA_signal_12648 ), .Q ( new_AGEMA_signal_14051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2555 ( .C ( clk ), .D ( new_AGEMA_signal_12650 ), .Q ( new_AGEMA_signal_14055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2561 ( .C ( clk ), .D ( new_AGEMA_signal_14060 ), .Q ( new_AGEMA_signal_14061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2567 ( .C ( clk ), .D ( new_AGEMA_signal_14066 ), .Q ( new_AGEMA_signal_14067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2573 ( .C ( clk ), .D ( new_AGEMA_signal_14072 ), .Q ( new_AGEMA_signal_14073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2579 ( .C ( clk ), .D ( new_AGEMA_signal_14078 ), .Q ( new_AGEMA_signal_14079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2583 ( .C ( clk ), .D ( new_AGEMA_signal_12932 ), .Q ( new_AGEMA_signal_14083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2587 ( .C ( clk ), .D ( new_AGEMA_signal_12934 ), .Q ( new_AGEMA_signal_14087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2591 ( .C ( clk ), .D ( new_AGEMA_signal_12936 ), .Q ( new_AGEMA_signal_14091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2595 ( .C ( clk ), .D ( new_AGEMA_signal_12938 ), .Q ( new_AGEMA_signal_14095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2599 ( .C ( clk ), .D ( new_AGEMA_signal_12988 ), .Q ( new_AGEMA_signal_14099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2603 ( .C ( clk ), .D ( new_AGEMA_signal_12990 ), .Q ( new_AGEMA_signal_14103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2607 ( .C ( clk ), .D ( new_AGEMA_signal_12992 ), .Q ( new_AGEMA_signal_14107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2611 ( .C ( clk ), .D ( new_AGEMA_signal_12994 ), .Q ( new_AGEMA_signal_14111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2647 ( .C ( clk ), .D ( n2245 ), .Q ( new_AGEMA_signal_14147 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2651 ( .C ( clk ), .D ( new_AGEMA_signal_1776 ), .Q ( new_AGEMA_signal_14151 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2655 ( .C ( clk ), .D ( new_AGEMA_signal_1777 ), .Q ( new_AGEMA_signal_14155 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2659 ( .C ( clk ), .D ( new_AGEMA_signal_1778 ), .Q ( new_AGEMA_signal_14159 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2665 ( .C ( clk ), .D ( new_AGEMA_signal_14164 ), .Q ( new_AGEMA_signal_14165 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2671 ( .C ( clk ), .D ( new_AGEMA_signal_14170 ), .Q ( new_AGEMA_signal_14171 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2677 ( .C ( clk ), .D ( new_AGEMA_signal_14176 ), .Q ( new_AGEMA_signal_14177 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2683 ( .C ( clk ), .D ( new_AGEMA_signal_14182 ), .Q ( new_AGEMA_signal_14183 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2687 ( .C ( clk ), .D ( n2262 ), .Q ( new_AGEMA_signal_14187 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2691 ( .C ( clk ), .D ( new_AGEMA_signal_1389 ), .Q ( new_AGEMA_signal_14191 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2695 ( .C ( clk ), .D ( new_AGEMA_signal_1390 ), .Q ( new_AGEMA_signal_14195 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2699 ( .C ( clk ), .D ( new_AGEMA_signal_1391 ), .Q ( new_AGEMA_signal_14199 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2727 ( .C ( clk ), .D ( n2343 ), .Q ( new_AGEMA_signal_14227 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2731 ( .C ( clk ), .D ( new_AGEMA_signal_1827 ), .Q ( new_AGEMA_signal_14231 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2735 ( .C ( clk ), .D ( new_AGEMA_signal_1828 ), .Q ( new_AGEMA_signal_14235 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2739 ( .C ( clk ), .D ( new_AGEMA_signal_1829 ), .Q ( new_AGEMA_signal_14239 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2759 ( .C ( clk ), .D ( new_AGEMA_signal_12940 ), .Q ( new_AGEMA_signal_14259 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2763 ( .C ( clk ), .D ( new_AGEMA_signal_12942 ), .Q ( new_AGEMA_signal_14263 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2767 ( .C ( clk ), .D ( new_AGEMA_signal_12944 ), .Q ( new_AGEMA_signal_14267 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2771 ( .C ( clk ), .D ( new_AGEMA_signal_12946 ), .Q ( new_AGEMA_signal_14271 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2775 ( .C ( clk ), .D ( new_AGEMA_signal_12908 ), .Q ( new_AGEMA_signal_14275 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2779 ( .C ( clk ), .D ( new_AGEMA_signal_12910 ), .Q ( new_AGEMA_signal_14279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2783 ( .C ( clk ), .D ( new_AGEMA_signal_12912 ), .Q ( new_AGEMA_signal_14283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2787 ( .C ( clk ), .D ( new_AGEMA_signal_12914 ), .Q ( new_AGEMA_signal_14287 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2791 ( .C ( clk ), .D ( new_AGEMA_signal_12628 ), .Q ( new_AGEMA_signal_14291 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2795 ( .C ( clk ), .D ( new_AGEMA_signal_12630 ), .Q ( new_AGEMA_signal_14295 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2799 ( .C ( clk ), .D ( new_AGEMA_signal_12632 ), .Q ( new_AGEMA_signal_14299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2803 ( .C ( clk ), .D ( new_AGEMA_signal_12634 ), .Q ( new_AGEMA_signal_14303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2807 ( .C ( clk ), .D ( new_AGEMA_signal_12732 ), .Q ( new_AGEMA_signal_14307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2811 ( .C ( clk ), .D ( new_AGEMA_signal_12734 ), .Q ( new_AGEMA_signal_14311 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2815 ( .C ( clk ), .D ( new_AGEMA_signal_12736 ), .Q ( new_AGEMA_signal_14315 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2819 ( .C ( clk ), .D ( new_AGEMA_signal_12738 ), .Q ( new_AGEMA_signal_14319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2823 ( .C ( clk ), .D ( n2417 ), .Q ( new_AGEMA_signal_14323 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2827 ( .C ( clk ), .D ( new_AGEMA_signal_2088 ), .Q ( new_AGEMA_signal_14327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2831 ( .C ( clk ), .D ( new_AGEMA_signal_2089 ), .Q ( new_AGEMA_signal_14331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2835 ( .C ( clk ), .D ( new_AGEMA_signal_2090 ), .Q ( new_AGEMA_signal_14335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2871 ( .C ( clk ), .D ( new_AGEMA_signal_13012 ), .Q ( new_AGEMA_signal_14371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2875 ( .C ( clk ), .D ( new_AGEMA_signal_13014 ), .Q ( new_AGEMA_signal_14375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2879 ( .C ( clk ), .D ( new_AGEMA_signal_13016 ), .Q ( new_AGEMA_signal_14379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2883 ( .C ( clk ), .D ( new_AGEMA_signal_13018 ), .Q ( new_AGEMA_signal_14383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2887 ( .C ( clk ), .D ( n2483 ), .Q ( new_AGEMA_signal_14387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2891 ( .C ( clk ), .D ( new_AGEMA_signal_1437 ), .Q ( new_AGEMA_signal_14391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2895 ( .C ( clk ), .D ( new_AGEMA_signal_1438 ), .Q ( new_AGEMA_signal_14395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2899 ( .C ( clk ), .D ( new_AGEMA_signal_1439 ), .Q ( new_AGEMA_signal_14399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2975 ( .C ( clk ), .D ( n2629 ), .Q ( new_AGEMA_signal_14475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2979 ( .C ( clk ), .D ( new_AGEMA_signal_1476 ), .Q ( new_AGEMA_signal_14479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2983 ( .C ( clk ), .D ( new_AGEMA_signal_1477 ), .Q ( new_AGEMA_signal_14483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2987 ( .C ( clk ), .D ( new_AGEMA_signal_1478 ), .Q ( new_AGEMA_signal_14487 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3031 ( .C ( clk ), .D ( n2736 ), .Q ( new_AGEMA_signal_14531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3035 ( .C ( clk ), .D ( new_AGEMA_signal_1269 ), .Q ( new_AGEMA_signal_14535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3039 ( .C ( clk ), .D ( new_AGEMA_signal_1270 ), .Q ( new_AGEMA_signal_14539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3043 ( .C ( clk ), .D ( new_AGEMA_signal_1271 ), .Q ( new_AGEMA_signal_14543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3047 ( .C ( clk ), .D ( new_AGEMA_signal_12836 ), .Q ( new_AGEMA_signal_14547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3051 ( .C ( clk ), .D ( new_AGEMA_signal_12838 ), .Q ( new_AGEMA_signal_14551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3055 ( .C ( clk ), .D ( new_AGEMA_signal_12840 ), .Q ( new_AGEMA_signal_14555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3059 ( .C ( clk ), .D ( new_AGEMA_signal_12842 ), .Q ( new_AGEMA_signal_14559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3063 ( .C ( clk ), .D ( new_AGEMA_signal_12724 ), .Q ( new_AGEMA_signal_14563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3067 ( .C ( clk ), .D ( new_AGEMA_signal_12726 ), .Q ( new_AGEMA_signal_14567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3071 ( .C ( clk ), .D ( new_AGEMA_signal_12728 ), .Q ( new_AGEMA_signal_14571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3075 ( .C ( clk ), .D ( new_AGEMA_signal_12730 ), .Q ( new_AGEMA_signal_14575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3079 ( .C ( clk ), .D ( n2787 ), .Q ( new_AGEMA_signal_14579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3083 ( .C ( clk ), .D ( new_AGEMA_signal_2025 ), .Q ( new_AGEMA_signal_14583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3087 ( .C ( clk ), .D ( new_AGEMA_signal_2026 ), .Q ( new_AGEMA_signal_14587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3091 ( .C ( clk ), .D ( new_AGEMA_signal_2027 ), .Q ( new_AGEMA_signal_14591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3129 ( .C ( clk ), .D ( new_AGEMA_signal_14628 ), .Q ( new_AGEMA_signal_14629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3137 ( .C ( clk ), .D ( new_AGEMA_signal_14636 ), .Q ( new_AGEMA_signal_14637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3145 ( .C ( clk ), .D ( new_AGEMA_signal_14644 ), .Q ( new_AGEMA_signal_14645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3153 ( .C ( clk ), .D ( new_AGEMA_signal_14652 ), .Q ( new_AGEMA_signal_14653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3169 ( .C ( clk ), .D ( new_AGEMA_signal_14668 ), .Q ( new_AGEMA_signal_14669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3177 ( .C ( clk ), .D ( new_AGEMA_signal_14676 ), .Q ( new_AGEMA_signal_14677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3185 ( .C ( clk ), .D ( new_AGEMA_signal_14684 ), .Q ( new_AGEMA_signal_14685 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3193 ( .C ( clk ), .D ( new_AGEMA_signal_14692 ), .Q ( new_AGEMA_signal_14693 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3199 ( .C ( clk ), .D ( n2009 ), .Q ( new_AGEMA_signal_14699 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3205 ( .C ( clk ), .D ( new_AGEMA_signal_1602 ), .Q ( new_AGEMA_signal_14705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3211 ( .C ( clk ), .D ( new_AGEMA_signal_1603 ), .Q ( new_AGEMA_signal_14711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3217 ( .C ( clk ), .D ( new_AGEMA_signal_1604 ), .Q ( new_AGEMA_signal_14717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3239 ( .C ( clk ), .D ( n2034 ), .Q ( new_AGEMA_signal_14739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3245 ( .C ( clk ), .D ( new_AGEMA_signal_1332 ), .Q ( new_AGEMA_signal_14745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3251 ( .C ( clk ), .D ( new_AGEMA_signal_1333 ), .Q ( new_AGEMA_signal_14751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3257 ( .C ( clk ), .D ( new_AGEMA_signal_1334 ), .Q ( new_AGEMA_signal_14757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3271 ( .C ( clk ), .D ( new_AGEMA_signal_13004 ), .Q ( new_AGEMA_signal_14771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3277 ( .C ( clk ), .D ( new_AGEMA_signal_13006 ), .Q ( new_AGEMA_signal_14777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3283 ( .C ( clk ), .D ( new_AGEMA_signal_13008 ), .Q ( new_AGEMA_signal_14783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3289 ( .C ( clk ), .D ( new_AGEMA_signal_13010 ), .Q ( new_AGEMA_signal_14789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3295 ( .C ( clk ), .D ( new_AGEMA_signal_13060 ), .Q ( new_AGEMA_signal_14795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3301 ( .C ( clk ), .D ( new_AGEMA_signal_13062 ), .Q ( new_AGEMA_signal_14801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3307 ( .C ( clk ), .D ( new_AGEMA_signal_13064 ), .Q ( new_AGEMA_signal_14807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3313 ( .C ( clk ), .D ( new_AGEMA_signal_13066 ), .Q ( new_AGEMA_signal_14813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3343 ( .C ( clk ), .D ( new_AGEMA_signal_12556 ), .Q ( new_AGEMA_signal_14843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3349 ( .C ( clk ), .D ( new_AGEMA_signal_12558 ), .Q ( new_AGEMA_signal_14849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3355 ( .C ( clk ), .D ( new_AGEMA_signal_12560 ), .Q ( new_AGEMA_signal_14855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3361 ( .C ( clk ), .D ( new_AGEMA_signal_12562 ), .Q ( new_AGEMA_signal_14861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3367 ( .C ( clk ), .D ( n2122 ), .Q ( new_AGEMA_signal_14867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3373 ( .C ( clk ), .D ( new_AGEMA_signal_1695 ), .Q ( new_AGEMA_signal_14873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3379 ( .C ( clk ), .D ( new_AGEMA_signal_1696 ), .Q ( new_AGEMA_signal_14879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3385 ( .C ( clk ), .D ( new_AGEMA_signal_1697 ), .Q ( new_AGEMA_signal_14885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3399 ( .C ( clk ), .D ( n2220 ), .Q ( new_AGEMA_signal_14899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3405 ( .C ( clk ), .D ( new_AGEMA_signal_1713 ), .Q ( new_AGEMA_signal_14905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3411 ( .C ( clk ), .D ( new_AGEMA_signal_1714 ), .Q ( new_AGEMA_signal_14911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3417 ( .C ( clk ), .D ( new_AGEMA_signal_1715 ), .Q ( new_AGEMA_signal_14917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3473 ( .C ( clk ), .D ( new_AGEMA_signal_14972 ), .Q ( new_AGEMA_signal_14973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3481 ( .C ( clk ), .D ( new_AGEMA_signal_14980 ), .Q ( new_AGEMA_signal_14981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3489 ( .C ( clk ), .D ( new_AGEMA_signal_14988 ), .Q ( new_AGEMA_signal_14989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3497 ( .C ( clk ), .D ( new_AGEMA_signal_14996 ), .Q ( new_AGEMA_signal_14997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3503 ( .C ( clk ), .D ( new_AGEMA_signal_12756 ), .Q ( new_AGEMA_signal_15003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3509 ( .C ( clk ), .D ( new_AGEMA_signal_12758 ), .Q ( new_AGEMA_signal_15009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3515 ( .C ( clk ), .D ( new_AGEMA_signal_12760 ), .Q ( new_AGEMA_signal_15015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3521 ( .C ( clk ), .D ( new_AGEMA_signal_12762 ), .Q ( new_AGEMA_signal_15021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3615 ( .C ( clk ), .D ( n2344 ), .Q ( new_AGEMA_signal_15115 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3621 ( .C ( clk ), .D ( new_AGEMA_signal_1833 ), .Q ( new_AGEMA_signal_15121 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3627 ( .C ( clk ), .D ( new_AGEMA_signal_1834 ), .Q ( new_AGEMA_signal_15127 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3633 ( .C ( clk ), .D ( new_AGEMA_signal_1835 ), .Q ( new_AGEMA_signal_15133 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3743 ( .C ( clk ), .D ( n2468 ), .Q ( new_AGEMA_signal_15243 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3749 ( .C ( clk ), .D ( new_AGEMA_signal_1446 ), .Q ( new_AGEMA_signal_15249 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3755 ( .C ( clk ), .D ( new_AGEMA_signal_1447 ), .Q ( new_AGEMA_signal_15255 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3761 ( .C ( clk ), .D ( new_AGEMA_signal_1448 ), .Q ( new_AGEMA_signal_15261 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3767 ( .C ( clk ), .D ( n2761 ), .Q ( new_AGEMA_signal_15267 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3773 ( .C ( clk ), .D ( new_AGEMA_signal_1548 ), .Q ( new_AGEMA_signal_15273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3779 ( .C ( clk ), .D ( new_AGEMA_signal_1549 ), .Q ( new_AGEMA_signal_15279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3785 ( .C ( clk ), .D ( new_AGEMA_signal_1550 ), .Q ( new_AGEMA_signal_15285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3817 ( .C ( clk ), .D ( new_AGEMA_signal_15316 ), .Q ( new_AGEMA_signal_15317 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3825 ( .C ( clk ), .D ( new_AGEMA_signal_15324 ), .Q ( new_AGEMA_signal_15325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3833 ( .C ( clk ), .D ( new_AGEMA_signal_15332 ), .Q ( new_AGEMA_signal_15333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3841 ( .C ( clk ), .D ( new_AGEMA_signal_15340 ), .Q ( new_AGEMA_signal_15341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3937 ( .C ( clk ), .D ( new_AGEMA_signal_15436 ), .Q ( new_AGEMA_signal_15437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3945 ( .C ( clk ), .D ( new_AGEMA_signal_15444 ), .Q ( new_AGEMA_signal_15445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3953 ( .C ( clk ), .D ( new_AGEMA_signal_15452 ), .Q ( new_AGEMA_signal_15453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3961 ( .C ( clk ), .D ( new_AGEMA_signal_15460 ), .Q ( new_AGEMA_signal_15461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3999 ( .C ( clk ), .D ( n2825 ), .Q ( new_AGEMA_signal_15499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4005 ( .C ( clk ), .D ( new_AGEMA_signal_2040 ), .Q ( new_AGEMA_signal_15505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4011 ( .C ( clk ), .D ( new_AGEMA_signal_2041 ), .Q ( new_AGEMA_signal_15511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4017 ( .C ( clk ), .D ( new_AGEMA_signal_2042 ), .Q ( new_AGEMA_signal_15517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4031 ( .C ( clk ), .D ( n1957 ), .Q ( new_AGEMA_signal_15531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4039 ( .C ( clk ), .D ( new_AGEMA_signal_1263 ), .Q ( new_AGEMA_signal_15539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4047 ( .C ( clk ), .D ( new_AGEMA_signal_1264 ), .Q ( new_AGEMA_signal_15547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4055 ( .C ( clk ), .D ( new_AGEMA_signal_1265 ), .Q ( new_AGEMA_signal_15555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4087 ( .C ( clk ), .D ( n2026 ), .Q ( new_AGEMA_signal_15587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4095 ( .C ( clk ), .D ( new_AGEMA_signal_1323 ), .Q ( new_AGEMA_signal_15595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4103 ( .C ( clk ), .D ( new_AGEMA_signal_1324 ), .Q ( new_AGEMA_signal_15603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4111 ( .C ( clk ), .D ( new_AGEMA_signal_1325 ), .Q ( new_AGEMA_signal_15611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4167 ( .C ( clk ), .D ( n2811 ), .Q ( new_AGEMA_signal_15667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4175 ( .C ( clk ), .D ( new_AGEMA_signal_1698 ), .Q ( new_AGEMA_signal_15675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4183 ( .C ( clk ), .D ( new_AGEMA_signal_1699 ), .Q ( new_AGEMA_signal_15683 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4191 ( .C ( clk ), .D ( new_AGEMA_signal_1700 ), .Q ( new_AGEMA_signal_15691 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4351 ( .C ( clk ), .D ( new_AGEMA_signal_13084 ), .Q ( new_AGEMA_signal_15851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4359 ( .C ( clk ), .D ( new_AGEMA_signal_13086 ), .Q ( new_AGEMA_signal_15859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4367 ( .C ( clk ), .D ( new_AGEMA_signal_13088 ), .Q ( new_AGEMA_signal_15867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4375 ( .C ( clk ), .D ( new_AGEMA_signal_13090 ), .Q ( new_AGEMA_signal_15875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4423 ( .C ( clk ), .D ( n2363 ), .Q ( new_AGEMA_signal_15923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4431 ( .C ( clk ), .D ( new_AGEMA_signal_1422 ), .Q ( new_AGEMA_signal_15931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4439 ( .C ( clk ), .D ( new_AGEMA_signal_1423 ), .Q ( new_AGEMA_signal_15939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4447 ( .C ( clk ), .D ( new_AGEMA_signal_1424 ), .Q ( new_AGEMA_signal_15947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4551 ( .C ( clk ), .D ( new_AGEMA_signal_12996 ), .Q ( new_AGEMA_signal_16051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4559 ( .C ( clk ), .D ( new_AGEMA_signal_12998 ), .Q ( new_AGEMA_signal_16059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4567 ( .C ( clk ), .D ( new_AGEMA_signal_13000 ), .Q ( new_AGEMA_signal_16067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4575 ( .C ( clk ), .D ( new_AGEMA_signal_13002 ), .Q ( new_AGEMA_signal_16075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4583 ( .C ( clk ), .D ( new_AGEMA_signal_12596 ), .Q ( new_AGEMA_signal_16083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4591 ( .C ( clk ), .D ( new_AGEMA_signal_12598 ), .Q ( new_AGEMA_signal_16091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4599 ( .C ( clk ), .D ( new_AGEMA_signal_12600 ), .Q ( new_AGEMA_signal_16099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4607 ( .C ( clk ), .D ( new_AGEMA_signal_12602 ), .Q ( new_AGEMA_signal_16107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4927 ( .C ( clk ), .D ( n2544 ), .Q ( new_AGEMA_signal_16427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4937 ( .C ( clk ), .D ( new_AGEMA_signal_1353 ), .Q ( new_AGEMA_signal_16437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4947 ( .C ( clk ), .D ( new_AGEMA_signal_1354 ), .Q ( new_AGEMA_signal_16447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4957 ( .C ( clk ), .D ( new_AGEMA_signal_1355 ), .Q ( new_AGEMA_signal_16457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5127 ( .C ( clk ), .D ( n2364 ), .Q ( new_AGEMA_signal_16627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5137 ( .C ( clk ), .D ( new_AGEMA_signal_1851 ), .Q ( new_AGEMA_signal_16637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5147 ( .C ( clk ), .D ( new_AGEMA_signal_1852 ), .Q ( new_AGEMA_signal_16647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5157 ( .C ( clk ), .D ( new_AGEMA_signal_1853 ), .Q ( new_AGEMA_signal_16657 ) ) ;

    /* cells in depth 6 */
    nor_HPC1 #(.security_order(3), .pipeline(1)) U1960 ( .ina ({new_AGEMA_signal_1499, new_AGEMA_signal_1498, new_AGEMA_signal_1497, n2575}), .inb ({new_AGEMA_signal_1502, new_AGEMA_signal_1501, new_AGEMA_signal_1500, n1962}), .clk ( clk ), .rnd ({Fresh[2389], Fresh[2388], Fresh[2387], Fresh[2386], Fresh[2385], Fresh[2384], Fresh[2383], Fresh[2382], Fresh[2381], Fresh[2380]}), .outt ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, new_AGEMA_signal_2043, n1924}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U1967 ( .ina ({new_AGEMA_signal_1505, new_AGEMA_signal_1504, new_AGEMA_signal_1503, n1922}), .inb ({new_AGEMA_signal_12554, new_AGEMA_signal_12552, new_AGEMA_signal_12550, new_AGEMA_signal_12548}), .clk ( clk ), .rnd ({Fresh[2399], Fresh[2398], Fresh[2397], Fresh[2396], Fresh[2395], Fresh[2394], Fresh[2393], Fresh[2392], Fresh[2391], Fresh[2390]}), .outt ({new_AGEMA_signal_2048, new_AGEMA_signal_2047, new_AGEMA_signal_2046, n1923}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U1981 ( .ina ({new_AGEMA_signal_1508, new_AGEMA_signal_1507, new_AGEMA_signal_1506, n1926}), .inb ({new_AGEMA_signal_1511, new_AGEMA_signal_1510, new_AGEMA_signal_1509, n1925}), .clk ( clk ), .rnd ({Fresh[2409], Fresh[2408], Fresh[2407], Fresh[2406], Fresh[2405], Fresh[2404], Fresh[2403], Fresh[2402], Fresh[2401], Fresh[2400]}), .outt ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, new_AGEMA_signal_2049, n1927}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U1993 ( .ina ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, new_AGEMA_signal_1515, n2734}), .inb ({new_AGEMA_signal_1520, new_AGEMA_signal_1519, new_AGEMA_signal_1518, n2763}), .clk ( clk ), .rnd ({Fresh[2419], Fresh[2418], Fresh[2417], Fresh[2416], Fresh[2415], Fresh[2414], Fresh[2413], Fresh[2412], Fresh[2411], Fresh[2410]}), .outt ({new_AGEMA_signal_2054, new_AGEMA_signal_2053, new_AGEMA_signal_2052, n1929}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2007 ( .ina ({new_AGEMA_signal_12562, new_AGEMA_signal_12560, new_AGEMA_signal_12558, new_AGEMA_signal_12556}), .inb ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, new_AGEMA_signal_1521, n2732}), .clk ( clk ), .rnd ({Fresh[2429], Fresh[2428], Fresh[2427], Fresh[2426], Fresh[2425], Fresh[2424], Fresh[2423], Fresh[2422], Fresh[2421], Fresh[2420]}), .outt ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, new_AGEMA_signal_2055, n2665}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2011 ( .ina ({new_AGEMA_signal_12570, new_AGEMA_signal_12568, new_AGEMA_signal_12566, new_AGEMA_signal_12564}), .inb ({new_AGEMA_signal_1526, new_AGEMA_signal_1525, new_AGEMA_signal_1524, n1937}), .clk ( clk ), .rnd ({Fresh[2439], Fresh[2438], Fresh[2437], Fresh[2436], Fresh[2435], Fresh[2434], Fresh[2433], Fresh[2432], Fresh[2431], Fresh[2430]}), .outt ({new_AGEMA_signal_2060, new_AGEMA_signal_2059, new_AGEMA_signal_2058, n1938}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2019 ( .ina ({new_AGEMA_signal_12578, new_AGEMA_signal_12576, new_AGEMA_signal_12574, new_AGEMA_signal_12572}), .inb ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, new_AGEMA_signal_1521, n2732}), .clk ( clk ), .rnd ({Fresh[2449], Fresh[2448], Fresh[2447], Fresh[2446], Fresh[2445], Fresh[2444], Fresh[2443], Fresh[2442], Fresh[2441], Fresh[2440]}), .outt ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, new_AGEMA_signal_2061, n2235}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2023 ( .ina ({new_AGEMA_signal_12586, new_AGEMA_signal_12584, new_AGEMA_signal_12582, new_AGEMA_signal_12580}), .inb ({new_AGEMA_signal_1244, new_AGEMA_signal_1243, new_AGEMA_signal_1242, n1942}), .clk ( clk ), .rnd ({Fresh[2459], Fresh[2458], Fresh[2457], Fresh[2456], Fresh[2455], Fresh[2454], Fresh[2453], Fresh[2452], Fresh[2451], Fresh[2450]}), .outt ({new_AGEMA_signal_1529, new_AGEMA_signal_1528, new_AGEMA_signal_1527, n1943}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2027 ( .ina ({new_AGEMA_signal_1247, new_AGEMA_signal_1246, new_AGEMA_signal_1245, n2676}), .inb ({new_AGEMA_signal_12594, new_AGEMA_signal_12592, new_AGEMA_signal_12590, new_AGEMA_signal_12588}), .clk ( clk ), .rnd ({Fresh[2469], Fresh[2468], Fresh[2467], Fresh[2466], Fresh[2465], Fresh[2464], Fresh[2463], Fresh[2462], Fresh[2461], Fresh[2460]}), .outt ({new_AGEMA_signal_1532, new_AGEMA_signal_1531, new_AGEMA_signal_1530, n1946}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2031 ( .ina ({new_AGEMA_signal_12602, new_AGEMA_signal_12600, new_AGEMA_signal_12598, new_AGEMA_signal_12596}), .inb ({new_AGEMA_signal_1535, new_AGEMA_signal_1534, new_AGEMA_signal_1533, n1944}), .clk ( clk ), .rnd ({Fresh[2479], Fresh[2478], Fresh[2477], Fresh[2476], Fresh[2475], Fresh[2474], Fresh[2473], Fresh[2472], Fresh[2471], Fresh[2470]}), .outt ({new_AGEMA_signal_2066, new_AGEMA_signal_2065, new_AGEMA_signal_2064, n1945}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2034 ( .ina ({new_AGEMA_signal_12610, new_AGEMA_signal_12608, new_AGEMA_signal_12606, new_AGEMA_signal_12604}), .inb ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, new_AGEMA_signal_1515, n2734}), .clk ( clk ), .rnd ({Fresh[2489], Fresh[2488], Fresh[2487], Fresh[2486], Fresh[2485], Fresh[2484], Fresh[2483], Fresh[2482], Fresh[2481], Fresh[2480]}), .outt ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, new_AGEMA_signal_2067, n1956}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2040 ( .ina ({new_AGEMA_signal_1538, new_AGEMA_signal_1537, new_AGEMA_signal_1536, n1950}), .inb ({new_AGEMA_signal_1256, new_AGEMA_signal_1255, new_AGEMA_signal_1254, n1949}), .clk ( clk ), .rnd ({Fresh[2499], Fresh[2498], Fresh[2497], Fresh[2496], Fresh[2495], Fresh[2494], Fresh[2493], Fresh[2492], Fresh[2491], Fresh[2490]}), .outt ({new_AGEMA_signal_2072, new_AGEMA_signal_2071, new_AGEMA_signal_2070, n1951}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2048 ( .ina ({new_AGEMA_signal_1541, new_AGEMA_signal_1540, new_AGEMA_signal_1539, n2662}), .inb ({new_AGEMA_signal_1262, new_AGEMA_signal_1261, new_AGEMA_signal_1260, n2627}), .clk ( clk ), .rnd ({Fresh[2509], Fresh[2508], Fresh[2507], Fresh[2506], Fresh[2505], Fresh[2504], Fresh[2503], Fresh[2502], Fresh[2501], Fresh[2500]}), .outt ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, new_AGEMA_signal_2073, n1952}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2057 ( .ina ({new_AGEMA_signal_12618, new_AGEMA_signal_12616, new_AGEMA_signal_12614, new_AGEMA_signal_12612}), .inb ({new_AGEMA_signal_1544, new_AGEMA_signal_1543, new_AGEMA_signal_1542, n2088}), .clk ( clk ), .rnd ({Fresh[2519], Fresh[2518], Fresh[2517], Fresh[2516], Fresh[2515], Fresh[2514], Fresh[2513], Fresh[2512], Fresh[2511], Fresh[2510]}), .outt ({new_AGEMA_signal_2078, new_AGEMA_signal_2077, new_AGEMA_signal_2076, n2687}) ) ;
    or_HPC1 #(.security_order(3), .pipeline(1)) U2061 ( .ina ({new_AGEMA_signal_1502, new_AGEMA_signal_1501, new_AGEMA_signal_1500, n1962}), .inb ({new_AGEMA_signal_12626, new_AGEMA_signal_12624, new_AGEMA_signal_12622, new_AGEMA_signal_12620}), .clk ( clk ), .rnd ({Fresh[2529], Fresh[2528], Fresh[2527], Fresh[2526], Fresh[2525], Fresh[2524], Fresh[2523], Fresh[2522], Fresh[2521], Fresh[2520]}), .outt ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, new_AGEMA_signal_2079, n1966}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2064 ( .ina ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, new_AGEMA_signal_1269, n2736}), .inb ({new_AGEMA_signal_12634, new_AGEMA_signal_12632, new_AGEMA_signal_12630, new_AGEMA_signal_12628}), .clk ( clk ), .rnd ({Fresh[2539], Fresh[2538], Fresh[2537], Fresh[2536], Fresh[2535], Fresh[2534], Fresh[2533], Fresh[2532], Fresh[2531], Fresh[2530]}), .outt ({new_AGEMA_signal_1547, new_AGEMA_signal_1546, new_AGEMA_signal_1545, n1963}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2077 ( .ina ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, new_AGEMA_signal_2085, n2720}), .inb ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, new_AGEMA_signal_2088, n2417}), .clk ( clk ), .rnd ({Fresh[2549], Fresh[2548], Fresh[2547], Fresh[2546], Fresh[2545], Fresh[2544], Fresh[2543], Fresh[2542], Fresh[2541], Fresh[2540]}), .outt ({new_AGEMA_signal_2558, new_AGEMA_signal_2557, new_AGEMA_signal_2556, n1968}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2082 ( .ina ({new_AGEMA_signal_1556, new_AGEMA_signal_1555, new_AGEMA_signal_1554, n2505}), .inb ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}), .clk ( clk ), .rnd ({Fresh[2559], Fresh[2558], Fresh[2557], Fresh[2556], Fresh[2555], Fresh[2554], Fresh[2553], Fresh[2552], Fresh[2551], Fresh[2550]}), .outt ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, new_AGEMA_signal_2091, n2684}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2088 ( .ina ({new_AGEMA_signal_12642, new_AGEMA_signal_12640, new_AGEMA_signal_12638, new_AGEMA_signal_12636}), .inb ({new_AGEMA_signal_1562, new_AGEMA_signal_1561, new_AGEMA_signal_1560, n2625}), .clk ( clk ), .rnd ({Fresh[2569], Fresh[2568], Fresh[2567], Fresh[2566], Fresh[2565], Fresh[2564], Fresh[2563], Fresh[2562], Fresh[2561], Fresh[2560]}), .outt ({new_AGEMA_signal_2096, new_AGEMA_signal_2095, new_AGEMA_signal_2094, n1972}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2092 ( .ina ({new_AGEMA_signal_12650, new_AGEMA_signal_12648, new_AGEMA_signal_12646, new_AGEMA_signal_12644}), .inb ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, new_AGEMA_signal_1293, n2190}), .clk ( clk ), .rnd ({Fresh[2579], Fresh[2578], Fresh[2577], Fresh[2576], Fresh[2575], Fresh[2574], Fresh[2573], Fresh[2572], Fresh[2571], Fresh[2570]}), .outt ({new_AGEMA_signal_1565, new_AGEMA_signal_1564, new_AGEMA_signal_1563, n1971}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2099 ( .ina ({new_AGEMA_signal_12658, new_AGEMA_signal_12656, new_AGEMA_signal_12654, new_AGEMA_signal_12652}), .inb ({new_AGEMA_signal_1568, new_AGEMA_signal_1567, new_AGEMA_signal_1566, n2535}), .clk ( clk ), .rnd ({Fresh[2589], Fresh[2588], Fresh[2587], Fresh[2586], Fresh[2585], Fresh[2584], Fresh[2583], Fresh[2582], Fresh[2581], Fresh[2580]}), .outt ({new_AGEMA_signal_2099, new_AGEMA_signal_2098, new_AGEMA_signal_2097, n1974}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2106 ( .ina ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, new_AGEMA_signal_1521, n2732}), .inb ({new_AGEMA_signal_12618, new_AGEMA_signal_12616, new_AGEMA_signal_12614, new_AGEMA_signal_12612}), .clk ( clk ), .rnd ({Fresh[2599], Fresh[2598], Fresh[2597], Fresh[2596], Fresh[2595], Fresh[2594], Fresh[2593], Fresh[2592], Fresh[2591], Fresh[2590]}), .outt ({new_AGEMA_signal_2102, new_AGEMA_signal_2101, new_AGEMA_signal_2100, n1979}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2112 ( .ina ({new_AGEMA_signal_12666, new_AGEMA_signal_12664, new_AGEMA_signal_12662, new_AGEMA_signal_12660}), .inb ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, new_AGEMA_signal_1302, n2817}), .clk ( clk ), .rnd ({Fresh[2609], Fresh[2608], Fresh[2607], Fresh[2606], Fresh[2605], Fresh[2604], Fresh[2603], Fresh[2602], Fresh[2601], Fresh[2600]}), .outt ({new_AGEMA_signal_1574, new_AGEMA_signal_1573, new_AGEMA_signal_1572, n1985}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2121 ( .ina ({new_AGEMA_signal_1580, new_AGEMA_signal_1579, new_AGEMA_signal_1578, n1992}), .inb ({new_AGEMA_signal_1583, new_AGEMA_signal_1582, new_AGEMA_signal_1581, n1991}), .clk ( clk ), .rnd ({Fresh[2619], Fresh[2618], Fresh[2617], Fresh[2616], Fresh[2615], Fresh[2614], Fresh[2613], Fresh[2612], Fresh[2611], Fresh[2610]}), .outt ({new_AGEMA_signal_2108, new_AGEMA_signal_2107, new_AGEMA_signal_2106, n1994}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2126 ( .ina ({new_AGEMA_signal_12674, new_AGEMA_signal_12672, new_AGEMA_signal_12670, new_AGEMA_signal_12668}), .inb ({new_AGEMA_signal_1586, new_AGEMA_signal_1585, new_AGEMA_signal_1584, n1995}), .clk ( clk ), .rnd ({Fresh[2629], Fresh[2628], Fresh[2627], Fresh[2626], Fresh[2625], Fresh[2624], Fresh[2623], Fresh[2622], Fresh[2621], Fresh[2620]}), .outt ({new_AGEMA_signal_2111, new_AGEMA_signal_2110, new_AGEMA_signal_2109, n1996}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2136 ( .ina ({new_AGEMA_signal_12682, new_AGEMA_signal_12680, new_AGEMA_signal_12678, new_AGEMA_signal_12676}), .inb ({new_AGEMA_signal_1592, new_AGEMA_signal_1591, new_AGEMA_signal_1590, n2003}), .clk ( clk ), .rnd ({Fresh[2639], Fresh[2638], Fresh[2637], Fresh[2636], Fresh[2635], Fresh[2634], Fresh[2633], Fresh[2632], Fresh[2631], Fresh[2630]}), .outt ({new_AGEMA_signal_2114, new_AGEMA_signal_2113, new_AGEMA_signal_2112, n2137}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2142 ( .ina ({new_AGEMA_signal_12690, new_AGEMA_signal_12688, new_AGEMA_signal_12686, new_AGEMA_signal_12684}), .inb ({new_AGEMA_signal_1598, new_AGEMA_signal_1597, new_AGEMA_signal_1596, n2572}), .clk ( clk ), .rnd ({Fresh[2649], Fresh[2648], Fresh[2647], Fresh[2646], Fresh[2645], Fresh[2644], Fresh[2643], Fresh[2642], Fresh[2641], Fresh[2640]}), .outt ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, new_AGEMA_signal_2115, n2006}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2144 ( .ina ({new_AGEMA_signal_12698, new_AGEMA_signal_12696, new_AGEMA_signal_12694, new_AGEMA_signal_12692}), .inb ({new_AGEMA_signal_1601, new_AGEMA_signal_1600, new_AGEMA_signal_1599, n2004}), .clk ( clk ), .rnd ({Fresh[2659], Fresh[2658], Fresh[2657], Fresh[2656], Fresh[2655], Fresh[2654], Fresh[2653], Fresh[2652], Fresh[2651], Fresh[2650]}), .outt ({new_AGEMA_signal_2120, new_AGEMA_signal_2119, new_AGEMA_signal_2118, n2005}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2152 ( .ina ({new_AGEMA_signal_12706, new_AGEMA_signal_12704, new_AGEMA_signal_12702, new_AGEMA_signal_12700}), .inb ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, new_AGEMA_signal_1605, n2533}), .clk ( clk ), .rnd ({Fresh[2669], Fresh[2668], Fresh[2667], Fresh[2666], Fresh[2665], Fresh[2664], Fresh[2663], Fresh[2662], Fresh[2661], Fresh[2660]}), .outt ({new_AGEMA_signal_2123, new_AGEMA_signal_2122, new_AGEMA_signal_2121, n2013}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2160 ( .ina ({new_AGEMA_signal_12714, new_AGEMA_signal_12712, new_AGEMA_signal_12710, new_AGEMA_signal_12708}), .inb ({new_AGEMA_signal_1328, new_AGEMA_signal_1327, new_AGEMA_signal_1326, n2227}), .clk ( clk ), .rnd ({Fresh[2679], Fresh[2678], Fresh[2677], Fresh[2676], Fresh[2675], Fresh[2674], Fresh[2673], Fresh[2672], Fresh[2671], Fresh[2670]}), .outt ({new_AGEMA_signal_1613, new_AGEMA_signal_1612, new_AGEMA_signal_1611, n2020}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2164 ( .ina ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, new_AGEMA_signal_1302, n2817}), .inb ({new_AGEMA_signal_12722, new_AGEMA_signal_12720, new_AGEMA_signal_12718, new_AGEMA_signal_12716}), .clk ( clk ), .rnd ({Fresh[2689], Fresh[2688], Fresh[2687], Fresh[2686], Fresh[2685], Fresh[2684], Fresh[2683], Fresh[2682], Fresh[2681], Fresh[2680]}), .outt ({new_AGEMA_signal_1616, new_AGEMA_signal_1615, new_AGEMA_signal_1614, n2023}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2168 ( .ina ({new_AGEMA_signal_1145, new_AGEMA_signal_1144, new_AGEMA_signal_1143, n2027}), .inb ({new_AGEMA_signal_12730, new_AGEMA_signal_12728, new_AGEMA_signal_12726, new_AGEMA_signal_12724}), .clk ( clk ), .rnd ({Fresh[2699], Fresh[2698], Fresh[2697], Fresh[2696], Fresh[2695], Fresh[2694], Fresh[2693], Fresh[2692], Fresh[2691], Fresh[2690]}), .outt ({new_AGEMA_signal_1331, new_AGEMA_signal_1330, new_AGEMA_signal_1329, n2028}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2172 ( .ina ({new_AGEMA_signal_1619, new_AGEMA_signal_1618, new_AGEMA_signal_1617, n2214}), .inb ({new_AGEMA_signal_12738, new_AGEMA_signal_12736, new_AGEMA_signal_12734, new_AGEMA_signal_12732}), .clk ( clk ), .rnd ({Fresh[2709], Fresh[2708], Fresh[2707], Fresh[2706], Fresh[2705], Fresh[2704], Fresh[2703], Fresh[2702], Fresh[2701], Fresh[2700]}), .outt ({new_AGEMA_signal_2129, new_AGEMA_signal_2128, new_AGEMA_signal_2127, n2033}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2175 ( .ina ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, new_AGEMA_signal_1623, n2376}), .inb ({new_AGEMA_signal_12746, new_AGEMA_signal_12744, new_AGEMA_signal_12742, new_AGEMA_signal_12740}), .clk ( clk ), .rnd ({Fresh[2719], Fresh[2718], Fresh[2717], Fresh[2716], Fresh[2715], Fresh[2714], Fresh[2713], Fresh[2712], Fresh[2711], Fresh[2710]}), .outt ({new_AGEMA_signal_2132, new_AGEMA_signal_2131, new_AGEMA_signal_2130, n2031}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2184 ( .ina ({new_AGEMA_signal_1262, new_AGEMA_signal_1261, new_AGEMA_signal_1260, n2627}), .inb ({new_AGEMA_signal_1628, new_AGEMA_signal_1627, new_AGEMA_signal_1626, n2039}), .clk ( clk ), .rnd ({Fresh[2729], Fresh[2728], Fresh[2727], Fresh[2726], Fresh[2725], Fresh[2724], Fresh[2723], Fresh[2722], Fresh[2721], Fresh[2720]}), .outt ({new_AGEMA_signal_2135, new_AGEMA_signal_2134, new_AGEMA_signal_2133, n2040}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2187 ( .ina ({new_AGEMA_signal_12754, new_AGEMA_signal_12752, new_AGEMA_signal_12750, new_AGEMA_signal_12748}), .inb ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}), .clk ( clk ), .rnd ({Fresh[2739], Fresh[2738], Fresh[2737], Fresh[2736], Fresh[2735], Fresh[2734], Fresh[2733], Fresh[2732], Fresh[2731], Fresh[2730]}), .outt ({new_AGEMA_signal_1631, new_AGEMA_signal_1630, new_AGEMA_signal_1629, n2050}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2193 ( .ina ({new_AGEMA_signal_12762, new_AGEMA_signal_12760, new_AGEMA_signal_12758, new_AGEMA_signal_12756}), .inb ({new_AGEMA_signal_1640, new_AGEMA_signal_1639, new_AGEMA_signal_1638, n2044}), .clk ( clk ), .rnd ({Fresh[2749], Fresh[2748], Fresh[2747], Fresh[2746], Fresh[2745], Fresh[2744], Fresh[2743], Fresh[2742], Fresh[2741], Fresh[2740]}), .outt ({new_AGEMA_signal_2138, new_AGEMA_signal_2137, new_AGEMA_signal_2136, n2045}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2199 ( .ina ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, new_AGEMA_signal_1641, n2654}), .inb ({new_AGEMA_signal_12618, new_AGEMA_signal_12616, new_AGEMA_signal_12614, new_AGEMA_signal_12612}), .clk ( clk ), .rnd ({Fresh[2759], Fresh[2758], Fresh[2757], Fresh[2756], Fresh[2755], Fresh[2754], Fresh[2753], Fresh[2752], Fresh[2751], Fresh[2750]}), .outt ({new_AGEMA_signal_2141, new_AGEMA_signal_2140, new_AGEMA_signal_2139, n2051}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2203 ( .ina ({new_AGEMA_signal_12770, new_AGEMA_signal_12768, new_AGEMA_signal_12766, new_AGEMA_signal_12764}), .inb ({new_AGEMA_signal_1646, new_AGEMA_signal_1645, new_AGEMA_signal_1644, n2055}), .clk ( clk ), .rnd ({Fresh[2769], Fresh[2768], Fresh[2767], Fresh[2766], Fresh[2765], Fresh[2764], Fresh[2763], Fresh[2762], Fresh[2761], Fresh[2760]}), .outt ({new_AGEMA_signal_2144, new_AGEMA_signal_2143, new_AGEMA_signal_2142, n2056}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2209 ( .ina ({new_AGEMA_signal_1652, new_AGEMA_signal_1651, new_AGEMA_signal_1650, n2407}), .inb ({new_AGEMA_signal_12778, new_AGEMA_signal_12776, new_AGEMA_signal_12774, new_AGEMA_signal_12772}), .clk ( clk ), .rnd ({Fresh[2779], Fresh[2778], Fresh[2777], Fresh[2776], Fresh[2775], Fresh[2774], Fresh[2773], Fresh[2772], Fresh[2771], Fresh[2770]}), .outt ({new_AGEMA_signal_2147, new_AGEMA_signal_2146, new_AGEMA_signal_2145, n2060}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2215 ( .ina ({new_AGEMA_signal_12786, new_AGEMA_signal_12784, new_AGEMA_signal_12782, new_AGEMA_signal_12780}), .inb ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, new_AGEMA_signal_1641, n2654}), .clk ( clk ), .rnd ({Fresh[2789], Fresh[2788], Fresh[2787], Fresh[2786], Fresh[2785], Fresh[2784], Fresh[2783], Fresh[2782], Fresh[2781], Fresh[2780]}), .outt ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, new_AGEMA_signal_2148, n2066}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2217 ( .ina ({new_AGEMA_signal_12730, new_AGEMA_signal_12728, new_AGEMA_signal_12726, new_AGEMA_signal_12724}), .inb ({new_AGEMA_signal_1658, new_AGEMA_signal_1657, new_AGEMA_signal_1656, n2731}), .clk ( clk ), .rnd ({Fresh[2799], Fresh[2798], Fresh[2797], Fresh[2796], Fresh[2795], Fresh[2794], Fresh[2793], Fresh[2792], Fresh[2791], Fresh[2790]}), .outt ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, new_AGEMA_signal_2151, n2065}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2221 ( .ina ({new_AGEMA_signal_1661, new_AGEMA_signal_1660, new_AGEMA_signal_1659, n2068}), .inb ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, new_AGEMA_signal_1302, n2817}), .clk ( clk ), .rnd ({Fresh[2809], Fresh[2808], Fresh[2807], Fresh[2806], Fresh[2805], Fresh[2804], Fresh[2803], Fresh[2802], Fresh[2801], Fresh[2800]}), .outt ({new_AGEMA_signal_2156, new_AGEMA_signal_2155, new_AGEMA_signal_2154, n2069}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2226 ( .ina ({new_AGEMA_signal_12794, new_AGEMA_signal_12792, new_AGEMA_signal_12790, new_AGEMA_signal_12788}), .inb ({new_AGEMA_signal_1664, new_AGEMA_signal_1663, new_AGEMA_signal_1662, n2252}), .clk ( clk ), .rnd ({Fresh[2819], Fresh[2818], Fresh[2817], Fresh[2816], Fresh[2815], Fresh[2814], Fresh[2813], Fresh[2812], Fresh[2811], Fresh[2810]}), .outt ({new_AGEMA_signal_2159, new_AGEMA_signal_2158, new_AGEMA_signal_2157, n2074}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2235 ( .ina ({new_AGEMA_signal_1346, new_AGEMA_signal_1345, new_AGEMA_signal_1344, n2081}), .inb ({new_AGEMA_signal_1667, new_AGEMA_signal_1666, new_AGEMA_signal_1665, n2080}), .clk ( clk ), .rnd ({Fresh[2829], Fresh[2828], Fresh[2827], Fresh[2826], Fresh[2825], Fresh[2824], Fresh[2823], Fresh[2822], Fresh[2821], Fresh[2820]}), .outt ({new_AGEMA_signal_2162, new_AGEMA_signal_2161, new_AGEMA_signal_2160, n2082}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2240 ( .ina ({new_AGEMA_signal_12698, new_AGEMA_signal_12696, new_AGEMA_signal_12694, new_AGEMA_signal_12692}), .inb ({new_AGEMA_signal_1673, new_AGEMA_signal_1672, new_AGEMA_signal_1671, n2083}), .clk ( clk ), .rnd ({Fresh[2839], Fresh[2838], Fresh[2837], Fresh[2836], Fresh[2835], Fresh[2834], Fresh[2833], Fresh[2832], Fresh[2831], Fresh[2830]}), .outt ({new_AGEMA_signal_2165, new_AGEMA_signal_2164, new_AGEMA_signal_2163, n2084}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2242 ( .ina ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, new_AGEMA_signal_1605, n2533}), .inb ({new_AGEMA_signal_12562, new_AGEMA_signal_12560, new_AGEMA_signal_12558, new_AGEMA_signal_12556}), .clk ( clk ), .rnd ({Fresh[2849], Fresh[2848], Fresh[2847], Fresh[2846], Fresh[2845], Fresh[2844], Fresh[2843], Fresh[2842], Fresh[2841], Fresh[2840]}), .outt ({new_AGEMA_signal_2168, new_AGEMA_signal_2167, new_AGEMA_signal_2166, n2085}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2245 ( .ina ({new_AGEMA_signal_12802, new_AGEMA_signal_12800, new_AGEMA_signal_12798, new_AGEMA_signal_12796}), .inb ({new_AGEMA_signal_1676, new_AGEMA_signal_1675, new_AGEMA_signal_1674, n2562}), .clk ( clk ), .rnd ({Fresh[2859], Fresh[2858], Fresh[2857], Fresh[2856], Fresh[2855], Fresh[2854], Fresh[2853], Fresh[2852], Fresh[2851], Fresh[2850]}), .outt ({new_AGEMA_signal_2171, new_AGEMA_signal_2170, new_AGEMA_signal_2169, n2131}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2248 ( .ina ({new_AGEMA_signal_1544, new_AGEMA_signal_1543, new_AGEMA_signal_1542, n2088}), .inb ({new_AGEMA_signal_1352, new_AGEMA_signal_1351, new_AGEMA_signal_1350, n2087}), .clk ( clk ), .rnd ({Fresh[2869], Fresh[2868], Fresh[2867], Fresh[2866], Fresh[2865], Fresh[2864], Fresh[2863], Fresh[2862], Fresh[2861], Fresh[2860]}), .outt ({new_AGEMA_signal_2174, new_AGEMA_signal_2173, new_AGEMA_signal_2172, n2089}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2252 ( .ina ({new_AGEMA_signal_12738, new_AGEMA_signal_12736, new_AGEMA_signal_12734, new_AGEMA_signal_12732}), .inb ({new_AGEMA_signal_1679, new_AGEMA_signal_1678, new_AGEMA_signal_1677, n2156}), .clk ( clk ), .rnd ({Fresh[2879], Fresh[2878], Fresh[2877], Fresh[2876], Fresh[2875], Fresh[2874], Fresh[2873], Fresh[2872], Fresh[2871], Fresh[2870]}), .outt ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, new_AGEMA_signal_2175, n2330}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2254 ( .ina ({new_AGEMA_signal_12810, new_AGEMA_signal_12808, new_AGEMA_signal_12806, new_AGEMA_signal_12804}), .inb ({new_AGEMA_signal_1514, new_AGEMA_signal_1513, new_AGEMA_signal_1512, n2151}), .clk ( clk ), .rnd ({Fresh[2889], Fresh[2888], Fresh[2887], Fresh[2886], Fresh[2885], Fresh[2884], Fresh[2883], Fresh[2882], Fresh[2881], Fresh[2880]}), .outt ({new_AGEMA_signal_2180, new_AGEMA_signal_2179, new_AGEMA_signal_2178, n2092}) ) ;
    or_HPC1 #(.security_order(3), .pipeline(1)) U2256 ( .ina ({new_AGEMA_signal_1550, new_AGEMA_signal_1549, new_AGEMA_signal_1548, n2761}), .inb ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, new_AGEMA_signal_1557, n2359}), .clk ( clk ), .rnd ({Fresh[2899], Fresh[2898], Fresh[2897], Fresh[2896], Fresh[2895], Fresh[2894], Fresh[2893], Fresh[2892], Fresh[2891], Fresh[2890]}), .outt ({new_AGEMA_signal_2183, new_AGEMA_signal_2182, new_AGEMA_signal_2181, n2094}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2261 ( .ina ({new_AGEMA_signal_1289, new_AGEMA_signal_1288, new_AGEMA_signal_1287, n2101}), .inb ({new_AGEMA_signal_1682, new_AGEMA_signal_1681, new_AGEMA_signal_1680, n2100}), .clk ( clk ), .rnd ({Fresh[2909], Fresh[2908], Fresh[2907], Fresh[2906], Fresh[2905], Fresh[2904], Fresh[2903], Fresh[2902], Fresh[2901], Fresh[2900]}), .outt ({new_AGEMA_signal_2186, new_AGEMA_signal_2185, new_AGEMA_signal_2184, n2160}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2265 ( .ina ({new_AGEMA_signal_1232, new_AGEMA_signal_1231, new_AGEMA_signal_1230, n2492}), .inb ({new_AGEMA_signal_12738, new_AGEMA_signal_12736, new_AGEMA_signal_12734, new_AGEMA_signal_12732}), .clk ( clk ), .rnd ({Fresh[2919], Fresh[2918], Fresh[2917], Fresh[2916], Fresh[2915], Fresh[2914], Fresh[2913], Fresh[2912], Fresh[2911], Fresh[2910]}), .outt ({new_AGEMA_signal_1685, new_AGEMA_signal_1684, new_AGEMA_signal_1683, n2504}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2271 ( .ina ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, new_AGEMA_signal_2088, n2417}), .inb ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}), .clk ( clk ), .rnd ({Fresh[2929], Fresh[2928], Fresh[2927], Fresh[2926], Fresh[2925], Fresh[2924], Fresh[2923], Fresh[2922], Fresh[2921], Fresh[2920]}), .outt ({new_AGEMA_signal_2630, new_AGEMA_signal_2629, new_AGEMA_signal_2628, n2114}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2273 ( .ina ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, new_AGEMA_signal_1257, n2677}), .inb ({new_AGEMA_signal_12698, new_AGEMA_signal_12696, new_AGEMA_signal_12694, new_AGEMA_signal_12692}), .clk ( clk ), .rnd ({Fresh[2939], Fresh[2938], Fresh[2937], Fresh[2936], Fresh[2935], Fresh[2934], Fresh[2933], Fresh[2932], Fresh[2931], Fresh[2930]}), .outt ({new_AGEMA_signal_1688, new_AGEMA_signal_1687, new_AGEMA_signal_1686, n2115}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2280 ( .ina ({new_AGEMA_signal_12818, new_AGEMA_signal_12816, new_AGEMA_signal_12814, new_AGEMA_signal_12812}), .inb ({new_AGEMA_signal_1658, new_AGEMA_signal_1657, new_AGEMA_signal_1656, n2731}), .clk ( clk ), .rnd ({Fresh[2949], Fresh[2948], Fresh[2947], Fresh[2946], Fresh[2945], Fresh[2944], Fresh[2943], Fresh[2942], Fresh[2941], Fresh[2940]}), .outt ({new_AGEMA_signal_2192, new_AGEMA_signal_2191, new_AGEMA_signal_2190, n2291}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2281 ( .ina ({new_AGEMA_signal_12562, new_AGEMA_signal_12560, new_AGEMA_signal_12558, new_AGEMA_signal_12556}), .inb ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, n2498}), .clk ( clk ), .rnd ({Fresh[2959], Fresh[2958], Fresh[2957], Fresh[2956], Fresh[2955], Fresh[2954], Fresh[2953], Fresh[2952], Fresh[2951], Fresh[2950]}), .outt ({new_AGEMA_signal_1694, new_AGEMA_signal_1693, new_AGEMA_signal_1692, n2119}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2291 ( .ina ({new_AGEMA_signal_12826, new_AGEMA_signal_12824, new_AGEMA_signal_12822, new_AGEMA_signal_12820}), .inb ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, n2498}), .clk ( clk ), .rnd ({Fresh[2969], Fresh[2968], Fresh[2967], Fresh[2966], Fresh[2965], Fresh[2964], Fresh[2963], Fresh[2962], Fresh[2961], Fresh[2960]}), .outt ({new_AGEMA_signal_1703, new_AGEMA_signal_1702, new_AGEMA_signal_1701, n2130}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2292 ( .ina ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, new_AGEMA_signal_1302, n2817}), .inb ({new_AGEMA_signal_1220, new_AGEMA_signal_1219, new_AGEMA_signal_1218, n2631}), .clk ( clk ), .rnd ({Fresh[2979], Fresh[2978], Fresh[2977], Fresh[2976], Fresh[2975], Fresh[2974], Fresh[2973], Fresh[2972], Fresh[2971], Fresh[2970]}), .outt ({new_AGEMA_signal_1706, new_AGEMA_signal_1705, new_AGEMA_signal_1704, n2129}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2295 ( .ina ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, new_AGEMA_signal_1359, n2647}), .inb ({new_AGEMA_signal_12834, new_AGEMA_signal_12832, new_AGEMA_signal_12830, new_AGEMA_signal_12828}), .clk ( clk ), .rnd ({Fresh[2989], Fresh[2988], Fresh[2987], Fresh[2986], Fresh[2985], Fresh[2984], Fresh[2983], Fresh[2982], Fresh[2981], Fresh[2980]}), .outt ({new_AGEMA_signal_1709, new_AGEMA_signal_1708, new_AGEMA_signal_1707, n2150}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2298 ( .ina ({new_AGEMA_signal_1232, new_AGEMA_signal_1231, new_AGEMA_signal_1230, n2492}), .inb ({new_AGEMA_signal_1364, new_AGEMA_signal_1363, new_AGEMA_signal_1362, n2132}), .clk ( clk ), .rnd ({Fresh[2999], Fresh[2998], Fresh[2997], Fresh[2996], Fresh[2995], Fresh[2994], Fresh[2993], Fresh[2992], Fresh[2991], Fresh[2990]}), .outt ({new_AGEMA_signal_1712, new_AGEMA_signal_1711, new_AGEMA_signal_1710, n2133}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2302 ( .ina ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, new_AGEMA_signal_1605, n2533}), .inb ({new_AGEMA_signal_12842, new_AGEMA_signal_12840, new_AGEMA_signal_12838, new_AGEMA_signal_12836}), .clk ( clk ), .rnd ({Fresh[3009], Fresh[3008], Fresh[3007], Fresh[3006], Fresh[3005], Fresh[3004], Fresh[3003], Fresh[3002], Fresh[3001], Fresh[3000]}), .outt ({new_AGEMA_signal_2201, new_AGEMA_signal_2200, new_AGEMA_signal_2199, n2136}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2306 ( .ina ({new_AGEMA_signal_1598, new_AGEMA_signal_1597, new_AGEMA_signal_1596, n2572}), .inb ({new_AGEMA_signal_1718, new_AGEMA_signal_1717, new_AGEMA_signal_1716, n2138}), .clk ( clk ), .rnd ({Fresh[3019], Fresh[3018], Fresh[3017], Fresh[3016], Fresh[3015], Fresh[3014], Fresh[3013], Fresh[3012], Fresh[3011], Fresh[3010]}), .outt ({new_AGEMA_signal_2204, new_AGEMA_signal_2203, new_AGEMA_signal_2202, n2139}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2313 ( .ina ({new_AGEMA_signal_12850, new_AGEMA_signal_12848, new_AGEMA_signal_12846, new_AGEMA_signal_12844}), .inb ({new_AGEMA_signal_1721, new_AGEMA_signal_1720, new_AGEMA_signal_1719, n2555}), .clk ( clk ), .rnd ({Fresh[3029], Fresh[3028], Fresh[3027], Fresh[3026], Fresh[3025], Fresh[3024], Fresh[3023], Fresh[3022], Fresh[3021], Fresh[3020]}), .outt ({new_AGEMA_signal_2207, new_AGEMA_signal_2206, new_AGEMA_signal_2205, n2144}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2318 ( .ina ({new_AGEMA_signal_1514, new_AGEMA_signal_1513, new_AGEMA_signal_1512, n2151}), .inb ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, new_AGEMA_signal_1605, n2533}), .clk ( clk ), .rnd ({Fresh[3039], Fresh[3038], Fresh[3037], Fresh[3036], Fresh[3035], Fresh[3034], Fresh[3033], Fresh[3032], Fresh[3031], Fresh[3030]}), .outt ({new_AGEMA_signal_2210, new_AGEMA_signal_2209, new_AGEMA_signal_2208, n2152}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2321 ( .ina ({new_AGEMA_signal_1262, new_AGEMA_signal_1261, new_AGEMA_signal_1260, n2627}), .inb ({new_AGEMA_signal_1679, new_AGEMA_signal_1678, new_AGEMA_signal_1677, n2156}), .clk ( clk ), .rnd ({Fresh[3049], Fresh[3048], Fresh[3047], Fresh[3046], Fresh[3045], Fresh[3044], Fresh[3043], Fresh[3042], Fresh[3041], Fresh[3040]}), .outt ({new_AGEMA_signal_2213, new_AGEMA_signal_2212, new_AGEMA_signal_2211, n2170}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2323 ( .ina ({new_AGEMA_signal_1724, new_AGEMA_signal_1723, new_AGEMA_signal_1722, n2429}), .inb ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, new_AGEMA_signal_1521, n2732}), .clk ( clk ), .rnd ({Fresh[3059], Fresh[3058], Fresh[3057], Fresh[3056], Fresh[3055], Fresh[3054], Fresh[3053], Fresh[3052], Fresh[3051], Fresh[3050]}), .outt ({new_AGEMA_signal_2216, new_AGEMA_signal_2215, new_AGEMA_signal_2214, n2157}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2329 ( .ina ({new_AGEMA_signal_12858, new_AGEMA_signal_12856, new_AGEMA_signal_12854, new_AGEMA_signal_12852}), .inb ({new_AGEMA_signal_1367, new_AGEMA_signal_1366, new_AGEMA_signal_1365, n2162}), .clk ( clk ), .rnd ({Fresh[3069], Fresh[3068], Fresh[3067], Fresh[3066], Fresh[3065], Fresh[3064], Fresh[3063], Fresh[3062], Fresh[3061], Fresh[3060]}), .outt ({new_AGEMA_signal_1727, new_AGEMA_signal_1726, new_AGEMA_signal_1725, n2163}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2335 ( .ina ({new_AGEMA_signal_1337, new_AGEMA_signal_1336, new_AGEMA_signal_1335, n2171}), .inb ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, new_AGEMA_signal_1623, n2376}), .clk ( clk ), .rnd ({Fresh[3079], Fresh[3078], Fresh[3077], Fresh[3076], Fresh[3075], Fresh[3074], Fresh[3073], Fresh[3072], Fresh[3071], Fresh[3070]}), .outt ({new_AGEMA_signal_2222, new_AGEMA_signal_2221, new_AGEMA_signal_2220, n2172}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2338 ( .ina ({new_AGEMA_signal_12562, new_AGEMA_signal_12560, new_AGEMA_signal_12558, new_AGEMA_signal_12556}), .inb ({new_AGEMA_signal_1160, new_AGEMA_signal_1159, new_AGEMA_signal_1158, n2545}), .clk ( clk ), .rnd ({Fresh[3089], Fresh[3088], Fresh[3087], Fresh[3086], Fresh[3085], Fresh[3084], Fresh[3083], Fresh[3082], Fresh[3081], Fresh[3080]}), .outt ({new_AGEMA_signal_1370, new_AGEMA_signal_1369, new_AGEMA_signal_1368, n2186}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2339 ( .ina ({new_AGEMA_signal_12658, new_AGEMA_signal_12656, new_AGEMA_signal_12654, new_AGEMA_signal_12652}), .inb ({new_AGEMA_signal_1622, new_AGEMA_signal_1621, new_AGEMA_signal_1620, n2290}), .clk ( clk ), .rnd ({Fresh[3099], Fresh[3098], Fresh[3097], Fresh[3096], Fresh[3095], Fresh[3094], Fresh[3093], Fresh[3092], Fresh[3091], Fresh[3090]}), .outt ({new_AGEMA_signal_2225, new_AGEMA_signal_2224, new_AGEMA_signal_2223, n2181}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2344 ( .ina ({new_AGEMA_signal_1730, new_AGEMA_signal_1729, new_AGEMA_signal_1728, n2176}), .inb ({new_AGEMA_signal_1733, new_AGEMA_signal_1732, new_AGEMA_signal_1731, n2175}), .clk ( clk ), .rnd ({Fresh[3109], Fresh[3108], Fresh[3107], Fresh[3106], Fresh[3105], Fresh[3104], Fresh[3103], Fresh[3102], Fresh[3101], Fresh[3100]}), .outt ({new_AGEMA_signal_2228, new_AGEMA_signal_2227, new_AGEMA_signal_2226, n2177}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2349 ( .ina ({new_AGEMA_signal_12618, new_AGEMA_signal_12616, new_AGEMA_signal_12614, new_AGEMA_signal_12612}), .inb ({new_AGEMA_signal_1166, new_AGEMA_signal_1165, new_AGEMA_signal_1164, n2182}), .clk ( clk ), .rnd ({Fresh[3119], Fresh[3118], Fresh[3117], Fresh[3116], Fresh[3115], Fresh[3114], Fresh[3113], Fresh[3112], Fresh[3111], Fresh[3110]}), .outt ({new_AGEMA_signal_1376, new_AGEMA_signal_1375, new_AGEMA_signal_1374, n2183}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2354 ( .ina ({new_AGEMA_signal_12866, new_AGEMA_signal_12864, new_AGEMA_signal_12862, new_AGEMA_signal_12860}), .inb ({new_AGEMA_signal_1736, new_AGEMA_signal_1735, new_AGEMA_signal_1734, n2188}), .clk ( clk ), .rnd ({Fresh[3129], Fresh[3128], Fresh[3127], Fresh[3126], Fresh[3125], Fresh[3124], Fresh[3123], Fresh[3122], Fresh[3121], Fresh[3120]}), .outt ({new_AGEMA_signal_2231, new_AGEMA_signal_2230, new_AGEMA_signal_2229, n2195}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2356 ( .ina ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, new_AGEMA_signal_1293, n2190}), .inb ({new_AGEMA_signal_1739, new_AGEMA_signal_1738, new_AGEMA_signal_1737, n2189}), .clk ( clk ), .rnd ({Fresh[3139], Fresh[3138], Fresh[3137], Fresh[3136], Fresh[3135], Fresh[3134], Fresh[3133], Fresh[3132], Fresh[3131], Fresh[3130]}), .outt ({new_AGEMA_signal_2234, new_AGEMA_signal_2233, new_AGEMA_signal_2232, n2193}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2358 ( .ina ({new_AGEMA_signal_12874, new_AGEMA_signal_12872, new_AGEMA_signal_12870, new_AGEMA_signal_12868}), .inb ({new_AGEMA_signal_1742, new_AGEMA_signal_1741, new_AGEMA_signal_1740, n2446}), .clk ( clk ), .rnd ({Fresh[3149], Fresh[3148], Fresh[3147], Fresh[3146], Fresh[3145], Fresh[3144], Fresh[3143], Fresh[3142], Fresh[3141], Fresh[3140]}), .outt ({new_AGEMA_signal_2237, new_AGEMA_signal_2236, new_AGEMA_signal_2235, n2191}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2364 ( .ina ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, new_AGEMA_signal_1377, n2576}), .inb ({new_AGEMA_signal_1382, new_AGEMA_signal_1381, new_AGEMA_signal_1380, n2748}), .clk ( clk ), .rnd ({Fresh[3159], Fresh[3158], Fresh[3157], Fresh[3156], Fresh[3155], Fresh[3154], Fresh[3153], Fresh[3152], Fresh[3151], Fresh[3150]}), .outt ({new_AGEMA_signal_1745, new_AGEMA_signal_1744, new_AGEMA_signal_1743, n2196}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2367 ( .ina ({new_AGEMA_signal_12594, new_AGEMA_signal_12592, new_AGEMA_signal_12590, new_AGEMA_signal_12588}), .inb ({new_AGEMA_signal_1556, new_AGEMA_signal_1555, new_AGEMA_signal_1554, n2505}), .clk ( clk ), .rnd ({Fresh[3169], Fresh[3168], Fresh[3167], Fresh[3166], Fresh[3165], Fresh[3164], Fresh[3163], Fresh[3162], Fresh[3161], Fresh[3160]}), .outt ({new_AGEMA_signal_2240, new_AGEMA_signal_2239, new_AGEMA_signal_2238, n2201}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2369 ( .ina ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, new_AGEMA_signal_2241, n2674}), .inb ({new_AGEMA_signal_12882, new_AGEMA_signal_12880, new_AGEMA_signal_12878, new_AGEMA_signal_12876}), .clk ( clk ), .rnd ({Fresh[3179], Fresh[3178], Fresh[3177], Fresh[3176], Fresh[3175], Fresh[3174], Fresh[3173], Fresh[3172], Fresh[3171], Fresh[3170]}), .outt ({new_AGEMA_signal_2663, new_AGEMA_signal_2662, new_AGEMA_signal_2661, n2200}) ) ;
    mux2_HPC1 #(.security_order(3), .pipeline(1)) U2371 ( .ins ({new_AGEMA_signal_12834, new_AGEMA_signal_12832, new_AGEMA_signal_12830, new_AGEMA_signal_12828}), .inb ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, new_AGEMA_signal_1515, n2734}), .ina ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, new_AGEMA_signal_2088, n2417}), .clk ( clk ), .rnd ({Fresh[3189], Fresh[3188], Fresh[3187], Fresh[3186], Fresh[3185], Fresh[3184], Fresh[3183], Fresh[3182], Fresh[3181], Fresh[3180]}), .outt ({new_AGEMA_signal_2666, new_AGEMA_signal_2665, new_AGEMA_signal_2664, n2202}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2379 ( .ina ({new_AGEMA_signal_1619, new_AGEMA_signal_1618, new_AGEMA_signal_1617, n2214}), .inb ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, new_AGEMA_signal_1383, n2213}), .clk ( clk ), .rnd ({Fresh[3199], Fresh[3198], Fresh[3197], Fresh[3196], Fresh[3195], Fresh[3194], Fresh[3193], Fresh[3192], Fresh[3191], Fresh[3190]}), .outt ({new_AGEMA_signal_2246, new_AGEMA_signal_2245, new_AGEMA_signal_2244, n2217}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2381 ( .ina ({new_AGEMA_signal_12890, new_AGEMA_signal_12888, new_AGEMA_signal_12886, new_AGEMA_signal_12884}), .inb ({new_AGEMA_signal_1388, new_AGEMA_signal_1387, new_AGEMA_signal_1386, n2215}), .clk ( clk ), .rnd ({Fresh[3209], Fresh[3208], Fresh[3207], Fresh[3206], Fresh[3205], Fresh[3204], Fresh[3203], Fresh[3202], Fresh[3201], Fresh[3200]}), .outt ({new_AGEMA_signal_1748, new_AGEMA_signal_1747, new_AGEMA_signal_1746, n2216}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2385 ( .ina ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, new_AGEMA_signal_1749, n2218}), .inb ({new_AGEMA_signal_12874, new_AGEMA_signal_12872, new_AGEMA_signal_12870, new_AGEMA_signal_12868}), .clk ( clk ), .rnd ({Fresh[3219], Fresh[3218], Fresh[3217], Fresh[3216], Fresh[3215], Fresh[3214], Fresh[3213], Fresh[3212], Fresh[3211], Fresh[3210]}), .outt ({new_AGEMA_signal_2249, new_AGEMA_signal_2248, new_AGEMA_signal_2247, n2222}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2387 ( .ina ({new_AGEMA_signal_1715, new_AGEMA_signal_1714, new_AGEMA_signal_1713, n2220}), .inb ({new_AGEMA_signal_1754, new_AGEMA_signal_1753, new_AGEMA_signal_1752, n2219}), .clk ( clk ), .rnd ({Fresh[3229], Fresh[3228], Fresh[3227], Fresh[3226], Fresh[3225], Fresh[3224], Fresh[3223], Fresh[3222], Fresh[3221], Fresh[3220]}), .outt ({new_AGEMA_signal_2252, new_AGEMA_signal_2251, new_AGEMA_signal_2250, n2221}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2391 ( .ina ({new_AGEMA_signal_1262, new_AGEMA_signal_1261, new_AGEMA_signal_1260, n2627}), .inb ({new_AGEMA_signal_12898, new_AGEMA_signal_12896, new_AGEMA_signal_12894, new_AGEMA_signal_12892}), .clk ( clk ), .rnd ({Fresh[3239], Fresh[3238], Fresh[3237], Fresh[3236], Fresh[3235], Fresh[3234], Fresh[3233], Fresh[3232], Fresh[3231], Fresh[3230]}), .outt ({new_AGEMA_signal_1757, new_AGEMA_signal_1756, new_AGEMA_signal_1755, n2226}) ) ;
    mux2_HPC1 #(.security_order(3), .pipeline(1)) U2393 ( .ins ({new_AGEMA_signal_12834, new_AGEMA_signal_12832, new_AGEMA_signal_12830, new_AGEMA_signal_12828}), .inb ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}), .ina ({new_AGEMA_signal_1328, new_AGEMA_signal_1327, new_AGEMA_signal_1326, n2227}), .clk ( clk ), .rnd ({Fresh[3249], Fresh[3248], Fresh[3247], Fresh[3246], Fresh[3245], Fresh[3244], Fresh[3243], Fresh[3242], Fresh[3241], Fresh[3240]}), .outt ({new_AGEMA_signal_1760, new_AGEMA_signal_1759, new_AGEMA_signal_1758, n2228}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2397 ( .ina ({new_AGEMA_signal_12714, new_AGEMA_signal_12712, new_AGEMA_signal_12710, new_AGEMA_signal_12708}), .inb ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}), .clk ( clk ), .rnd ({Fresh[3259], Fresh[3258], Fresh[3257], Fresh[3256], Fresh[3255], Fresh[3254], Fresh[3253], Fresh[3252], Fresh[3251], Fresh[3250]}), .outt ({new_AGEMA_signal_1763, new_AGEMA_signal_1762, new_AGEMA_signal_1761, n2237}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2398 ( .ina ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, new_AGEMA_signal_2088, n2417}), .inb ({new_AGEMA_signal_12834, new_AGEMA_signal_12832, new_AGEMA_signal_12830, new_AGEMA_signal_12828}), .clk ( clk ), .rnd ({Fresh[3269], Fresh[3268], Fresh[3267], Fresh[3266], Fresh[3265], Fresh[3264], Fresh[3263], Fresh[3262], Fresh[3261], Fresh[3260]}), .outt ({new_AGEMA_signal_2678, new_AGEMA_signal_2677, new_AGEMA_signal_2676, n2233}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2403 ( .ina ({new_AGEMA_signal_12906, new_AGEMA_signal_12904, new_AGEMA_signal_12902, new_AGEMA_signal_12900}), .inb ({new_AGEMA_signal_1220, new_AGEMA_signal_1219, new_AGEMA_signal_1218, n2631}), .clk ( clk ), .rnd ({Fresh[3279], Fresh[3278], Fresh[3277], Fresh[3276], Fresh[3275], Fresh[3274], Fresh[3273], Fresh[3272], Fresh[3271], Fresh[3270]}), .outt ({new_AGEMA_signal_1766, new_AGEMA_signal_1765, new_AGEMA_signal_1764, n2238}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2406 ( .ina ({new_AGEMA_signal_1589, new_AGEMA_signal_1588, new_AGEMA_signal_1587, n2241}), .inb ({new_AGEMA_signal_1769, new_AGEMA_signal_1768, new_AGEMA_signal_1767, n2240}), .clk ( clk ), .rnd ({Fresh[3289], Fresh[3288], Fresh[3287], Fresh[3286], Fresh[3285], Fresh[3284], Fresh[3283], Fresh[3282], Fresh[3281], Fresh[3280]}), .outt ({new_AGEMA_signal_2258, new_AGEMA_signal_2257, new_AGEMA_signal_2256, n2248}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2409 ( .ina ({new_AGEMA_signal_1772, new_AGEMA_signal_1771, new_AGEMA_signal_1770, n2561}), .inb ({new_AGEMA_signal_1775, new_AGEMA_signal_1774, new_AGEMA_signal_1773, n2243}), .clk ( clk ), .rnd ({Fresh[3299], Fresh[3298], Fresh[3297], Fresh[3296], Fresh[3295], Fresh[3294], Fresh[3293], Fresh[3292], Fresh[3291], Fresh[3290]}), .outt ({new_AGEMA_signal_2261, new_AGEMA_signal_2260, new_AGEMA_signal_2259, n2244}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2414 ( .ina ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, new_AGEMA_signal_1623, n2376}), .inb ({new_AGEMA_signal_12554, new_AGEMA_signal_12552, new_AGEMA_signal_12550, new_AGEMA_signal_12548}), .clk ( clk ), .rnd ({Fresh[3309], Fresh[3308], Fresh[3307], Fresh[3306], Fresh[3305], Fresh[3304], Fresh[3303], Fresh[3302], Fresh[3301], Fresh[3300]}), .outt ({new_AGEMA_signal_2264, new_AGEMA_signal_2263, new_AGEMA_signal_2262, n2249}) ) ;
    mux2_HPC1 #(.security_order(3), .pipeline(1)) U2417 ( .ins ({new_AGEMA_signal_12834, new_AGEMA_signal_12832, new_AGEMA_signal_12830, new_AGEMA_signal_12828}), .inb ({new_AGEMA_signal_1664, new_AGEMA_signal_1663, new_AGEMA_signal_1662, n2252}), .ina ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}), .clk ( clk ), .rnd ({Fresh[3319], Fresh[3318], Fresh[3317], Fresh[3316], Fresh[3315], Fresh[3314], Fresh[3313], Fresh[3312], Fresh[3311], Fresh[3310]}), .outt ({new_AGEMA_signal_2267, new_AGEMA_signal_2266, new_AGEMA_signal_2265, n2253}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2424 ( .ina ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, new_AGEMA_signal_1605, n2533}), .inb ({new_AGEMA_signal_1784, new_AGEMA_signal_1783, new_AGEMA_signal_1782, n2259}), .clk ( clk ), .rnd ({Fresh[3329], Fresh[3328], Fresh[3327], Fresh[3326], Fresh[3325], Fresh[3324], Fresh[3323], Fresh[3322], Fresh[3321], Fresh[3320]}), .outt ({new_AGEMA_signal_2270, new_AGEMA_signal_2269, new_AGEMA_signal_2268, n2260}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2429 ( .ina ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, new_AGEMA_signal_2088, n2417}), .inb ({new_AGEMA_signal_12914, new_AGEMA_signal_12912, new_AGEMA_signal_12910, new_AGEMA_signal_12908}), .clk ( clk ), .rnd ({Fresh[3339], Fresh[3338], Fresh[3337], Fresh[3336], Fresh[3335], Fresh[3334], Fresh[3333], Fresh[3332], Fresh[3331], Fresh[3330]}), .outt ({new_AGEMA_signal_2690, new_AGEMA_signal_2689, new_AGEMA_signal_2688, n2273}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2430 ( .ina ({new_AGEMA_signal_12922, new_AGEMA_signal_12920, new_AGEMA_signal_12918, new_AGEMA_signal_12916}), .inb ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, new_AGEMA_signal_2085, n2720}), .clk ( clk ), .rnd ({Fresh[3349], Fresh[3348], Fresh[3347], Fresh[3346], Fresh[3345], Fresh[3344], Fresh[3343], Fresh[3342], Fresh[3341], Fresh[3340]}), .outt ({new_AGEMA_signal_2693, new_AGEMA_signal_2692, new_AGEMA_signal_2691, n2752}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2433 ( .ina ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, new_AGEMA_signal_1395, n2645}), .inb ({new_AGEMA_signal_12818, new_AGEMA_signal_12816, new_AGEMA_signal_12814, new_AGEMA_signal_12812}), .clk ( clk ), .rnd ({Fresh[3359], Fresh[3358], Fresh[3357], Fresh[3356], Fresh[3355], Fresh[3354], Fresh[3353], Fresh[3352], Fresh[3351], Fresh[3350]}), .outt ({new_AGEMA_signal_1787, new_AGEMA_signal_1786, new_AGEMA_signal_1785, n2265}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2437 ( .ina ({new_AGEMA_signal_12930, new_AGEMA_signal_12928, new_AGEMA_signal_12926, new_AGEMA_signal_12924}), .inb ({new_AGEMA_signal_1400, new_AGEMA_signal_1399, new_AGEMA_signal_1398, n2268}), .clk ( clk ), .rnd ({Fresh[3369], Fresh[3368], Fresh[3367], Fresh[3366], Fresh[3365], Fresh[3364], Fresh[3363], Fresh[3362], Fresh[3361], Fresh[3360]}), .outt ({new_AGEMA_signal_1790, new_AGEMA_signal_1789, new_AGEMA_signal_1788, n2269}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2444 ( .ina ({new_AGEMA_signal_12634, new_AGEMA_signal_12632, new_AGEMA_signal_12630, new_AGEMA_signal_12628}), .inb ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, new_AGEMA_signal_1302, n2817}), .clk ( clk ), .rnd ({Fresh[3379], Fresh[3378], Fresh[3377], Fresh[3376], Fresh[3375], Fresh[3374], Fresh[3373], Fresh[3372], Fresh[3371], Fresh[3370]}), .outt ({new_AGEMA_signal_1796, new_AGEMA_signal_1795, new_AGEMA_signal_1794, n2277}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2449 ( .ina ({new_AGEMA_signal_12938, new_AGEMA_signal_12936, new_AGEMA_signal_12934, new_AGEMA_signal_12932}), .inb ({new_AGEMA_signal_1403, new_AGEMA_signal_1402, new_AGEMA_signal_1401, n2383}), .clk ( clk ), .rnd ({Fresh[3389], Fresh[3388], Fresh[3387], Fresh[3386], Fresh[3385], Fresh[3384], Fresh[3383], Fresh[3382], Fresh[3381], Fresh[3380]}), .outt ({new_AGEMA_signal_1799, new_AGEMA_signal_1798, new_AGEMA_signal_1797, n2282}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2452 ( .ina ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, new_AGEMA_signal_1269, n2736}), .inb ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, new_AGEMA_signal_1605, n2533}), .clk ( clk ), .rnd ({Fresh[3399], Fresh[3398], Fresh[3397], Fresh[3396], Fresh[3395], Fresh[3394], Fresh[3393], Fresh[3392], Fresh[3391], Fresh[3390]}), .outt ({new_AGEMA_signal_2285, new_AGEMA_signal_2284, new_AGEMA_signal_2283, n2284}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2456 ( .ina ({new_AGEMA_signal_1802, new_AGEMA_signal_1801, new_AGEMA_signal_1800, n2774}), .inb ({new_AGEMA_signal_12946, new_AGEMA_signal_12944, new_AGEMA_signal_12942, new_AGEMA_signal_12940}), .clk ( clk ), .rnd ({Fresh[3409], Fresh[3408], Fresh[3407], Fresh[3406], Fresh[3405], Fresh[3404], Fresh[3403], Fresh[3402], Fresh[3401], Fresh[3400]}), .outt ({new_AGEMA_signal_2288, new_AGEMA_signal_2287, new_AGEMA_signal_2286, n2459}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2459 ( .ina ({new_AGEMA_signal_12570, new_AGEMA_signal_12568, new_AGEMA_signal_12566, new_AGEMA_signal_12564}), .inb ({new_AGEMA_signal_1805, new_AGEMA_signal_1804, new_AGEMA_signal_1803, n2287}), .clk ( clk ), .rnd ({Fresh[3419], Fresh[3418], Fresh[3417], Fresh[3416], Fresh[3415], Fresh[3414], Fresh[3413], Fresh[3412], Fresh[3411], Fresh[3410]}), .outt ({new_AGEMA_signal_2291, new_AGEMA_signal_2290, new_AGEMA_signal_2289, n2288}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2462 ( .ina ({new_AGEMA_signal_12562, new_AGEMA_signal_12560, new_AGEMA_signal_12558, new_AGEMA_signal_12556}), .inb ({new_AGEMA_signal_1550, new_AGEMA_signal_1549, new_AGEMA_signal_1548, n2761}), .clk ( clk ), .rnd ({Fresh[3429], Fresh[3428], Fresh[3427], Fresh[3426], Fresh[3425], Fresh[3424], Fresh[3423], Fresh[3422], Fresh[3421], Fresh[3420]}), .outt ({new_AGEMA_signal_2294, new_AGEMA_signal_2293, new_AGEMA_signal_2292, n2458}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2464 ( .ina ({new_AGEMA_signal_12858, new_AGEMA_signal_12856, new_AGEMA_signal_12854, new_AGEMA_signal_12852}), .inb ({new_AGEMA_signal_1622, new_AGEMA_signal_1621, new_AGEMA_signal_1620, n2290}), .clk ( clk ), .rnd ({Fresh[3439], Fresh[3438], Fresh[3437], Fresh[3436], Fresh[3435], Fresh[3434], Fresh[3433], Fresh[3432], Fresh[3431], Fresh[3430]}), .outt ({new_AGEMA_signal_2297, new_AGEMA_signal_2296, new_AGEMA_signal_2295, n2293}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2467 ( .ina ({new_AGEMA_signal_12810, new_AGEMA_signal_12808, new_AGEMA_signal_12806, new_AGEMA_signal_12804}), .inb ({new_AGEMA_signal_1340, new_AGEMA_signal_1339, new_AGEMA_signal_1338, n2642}), .clk ( clk ), .rnd ({Fresh[3449], Fresh[3448], Fresh[3447], Fresh[3446], Fresh[3445], Fresh[3444], Fresh[3443], Fresh[3442], Fresh[3441], Fresh[3440]}), .outt ({new_AGEMA_signal_1808, new_AGEMA_signal_1807, new_AGEMA_signal_1806, n2294}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2472 ( .ina ({new_AGEMA_signal_1811, new_AGEMA_signal_1810, new_AGEMA_signal_1809, n2438}), .inb ({new_AGEMA_signal_1406, new_AGEMA_signal_1405, new_AGEMA_signal_1404, n2299}), .clk ( clk ), .rnd ({Fresh[3459], Fresh[3458], Fresh[3457], Fresh[3456], Fresh[3455], Fresh[3454], Fresh[3453], Fresh[3452], Fresh[3451], Fresh[3450]}), .outt ({new_AGEMA_signal_2300, new_AGEMA_signal_2299, new_AGEMA_signal_2298, n2300}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2480 ( .ina ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, new_AGEMA_signal_1515, n2734}), .inb ({new_AGEMA_signal_12874, new_AGEMA_signal_12872, new_AGEMA_signal_12870, new_AGEMA_signal_12868}), .clk ( clk ), .rnd ({Fresh[3469], Fresh[3468], Fresh[3467], Fresh[3466], Fresh[3465], Fresh[3464], Fresh[3463], Fresh[3462], Fresh[3461], Fresh[3460]}), .outt ({new_AGEMA_signal_2303, new_AGEMA_signal_2302, new_AGEMA_signal_2301, n2323}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) U2482 ( .ina ({new_AGEMA_signal_1283, new_AGEMA_signal_1282, new_AGEMA_signal_1281, n2571}), .inb ({new_AGEMA_signal_1814, new_AGEMA_signal_1813, new_AGEMA_signal_1812, n2371}), .clk ( clk ), .rnd ({Fresh[3479], Fresh[3478], Fresh[3477], Fresh[3476], Fresh[3475], Fresh[3474], Fresh[3473], Fresh[3472], Fresh[3471], Fresh[3470]}), .outt ({new_AGEMA_signal_2306, new_AGEMA_signal_2305, new_AGEMA_signal_2304, n2314}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2485 ( .ina ({new_AGEMA_signal_1172, new_AGEMA_signal_1171, new_AGEMA_signal_1170, n2316}), .inb ({new_AGEMA_signal_12954, new_AGEMA_signal_12952, new_AGEMA_signal_12950, new_AGEMA_signal_12948}), .clk ( clk ), .rnd ({Fresh[3489], Fresh[3488], Fresh[3487], Fresh[3486], Fresh[3485], Fresh[3484], Fresh[3483], Fresh[3482], Fresh[3481], Fresh[3480]}), .outt ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, new_AGEMA_signal_1407, n2319}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2491 ( .ina ({new_AGEMA_signal_1340, new_AGEMA_signal_1339, new_AGEMA_signal_1338, n2642}), .inb ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, n2498}), .clk ( clk ), .rnd ({Fresh[3499], Fresh[3498], Fresh[3497], Fresh[3496], Fresh[3495], Fresh[3494], Fresh[3493], Fresh[3492], Fresh[3491], Fresh[3490]}), .outt ({new_AGEMA_signal_1820, new_AGEMA_signal_1819, new_AGEMA_signal_1818, n2326}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2496 ( .ina ({new_AGEMA_signal_1826, new_AGEMA_signal_1825, new_AGEMA_signal_1824, n2328}), .inb ({new_AGEMA_signal_1415, new_AGEMA_signal_1414, new_AGEMA_signal_1413, n2327}), .clk ( clk ), .rnd ({Fresh[3509], Fresh[3508], Fresh[3507], Fresh[3506], Fresh[3505], Fresh[3504], Fresh[3503], Fresh[3502], Fresh[3501], Fresh[3500]}), .outt ({new_AGEMA_signal_2312, new_AGEMA_signal_2311, new_AGEMA_signal_2310, n2329}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2501 ( .ina ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, new_AGEMA_signal_2088, n2417}), .inb ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, new_AGEMA_signal_2241, n2674}), .clk ( clk ), .rnd ({Fresh[3519], Fresh[3518], Fresh[3517], Fresh[3516], Fresh[3515], Fresh[3514], Fresh[3513], Fresh[3512], Fresh[3511], Fresh[3510]}), .outt ({new_AGEMA_signal_2729, new_AGEMA_signal_2728, new_AGEMA_signal_2727, n2335}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2506 ( .ina ({new_AGEMA_signal_12706, new_AGEMA_signal_12704, new_AGEMA_signal_12702, new_AGEMA_signal_12700}), .inb ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, new_AGEMA_signal_1623, n2376}), .clk ( clk ), .rnd ({Fresh[3529], Fresh[3528], Fresh[3527], Fresh[3526], Fresh[3525], Fresh[3524], Fresh[3523], Fresh[3522], Fresh[3521], Fresh[3520]}), .outt ({new_AGEMA_signal_2315, new_AGEMA_signal_2314, new_AGEMA_signal_2313, n2341}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2507 ( .ina ({new_AGEMA_signal_12962, new_AGEMA_signal_12960, new_AGEMA_signal_12958, new_AGEMA_signal_12956}), .inb ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, new_AGEMA_signal_1269, n2736}), .clk ( clk ), .rnd ({Fresh[3539], Fresh[3538], Fresh[3537], Fresh[3536], Fresh[3535], Fresh[3534], Fresh[3533], Fresh[3532], Fresh[3531], Fresh[3530]}), .outt ({new_AGEMA_signal_1832, new_AGEMA_signal_1831, new_AGEMA_signal_1830, n2340}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2514 ( .ina ({new_AGEMA_signal_1418, new_AGEMA_signal_1417, new_AGEMA_signal_1416, n2348}), .inb ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, new_AGEMA_signal_1419, n2347}), .clk ( clk ), .rnd ({Fresh[3549], Fresh[3548], Fresh[3547], Fresh[3546], Fresh[3545], Fresh[3544], Fresh[3543], Fresh[3542], Fresh[3541], Fresh[3540]}), .outt ({new_AGEMA_signal_1838, new_AGEMA_signal_1837, new_AGEMA_signal_1836, n2349}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2517 ( .ina ({new_AGEMA_signal_12970, new_AGEMA_signal_12968, new_AGEMA_signal_12966, new_AGEMA_signal_12964}), .inb ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, new_AGEMA_signal_1299, n2690}), .clk ( clk ), .rnd ({Fresh[3559], Fresh[3558], Fresh[3557], Fresh[3556], Fresh[3555], Fresh[3554], Fresh[3553], Fresh[3552], Fresh[3551], Fresh[3550]}), .outt ({new_AGEMA_signal_1841, new_AGEMA_signal_1840, new_AGEMA_signal_1839, n2375}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2518 ( .ina ({new_AGEMA_signal_12850, new_AGEMA_signal_12848, new_AGEMA_signal_12846, new_AGEMA_signal_12844}), .inb ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, new_AGEMA_signal_1269, n2736}), .clk ( clk ), .rnd ({Fresh[3569], Fresh[3568], Fresh[3567], Fresh[3566], Fresh[3565], Fresh[3564], Fresh[3563], Fresh[3562], Fresh[3561], Fresh[3560]}), .outt ({new_AGEMA_signal_1844, new_AGEMA_signal_1843, new_AGEMA_signal_1842, n2352}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2522 ( .ina ({new_AGEMA_signal_1847, new_AGEMA_signal_1846, new_AGEMA_signal_1845, n2353}), .inb ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, new_AGEMA_signal_1605, n2533}), .clk ( clk ), .rnd ({Fresh[3579], Fresh[3578], Fresh[3577], Fresh[3576], Fresh[3575], Fresh[3574], Fresh[3573], Fresh[3572], Fresh[3571], Fresh[3570]}), .outt ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, new_AGEMA_signal_2319, n2354}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2525 ( .ina ({new_AGEMA_signal_12978, new_AGEMA_signal_12976, new_AGEMA_signal_12974, new_AGEMA_signal_12972}), .inb ({new_AGEMA_signal_1850, new_AGEMA_signal_1849, new_AGEMA_signal_1848, n2355}), .clk ( clk ), .rnd ({Fresh[3589], Fresh[3588], Fresh[3587], Fresh[3586], Fresh[3585], Fresh[3584], Fresh[3583], Fresh[3582], Fresh[3581], Fresh[3580]}), .outt ({new_AGEMA_signal_2324, new_AGEMA_signal_2323, new_AGEMA_signal_2322, n2357}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2527 ( .ina ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, new_AGEMA_signal_1557, n2359}), .inb ({new_AGEMA_signal_12986, new_AGEMA_signal_12984, new_AGEMA_signal_12982, new_AGEMA_signal_12980}), .clk ( clk ), .rnd ({Fresh[3599], Fresh[3598], Fresh[3597], Fresh[3596], Fresh[3595], Fresh[3594], Fresh[3593], Fresh[3592], Fresh[3591], Fresh[3590]}), .outt ({new_AGEMA_signal_2327, new_AGEMA_signal_2326, new_AGEMA_signal_2325, n2360}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2534 ( .ina ({new_AGEMA_signal_12562, new_AGEMA_signal_12560, new_AGEMA_signal_12558, new_AGEMA_signal_12556}), .inb ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, new_AGEMA_signal_2241, n2674}), .clk ( clk ), .rnd ({Fresh[3609], Fresh[3608], Fresh[3607], Fresh[3606], Fresh[3605], Fresh[3604], Fresh[3603], Fresh[3602], Fresh[3601], Fresh[3600]}), .outt ({new_AGEMA_signal_2738, new_AGEMA_signal_2737, new_AGEMA_signal_2736, n2369}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2536 ( .ina ({new_AGEMA_signal_1814, new_AGEMA_signal_1813, new_AGEMA_signal_1812, n2371}), .inb ({new_AGEMA_signal_12898, new_AGEMA_signal_12896, new_AGEMA_signal_12894, new_AGEMA_signal_12892}), .clk ( clk ), .rnd ({Fresh[3619], Fresh[3618], Fresh[3617], Fresh[3616], Fresh[3615], Fresh[3614], Fresh[3613], Fresh[3612], Fresh[3611], Fresh[3610]}), .outt ({new_AGEMA_signal_2330, new_AGEMA_signal_2329, new_AGEMA_signal_2328, n2372}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2539 ( .ina ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, new_AGEMA_signal_1377, n2576}), .inb ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, new_AGEMA_signal_1623, n2376}), .clk ( clk ), .rnd ({Fresh[3629], Fresh[3628], Fresh[3627], Fresh[3626], Fresh[3625], Fresh[3624], Fresh[3623], Fresh[3622], Fresh[3621], Fresh[3620]}), .outt ({new_AGEMA_signal_2333, new_AGEMA_signal_2332, new_AGEMA_signal_2331, n2377}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2544 ( .ina ({new_AGEMA_signal_12874, new_AGEMA_signal_12872, new_AGEMA_signal_12870, new_AGEMA_signal_12868}), .inb ({new_AGEMA_signal_1427, new_AGEMA_signal_1426, new_AGEMA_signal_1425, n2415}), .clk ( clk ), .rnd ({Fresh[3639], Fresh[3638], Fresh[3637], Fresh[3636], Fresh[3635], Fresh[3634], Fresh[3633], Fresh[3632], Fresh[3631], Fresh[3630]}), .outt ({new_AGEMA_signal_1856, new_AGEMA_signal_1855, new_AGEMA_signal_1854, n2467}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2545 ( .ina ({new_AGEMA_signal_12994, new_AGEMA_signal_12992, new_AGEMA_signal_12990, new_AGEMA_signal_12988}), .inb ({new_AGEMA_signal_1403, new_AGEMA_signal_1402, new_AGEMA_signal_1401, n2383}), .clk ( clk ), .rnd ({Fresh[3649], Fresh[3648], Fresh[3647], Fresh[3646], Fresh[3645], Fresh[3644], Fresh[3643], Fresh[3642], Fresh[3641], Fresh[3640]}), .outt ({new_AGEMA_signal_1859, new_AGEMA_signal_1858, new_AGEMA_signal_1857, n2385}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2546 ( .ina ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}), .inb ({new_AGEMA_signal_12738, new_AGEMA_signal_12736, new_AGEMA_signal_12734, new_AGEMA_signal_12732}), .clk ( clk ), .rnd ({Fresh[3659], Fresh[3658], Fresh[3657], Fresh[3656], Fresh[3655], Fresh[3654], Fresh[3653], Fresh[3652], Fresh[3651], Fresh[3650]}), .outt ({new_AGEMA_signal_1862, new_AGEMA_signal_1861, new_AGEMA_signal_1860, n2384}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2548 ( .ina ({new_AGEMA_signal_12698, new_AGEMA_signal_12696, new_AGEMA_signal_12694, new_AGEMA_signal_12692}), .inb ({new_AGEMA_signal_1724, new_AGEMA_signal_1723, new_AGEMA_signal_1722, n2429}), .clk ( clk ), .rnd ({Fresh[3669], Fresh[3668], Fresh[3667], Fresh[3666], Fresh[3665], Fresh[3664], Fresh[3663], Fresh[3662], Fresh[3661], Fresh[3660]}), .outt ({new_AGEMA_signal_2339, new_AGEMA_signal_2338, new_AGEMA_signal_2337, n2386}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2552 ( .ina ({new_AGEMA_signal_12866, new_AGEMA_signal_12864, new_AGEMA_signal_12862, new_AGEMA_signal_12860}), .inb ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, new_AGEMA_signal_1359, n2647}), .clk ( clk ), .rnd ({Fresh[3679], Fresh[3678], Fresh[3677], Fresh[3676], Fresh[3675], Fresh[3674], Fresh[3673], Fresh[3672], Fresh[3671], Fresh[3670]}), .outt ({new_AGEMA_signal_1865, new_AGEMA_signal_1864, new_AGEMA_signal_1863, n2394}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2553 ( .ina ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}), .inb ({new_AGEMA_signal_12874, new_AGEMA_signal_12872, new_AGEMA_signal_12870, new_AGEMA_signal_12868}), .clk ( clk ), .rnd ({Fresh[3689], Fresh[3688], Fresh[3687], Fresh[3686], Fresh[3685], Fresh[3684], Fresh[3683], Fresh[3682], Fresh[3681], Fresh[3680]}), .outt ({new_AGEMA_signal_1868, new_AGEMA_signal_1867, new_AGEMA_signal_1866, n2391}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2554 ( .ina ({new_AGEMA_signal_1556, new_AGEMA_signal_1555, new_AGEMA_signal_1554, n2505}), .inb ({new_AGEMA_signal_12738, new_AGEMA_signal_12736, new_AGEMA_signal_12734, new_AGEMA_signal_12732}), .clk ( clk ), .rnd ({Fresh[3699], Fresh[3698], Fresh[3697], Fresh[3696], Fresh[3695], Fresh[3694], Fresh[3693], Fresh[3692], Fresh[3691], Fresh[3690]}), .outt ({new_AGEMA_signal_2342, new_AGEMA_signal_2341, new_AGEMA_signal_2340, n2390}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2559 ( .ina ({new_AGEMA_signal_12810, new_AGEMA_signal_12808, new_AGEMA_signal_12806, new_AGEMA_signal_12804}), .inb ({new_AGEMA_signal_1430, new_AGEMA_signal_1429, new_AGEMA_signal_1428, n2700}), .clk ( clk ), .rnd ({Fresh[3709], Fresh[3708], Fresh[3707], Fresh[3706], Fresh[3705], Fresh[3704], Fresh[3703], Fresh[3702], Fresh[3701], Fresh[3700]}), .outt ({new_AGEMA_signal_1871, new_AGEMA_signal_1870, new_AGEMA_signal_1869, n2396}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2562 ( .ina ({new_AGEMA_signal_13002, new_AGEMA_signal_13000, new_AGEMA_signal_12998, new_AGEMA_signal_12996}), .inb ({new_AGEMA_signal_1811, new_AGEMA_signal_1810, new_AGEMA_signal_1809, n2438}), .clk ( clk ), .rnd ({Fresh[3719], Fresh[3718], Fresh[3717], Fresh[3716], Fresh[3715], Fresh[3714], Fresh[3713], Fresh[3712], Fresh[3711], Fresh[3710]}), .outt ({new_AGEMA_signal_2345, new_AGEMA_signal_2344, new_AGEMA_signal_2343, n2406}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2565 ( .ina ({new_AGEMA_signal_1433, new_AGEMA_signal_1432, new_AGEMA_signal_1431, n2594}), .inb ({new_AGEMA_signal_1436, new_AGEMA_signal_1435, new_AGEMA_signal_1434, n2402}), .clk ( clk ), .rnd ({Fresh[3729], Fresh[3728], Fresh[3727], Fresh[3726], Fresh[3725], Fresh[3724], Fresh[3723], Fresh[3722], Fresh[3721], Fresh[3720]}), .outt ({new_AGEMA_signal_1874, new_AGEMA_signal_1873, new_AGEMA_signal_1872, n2403}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2569 ( .ina ({new_AGEMA_signal_1652, new_AGEMA_signal_1651, new_AGEMA_signal_1650, n2407}), .inb ({new_AGEMA_signal_12842, new_AGEMA_signal_12840, new_AGEMA_signal_12838, new_AGEMA_signal_12836}), .clk ( clk ), .rnd ({Fresh[3739], Fresh[3738], Fresh[3737], Fresh[3736], Fresh[3735], Fresh[3734], Fresh[3733], Fresh[3732], Fresh[3731], Fresh[3730]}), .outt ({new_AGEMA_signal_2351, new_AGEMA_signal_2350, new_AGEMA_signal_2349, n2408}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2573 ( .ina ({new_AGEMA_signal_1553, new_AGEMA_signal_1552, new_AGEMA_signal_1551, n2412}), .inb ({new_AGEMA_signal_12906, new_AGEMA_signal_12904, new_AGEMA_signal_12902, new_AGEMA_signal_12900}), .clk ( clk ), .rnd ({Fresh[3749], Fresh[3748], Fresh[3747], Fresh[3746], Fresh[3745], Fresh[3744], Fresh[3743], Fresh[3742], Fresh[3741], Fresh[3740]}), .outt ({new_AGEMA_signal_2354, new_AGEMA_signal_2353, new_AGEMA_signal_2352, n2574}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2574 ( .ina ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, n2498}), .inb ({new_AGEMA_signal_12762, new_AGEMA_signal_12760, new_AGEMA_signal_12758, new_AGEMA_signal_12756}), .clk ( clk ), .rnd ({Fresh[3759], Fresh[3758], Fresh[3757], Fresh[3756], Fresh[3755], Fresh[3754], Fresh[3753], Fresh[3752], Fresh[3751], Fresh[3750]}), .outt ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, new_AGEMA_signal_1875, n2413}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2577 ( .ina ({new_AGEMA_signal_1427, new_AGEMA_signal_1426, new_AGEMA_signal_1425, n2415}), .inb ({new_AGEMA_signal_12738, new_AGEMA_signal_12736, new_AGEMA_signal_12734, new_AGEMA_signal_12732}), .clk ( clk ), .rnd ({Fresh[3769], Fresh[3768], Fresh[3767], Fresh[3766], Fresh[3765], Fresh[3764], Fresh[3763], Fresh[3762], Fresh[3761], Fresh[3760]}), .outt ({new_AGEMA_signal_1880, new_AGEMA_signal_1879, new_AGEMA_signal_1878, n2416}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2586 ( .ina ({new_AGEMA_signal_1883, new_AGEMA_signal_1882, new_AGEMA_signal_1881, n2428}), .inb ({new_AGEMA_signal_13010, new_AGEMA_signal_13008, new_AGEMA_signal_13006, new_AGEMA_signal_13004}), .clk ( clk ), .rnd ({Fresh[3779], Fresh[3778], Fresh[3777], Fresh[3776], Fresh[3775], Fresh[3774], Fresh[3773], Fresh[3772], Fresh[3771], Fresh[3770]}), .outt ({new_AGEMA_signal_2360, new_AGEMA_signal_2359, new_AGEMA_signal_2358, n2433}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2587 ( .ina ({new_AGEMA_signal_12562, new_AGEMA_signal_12560, new_AGEMA_signal_12558, new_AGEMA_signal_12556}), .inb ({new_AGEMA_signal_1724, new_AGEMA_signal_1723, new_AGEMA_signal_1722, n2429}), .clk ( clk ), .rnd ({Fresh[3789], Fresh[3788], Fresh[3787], Fresh[3786], Fresh[3785], Fresh[3784], Fresh[3783], Fresh[3782], Fresh[3781], Fresh[3780]}), .outt ({new_AGEMA_signal_2363, new_AGEMA_signal_2362, new_AGEMA_signal_2361, n2689}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2591 ( .ina ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, new_AGEMA_signal_1359, n2647}), .inb ({new_AGEMA_signal_1232, new_AGEMA_signal_1231, new_AGEMA_signal_1230, n2492}), .clk ( clk ), .rnd ({Fresh[3799], Fresh[3798], Fresh[3797], Fresh[3796], Fresh[3795], Fresh[3794], Fresh[3793], Fresh[3792], Fresh[3791], Fresh[3790]}), .outt ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, new_AGEMA_signal_1887, n2434}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2595 ( .ina ({new_AGEMA_signal_1811, new_AGEMA_signal_1810, new_AGEMA_signal_1809, n2438}), .inb ({new_AGEMA_signal_1439, new_AGEMA_signal_1438, new_AGEMA_signal_1437, n2483}), .clk ( clk ), .rnd ({Fresh[3809], Fresh[3808], Fresh[3807], Fresh[3806], Fresh[3805], Fresh[3804], Fresh[3803], Fresh[3802], Fresh[3801], Fresh[3800]}), .outt ({new_AGEMA_signal_2369, new_AGEMA_signal_2368, new_AGEMA_signal_2367, n2439}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2598 ( .ina ({new_AGEMA_signal_12994, new_AGEMA_signal_12992, new_AGEMA_signal_12990, new_AGEMA_signal_12988}), .inb ({new_AGEMA_signal_1781, new_AGEMA_signal_1780, new_AGEMA_signal_1779, n2540}), .clk ( clk ), .rnd ({Fresh[3819], Fresh[3818], Fresh[3817], Fresh[3816], Fresh[3815], Fresh[3814], Fresh[3813], Fresh[3812], Fresh[3811], Fresh[3810]}), .outt ({new_AGEMA_signal_2372, new_AGEMA_signal_2371, new_AGEMA_signal_2370, n2445}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2600 ( .ina ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, new_AGEMA_signal_1299, n2690}), .inb ({new_AGEMA_signal_1892, new_AGEMA_signal_1891, new_AGEMA_signal_1890, n2443}), .clk ( clk ), .rnd ({Fresh[3829], Fresh[3828], Fresh[3827], Fresh[3826], Fresh[3825], Fresh[3824], Fresh[3823], Fresh[3822], Fresh[3821], Fresh[3820]}), .outt ({new_AGEMA_signal_2375, new_AGEMA_signal_2374, new_AGEMA_signal_2373, n2444}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2602 ( .ina ({new_AGEMA_signal_12658, new_AGEMA_signal_12656, new_AGEMA_signal_12654, new_AGEMA_signal_12652}), .inb ({new_AGEMA_signal_1742, new_AGEMA_signal_1741, new_AGEMA_signal_1740, n2446}), .clk ( clk ), .rnd ({Fresh[3839], Fresh[3838], Fresh[3837], Fresh[3836], Fresh[3835], Fresh[3834], Fresh[3833], Fresh[3832], Fresh[3831], Fresh[3830]}), .outt ({new_AGEMA_signal_2378, new_AGEMA_signal_2377, new_AGEMA_signal_2376, n2447}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2607 ( .ina ({new_AGEMA_signal_1550, new_AGEMA_signal_1549, new_AGEMA_signal_1548, n2761}), .inb ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, new_AGEMA_signal_1893, n2693}), .clk ( clk ), .rnd ({Fresh[3849], Fresh[3848], Fresh[3847], Fresh[3846], Fresh[3845], Fresh[3844], Fresh[3843], Fresh[3842], Fresh[3841], Fresh[3840]}), .outt ({new_AGEMA_signal_2381, new_AGEMA_signal_2380, new_AGEMA_signal_2379, n2454}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2617 ( .ina ({new_AGEMA_signal_12818, new_AGEMA_signal_12816, new_AGEMA_signal_12814, new_AGEMA_signal_12812}), .inb ({new_AGEMA_signal_1445, new_AGEMA_signal_1444, new_AGEMA_signal_1443, n2464}), .clk ( clk ), .rnd ({Fresh[3859], Fresh[3858], Fresh[3857], Fresh[3856], Fresh[3855], Fresh[3854], Fresh[3853], Fresh[3852], Fresh[3851], Fresh[3850]}), .outt ({new_AGEMA_signal_1898, new_AGEMA_signal_1897, new_AGEMA_signal_1896, n2465}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2622 ( .ina ({new_AGEMA_signal_12834, new_AGEMA_signal_12832, new_AGEMA_signal_12830, new_AGEMA_signal_12828}), .inb ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, new_AGEMA_signal_1377, n2576}), .clk ( clk ), .rnd ({Fresh[3869], Fresh[3868], Fresh[3867], Fresh[3866], Fresh[3865], Fresh[3864], Fresh[3863], Fresh[3862], Fresh[3861], Fresh[3860]}), .outt ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, new_AGEMA_signal_1899, n2470}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2626 ( .ina ({new_AGEMA_signal_1451, new_AGEMA_signal_1450, new_AGEMA_signal_1449, n2473}), .inb ({new_AGEMA_signal_1454, new_AGEMA_signal_1453, new_AGEMA_signal_1452, n2472}), .clk ( clk ), .rnd ({Fresh[3879], Fresh[3878], Fresh[3877], Fresh[3876], Fresh[3875], Fresh[3874], Fresh[3873], Fresh[3872], Fresh[3871], Fresh[3870]}), .outt ({new_AGEMA_signal_1904, new_AGEMA_signal_1903, new_AGEMA_signal_1902, n2476}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2633 ( .ina ({new_AGEMA_signal_13018, new_AGEMA_signal_13016, new_AGEMA_signal_13014, new_AGEMA_signal_13012}), .inb ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, new_AGEMA_signal_1905, n2480}), .clk ( clk ), .rnd ({Fresh[3889], Fresh[3888], Fresh[3887], Fresh[3886], Fresh[3885], Fresh[3884], Fresh[3883], Fresh[3882], Fresh[3881], Fresh[3880]}), .outt ({new_AGEMA_signal_2390, new_AGEMA_signal_2389, new_AGEMA_signal_2388, n2481}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2639 ( .ina ({new_AGEMA_signal_13026, new_AGEMA_signal_13024, new_AGEMA_signal_13022, new_AGEMA_signal_13020}), .inb ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, new_AGEMA_signal_1302, n2817}), .clk ( clk ), .rnd ({Fresh[3899], Fresh[3898], Fresh[3897], Fresh[3896], Fresh[3895], Fresh[3894], Fresh[3893], Fresh[3892], Fresh[3891], Fresh[3890]}), .outt ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, new_AGEMA_signal_1911, n2486}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2642 ( .ina ({new_AGEMA_signal_12922, new_AGEMA_signal_12920, new_AGEMA_signal_12918, new_AGEMA_signal_12916}), .inb ({new_AGEMA_signal_1460, new_AGEMA_signal_1459, new_AGEMA_signal_1458, n2488}), .clk ( clk ), .rnd ({Fresh[3909], Fresh[3908], Fresh[3907], Fresh[3906], Fresh[3905], Fresh[3904], Fresh[3903], Fresh[3902], Fresh[3901], Fresh[3900]}), .outt ({new_AGEMA_signal_1916, new_AGEMA_signal_1915, new_AGEMA_signal_1914, n2489}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2645 ( .ina ({new_AGEMA_signal_13034, new_AGEMA_signal_13032, new_AGEMA_signal_13030, new_AGEMA_signal_13028}), .inb ({new_AGEMA_signal_1232, new_AGEMA_signal_1231, new_AGEMA_signal_1230, n2492}), .clk ( clk ), .rnd ({Fresh[3919], Fresh[3918], Fresh[3917], Fresh[3916], Fresh[3915], Fresh[3914], Fresh[3913], Fresh[3912], Fresh[3911], Fresh[3910]}), .outt ({new_AGEMA_signal_1919, new_AGEMA_signal_1918, new_AGEMA_signal_1917, n2497}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2646 ( .ina ({new_AGEMA_signal_13042, new_AGEMA_signal_13040, new_AGEMA_signal_13038, new_AGEMA_signal_13036}), .inb ({new_AGEMA_signal_1430, new_AGEMA_signal_1429, new_AGEMA_signal_1428, n2700}), .clk ( clk ), .rnd ({Fresh[3929], Fresh[3928], Fresh[3927], Fresh[3926], Fresh[3925], Fresh[3924], Fresh[3923], Fresh[3922], Fresh[3921], Fresh[3920]}), .outt ({new_AGEMA_signal_1922, new_AGEMA_signal_1921, new_AGEMA_signal_1920, n2495}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2647 ( .ina ({new_AGEMA_signal_12826, new_AGEMA_signal_12824, new_AGEMA_signal_12822, new_AGEMA_signal_12820}), .inb ({new_AGEMA_signal_1562, new_AGEMA_signal_1561, new_AGEMA_signal_1560, n2625}), .clk ( clk ), .rnd ({Fresh[3939], Fresh[3938], Fresh[3937], Fresh[3936], Fresh[3935], Fresh[3934], Fresh[3933], Fresh[3932], Fresh[3931], Fresh[3930]}), .outt ({new_AGEMA_signal_2396, new_AGEMA_signal_2395, new_AGEMA_signal_2394, n2494}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2650 ( .ina ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, n2498}), .inb ({new_AGEMA_signal_12594, new_AGEMA_signal_12592, new_AGEMA_signal_12590, new_AGEMA_signal_12588}), .clk ( clk ), .rnd ({Fresh[3949], Fresh[3948], Fresh[3947], Fresh[3946], Fresh[3945], Fresh[3944], Fresh[3943], Fresh[3942], Fresh[3941], Fresh[3940]}), .outt ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, new_AGEMA_signal_1923, n2499}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2653 ( .ina ({new_AGEMA_signal_12594, new_AGEMA_signal_12592, new_AGEMA_signal_12590, new_AGEMA_signal_12588}), .inb ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, new_AGEMA_signal_2241, n2674}), .clk ( clk ), .rnd ({Fresh[3959], Fresh[3958], Fresh[3957], Fresh[3956], Fresh[3955], Fresh[3954], Fresh[3953], Fresh[3952], Fresh[3951], Fresh[3950]}), .outt ({new_AGEMA_signal_2789, new_AGEMA_signal_2788, new_AGEMA_signal_2787, n2503}) ) ;
    mux2_HPC1 #(.security_order(3), .pipeline(1)) U2655 ( .ins ({new_AGEMA_signal_12834, new_AGEMA_signal_12832, new_AGEMA_signal_12830, new_AGEMA_signal_12828}), .inb ({new_AGEMA_signal_1556, new_AGEMA_signal_1555, new_AGEMA_signal_1554, n2505}), .ina ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}), .clk ( clk ), .rnd ({Fresh[3969], Fresh[3968], Fresh[3967], Fresh[3966], Fresh[3965], Fresh[3964], Fresh[3963], Fresh[3962], Fresh[3961], Fresh[3960]}), .outt ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, new_AGEMA_signal_2397, n2506}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2662 ( .ina ({new_AGEMA_signal_1541, new_AGEMA_signal_1540, new_AGEMA_signal_1539, n2662}), .inb ({new_AGEMA_signal_12682, new_AGEMA_signal_12680, new_AGEMA_signal_12678, new_AGEMA_signal_12676}), .clk ( clk ), .rnd ({Fresh[3979], Fresh[3978], Fresh[3977], Fresh[3976], Fresh[3975], Fresh[3974], Fresh[3973], Fresh[3972], Fresh[3971], Fresh[3970]}), .outt ({new_AGEMA_signal_2402, new_AGEMA_signal_2401, new_AGEMA_signal_2400, n2518}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2663 ( .ina ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, new_AGEMA_signal_2085, n2720}), .inb ({new_AGEMA_signal_12738, new_AGEMA_signal_12736, new_AGEMA_signal_12734, new_AGEMA_signal_12732}), .clk ( clk ), .rnd ({Fresh[3989], Fresh[3988], Fresh[3987], Fresh[3986], Fresh[3985], Fresh[3984], Fresh[3983], Fresh[3982], Fresh[3981], Fresh[3980]}), .outt ({new_AGEMA_signal_2792, new_AGEMA_signal_2791, new_AGEMA_signal_2790, n2517}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2666 ( .ina ({new_AGEMA_signal_1928, new_AGEMA_signal_1927, new_AGEMA_signal_1926, n2520}), .inb ({new_AGEMA_signal_12874, new_AGEMA_signal_12872, new_AGEMA_signal_12870, new_AGEMA_signal_12868}), .clk ( clk ), .rnd ({Fresh[3999], Fresh[3998], Fresh[3997], Fresh[3996], Fresh[3995], Fresh[3994], Fresh[3993], Fresh[3992], Fresh[3991], Fresh[3990]}), .outt ({new_AGEMA_signal_2405, new_AGEMA_signal_2404, new_AGEMA_signal_2403, n2523}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2668 ( .ina ({new_AGEMA_signal_1802, new_AGEMA_signal_1801, new_AGEMA_signal_1800, n2774}), .inb ({new_AGEMA_signal_1463, new_AGEMA_signal_1462, new_AGEMA_signal_1461, n2521}), .clk ( clk ), .rnd ({Fresh[4009], Fresh[4008], Fresh[4007], Fresh[4006], Fresh[4005], Fresh[4004], Fresh[4003], Fresh[4002], Fresh[4001], Fresh[4000]}), .outt ({new_AGEMA_signal_2408, new_AGEMA_signal_2407, new_AGEMA_signal_2406, n2522}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2675 ( .ina ({new_AGEMA_signal_12682, new_AGEMA_signal_12680, new_AGEMA_signal_12678, new_AGEMA_signal_12676}), .inb ({new_AGEMA_signal_1931, new_AGEMA_signal_1930, new_AGEMA_signal_1929, n2531}), .clk ( clk ), .rnd ({Fresh[4019], Fresh[4018], Fresh[4017], Fresh[4016], Fresh[4015], Fresh[4014], Fresh[4013], Fresh[4012], Fresh[4011], Fresh[4010]}), .outt ({new_AGEMA_signal_2411, new_AGEMA_signal_2410, new_AGEMA_signal_2409, n2532}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2677 ( .ina ({new_AGEMA_signal_12554, new_AGEMA_signal_12552, new_AGEMA_signal_12550, new_AGEMA_signal_12548}), .inb ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, new_AGEMA_signal_1605, n2533}), .clk ( clk ), .rnd ({Fresh[4029], Fresh[4028], Fresh[4027], Fresh[4026], Fresh[4025], Fresh[4024], Fresh[4023], Fresh[4022], Fresh[4021], Fresh[4020]}), .outt ({new_AGEMA_signal_2414, new_AGEMA_signal_2413, new_AGEMA_signal_2412, n2534}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2681 ( .ina ({new_AGEMA_signal_13050, new_AGEMA_signal_13048, new_AGEMA_signal_13046, new_AGEMA_signal_13044}), .inb ({new_AGEMA_signal_1781, new_AGEMA_signal_1780, new_AGEMA_signal_1779, n2540}), .clk ( clk ), .rnd ({Fresh[4039], Fresh[4038], Fresh[4037], Fresh[4036], Fresh[4035], Fresh[4034], Fresh[4033], Fresh[4032], Fresh[4031], Fresh[4030]}), .outt ({new_AGEMA_signal_2417, new_AGEMA_signal_2416, new_AGEMA_signal_2415, n2542}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2683 ( .ina ({new_AGEMA_signal_1160, new_AGEMA_signal_1159, new_AGEMA_signal_1158, n2545}), .inb ({new_AGEMA_signal_1355, new_AGEMA_signal_1354, new_AGEMA_signal_1353, n2544}), .clk ( clk ), .rnd ({Fresh[4049], Fresh[4048], Fresh[4047], Fresh[4046], Fresh[4045], Fresh[4044], Fresh[4043], Fresh[4042], Fresh[4041], Fresh[4040]}), .outt ({new_AGEMA_signal_1934, new_AGEMA_signal_1933, new_AGEMA_signal_1932, n2546}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2687 ( .ina ({new_AGEMA_signal_1274, new_AGEMA_signal_1273, new_AGEMA_signal_1272, n2673}), .inb ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, new_AGEMA_signal_1521, n2732}), .clk ( clk ), .rnd ({Fresh[4059], Fresh[4058], Fresh[4057], Fresh[4056], Fresh[4055], Fresh[4054], Fresh[4053], Fresh[4052], Fresh[4051], Fresh[4050]}), .outt ({new_AGEMA_signal_2423, new_AGEMA_signal_2422, new_AGEMA_signal_2421, n2551}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2690 ( .ina ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, new_AGEMA_signal_1935, n2553}), .inb ({new_AGEMA_signal_13058, new_AGEMA_signal_13056, new_AGEMA_signal_13054, new_AGEMA_signal_13052}), .clk ( clk ), .rnd ({Fresh[4069], Fresh[4068], Fresh[4067], Fresh[4066], Fresh[4065], Fresh[4064], Fresh[4063], Fresh[4062], Fresh[4061], Fresh[4060]}), .outt ({new_AGEMA_signal_2426, new_AGEMA_signal_2425, new_AGEMA_signal_2424, n2558}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2692 ( .ina ({new_AGEMA_signal_1721, new_AGEMA_signal_1720, new_AGEMA_signal_1719, n2555}), .inb ({new_AGEMA_signal_1940, new_AGEMA_signal_1939, new_AGEMA_signal_1938, n2554}), .clk ( clk ), .rnd ({Fresh[4079], Fresh[4078], Fresh[4077], Fresh[4076], Fresh[4075], Fresh[4074], Fresh[4073], Fresh[4072], Fresh[4071], Fresh[4070]}), .outt ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, new_AGEMA_signal_2427, n2556}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2696 ( .ina ({new_AGEMA_signal_1772, new_AGEMA_signal_1771, new_AGEMA_signal_1770, n2561}), .inb ({new_AGEMA_signal_1466, new_AGEMA_signal_1465, new_AGEMA_signal_1464, n2560}), .clk ( clk ), .rnd ({Fresh[4089], Fresh[4088], Fresh[4087], Fresh[4086], Fresh[4085], Fresh[4084], Fresh[4083], Fresh[4082], Fresh[4081], Fresh[4080]}), .outt ({new_AGEMA_signal_2432, new_AGEMA_signal_2431, new_AGEMA_signal_2430, n2566}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2697 ( .ina ({new_AGEMA_signal_13066, new_AGEMA_signal_13064, new_AGEMA_signal_13062, new_AGEMA_signal_13060}), .inb ({new_AGEMA_signal_1676, new_AGEMA_signal_1675, new_AGEMA_signal_1674, n2562}), .clk ( clk ), .rnd ({Fresh[4099], Fresh[4098], Fresh[4097], Fresh[4096], Fresh[4095], Fresh[4094], Fresh[4093], Fresh[4092], Fresh[4091], Fresh[4090]}), .outt ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, new_AGEMA_signal_2433, n2715}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2703 ( .ina ({new_AGEMA_signal_1598, new_AGEMA_signal_1597, new_AGEMA_signal_1596, n2572}), .inb ({new_AGEMA_signal_1283, new_AGEMA_signal_1282, new_AGEMA_signal_1281, n2571}), .clk ( clk ), .rnd ({Fresh[4109], Fresh[4108], Fresh[4107], Fresh[4106], Fresh[4105], Fresh[4104], Fresh[4103], Fresh[4102], Fresh[4101], Fresh[4100]}), .outt ({new_AGEMA_signal_2438, new_AGEMA_signal_2437, new_AGEMA_signal_2436, n2573}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2705 ( .ina ({new_AGEMA_signal_13002, new_AGEMA_signal_13000, new_AGEMA_signal_12998, new_AGEMA_signal_12996}), .inb ({new_AGEMA_signal_1637, new_AGEMA_signal_1636, new_AGEMA_signal_1635, n2754}), .clk ( clk ), .rnd ({Fresh[4119], Fresh[4118], Fresh[4117], Fresh[4116], Fresh[4115], Fresh[4114], Fresh[4113], Fresh[4112], Fresh[4111], Fresh[4110]}), .outt ({new_AGEMA_signal_2441, new_AGEMA_signal_2440, new_AGEMA_signal_2439, n2585}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2706 ( .ina ({new_AGEMA_signal_12914, new_AGEMA_signal_12912, new_AGEMA_signal_12910, new_AGEMA_signal_12908}), .inb ({new_AGEMA_signal_1262, new_AGEMA_signal_1261, new_AGEMA_signal_1260, n2627}), .clk ( clk ), .rnd ({Fresh[4129], Fresh[4128], Fresh[4127], Fresh[4126], Fresh[4125], Fresh[4124], Fresh[4123], Fresh[4122], Fresh[4121], Fresh[4120]}), .outt ({new_AGEMA_signal_1946, new_AGEMA_signal_1945, new_AGEMA_signal_1944, n2581}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2707 ( .ina ({new_AGEMA_signal_1499, new_AGEMA_signal_1498, new_AGEMA_signal_1497, n2575}), .inb ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, new_AGEMA_signal_1302, n2817}), .clk ( clk ), .rnd ({Fresh[4139], Fresh[4138], Fresh[4137], Fresh[4136], Fresh[4135], Fresh[4134], Fresh[4133], Fresh[4132], Fresh[4131], Fresh[4130]}), .outt ({new_AGEMA_signal_2444, new_AGEMA_signal_2443, new_AGEMA_signal_2442, n2579}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2708 ( .ina ({new_AGEMA_signal_13042, new_AGEMA_signal_13040, new_AGEMA_signal_13038, new_AGEMA_signal_13036}), .inb ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, new_AGEMA_signal_1377, n2576}), .clk ( clk ), .rnd ({Fresh[4149], Fresh[4148], Fresh[4147], Fresh[4146], Fresh[4145], Fresh[4144], Fresh[4143], Fresh[4142], Fresh[4141], Fresh[4140]}), .outt ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, new_AGEMA_signal_1947, n2578}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2711 ( .ina ({new_AGEMA_signal_1562, new_AGEMA_signal_1561, new_AGEMA_signal_1560, n2625}), .inb ({new_AGEMA_signal_12882, new_AGEMA_signal_12880, new_AGEMA_signal_12878, new_AGEMA_signal_12876}), .clk ( clk ), .rnd ({Fresh[4159], Fresh[4158], Fresh[4157], Fresh[4156], Fresh[4155], Fresh[4154], Fresh[4153], Fresh[4152], Fresh[4151], Fresh[4150]}), .outt ({new_AGEMA_signal_2447, new_AGEMA_signal_2446, new_AGEMA_signal_2445, n2582}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2715 ( .ina ({new_AGEMA_signal_12626, new_AGEMA_signal_12624, new_AGEMA_signal_12622, new_AGEMA_signal_12620}), .inb ({new_AGEMA_signal_1952, new_AGEMA_signal_1951, new_AGEMA_signal_1950, n2586}), .clk ( clk ), .rnd ({Fresh[4169], Fresh[4168], Fresh[4167], Fresh[4166], Fresh[4165], Fresh[4164], Fresh[4163], Fresh[4162], Fresh[4161], Fresh[4160]}), .outt ({new_AGEMA_signal_2450, new_AGEMA_signal_2449, new_AGEMA_signal_2448, n2588}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2719 ( .ina ({new_AGEMA_signal_1433, new_AGEMA_signal_1432, new_AGEMA_signal_1431, n2594}), .inb ({new_AGEMA_signal_13002, new_AGEMA_signal_13000, new_AGEMA_signal_12998, new_AGEMA_signal_12996}), .clk ( clk ), .rnd ({Fresh[4179], Fresh[4178], Fresh[4177], Fresh[4176], Fresh[4175], Fresh[4174], Fresh[4173], Fresh[4172], Fresh[4171], Fresh[4170]}), .outt ({new_AGEMA_signal_1955, new_AGEMA_signal_1954, new_AGEMA_signal_1953, n2607}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2722 ( .ina ({new_AGEMA_signal_1469, new_AGEMA_signal_1468, new_AGEMA_signal_1467, n2597}), .inb ({new_AGEMA_signal_1958, new_AGEMA_signal_1957, new_AGEMA_signal_1956, n2596}), .clk ( clk ), .rnd ({Fresh[4189], Fresh[4188], Fresh[4187], Fresh[4186], Fresh[4185], Fresh[4184], Fresh[4183], Fresh[4182], Fresh[4181], Fresh[4180]}), .outt ({new_AGEMA_signal_2453, new_AGEMA_signal_2452, new_AGEMA_signal_2451, n2605}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2724 ( .ina ({new_AGEMA_signal_1961, new_AGEMA_signal_1960, new_AGEMA_signal_1959, n2598}), .inb ({new_AGEMA_signal_13074, new_AGEMA_signal_13072, new_AGEMA_signal_13070, new_AGEMA_signal_13068}), .clk ( clk ), .rnd ({Fresh[4199], Fresh[4198], Fresh[4197], Fresh[4196], Fresh[4195], Fresh[4194], Fresh[4193], Fresh[4192], Fresh[4191], Fresh[4190]}), .outt ({new_AGEMA_signal_2456, new_AGEMA_signal_2455, new_AGEMA_signal_2454, n2603}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2726 ( .ina ({new_AGEMA_signal_1181, new_AGEMA_signal_1180, new_AGEMA_signal_1179, n2599}), .inb ({new_AGEMA_signal_12906, new_AGEMA_signal_12904, new_AGEMA_signal_12902, new_AGEMA_signal_12900}), .clk ( clk ), .rnd ({Fresh[4209], Fresh[4208], Fresh[4207], Fresh[4206], Fresh[4205], Fresh[4204], Fresh[4203], Fresh[4202], Fresh[4201], Fresh[4200]}), .outt ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, new_AGEMA_signal_1470, n2601}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2733 ( .ina ({new_AGEMA_signal_1967, new_AGEMA_signal_1966, new_AGEMA_signal_1965, n2610}), .inb ({new_AGEMA_signal_12874, new_AGEMA_signal_12872, new_AGEMA_signal_12870, new_AGEMA_signal_12868}), .clk ( clk ), .rnd ({Fresh[4219], Fresh[4218], Fresh[4217], Fresh[4216], Fresh[4215], Fresh[4214], Fresh[4213], Fresh[4212], Fresh[4211], Fresh[4210]}), .outt ({new_AGEMA_signal_2459, new_AGEMA_signal_2458, new_AGEMA_signal_2457, n2620}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2736 ( .ina ({new_AGEMA_signal_1970, new_AGEMA_signal_1969, new_AGEMA_signal_1968, n2614}), .inb ({new_AGEMA_signal_1973, new_AGEMA_signal_1972, new_AGEMA_signal_1971, n2613}), .clk ( clk ), .rnd ({Fresh[4229], Fresh[4228], Fresh[4227], Fresh[4226], Fresh[4225], Fresh[4224], Fresh[4223], Fresh[4222], Fresh[4221], Fresh[4220]}), .outt ({new_AGEMA_signal_2462, new_AGEMA_signal_2461, new_AGEMA_signal_2460, n2618}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2743 ( .ina ({new_AGEMA_signal_12834, new_AGEMA_signal_12832, new_AGEMA_signal_12830, new_AGEMA_signal_12828}), .inb ({new_AGEMA_signal_1562, new_AGEMA_signal_1561, new_AGEMA_signal_1560, n2625}), .clk ( clk ), .rnd ({Fresh[4239], Fresh[4238], Fresh[4237], Fresh[4236], Fresh[4235], Fresh[4234], Fresh[4233], Fresh[4232], Fresh[4231], Fresh[4230]}), .outt ({new_AGEMA_signal_2465, new_AGEMA_signal_2464, new_AGEMA_signal_2463, n2626}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2746 ( .ina ({new_AGEMA_signal_1220, new_AGEMA_signal_1219, new_AGEMA_signal_1218, n2631}), .inb ({new_AGEMA_signal_12738, new_AGEMA_signal_12736, new_AGEMA_signal_12734, new_AGEMA_signal_12732}), .clk ( clk ), .rnd ({Fresh[4249], Fresh[4248], Fresh[4247], Fresh[4246], Fresh[4245], Fresh[4244], Fresh[4243], Fresh[4242], Fresh[4241], Fresh[4240]}), .outt ({new_AGEMA_signal_1976, new_AGEMA_signal_1975, new_AGEMA_signal_1974, n2632}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2752 ( .ina ({new_AGEMA_signal_1979, new_AGEMA_signal_1978, new_AGEMA_signal_1977, n2784}), .inb ({new_AGEMA_signal_1340, new_AGEMA_signal_1339, new_AGEMA_signal_1338, n2642}), .clk ( clk ), .rnd ({Fresh[4259], Fresh[4258], Fresh[4257], Fresh[4256], Fresh[4255], Fresh[4254], Fresh[4253], Fresh[4252], Fresh[4251], Fresh[4250]}), .outt ({new_AGEMA_signal_2468, new_AGEMA_signal_2467, new_AGEMA_signal_2466, n2644}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2754 ( .ina ({new_AGEMA_signal_12586, new_AGEMA_signal_12584, new_AGEMA_signal_12582, new_AGEMA_signal_12580}), .inb ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, new_AGEMA_signal_1395, n2645}), .clk ( clk ), .rnd ({Fresh[4269], Fresh[4268], Fresh[4267], Fresh[4266], Fresh[4265], Fresh[4264], Fresh[4263], Fresh[4262], Fresh[4261], Fresh[4260]}), .outt ({new_AGEMA_signal_1982, new_AGEMA_signal_1981, new_AGEMA_signal_1980, n2646}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2758 ( .ina ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}), .inb ({new_AGEMA_signal_1481, new_AGEMA_signal_1480, new_AGEMA_signal_1479, n2650}), .clk ( clk ), .rnd ({Fresh[4279], Fresh[4278], Fresh[4277], Fresh[4276], Fresh[4275], Fresh[4274], Fresh[4273], Fresh[4272], Fresh[4271], Fresh[4270]}), .outt ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, new_AGEMA_signal_1983, n2653}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2760 ( .ina ({new_AGEMA_signal_12906, new_AGEMA_signal_12904, new_AGEMA_signal_12902, new_AGEMA_signal_12900}), .inb ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, new_AGEMA_signal_1641, n2654}), .clk ( clk ), .rnd ({Fresh[4289], Fresh[4288], Fresh[4287], Fresh[4286], Fresh[4285], Fresh[4284], Fresh[4283], Fresh[4282], Fresh[4281], Fresh[4280]}), .outt ({new_AGEMA_signal_2474, new_AGEMA_signal_2473, new_AGEMA_signal_2472, n2655}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2764 ( .ina ({new_AGEMA_signal_1541, new_AGEMA_signal_1540, new_AGEMA_signal_1539, n2662}), .inb ({new_AGEMA_signal_12922, new_AGEMA_signal_12920, new_AGEMA_signal_12918, new_AGEMA_signal_12916}), .clk ( clk ), .rnd ({Fresh[4299], Fresh[4298], Fresh[4297], Fresh[4296], Fresh[4295], Fresh[4294], Fresh[4293], Fresh[4292], Fresh[4291], Fresh[4290]}), .outt ({new_AGEMA_signal_2477, new_AGEMA_signal_2476, new_AGEMA_signal_2475, n2663}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2770 ( .ina ({new_AGEMA_signal_1274, new_AGEMA_signal_1273, new_AGEMA_signal_1272, n2673}), .inb ({new_AGEMA_signal_12882, new_AGEMA_signal_12880, new_AGEMA_signal_12878, new_AGEMA_signal_12876}), .clk ( clk ), .rnd ({Fresh[4309], Fresh[4308], Fresh[4307], Fresh[4306], Fresh[4305], Fresh[4304], Fresh[4303], Fresh[4302], Fresh[4301], Fresh[4300]}), .outt ({new_AGEMA_signal_1988, new_AGEMA_signal_1987, new_AGEMA_signal_1986, n2675}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2772 ( .ina ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, new_AGEMA_signal_1257, n2677}), .inb ({new_AGEMA_signal_1247, new_AGEMA_signal_1246, new_AGEMA_signal_1245, n2676}), .clk ( clk ), .rnd ({Fresh[4319], Fresh[4318], Fresh[4317], Fresh[4316], Fresh[4315], Fresh[4314], Fresh[4313], Fresh[4312], Fresh[4311], Fresh[4310]}), .outt ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, new_AGEMA_signal_1989, n2678}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2780 ( .ina ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, new_AGEMA_signal_1299, n2690}), .inb ({new_AGEMA_signal_12914, new_AGEMA_signal_12912, new_AGEMA_signal_12910, new_AGEMA_signal_12908}), .clk ( clk ), .rnd ({Fresh[4329], Fresh[4328], Fresh[4327], Fresh[4326], Fresh[4325], Fresh[4324], Fresh[4323], Fresh[4322], Fresh[4321], Fresh[4320]}), .outt ({new_AGEMA_signal_1994, new_AGEMA_signal_1993, new_AGEMA_signal_1992, n2691}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2782 ( .ina ({new_AGEMA_signal_12938, new_AGEMA_signal_12936, new_AGEMA_signal_12934, new_AGEMA_signal_12932}), .inb ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, new_AGEMA_signal_1893, n2693}), .clk ( clk ), .rnd ({Fresh[4339], Fresh[4338], Fresh[4337], Fresh[4336], Fresh[4335], Fresh[4334], Fresh[4333], Fresh[4332], Fresh[4331], Fresh[4330]}), .outt ({new_AGEMA_signal_2483, new_AGEMA_signal_2482, new_AGEMA_signal_2481, n2695}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2785 ( .ina ({new_AGEMA_signal_1430, new_AGEMA_signal_1429, new_AGEMA_signal_1428, n2700}), .inb ({new_AGEMA_signal_13066, new_AGEMA_signal_13064, new_AGEMA_signal_13062, new_AGEMA_signal_13060}), .clk ( clk ), .rnd ({Fresh[4349], Fresh[4348], Fresh[4347], Fresh[4346], Fresh[4345], Fresh[4344], Fresh[4343], Fresh[4342], Fresh[4341], Fresh[4340]}), .outt ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, new_AGEMA_signal_1995, n2701}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2791 ( .ina ({new_AGEMA_signal_2000, new_AGEMA_signal_1999, new_AGEMA_signal_1998, n2711}), .inb ({new_AGEMA_signal_2003, new_AGEMA_signal_2002, new_AGEMA_signal_2001, n2710}), .clk ( clk ), .rnd ({Fresh[4359], Fresh[4358], Fresh[4357], Fresh[4356], Fresh[4355], Fresh[4354], Fresh[4353], Fresh[4352], Fresh[4351], Fresh[4350]}), .outt ({new_AGEMA_signal_2486, new_AGEMA_signal_2485, new_AGEMA_signal_2484, n2717}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2796 ( .ina ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, new_AGEMA_signal_2085, n2720}), .inb ({new_AGEMA_signal_12834, new_AGEMA_signal_12832, new_AGEMA_signal_12830, new_AGEMA_signal_12828}), .clk ( clk ), .rnd ({Fresh[4369], Fresh[4368], Fresh[4367], Fresh[4366], Fresh[4365], Fresh[4364], Fresh[4363], Fresh[4362], Fresh[4361], Fresh[4360]}), .outt ({new_AGEMA_signal_2846, new_AGEMA_signal_2845, new_AGEMA_signal_2844, n2729}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2798 ( .ina ({new_AGEMA_signal_12698, new_AGEMA_signal_12696, new_AGEMA_signal_12694, new_AGEMA_signal_12692}), .inb ({new_AGEMA_signal_1487, new_AGEMA_signal_1486, new_AGEMA_signal_1485, n2722}), .clk ( clk ), .rnd ({Fresh[4379], Fresh[4378], Fresh[4377], Fresh[4376], Fresh[4375], Fresh[4374], Fresh[4373], Fresh[4372], Fresh[4371], Fresh[4370]}), .outt ({new_AGEMA_signal_2006, new_AGEMA_signal_2005, new_AGEMA_signal_2004, n2727}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2803 ( .ina ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, new_AGEMA_signal_1521, n2732}), .inb ({new_AGEMA_signal_1658, new_AGEMA_signal_1657, new_AGEMA_signal_1656, n2731}), .clk ( clk ), .rnd ({Fresh[4389], Fresh[4388], Fresh[4387], Fresh[4386], Fresh[4385], Fresh[4384], Fresh[4383], Fresh[4382], Fresh[4381], Fresh[4380]}), .outt ({new_AGEMA_signal_2492, new_AGEMA_signal_2491, new_AGEMA_signal_2490, n2733}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2807 ( .ina ({new_AGEMA_signal_13082, new_AGEMA_signal_13080, new_AGEMA_signal_13078, new_AGEMA_signal_13076}), .inb ({new_AGEMA_signal_2012, new_AGEMA_signal_2011, new_AGEMA_signal_2010, n2738}), .clk ( clk ), .rnd ({Fresh[4399], Fresh[4398], Fresh[4397], Fresh[4396], Fresh[4395], Fresh[4394], Fresh[4393], Fresh[4392], Fresh[4391], Fresh[4390]}), .outt ({new_AGEMA_signal_2495, new_AGEMA_signal_2494, new_AGEMA_signal_2493, n2740}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2812 ( .ina ({new_AGEMA_signal_1382, new_AGEMA_signal_1381, new_AGEMA_signal_1380, n2748}), .inb ({new_AGEMA_signal_12554, new_AGEMA_signal_12552, new_AGEMA_signal_12550, new_AGEMA_signal_12548}), .clk ( clk ), .rnd ({Fresh[4409], Fresh[4408], Fresh[4407], Fresh[4406], Fresh[4405], Fresh[4404], Fresh[4403], Fresh[4402], Fresh[4401], Fresh[4400]}), .outt ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, new_AGEMA_signal_2013, n2749}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2815 ( .ina ({new_AGEMA_signal_1637, new_AGEMA_signal_1636, new_AGEMA_signal_1635, n2754}), .inb ({new_AGEMA_signal_12714, new_AGEMA_signal_12712, new_AGEMA_signal_12710, new_AGEMA_signal_12708}), .clk ( clk ), .rnd ({Fresh[4419], Fresh[4418], Fresh[4417], Fresh[4416], Fresh[4415], Fresh[4414], Fresh[4413], Fresh[4412], Fresh[4411], Fresh[4410]}), .outt ({new_AGEMA_signal_2501, new_AGEMA_signal_2500, new_AGEMA_signal_2499, n2757}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2816 ( .ina ({new_AGEMA_signal_1208, new_AGEMA_signal_1207, new_AGEMA_signal_1206, n2755}), .inb ({new_AGEMA_signal_13090, new_AGEMA_signal_13088, new_AGEMA_signal_13086, new_AGEMA_signal_13084}), .clk ( clk ), .rnd ({Fresh[4429], Fresh[4428], Fresh[4427], Fresh[4426], Fresh[4425], Fresh[4424], Fresh[4423], Fresh[4422], Fresh[4421], Fresh[4420]}), .outt ({new_AGEMA_signal_2018, new_AGEMA_signal_2017, new_AGEMA_signal_2016, n2756}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2819 ( .ina ({new_AGEMA_signal_1550, new_AGEMA_signal_1549, new_AGEMA_signal_1548, n2761}), .inb ({new_AGEMA_signal_12946, new_AGEMA_signal_12944, new_AGEMA_signal_12942, new_AGEMA_signal_12940}), .clk ( clk ), .rnd ({Fresh[4439], Fresh[4438], Fresh[4437], Fresh[4436], Fresh[4435], Fresh[4434], Fresh[4433], Fresh[4432], Fresh[4431], Fresh[4430]}), .outt ({new_AGEMA_signal_2504, new_AGEMA_signal_2503, new_AGEMA_signal_2502, n2762}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2823 ( .ina ({new_AGEMA_signal_12554, new_AGEMA_signal_12552, new_AGEMA_signal_12550, new_AGEMA_signal_12548}), .inb ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, new_AGEMA_signal_2019, n2768}), .clk ( clk ), .rnd ({Fresh[4449], Fresh[4448], Fresh[4447], Fresh[4446], Fresh[4445], Fresh[4444], Fresh[4443], Fresh[4442], Fresh[4441], Fresh[4440]}), .outt ({new_AGEMA_signal_2507, new_AGEMA_signal_2506, new_AGEMA_signal_2505, n2770}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2825 ( .ina ({new_AGEMA_signal_1670, new_AGEMA_signal_1669, new_AGEMA_signal_1668, n2773}), .inb ({new_AGEMA_signal_13090, new_AGEMA_signal_13088, new_AGEMA_signal_13086, new_AGEMA_signal_13084}), .clk ( clk ), .rnd ({Fresh[4459], Fresh[4458], Fresh[4457], Fresh[4456], Fresh[4455], Fresh[4454], Fresh[4453], Fresh[4452], Fresh[4451], Fresh[4450]}), .outt ({new_AGEMA_signal_2510, new_AGEMA_signal_2509, new_AGEMA_signal_2508, n2776}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2826 ( .ina ({new_AGEMA_signal_1802, new_AGEMA_signal_1801, new_AGEMA_signal_1800, n2774}), .inb ({new_AGEMA_signal_12562, new_AGEMA_signal_12560, new_AGEMA_signal_12558, new_AGEMA_signal_12556}), .clk ( clk ), .rnd ({Fresh[4469], Fresh[4468], Fresh[4467], Fresh[4466], Fresh[4465], Fresh[4464], Fresh[4463], Fresh[4462], Fresh[4461], Fresh[4460]}), .outt ({new_AGEMA_signal_2513, new_AGEMA_signal_2512, new_AGEMA_signal_2511, n2775}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2830 ( .ina ({new_AGEMA_signal_1490, new_AGEMA_signal_1489, new_AGEMA_signal_1488, n2782}), .inb ({new_AGEMA_signal_1493, new_AGEMA_signal_1492, new_AGEMA_signal_1491, n2781}), .clk ( clk ), .rnd ({Fresh[4479], Fresh[4478], Fresh[4477], Fresh[4476], Fresh[4475], Fresh[4474], Fresh[4473], Fresh[4472], Fresh[4471], Fresh[4470]}), .outt ({new_AGEMA_signal_2024, new_AGEMA_signal_2023, new_AGEMA_signal_2022, n2783}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2836 ( .ina ({new_AGEMA_signal_2030, new_AGEMA_signal_2029, new_AGEMA_signal_2028, n2794}), .inb ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, new_AGEMA_signal_2031, n2793}), .clk ( clk ), .rnd ({Fresh[4489], Fresh[4488], Fresh[4487], Fresh[4486], Fresh[4485], Fresh[4484], Fresh[4483], Fresh[4482], Fresh[4481], Fresh[4480]}), .outt ({new_AGEMA_signal_2519, new_AGEMA_signal_2518, new_AGEMA_signal_2517, n2795}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2845 ( .ina ({new_AGEMA_signal_2036, new_AGEMA_signal_2035, new_AGEMA_signal_2034, n2812}), .inb ({new_AGEMA_signal_1700, new_AGEMA_signal_1699, new_AGEMA_signal_1698, n2811}), .clk ( clk ), .rnd ({Fresh[4499], Fresh[4498], Fresh[4497], Fresh[4496], Fresh[4495], Fresh[4494], Fresh[4493], Fresh[4492], Fresh[4491], Fresh[4490]}), .outt ({new_AGEMA_signal_2522, new_AGEMA_signal_2521, new_AGEMA_signal_2520, n2814}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2848 ( .ina ({new_AGEMA_signal_12650, new_AGEMA_signal_12648, new_AGEMA_signal_12646, new_AGEMA_signal_12644}), .inb ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, new_AGEMA_signal_1302, n2817}), .clk ( clk ), .rnd ({Fresh[4509], Fresh[4508], Fresh[4507], Fresh[4506], Fresh[4505], Fresh[4504], Fresh[4503], Fresh[4502], Fresh[4501], Fresh[4500]}), .outt ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, new_AGEMA_signal_2037, n2819}) ) ;
    buf_clk new_AGEMA_reg_buffer_1592 ( .C ( clk ), .D ( new_AGEMA_signal_13091 ), .Q ( new_AGEMA_signal_13092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1594 ( .C ( clk ), .D ( new_AGEMA_signal_13093 ), .Q ( new_AGEMA_signal_13094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1596 ( .C ( clk ), .D ( new_AGEMA_signal_13095 ), .Q ( new_AGEMA_signal_13096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1598 ( .C ( clk ), .D ( new_AGEMA_signal_13097 ), .Q ( new_AGEMA_signal_13098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1600 ( .C ( clk ), .D ( new_AGEMA_signal_13099 ), .Q ( new_AGEMA_signal_13100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1602 ( .C ( clk ), .D ( new_AGEMA_signal_13101 ), .Q ( new_AGEMA_signal_13102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1604 ( .C ( clk ), .D ( new_AGEMA_signal_13103 ), .Q ( new_AGEMA_signal_13104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1606 ( .C ( clk ), .D ( new_AGEMA_signal_13105 ), .Q ( new_AGEMA_signal_13106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1610 ( .C ( clk ), .D ( new_AGEMA_signal_13109 ), .Q ( new_AGEMA_signal_13110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1614 ( .C ( clk ), .D ( new_AGEMA_signal_13113 ), .Q ( new_AGEMA_signal_13114 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1618 ( .C ( clk ), .D ( new_AGEMA_signal_13117 ), .Q ( new_AGEMA_signal_13118 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1622 ( .C ( clk ), .D ( new_AGEMA_signal_13121 ), .Q ( new_AGEMA_signal_13122 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1624 ( .C ( clk ), .D ( new_AGEMA_signal_13123 ), .Q ( new_AGEMA_signal_13124 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1626 ( .C ( clk ), .D ( new_AGEMA_signal_13125 ), .Q ( new_AGEMA_signal_13126 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1628 ( .C ( clk ), .D ( new_AGEMA_signal_13127 ), .Q ( new_AGEMA_signal_13128 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1630 ( .C ( clk ), .D ( new_AGEMA_signal_13129 ), .Q ( new_AGEMA_signal_13130 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1632 ( .C ( clk ), .D ( new_AGEMA_signal_13131 ), .Q ( new_AGEMA_signal_13132 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1634 ( .C ( clk ), .D ( new_AGEMA_signal_13133 ), .Q ( new_AGEMA_signal_13134 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1636 ( .C ( clk ), .D ( new_AGEMA_signal_13135 ), .Q ( new_AGEMA_signal_13136 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1638 ( .C ( clk ), .D ( new_AGEMA_signal_13137 ), .Q ( new_AGEMA_signal_13138 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1640 ( .C ( clk ), .D ( new_AGEMA_signal_13139 ), .Q ( new_AGEMA_signal_13140 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1642 ( .C ( clk ), .D ( new_AGEMA_signal_13141 ), .Q ( new_AGEMA_signal_13142 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1644 ( .C ( clk ), .D ( new_AGEMA_signal_13143 ), .Q ( new_AGEMA_signal_13144 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1646 ( .C ( clk ), .D ( new_AGEMA_signal_13145 ), .Q ( new_AGEMA_signal_13146 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1648 ( .C ( clk ), .D ( new_AGEMA_signal_13147 ), .Q ( new_AGEMA_signal_13148 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1650 ( .C ( clk ), .D ( new_AGEMA_signal_13149 ), .Q ( new_AGEMA_signal_13150 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1652 ( .C ( clk ), .D ( new_AGEMA_signal_13151 ), .Q ( new_AGEMA_signal_13152 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1654 ( .C ( clk ), .D ( new_AGEMA_signal_13153 ), .Q ( new_AGEMA_signal_13154 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1656 ( .C ( clk ), .D ( new_AGEMA_signal_13155 ), .Q ( new_AGEMA_signal_13156 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1658 ( .C ( clk ), .D ( new_AGEMA_signal_13157 ), .Q ( new_AGEMA_signal_13158 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1660 ( .C ( clk ), .D ( new_AGEMA_signal_13159 ), .Q ( new_AGEMA_signal_13160 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1662 ( .C ( clk ), .D ( new_AGEMA_signal_13161 ), .Q ( new_AGEMA_signal_13162 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1664 ( .C ( clk ), .D ( new_AGEMA_signal_13163 ), .Q ( new_AGEMA_signal_13164 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1666 ( .C ( clk ), .D ( new_AGEMA_signal_13165 ), .Q ( new_AGEMA_signal_13166 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1668 ( .C ( clk ), .D ( new_AGEMA_signal_13167 ), .Q ( new_AGEMA_signal_13168 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1670 ( .C ( clk ), .D ( new_AGEMA_signal_13169 ), .Q ( new_AGEMA_signal_13170 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1672 ( .C ( clk ), .D ( new_AGEMA_signal_13171 ), .Q ( new_AGEMA_signal_13172 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1674 ( .C ( clk ), .D ( new_AGEMA_signal_13173 ), .Q ( new_AGEMA_signal_13174 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1676 ( .C ( clk ), .D ( new_AGEMA_signal_13175 ), .Q ( new_AGEMA_signal_13176 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1678 ( .C ( clk ), .D ( new_AGEMA_signal_13177 ), .Q ( new_AGEMA_signal_13178 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1680 ( .C ( clk ), .D ( new_AGEMA_signal_13179 ), .Q ( new_AGEMA_signal_13180 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1682 ( .C ( clk ), .D ( new_AGEMA_signal_13181 ), .Q ( new_AGEMA_signal_13182 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1684 ( .C ( clk ), .D ( new_AGEMA_signal_13183 ), .Q ( new_AGEMA_signal_13184 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1686 ( .C ( clk ), .D ( new_AGEMA_signal_13185 ), .Q ( new_AGEMA_signal_13186 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1688 ( .C ( clk ), .D ( new_AGEMA_signal_13187 ), .Q ( new_AGEMA_signal_13188 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1690 ( .C ( clk ), .D ( new_AGEMA_signal_13189 ), .Q ( new_AGEMA_signal_13190 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1692 ( .C ( clk ), .D ( new_AGEMA_signal_13191 ), .Q ( new_AGEMA_signal_13192 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1694 ( .C ( clk ), .D ( new_AGEMA_signal_13193 ), .Q ( new_AGEMA_signal_13194 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1696 ( .C ( clk ), .D ( new_AGEMA_signal_13195 ), .Q ( new_AGEMA_signal_13196 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1698 ( .C ( clk ), .D ( new_AGEMA_signal_13197 ), .Q ( new_AGEMA_signal_13198 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1700 ( .C ( clk ), .D ( new_AGEMA_signal_13199 ), .Q ( new_AGEMA_signal_13200 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1702 ( .C ( clk ), .D ( new_AGEMA_signal_13201 ), .Q ( new_AGEMA_signal_13202 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1704 ( .C ( clk ), .D ( new_AGEMA_signal_13203 ), .Q ( new_AGEMA_signal_13204 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1706 ( .C ( clk ), .D ( new_AGEMA_signal_13205 ), .Q ( new_AGEMA_signal_13206 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1708 ( .C ( clk ), .D ( new_AGEMA_signal_13207 ), .Q ( new_AGEMA_signal_13208 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1710 ( .C ( clk ), .D ( new_AGEMA_signal_13209 ), .Q ( new_AGEMA_signal_13210 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1714 ( .C ( clk ), .D ( new_AGEMA_signal_13213 ), .Q ( new_AGEMA_signal_13214 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1718 ( .C ( clk ), .D ( new_AGEMA_signal_13217 ), .Q ( new_AGEMA_signal_13218 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1722 ( .C ( clk ), .D ( new_AGEMA_signal_13221 ), .Q ( new_AGEMA_signal_13222 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1726 ( .C ( clk ), .D ( new_AGEMA_signal_13225 ), .Q ( new_AGEMA_signal_13226 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1728 ( .C ( clk ), .D ( new_AGEMA_signal_13227 ), .Q ( new_AGEMA_signal_13228 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1730 ( .C ( clk ), .D ( new_AGEMA_signal_13229 ), .Q ( new_AGEMA_signal_13230 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1732 ( .C ( clk ), .D ( new_AGEMA_signal_13231 ), .Q ( new_AGEMA_signal_13232 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1734 ( .C ( clk ), .D ( new_AGEMA_signal_13233 ), .Q ( new_AGEMA_signal_13234 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1736 ( .C ( clk ), .D ( new_AGEMA_signal_13235 ), .Q ( new_AGEMA_signal_13236 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1738 ( .C ( clk ), .D ( new_AGEMA_signal_13237 ), .Q ( new_AGEMA_signal_13238 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1740 ( .C ( clk ), .D ( new_AGEMA_signal_13239 ), .Q ( new_AGEMA_signal_13240 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1742 ( .C ( clk ), .D ( new_AGEMA_signal_13241 ), .Q ( new_AGEMA_signal_13242 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1744 ( .C ( clk ), .D ( new_AGEMA_signal_13243 ), .Q ( new_AGEMA_signal_13244 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1746 ( .C ( clk ), .D ( new_AGEMA_signal_13245 ), .Q ( new_AGEMA_signal_13246 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1748 ( .C ( clk ), .D ( new_AGEMA_signal_13247 ), .Q ( new_AGEMA_signal_13248 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1750 ( .C ( clk ), .D ( new_AGEMA_signal_13249 ), .Q ( new_AGEMA_signal_13250 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1752 ( .C ( clk ), .D ( new_AGEMA_signal_13251 ), .Q ( new_AGEMA_signal_13252 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1754 ( .C ( clk ), .D ( new_AGEMA_signal_13253 ), .Q ( new_AGEMA_signal_13254 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1756 ( .C ( clk ), .D ( new_AGEMA_signal_13255 ), .Q ( new_AGEMA_signal_13256 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1758 ( .C ( clk ), .D ( new_AGEMA_signal_13257 ), .Q ( new_AGEMA_signal_13258 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1760 ( .C ( clk ), .D ( new_AGEMA_signal_13259 ), .Q ( new_AGEMA_signal_13260 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1762 ( .C ( clk ), .D ( new_AGEMA_signal_13261 ), .Q ( new_AGEMA_signal_13262 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1764 ( .C ( clk ), .D ( new_AGEMA_signal_13263 ), .Q ( new_AGEMA_signal_13264 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1766 ( .C ( clk ), .D ( new_AGEMA_signal_13265 ), .Q ( new_AGEMA_signal_13266 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1768 ( .C ( clk ), .D ( new_AGEMA_signal_13267 ), .Q ( new_AGEMA_signal_13268 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1770 ( .C ( clk ), .D ( new_AGEMA_signal_13269 ), .Q ( new_AGEMA_signal_13270 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1772 ( .C ( clk ), .D ( new_AGEMA_signal_13271 ), .Q ( new_AGEMA_signal_13272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1774 ( .C ( clk ), .D ( new_AGEMA_signal_13273 ), .Q ( new_AGEMA_signal_13274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1776 ( .C ( clk ), .D ( new_AGEMA_signal_13275 ), .Q ( new_AGEMA_signal_13276 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1778 ( .C ( clk ), .D ( new_AGEMA_signal_13277 ), .Q ( new_AGEMA_signal_13278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1780 ( .C ( clk ), .D ( new_AGEMA_signal_13279 ), .Q ( new_AGEMA_signal_13280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1782 ( .C ( clk ), .D ( new_AGEMA_signal_13281 ), .Q ( new_AGEMA_signal_13282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1786 ( .C ( clk ), .D ( new_AGEMA_signal_13285 ), .Q ( new_AGEMA_signal_13286 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1790 ( .C ( clk ), .D ( new_AGEMA_signal_13289 ), .Q ( new_AGEMA_signal_13290 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1794 ( .C ( clk ), .D ( new_AGEMA_signal_13293 ), .Q ( new_AGEMA_signal_13294 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1798 ( .C ( clk ), .D ( new_AGEMA_signal_13297 ), .Q ( new_AGEMA_signal_13298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1800 ( .C ( clk ), .D ( new_AGEMA_signal_13299 ), .Q ( new_AGEMA_signal_13300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1802 ( .C ( clk ), .D ( new_AGEMA_signal_13301 ), .Q ( new_AGEMA_signal_13302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1804 ( .C ( clk ), .D ( new_AGEMA_signal_13303 ), .Q ( new_AGEMA_signal_13304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1806 ( .C ( clk ), .D ( new_AGEMA_signal_13305 ), .Q ( new_AGEMA_signal_13306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1808 ( .C ( clk ), .D ( new_AGEMA_signal_13307 ), .Q ( new_AGEMA_signal_13308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1810 ( .C ( clk ), .D ( new_AGEMA_signal_13309 ), .Q ( new_AGEMA_signal_13310 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1812 ( .C ( clk ), .D ( new_AGEMA_signal_13311 ), .Q ( new_AGEMA_signal_13312 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1814 ( .C ( clk ), .D ( new_AGEMA_signal_13313 ), .Q ( new_AGEMA_signal_13314 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1816 ( .C ( clk ), .D ( new_AGEMA_signal_13315 ), .Q ( new_AGEMA_signal_13316 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1818 ( .C ( clk ), .D ( new_AGEMA_signal_13317 ), .Q ( new_AGEMA_signal_13318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1820 ( .C ( clk ), .D ( new_AGEMA_signal_13319 ), .Q ( new_AGEMA_signal_13320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1822 ( .C ( clk ), .D ( new_AGEMA_signal_13321 ), .Q ( new_AGEMA_signal_13322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1824 ( .C ( clk ), .D ( new_AGEMA_signal_13323 ), .Q ( new_AGEMA_signal_13324 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1826 ( .C ( clk ), .D ( new_AGEMA_signal_13325 ), .Q ( new_AGEMA_signal_13326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1828 ( .C ( clk ), .D ( new_AGEMA_signal_13327 ), .Q ( new_AGEMA_signal_13328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1830 ( .C ( clk ), .D ( new_AGEMA_signal_13329 ), .Q ( new_AGEMA_signal_13330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1832 ( .C ( clk ), .D ( new_AGEMA_signal_13331 ), .Q ( new_AGEMA_signal_13332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1834 ( .C ( clk ), .D ( new_AGEMA_signal_13333 ), .Q ( new_AGEMA_signal_13334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1836 ( .C ( clk ), .D ( new_AGEMA_signal_13335 ), .Q ( new_AGEMA_signal_13336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1838 ( .C ( clk ), .D ( new_AGEMA_signal_13337 ), .Q ( new_AGEMA_signal_13338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1842 ( .C ( clk ), .D ( new_AGEMA_signal_13341 ), .Q ( new_AGEMA_signal_13342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1846 ( .C ( clk ), .D ( new_AGEMA_signal_13345 ), .Q ( new_AGEMA_signal_13346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1850 ( .C ( clk ), .D ( new_AGEMA_signal_13349 ), .Q ( new_AGEMA_signal_13350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1854 ( .C ( clk ), .D ( new_AGEMA_signal_13353 ), .Q ( new_AGEMA_signal_13354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1856 ( .C ( clk ), .D ( new_AGEMA_signal_13355 ), .Q ( new_AGEMA_signal_13356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1858 ( .C ( clk ), .D ( new_AGEMA_signal_13357 ), .Q ( new_AGEMA_signal_13358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1860 ( .C ( clk ), .D ( new_AGEMA_signal_13359 ), .Q ( new_AGEMA_signal_13360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1862 ( .C ( clk ), .D ( new_AGEMA_signal_13361 ), .Q ( new_AGEMA_signal_13362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1864 ( .C ( clk ), .D ( new_AGEMA_signal_13363 ), .Q ( new_AGEMA_signal_13364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1866 ( .C ( clk ), .D ( new_AGEMA_signal_13365 ), .Q ( new_AGEMA_signal_13366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1868 ( .C ( clk ), .D ( new_AGEMA_signal_13367 ), .Q ( new_AGEMA_signal_13368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1870 ( .C ( clk ), .D ( new_AGEMA_signal_13369 ), .Q ( new_AGEMA_signal_13370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1872 ( .C ( clk ), .D ( new_AGEMA_signal_13371 ), .Q ( new_AGEMA_signal_13372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1874 ( .C ( clk ), .D ( new_AGEMA_signal_13373 ), .Q ( new_AGEMA_signal_13374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1876 ( .C ( clk ), .D ( new_AGEMA_signal_13375 ), .Q ( new_AGEMA_signal_13376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1878 ( .C ( clk ), .D ( new_AGEMA_signal_13377 ), .Q ( new_AGEMA_signal_13378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1882 ( .C ( clk ), .D ( new_AGEMA_signal_13381 ), .Q ( new_AGEMA_signal_13382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1886 ( .C ( clk ), .D ( new_AGEMA_signal_13385 ), .Q ( new_AGEMA_signal_13386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1890 ( .C ( clk ), .D ( new_AGEMA_signal_13389 ), .Q ( new_AGEMA_signal_13390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1894 ( .C ( clk ), .D ( new_AGEMA_signal_13393 ), .Q ( new_AGEMA_signal_13394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1896 ( .C ( clk ), .D ( new_AGEMA_signal_13395 ), .Q ( new_AGEMA_signal_13396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1898 ( .C ( clk ), .D ( new_AGEMA_signal_13397 ), .Q ( new_AGEMA_signal_13398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1900 ( .C ( clk ), .D ( new_AGEMA_signal_13399 ), .Q ( new_AGEMA_signal_13400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1902 ( .C ( clk ), .D ( new_AGEMA_signal_13401 ), .Q ( new_AGEMA_signal_13402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1904 ( .C ( clk ), .D ( new_AGEMA_signal_13403 ), .Q ( new_AGEMA_signal_13404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1906 ( .C ( clk ), .D ( new_AGEMA_signal_13405 ), .Q ( new_AGEMA_signal_13406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1908 ( .C ( clk ), .D ( new_AGEMA_signal_13407 ), .Q ( new_AGEMA_signal_13408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1910 ( .C ( clk ), .D ( new_AGEMA_signal_13409 ), .Q ( new_AGEMA_signal_13410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1912 ( .C ( clk ), .D ( new_AGEMA_signal_13411 ), .Q ( new_AGEMA_signal_13412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1914 ( .C ( clk ), .D ( new_AGEMA_signal_13413 ), .Q ( new_AGEMA_signal_13414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1916 ( .C ( clk ), .D ( new_AGEMA_signal_13415 ), .Q ( new_AGEMA_signal_13416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1918 ( .C ( clk ), .D ( new_AGEMA_signal_13417 ), .Q ( new_AGEMA_signal_13418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1922 ( .C ( clk ), .D ( new_AGEMA_signal_13421 ), .Q ( new_AGEMA_signal_13422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1926 ( .C ( clk ), .D ( new_AGEMA_signal_13425 ), .Q ( new_AGEMA_signal_13426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1930 ( .C ( clk ), .D ( new_AGEMA_signal_13429 ), .Q ( new_AGEMA_signal_13430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1934 ( .C ( clk ), .D ( new_AGEMA_signal_13433 ), .Q ( new_AGEMA_signal_13434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1936 ( .C ( clk ), .D ( new_AGEMA_signal_13435 ), .Q ( new_AGEMA_signal_13436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1938 ( .C ( clk ), .D ( new_AGEMA_signal_13437 ), .Q ( new_AGEMA_signal_13438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1940 ( .C ( clk ), .D ( new_AGEMA_signal_13439 ), .Q ( new_AGEMA_signal_13440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1942 ( .C ( clk ), .D ( new_AGEMA_signal_13441 ), .Q ( new_AGEMA_signal_13442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1944 ( .C ( clk ), .D ( new_AGEMA_signal_13443 ), .Q ( new_AGEMA_signal_13444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1946 ( .C ( clk ), .D ( new_AGEMA_signal_13445 ), .Q ( new_AGEMA_signal_13446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1948 ( .C ( clk ), .D ( new_AGEMA_signal_13447 ), .Q ( new_AGEMA_signal_13448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1950 ( .C ( clk ), .D ( new_AGEMA_signal_13449 ), .Q ( new_AGEMA_signal_13450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1952 ( .C ( clk ), .D ( new_AGEMA_signal_13451 ), .Q ( new_AGEMA_signal_13452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1954 ( .C ( clk ), .D ( new_AGEMA_signal_13453 ), .Q ( new_AGEMA_signal_13454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1956 ( .C ( clk ), .D ( new_AGEMA_signal_13455 ), .Q ( new_AGEMA_signal_13456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1958 ( .C ( clk ), .D ( new_AGEMA_signal_13457 ), .Q ( new_AGEMA_signal_13458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1960 ( .C ( clk ), .D ( new_AGEMA_signal_13459 ), .Q ( new_AGEMA_signal_13460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1962 ( .C ( clk ), .D ( new_AGEMA_signal_13461 ), .Q ( new_AGEMA_signal_13462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1964 ( .C ( clk ), .D ( new_AGEMA_signal_13463 ), .Q ( new_AGEMA_signal_13464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1966 ( .C ( clk ), .D ( new_AGEMA_signal_13465 ), .Q ( new_AGEMA_signal_13466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1968 ( .C ( clk ), .D ( new_AGEMA_signal_13467 ), .Q ( new_AGEMA_signal_13468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1970 ( .C ( clk ), .D ( new_AGEMA_signal_13469 ), .Q ( new_AGEMA_signal_13470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1972 ( .C ( clk ), .D ( new_AGEMA_signal_13471 ), .Q ( new_AGEMA_signal_13472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1974 ( .C ( clk ), .D ( new_AGEMA_signal_13473 ), .Q ( new_AGEMA_signal_13474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1976 ( .C ( clk ), .D ( new_AGEMA_signal_13475 ), .Q ( new_AGEMA_signal_13476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1978 ( .C ( clk ), .D ( new_AGEMA_signal_13477 ), .Q ( new_AGEMA_signal_13478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1980 ( .C ( clk ), .D ( new_AGEMA_signal_13479 ), .Q ( new_AGEMA_signal_13480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1982 ( .C ( clk ), .D ( new_AGEMA_signal_13481 ), .Q ( new_AGEMA_signal_13482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1984 ( .C ( clk ), .D ( new_AGEMA_signal_13483 ), .Q ( new_AGEMA_signal_13484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1986 ( .C ( clk ), .D ( new_AGEMA_signal_13485 ), .Q ( new_AGEMA_signal_13486 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1988 ( .C ( clk ), .D ( new_AGEMA_signal_13487 ), .Q ( new_AGEMA_signal_13488 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1990 ( .C ( clk ), .D ( new_AGEMA_signal_13489 ), .Q ( new_AGEMA_signal_13490 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1992 ( .C ( clk ), .D ( new_AGEMA_signal_13491 ), .Q ( new_AGEMA_signal_13492 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1994 ( .C ( clk ), .D ( new_AGEMA_signal_13493 ), .Q ( new_AGEMA_signal_13494 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1996 ( .C ( clk ), .D ( new_AGEMA_signal_13495 ), .Q ( new_AGEMA_signal_13496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1998 ( .C ( clk ), .D ( new_AGEMA_signal_13497 ), .Q ( new_AGEMA_signal_13498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2000 ( .C ( clk ), .D ( new_AGEMA_signal_13499 ), .Q ( new_AGEMA_signal_13500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2002 ( .C ( clk ), .D ( new_AGEMA_signal_13501 ), .Q ( new_AGEMA_signal_13502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2004 ( .C ( clk ), .D ( new_AGEMA_signal_13503 ), .Q ( new_AGEMA_signal_13504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2006 ( .C ( clk ), .D ( new_AGEMA_signal_13505 ), .Q ( new_AGEMA_signal_13506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2008 ( .C ( clk ), .D ( new_AGEMA_signal_13507 ), .Q ( new_AGEMA_signal_13508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2010 ( .C ( clk ), .D ( new_AGEMA_signal_13509 ), .Q ( new_AGEMA_signal_13510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2012 ( .C ( clk ), .D ( new_AGEMA_signal_13511 ), .Q ( new_AGEMA_signal_13512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2014 ( .C ( clk ), .D ( new_AGEMA_signal_13513 ), .Q ( new_AGEMA_signal_13514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2016 ( .C ( clk ), .D ( new_AGEMA_signal_13515 ), .Q ( new_AGEMA_signal_13516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2018 ( .C ( clk ), .D ( new_AGEMA_signal_13517 ), .Q ( new_AGEMA_signal_13518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2020 ( .C ( clk ), .D ( new_AGEMA_signal_13519 ), .Q ( new_AGEMA_signal_13520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2022 ( .C ( clk ), .D ( new_AGEMA_signal_13521 ), .Q ( new_AGEMA_signal_13522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2024 ( .C ( clk ), .D ( new_AGEMA_signal_13523 ), .Q ( new_AGEMA_signal_13524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2026 ( .C ( clk ), .D ( new_AGEMA_signal_13525 ), .Q ( new_AGEMA_signal_13526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2028 ( .C ( clk ), .D ( new_AGEMA_signal_13527 ), .Q ( new_AGEMA_signal_13528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2030 ( .C ( clk ), .D ( new_AGEMA_signal_13529 ), .Q ( new_AGEMA_signal_13530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2032 ( .C ( clk ), .D ( new_AGEMA_signal_13531 ), .Q ( new_AGEMA_signal_13532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2034 ( .C ( clk ), .D ( new_AGEMA_signal_13533 ), .Q ( new_AGEMA_signal_13534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2036 ( .C ( clk ), .D ( new_AGEMA_signal_13535 ), .Q ( new_AGEMA_signal_13536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2038 ( .C ( clk ), .D ( new_AGEMA_signal_13537 ), .Q ( new_AGEMA_signal_13538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2040 ( .C ( clk ), .D ( new_AGEMA_signal_13539 ), .Q ( new_AGEMA_signal_13540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2042 ( .C ( clk ), .D ( new_AGEMA_signal_13541 ), .Q ( new_AGEMA_signal_13542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2044 ( .C ( clk ), .D ( new_AGEMA_signal_13543 ), .Q ( new_AGEMA_signal_13544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2046 ( .C ( clk ), .D ( new_AGEMA_signal_13545 ), .Q ( new_AGEMA_signal_13546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2048 ( .C ( clk ), .D ( new_AGEMA_signal_13547 ), .Q ( new_AGEMA_signal_13548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2050 ( .C ( clk ), .D ( new_AGEMA_signal_13549 ), .Q ( new_AGEMA_signal_13550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2052 ( .C ( clk ), .D ( new_AGEMA_signal_13551 ), .Q ( new_AGEMA_signal_13552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2054 ( .C ( clk ), .D ( new_AGEMA_signal_13553 ), .Q ( new_AGEMA_signal_13554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2056 ( .C ( clk ), .D ( new_AGEMA_signal_13555 ), .Q ( new_AGEMA_signal_13556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2058 ( .C ( clk ), .D ( new_AGEMA_signal_13557 ), .Q ( new_AGEMA_signal_13558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2060 ( .C ( clk ), .D ( new_AGEMA_signal_13559 ), .Q ( new_AGEMA_signal_13560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2062 ( .C ( clk ), .D ( new_AGEMA_signal_13561 ), .Q ( new_AGEMA_signal_13562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2064 ( .C ( clk ), .D ( new_AGEMA_signal_13563 ), .Q ( new_AGEMA_signal_13564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2066 ( .C ( clk ), .D ( new_AGEMA_signal_13565 ), .Q ( new_AGEMA_signal_13566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2068 ( .C ( clk ), .D ( new_AGEMA_signal_13567 ), .Q ( new_AGEMA_signal_13568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2070 ( .C ( clk ), .D ( new_AGEMA_signal_13569 ), .Q ( new_AGEMA_signal_13570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2076 ( .C ( clk ), .D ( new_AGEMA_signal_13575 ), .Q ( new_AGEMA_signal_13576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2082 ( .C ( clk ), .D ( new_AGEMA_signal_13581 ), .Q ( new_AGEMA_signal_13582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2088 ( .C ( clk ), .D ( new_AGEMA_signal_13587 ), .Q ( new_AGEMA_signal_13588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2094 ( .C ( clk ), .D ( new_AGEMA_signal_13593 ), .Q ( new_AGEMA_signal_13594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2096 ( .C ( clk ), .D ( new_AGEMA_signal_13595 ), .Q ( new_AGEMA_signal_13596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2098 ( .C ( clk ), .D ( new_AGEMA_signal_13597 ), .Q ( new_AGEMA_signal_13598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2100 ( .C ( clk ), .D ( new_AGEMA_signal_13599 ), .Q ( new_AGEMA_signal_13600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2102 ( .C ( clk ), .D ( new_AGEMA_signal_13601 ), .Q ( new_AGEMA_signal_13602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2104 ( .C ( clk ), .D ( new_AGEMA_signal_13603 ), .Q ( new_AGEMA_signal_13604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2106 ( .C ( clk ), .D ( new_AGEMA_signal_13605 ), .Q ( new_AGEMA_signal_13606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2108 ( .C ( clk ), .D ( new_AGEMA_signal_13607 ), .Q ( new_AGEMA_signal_13608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2110 ( .C ( clk ), .D ( new_AGEMA_signal_13609 ), .Q ( new_AGEMA_signal_13610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2112 ( .C ( clk ), .D ( new_AGEMA_signal_13611 ), .Q ( new_AGEMA_signal_13612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2114 ( .C ( clk ), .D ( new_AGEMA_signal_13613 ), .Q ( new_AGEMA_signal_13614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2116 ( .C ( clk ), .D ( new_AGEMA_signal_13615 ), .Q ( new_AGEMA_signal_13616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2118 ( .C ( clk ), .D ( new_AGEMA_signal_13617 ), .Q ( new_AGEMA_signal_13618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2122 ( .C ( clk ), .D ( new_AGEMA_signal_13621 ), .Q ( new_AGEMA_signal_13622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2126 ( .C ( clk ), .D ( new_AGEMA_signal_13625 ), .Q ( new_AGEMA_signal_13626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2130 ( .C ( clk ), .D ( new_AGEMA_signal_13629 ), .Q ( new_AGEMA_signal_13630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2134 ( .C ( clk ), .D ( new_AGEMA_signal_13633 ), .Q ( new_AGEMA_signal_13634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2136 ( .C ( clk ), .D ( new_AGEMA_signal_13635 ), .Q ( new_AGEMA_signal_13636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2138 ( .C ( clk ), .D ( new_AGEMA_signal_13637 ), .Q ( new_AGEMA_signal_13638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2140 ( .C ( clk ), .D ( new_AGEMA_signal_13639 ), .Q ( new_AGEMA_signal_13640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2142 ( .C ( clk ), .D ( new_AGEMA_signal_13641 ), .Q ( new_AGEMA_signal_13642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2144 ( .C ( clk ), .D ( new_AGEMA_signal_13643 ), .Q ( new_AGEMA_signal_13644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2146 ( .C ( clk ), .D ( new_AGEMA_signal_13645 ), .Q ( new_AGEMA_signal_13646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2148 ( .C ( clk ), .D ( new_AGEMA_signal_13647 ), .Q ( new_AGEMA_signal_13648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2150 ( .C ( clk ), .D ( new_AGEMA_signal_13649 ), .Q ( new_AGEMA_signal_13650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2152 ( .C ( clk ), .D ( new_AGEMA_signal_13651 ), .Q ( new_AGEMA_signal_13652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2154 ( .C ( clk ), .D ( new_AGEMA_signal_13653 ), .Q ( new_AGEMA_signal_13654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2156 ( .C ( clk ), .D ( new_AGEMA_signal_13655 ), .Q ( new_AGEMA_signal_13656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2158 ( .C ( clk ), .D ( new_AGEMA_signal_13657 ), .Q ( new_AGEMA_signal_13658 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2162 ( .C ( clk ), .D ( new_AGEMA_signal_13661 ), .Q ( new_AGEMA_signal_13662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2166 ( .C ( clk ), .D ( new_AGEMA_signal_13665 ), .Q ( new_AGEMA_signal_13666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2170 ( .C ( clk ), .D ( new_AGEMA_signal_13669 ), .Q ( new_AGEMA_signal_13670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2174 ( .C ( clk ), .D ( new_AGEMA_signal_13673 ), .Q ( new_AGEMA_signal_13674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2176 ( .C ( clk ), .D ( new_AGEMA_signal_13675 ), .Q ( new_AGEMA_signal_13676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2178 ( .C ( clk ), .D ( new_AGEMA_signal_13677 ), .Q ( new_AGEMA_signal_13678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2180 ( .C ( clk ), .D ( new_AGEMA_signal_13679 ), .Q ( new_AGEMA_signal_13680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2182 ( .C ( clk ), .D ( new_AGEMA_signal_13681 ), .Q ( new_AGEMA_signal_13682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2184 ( .C ( clk ), .D ( new_AGEMA_signal_13683 ), .Q ( new_AGEMA_signal_13684 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2186 ( .C ( clk ), .D ( new_AGEMA_signal_13685 ), .Q ( new_AGEMA_signal_13686 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2188 ( .C ( clk ), .D ( new_AGEMA_signal_13687 ), .Q ( new_AGEMA_signal_13688 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2190 ( .C ( clk ), .D ( new_AGEMA_signal_13689 ), .Q ( new_AGEMA_signal_13690 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2192 ( .C ( clk ), .D ( new_AGEMA_signal_13691 ), .Q ( new_AGEMA_signal_13692 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2194 ( .C ( clk ), .D ( new_AGEMA_signal_13693 ), .Q ( new_AGEMA_signal_13694 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2196 ( .C ( clk ), .D ( new_AGEMA_signal_13695 ), .Q ( new_AGEMA_signal_13696 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2198 ( .C ( clk ), .D ( new_AGEMA_signal_13697 ), .Q ( new_AGEMA_signal_13698 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2200 ( .C ( clk ), .D ( new_AGEMA_signal_13699 ), .Q ( new_AGEMA_signal_13700 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2202 ( .C ( clk ), .D ( new_AGEMA_signal_13701 ), .Q ( new_AGEMA_signal_13702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2204 ( .C ( clk ), .D ( new_AGEMA_signal_13703 ), .Q ( new_AGEMA_signal_13704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2206 ( .C ( clk ), .D ( new_AGEMA_signal_13705 ), .Q ( new_AGEMA_signal_13706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2208 ( .C ( clk ), .D ( new_AGEMA_signal_13707 ), .Q ( new_AGEMA_signal_13708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2210 ( .C ( clk ), .D ( new_AGEMA_signal_13709 ), .Q ( new_AGEMA_signal_13710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2212 ( .C ( clk ), .D ( new_AGEMA_signal_13711 ), .Q ( new_AGEMA_signal_13712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2214 ( .C ( clk ), .D ( new_AGEMA_signal_13713 ), .Q ( new_AGEMA_signal_13714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2216 ( .C ( clk ), .D ( new_AGEMA_signal_13715 ), .Q ( new_AGEMA_signal_13716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2218 ( .C ( clk ), .D ( new_AGEMA_signal_13717 ), .Q ( new_AGEMA_signal_13718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2220 ( .C ( clk ), .D ( new_AGEMA_signal_13719 ), .Q ( new_AGEMA_signal_13720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2222 ( .C ( clk ), .D ( new_AGEMA_signal_13721 ), .Q ( new_AGEMA_signal_13722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2224 ( .C ( clk ), .D ( new_AGEMA_signal_13723 ), .Q ( new_AGEMA_signal_13724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2226 ( .C ( clk ), .D ( new_AGEMA_signal_13725 ), .Q ( new_AGEMA_signal_13726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2228 ( .C ( clk ), .D ( new_AGEMA_signal_13727 ), .Q ( new_AGEMA_signal_13728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2230 ( .C ( clk ), .D ( new_AGEMA_signal_13729 ), .Q ( new_AGEMA_signal_13730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2234 ( .C ( clk ), .D ( new_AGEMA_signal_13733 ), .Q ( new_AGEMA_signal_13734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2238 ( .C ( clk ), .D ( new_AGEMA_signal_13737 ), .Q ( new_AGEMA_signal_13738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2242 ( .C ( clk ), .D ( new_AGEMA_signal_13741 ), .Q ( new_AGEMA_signal_13742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2246 ( .C ( clk ), .D ( new_AGEMA_signal_13745 ), .Q ( new_AGEMA_signal_13746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2248 ( .C ( clk ), .D ( new_AGEMA_signal_13747 ), .Q ( new_AGEMA_signal_13748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2250 ( .C ( clk ), .D ( new_AGEMA_signal_13749 ), .Q ( new_AGEMA_signal_13750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2252 ( .C ( clk ), .D ( new_AGEMA_signal_13751 ), .Q ( new_AGEMA_signal_13752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2254 ( .C ( clk ), .D ( new_AGEMA_signal_13753 ), .Q ( new_AGEMA_signal_13754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2256 ( .C ( clk ), .D ( new_AGEMA_signal_13755 ), .Q ( new_AGEMA_signal_13756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2258 ( .C ( clk ), .D ( new_AGEMA_signal_13757 ), .Q ( new_AGEMA_signal_13758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2260 ( .C ( clk ), .D ( new_AGEMA_signal_13759 ), .Q ( new_AGEMA_signal_13760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2262 ( .C ( clk ), .D ( new_AGEMA_signal_13761 ), .Q ( new_AGEMA_signal_13762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2266 ( .C ( clk ), .D ( new_AGEMA_signal_13765 ), .Q ( new_AGEMA_signal_13766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2270 ( .C ( clk ), .D ( new_AGEMA_signal_13769 ), .Q ( new_AGEMA_signal_13770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2274 ( .C ( clk ), .D ( new_AGEMA_signal_13773 ), .Q ( new_AGEMA_signal_13774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2278 ( .C ( clk ), .D ( new_AGEMA_signal_13777 ), .Q ( new_AGEMA_signal_13778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2280 ( .C ( clk ), .D ( new_AGEMA_signal_13779 ), .Q ( new_AGEMA_signal_13780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2282 ( .C ( clk ), .D ( new_AGEMA_signal_13781 ), .Q ( new_AGEMA_signal_13782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2284 ( .C ( clk ), .D ( new_AGEMA_signal_13783 ), .Q ( new_AGEMA_signal_13784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2286 ( .C ( clk ), .D ( new_AGEMA_signal_13785 ), .Q ( new_AGEMA_signal_13786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2288 ( .C ( clk ), .D ( new_AGEMA_signal_13787 ), .Q ( new_AGEMA_signal_13788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2292 ( .C ( clk ), .D ( new_AGEMA_signal_13791 ), .Q ( new_AGEMA_signal_13792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2296 ( .C ( clk ), .D ( new_AGEMA_signal_13795 ), .Q ( new_AGEMA_signal_13796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2300 ( .C ( clk ), .D ( new_AGEMA_signal_13799 ), .Q ( new_AGEMA_signal_13800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2304 ( .C ( clk ), .D ( new_AGEMA_signal_13803 ), .Q ( new_AGEMA_signal_13804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2308 ( .C ( clk ), .D ( new_AGEMA_signal_13807 ), .Q ( new_AGEMA_signal_13808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2312 ( .C ( clk ), .D ( new_AGEMA_signal_13811 ), .Q ( new_AGEMA_signal_13812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2316 ( .C ( clk ), .D ( new_AGEMA_signal_13815 ), .Q ( new_AGEMA_signal_13816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2336 ( .C ( clk ), .D ( new_AGEMA_signal_13835 ), .Q ( new_AGEMA_signal_13836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2340 ( .C ( clk ), .D ( new_AGEMA_signal_13839 ), .Q ( new_AGEMA_signal_13840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2344 ( .C ( clk ), .D ( new_AGEMA_signal_13843 ), .Q ( new_AGEMA_signal_13844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2348 ( .C ( clk ), .D ( new_AGEMA_signal_13847 ), .Q ( new_AGEMA_signal_13848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2360 ( .C ( clk ), .D ( new_AGEMA_signal_13859 ), .Q ( new_AGEMA_signal_13860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2364 ( .C ( clk ), .D ( new_AGEMA_signal_13863 ), .Q ( new_AGEMA_signal_13864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2368 ( .C ( clk ), .D ( new_AGEMA_signal_13867 ), .Q ( new_AGEMA_signal_13868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2372 ( .C ( clk ), .D ( new_AGEMA_signal_13871 ), .Q ( new_AGEMA_signal_13872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2384 ( .C ( clk ), .D ( new_AGEMA_signal_13883 ), .Q ( new_AGEMA_signal_13884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2388 ( .C ( clk ), .D ( new_AGEMA_signal_13887 ), .Q ( new_AGEMA_signal_13888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2392 ( .C ( clk ), .D ( new_AGEMA_signal_13891 ), .Q ( new_AGEMA_signal_13892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2396 ( .C ( clk ), .D ( new_AGEMA_signal_13895 ), .Q ( new_AGEMA_signal_13896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2400 ( .C ( clk ), .D ( new_AGEMA_signal_13899 ), .Q ( new_AGEMA_signal_13900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2404 ( .C ( clk ), .D ( new_AGEMA_signal_13903 ), .Q ( new_AGEMA_signal_13904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2408 ( .C ( clk ), .D ( new_AGEMA_signal_13907 ), .Q ( new_AGEMA_signal_13908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2412 ( .C ( clk ), .D ( new_AGEMA_signal_13911 ), .Q ( new_AGEMA_signal_13912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2448 ( .C ( clk ), .D ( new_AGEMA_signal_13947 ), .Q ( new_AGEMA_signal_13948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2452 ( .C ( clk ), .D ( new_AGEMA_signal_13951 ), .Q ( new_AGEMA_signal_13952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2456 ( .C ( clk ), .D ( new_AGEMA_signal_13955 ), .Q ( new_AGEMA_signal_13956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2460 ( .C ( clk ), .D ( new_AGEMA_signal_13959 ), .Q ( new_AGEMA_signal_13960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2464 ( .C ( clk ), .D ( new_AGEMA_signal_13963 ), .Q ( new_AGEMA_signal_13964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2468 ( .C ( clk ), .D ( new_AGEMA_signal_13967 ), .Q ( new_AGEMA_signal_13968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2472 ( .C ( clk ), .D ( new_AGEMA_signal_13971 ), .Q ( new_AGEMA_signal_13972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2476 ( .C ( clk ), .D ( new_AGEMA_signal_13975 ), .Q ( new_AGEMA_signal_13976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2480 ( .C ( clk ), .D ( new_AGEMA_signal_13979 ), .Q ( new_AGEMA_signal_13980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2484 ( .C ( clk ), .D ( new_AGEMA_signal_13983 ), .Q ( new_AGEMA_signal_13984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2488 ( .C ( clk ), .D ( new_AGEMA_signal_13987 ), .Q ( new_AGEMA_signal_13988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2492 ( .C ( clk ), .D ( new_AGEMA_signal_13991 ), .Q ( new_AGEMA_signal_13992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2520 ( .C ( clk ), .D ( new_AGEMA_signal_14019 ), .Q ( new_AGEMA_signal_14020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2524 ( .C ( clk ), .D ( new_AGEMA_signal_14023 ), .Q ( new_AGEMA_signal_14024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2528 ( .C ( clk ), .D ( new_AGEMA_signal_14027 ), .Q ( new_AGEMA_signal_14028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2532 ( .C ( clk ), .D ( new_AGEMA_signal_14031 ), .Q ( new_AGEMA_signal_14032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2544 ( .C ( clk ), .D ( new_AGEMA_signal_14043 ), .Q ( new_AGEMA_signal_14044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2548 ( .C ( clk ), .D ( new_AGEMA_signal_14047 ), .Q ( new_AGEMA_signal_14048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2552 ( .C ( clk ), .D ( new_AGEMA_signal_14051 ), .Q ( new_AGEMA_signal_14052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2556 ( .C ( clk ), .D ( new_AGEMA_signal_14055 ), .Q ( new_AGEMA_signal_14056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2562 ( .C ( clk ), .D ( new_AGEMA_signal_14061 ), .Q ( new_AGEMA_signal_14062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2568 ( .C ( clk ), .D ( new_AGEMA_signal_14067 ), .Q ( new_AGEMA_signal_14068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2574 ( .C ( clk ), .D ( new_AGEMA_signal_14073 ), .Q ( new_AGEMA_signal_14074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2580 ( .C ( clk ), .D ( new_AGEMA_signal_14079 ), .Q ( new_AGEMA_signal_14080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2584 ( .C ( clk ), .D ( new_AGEMA_signal_14083 ), .Q ( new_AGEMA_signal_14084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2588 ( .C ( clk ), .D ( new_AGEMA_signal_14087 ), .Q ( new_AGEMA_signal_14088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2592 ( .C ( clk ), .D ( new_AGEMA_signal_14091 ), .Q ( new_AGEMA_signal_14092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2596 ( .C ( clk ), .D ( new_AGEMA_signal_14095 ), .Q ( new_AGEMA_signal_14096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2600 ( .C ( clk ), .D ( new_AGEMA_signal_14099 ), .Q ( new_AGEMA_signal_14100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2604 ( .C ( clk ), .D ( new_AGEMA_signal_14103 ), .Q ( new_AGEMA_signal_14104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2608 ( .C ( clk ), .D ( new_AGEMA_signal_14107 ), .Q ( new_AGEMA_signal_14108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2612 ( .C ( clk ), .D ( new_AGEMA_signal_14111 ), .Q ( new_AGEMA_signal_14112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2648 ( .C ( clk ), .D ( new_AGEMA_signal_14147 ), .Q ( new_AGEMA_signal_14148 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2652 ( .C ( clk ), .D ( new_AGEMA_signal_14151 ), .Q ( new_AGEMA_signal_14152 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2656 ( .C ( clk ), .D ( new_AGEMA_signal_14155 ), .Q ( new_AGEMA_signal_14156 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2660 ( .C ( clk ), .D ( new_AGEMA_signal_14159 ), .Q ( new_AGEMA_signal_14160 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2666 ( .C ( clk ), .D ( new_AGEMA_signal_14165 ), .Q ( new_AGEMA_signal_14166 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2672 ( .C ( clk ), .D ( new_AGEMA_signal_14171 ), .Q ( new_AGEMA_signal_14172 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2678 ( .C ( clk ), .D ( new_AGEMA_signal_14177 ), .Q ( new_AGEMA_signal_14178 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2684 ( .C ( clk ), .D ( new_AGEMA_signal_14183 ), .Q ( new_AGEMA_signal_14184 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2688 ( .C ( clk ), .D ( new_AGEMA_signal_14187 ), .Q ( new_AGEMA_signal_14188 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2692 ( .C ( clk ), .D ( new_AGEMA_signal_14191 ), .Q ( new_AGEMA_signal_14192 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2696 ( .C ( clk ), .D ( new_AGEMA_signal_14195 ), .Q ( new_AGEMA_signal_14196 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2700 ( .C ( clk ), .D ( new_AGEMA_signal_14199 ), .Q ( new_AGEMA_signal_14200 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2728 ( .C ( clk ), .D ( new_AGEMA_signal_14227 ), .Q ( new_AGEMA_signal_14228 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2732 ( .C ( clk ), .D ( new_AGEMA_signal_14231 ), .Q ( new_AGEMA_signal_14232 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2736 ( .C ( clk ), .D ( new_AGEMA_signal_14235 ), .Q ( new_AGEMA_signal_14236 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2740 ( .C ( clk ), .D ( new_AGEMA_signal_14239 ), .Q ( new_AGEMA_signal_14240 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2760 ( .C ( clk ), .D ( new_AGEMA_signal_14259 ), .Q ( new_AGEMA_signal_14260 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2764 ( .C ( clk ), .D ( new_AGEMA_signal_14263 ), .Q ( new_AGEMA_signal_14264 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2768 ( .C ( clk ), .D ( new_AGEMA_signal_14267 ), .Q ( new_AGEMA_signal_14268 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2772 ( .C ( clk ), .D ( new_AGEMA_signal_14271 ), .Q ( new_AGEMA_signal_14272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2776 ( .C ( clk ), .D ( new_AGEMA_signal_14275 ), .Q ( new_AGEMA_signal_14276 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2780 ( .C ( clk ), .D ( new_AGEMA_signal_14279 ), .Q ( new_AGEMA_signal_14280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2784 ( .C ( clk ), .D ( new_AGEMA_signal_14283 ), .Q ( new_AGEMA_signal_14284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2788 ( .C ( clk ), .D ( new_AGEMA_signal_14287 ), .Q ( new_AGEMA_signal_14288 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2792 ( .C ( clk ), .D ( new_AGEMA_signal_14291 ), .Q ( new_AGEMA_signal_14292 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2796 ( .C ( clk ), .D ( new_AGEMA_signal_14295 ), .Q ( new_AGEMA_signal_14296 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2800 ( .C ( clk ), .D ( new_AGEMA_signal_14299 ), .Q ( new_AGEMA_signal_14300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2804 ( .C ( clk ), .D ( new_AGEMA_signal_14303 ), .Q ( new_AGEMA_signal_14304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2808 ( .C ( clk ), .D ( new_AGEMA_signal_14307 ), .Q ( new_AGEMA_signal_14308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2812 ( .C ( clk ), .D ( new_AGEMA_signal_14311 ), .Q ( new_AGEMA_signal_14312 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2816 ( .C ( clk ), .D ( new_AGEMA_signal_14315 ), .Q ( new_AGEMA_signal_14316 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2820 ( .C ( clk ), .D ( new_AGEMA_signal_14319 ), .Q ( new_AGEMA_signal_14320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2824 ( .C ( clk ), .D ( new_AGEMA_signal_14323 ), .Q ( new_AGEMA_signal_14324 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2828 ( .C ( clk ), .D ( new_AGEMA_signal_14327 ), .Q ( new_AGEMA_signal_14328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2832 ( .C ( clk ), .D ( new_AGEMA_signal_14331 ), .Q ( new_AGEMA_signal_14332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2836 ( .C ( clk ), .D ( new_AGEMA_signal_14335 ), .Q ( new_AGEMA_signal_14336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2872 ( .C ( clk ), .D ( new_AGEMA_signal_14371 ), .Q ( new_AGEMA_signal_14372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2876 ( .C ( clk ), .D ( new_AGEMA_signal_14375 ), .Q ( new_AGEMA_signal_14376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2880 ( .C ( clk ), .D ( new_AGEMA_signal_14379 ), .Q ( new_AGEMA_signal_14380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2884 ( .C ( clk ), .D ( new_AGEMA_signal_14383 ), .Q ( new_AGEMA_signal_14384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2888 ( .C ( clk ), .D ( new_AGEMA_signal_14387 ), .Q ( new_AGEMA_signal_14388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2892 ( .C ( clk ), .D ( new_AGEMA_signal_14391 ), .Q ( new_AGEMA_signal_14392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2896 ( .C ( clk ), .D ( new_AGEMA_signal_14395 ), .Q ( new_AGEMA_signal_14396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2900 ( .C ( clk ), .D ( new_AGEMA_signal_14399 ), .Q ( new_AGEMA_signal_14400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2976 ( .C ( clk ), .D ( new_AGEMA_signal_14475 ), .Q ( new_AGEMA_signal_14476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2980 ( .C ( clk ), .D ( new_AGEMA_signal_14479 ), .Q ( new_AGEMA_signal_14480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2984 ( .C ( clk ), .D ( new_AGEMA_signal_14483 ), .Q ( new_AGEMA_signal_14484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2988 ( .C ( clk ), .D ( new_AGEMA_signal_14487 ), .Q ( new_AGEMA_signal_14488 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3032 ( .C ( clk ), .D ( new_AGEMA_signal_14531 ), .Q ( new_AGEMA_signal_14532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3036 ( .C ( clk ), .D ( new_AGEMA_signal_14535 ), .Q ( new_AGEMA_signal_14536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3040 ( .C ( clk ), .D ( new_AGEMA_signal_14539 ), .Q ( new_AGEMA_signal_14540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3044 ( .C ( clk ), .D ( new_AGEMA_signal_14543 ), .Q ( new_AGEMA_signal_14544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3048 ( .C ( clk ), .D ( new_AGEMA_signal_14547 ), .Q ( new_AGEMA_signal_14548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3052 ( .C ( clk ), .D ( new_AGEMA_signal_14551 ), .Q ( new_AGEMA_signal_14552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3056 ( .C ( clk ), .D ( new_AGEMA_signal_14555 ), .Q ( new_AGEMA_signal_14556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3060 ( .C ( clk ), .D ( new_AGEMA_signal_14559 ), .Q ( new_AGEMA_signal_14560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3064 ( .C ( clk ), .D ( new_AGEMA_signal_14563 ), .Q ( new_AGEMA_signal_14564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3068 ( .C ( clk ), .D ( new_AGEMA_signal_14567 ), .Q ( new_AGEMA_signal_14568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3072 ( .C ( clk ), .D ( new_AGEMA_signal_14571 ), .Q ( new_AGEMA_signal_14572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3076 ( .C ( clk ), .D ( new_AGEMA_signal_14575 ), .Q ( new_AGEMA_signal_14576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3080 ( .C ( clk ), .D ( new_AGEMA_signal_14579 ), .Q ( new_AGEMA_signal_14580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3084 ( .C ( clk ), .D ( new_AGEMA_signal_14583 ), .Q ( new_AGEMA_signal_14584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3088 ( .C ( clk ), .D ( new_AGEMA_signal_14587 ), .Q ( new_AGEMA_signal_14588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3092 ( .C ( clk ), .D ( new_AGEMA_signal_14591 ), .Q ( new_AGEMA_signal_14592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3130 ( .C ( clk ), .D ( new_AGEMA_signal_14629 ), .Q ( new_AGEMA_signal_14630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3138 ( .C ( clk ), .D ( new_AGEMA_signal_14637 ), .Q ( new_AGEMA_signal_14638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3146 ( .C ( clk ), .D ( new_AGEMA_signal_14645 ), .Q ( new_AGEMA_signal_14646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3154 ( .C ( clk ), .D ( new_AGEMA_signal_14653 ), .Q ( new_AGEMA_signal_14654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3170 ( .C ( clk ), .D ( new_AGEMA_signal_14669 ), .Q ( new_AGEMA_signal_14670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3178 ( .C ( clk ), .D ( new_AGEMA_signal_14677 ), .Q ( new_AGEMA_signal_14678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3186 ( .C ( clk ), .D ( new_AGEMA_signal_14685 ), .Q ( new_AGEMA_signal_14686 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3194 ( .C ( clk ), .D ( new_AGEMA_signal_14693 ), .Q ( new_AGEMA_signal_14694 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3200 ( .C ( clk ), .D ( new_AGEMA_signal_14699 ), .Q ( new_AGEMA_signal_14700 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3206 ( .C ( clk ), .D ( new_AGEMA_signal_14705 ), .Q ( new_AGEMA_signal_14706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3212 ( .C ( clk ), .D ( new_AGEMA_signal_14711 ), .Q ( new_AGEMA_signal_14712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3218 ( .C ( clk ), .D ( new_AGEMA_signal_14717 ), .Q ( new_AGEMA_signal_14718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3240 ( .C ( clk ), .D ( new_AGEMA_signal_14739 ), .Q ( new_AGEMA_signal_14740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3246 ( .C ( clk ), .D ( new_AGEMA_signal_14745 ), .Q ( new_AGEMA_signal_14746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3252 ( .C ( clk ), .D ( new_AGEMA_signal_14751 ), .Q ( new_AGEMA_signal_14752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3258 ( .C ( clk ), .D ( new_AGEMA_signal_14757 ), .Q ( new_AGEMA_signal_14758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3272 ( .C ( clk ), .D ( new_AGEMA_signal_14771 ), .Q ( new_AGEMA_signal_14772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3278 ( .C ( clk ), .D ( new_AGEMA_signal_14777 ), .Q ( new_AGEMA_signal_14778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3284 ( .C ( clk ), .D ( new_AGEMA_signal_14783 ), .Q ( new_AGEMA_signal_14784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3290 ( .C ( clk ), .D ( new_AGEMA_signal_14789 ), .Q ( new_AGEMA_signal_14790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3296 ( .C ( clk ), .D ( new_AGEMA_signal_14795 ), .Q ( new_AGEMA_signal_14796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3302 ( .C ( clk ), .D ( new_AGEMA_signal_14801 ), .Q ( new_AGEMA_signal_14802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3308 ( .C ( clk ), .D ( new_AGEMA_signal_14807 ), .Q ( new_AGEMA_signal_14808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3314 ( .C ( clk ), .D ( new_AGEMA_signal_14813 ), .Q ( new_AGEMA_signal_14814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3344 ( .C ( clk ), .D ( new_AGEMA_signal_14843 ), .Q ( new_AGEMA_signal_14844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3350 ( .C ( clk ), .D ( new_AGEMA_signal_14849 ), .Q ( new_AGEMA_signal_14850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3356 ( .C ( clk ), .D ( new_AGEMA_signal_14855 ), .Q ( new_AGEMA_signal_14856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3362 ( .C ( clk ), .D ( new_AGEMA_signal_14861 ), .Q ( new_AGEMA_signal_14862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3368 ( .C ( clk ), .D ( new_AGEMA_signal_14867 ), .Q ( new_AGEMA_signal_14868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3374 ( .C ( clk ), .D ( new_AGEMA_signal_14873 ), .Q ( new_AGEMA_signal_14874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3380 ( .C ( clk ), .D ( new_AGEMA_signal_14879 ), .Q ( new_AGEMA_signal_14880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3386 ( .C ( clk ), .D ( new_AGEMA_signal_14885 ), .Q ( new_AGEMA_signal_14886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3400 ( .C ( clk ), .D ( new_AGEMA_signal_14899 ), .Q ( new_AGEMA_signal_14900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3406 ( .C ( clk ), .D ( new_AGEMA_signal_14905 ), .Q ( new_AGEMA_signal_14906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3412 ( .C ( clk ), .D ( new_AGEMA_signal_14911 ), .Q ( new_AGEMA_signal_14912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3418 ( .C ( clk ), .D ( new_AGEMA_signal_14917 ), .Q ( new_AGEMA_signal_14918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3474 ( .C ( clk ), .D ( new_AGEMA_signal_14973 ), .Q ( new_AGEMA_signal_14974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3482 ( .C ( clk ), .D ( new_AGEMA_signal_14981 ), .Q ( new_AGEMA_signal_14982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3490 ( .C ( clk ), .D ( new_AGEMA_signal_14989 ), .Q ( new_AGEMA_signal_14990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3498 ( .C ( clk ), .D ( new_AGEMA_signal_14997 ), .Q ( new_AGEMA_signal_14998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3504 ( .C ( clk ), .D ( new_AGEMA_signal_15003 ), .Q ( new_AGEMA_signal_15004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3510 ( .C ( clk ), .D ( new_AGEMA_signal_15009 ), .Q ( new_AGEMA_signal_15010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3516 ( .C ( clk ), .D ( new_AGEMA_signal_15015 ), .Q ( new_AGEMA_signal_15016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3522 ( .C ( clk ), .D ( new_AGEMA_signal_15021 ), .Q ( new_AGEMA_signal_15022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3616 ( .C ( clk ), .D ( new_AGEMA_signal_15115 ), .Q ( new_AGEMA_signal_15116 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3622 ( .C ( clk ), .D ( new_AGEMA_signal_15121 ), .Q ( new_AGEMA_signal_15122 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3628 ( .C ( clk ), .D ( new_AGEMA_signal_15127 ), .Q ( new_AGEMA_signal_15128 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3634 ( .C ( clk ), .D ( new_AGEMA_signal_15133 ), .Q ( new_AGEMA_signal_15134 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3744 ( .C ( clk ), .D ( new_AGEMA_signal_15243 ), .Q ( new_AGEMA_signal_15244 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3750 ( .C ( clk ), .D ( new_AGEMA_signal_15249 ), .Q ( new_AGEMA_signal_15250 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3756 ( .C ( clk ), .D ( new_AGEMA_signal_15255 ), .Q ( new_AGEMA_signal_15256 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3762 ( .C ( clk ), .D ( new_AGEMA_signal_15261 ), .Q ( new_AGEMA_signal_15262 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3768 ( .C ( clk ), .D ( new_AGEMA_signal_15267 ), .Q ( new_AGEMA_signal_15268 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3774 ( .C ( clk ), .D ( new_AGEMA_signal_15273 ), .Q ( new_AGEMA_signal_15274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3780 ( .C ( clk ), .D ( new_AGEMA_signal_15279 ), .Q ( new_AGEMA_signal_15280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3786 ( .C ( clk ), .D ( new_AGEMA_signal_15285 ), .Q ( new_AGEMA_signal_15286 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3818 ( .C ( clk ), .D ( new_AGEMA_signal_15317 ), .Q ( new_AGEMA_signal_15318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3826 ( .C ( clk ), .D ( new_AGEMA_signal_15325 ), .Q ( new_AGEMA_signal_15326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3834 ( .C ( clk ), .D ( new_AGEMA_signal_15333 ), .Q ( new_AGEMA_signal_15334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3842 ( .C ( clk ), .D ( new_AGEMA_signal_15341 ), .Q ( new_AGEMA_signal_15342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3938 ( .C ( clk ), .D ( new_AGEMA_signal_15437 ), .Q ( new_AGEMA_signal_15438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3946 ( .C ( clk ), .D ( new_AGEMA_signal_15445 ), .Q ( new_AGEMA_signal_15446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3954 ( .C ( clk ), .D ( new_AGEMA_signal_15453 ), .Q ( new_AGEMA_signal_15454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3962 ( .C ( clk ), .D ( new_AGEMA_signal_15461 ), .Q ( new_AGEMA_signal_15462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4000 ( .C ( clk ), .D ( new_AGEMA_signal_15499 ), .Q ( new_AGEMA_signal_15500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4006 ( .C ( clk ), .D ( new_AGEMA_signal_15505 ), .Q ( new_AGEMA_signal_15506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4012 ( .C ( clk ), .D ( new_AGEMA_signal_15511 ), .Q ( new_AGEMA_signal_15512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4018 ( .C ( clk ), .D ( new_AGEMA_signal_15517 ), .Q ( new_AGEMA_signal_15518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4032 ( .C ( clk ), .D ( new_AGEMA_signal_15531 ), .Q ( new_AGEMA_signal_15532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4040 ( .C ( clk ), .D ( new_AGEMA_signal_15539 ), .Q ( new_AGEMA_signal_15540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4048 ( .C ( clk ), .D ( new_AGEMA_signal_15547 ), .Q ( new_AGEMA_signal_15548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4056 ( .C ( clk ), .D ( new_AGEMA_signal_15555 ), .Q ( new_AGEMA_signal_15556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4088 ( .C ( clk ), .D ( new_AGEMA_signal_15587 ), .Q ( new_AGEMA_signal_15588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4096 ( .C ( clk ), .D ( new_AGEMA_signal_15595 ), .Q ( new_AGEMA_signal_15596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4104 ( .C ( clk ), .D ( new_AGEMA_signal_15603 ), .Q ( new_AGEMA_signal_15604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4112 ( .C ( clk ), .D ( new_AGEMA_signal_15611 ), .Q ( new_AGEMA_signal_15612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4168 ( .C ( clk ), .D ( new_AGEMA_signal_15667 ), .Q ( new_AGEMA_signal_15668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4176 ( .C ( clk ), .D ( new_AGEMA_signal_15675 ), .Q ( new_AGEMA_signal_15676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4184 ( .C ( clk ), .D ( new_AGEMA_signal_15683 ), .Q ( new_AGEMA_signal_15684 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4192 ( .C ( clk ), .D ( new_AGEMA_signal_15691 ), .Q ( new_AGEMA_signal_15692 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4352 ( .C ( clk ), .D ( new_AGEMA_signal_15851 ), .Q ( new_AGEMA_signal_15852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4360 ( .C ( clk ), .D ( new_AGEMA_signal_15859 ), .Q ( new_AGEMA_signal_15860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4368 ( .C ( clk ), .D ( new_AGEMA_signal_15867 ), .Q ( new_AGEMA_signal_15868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4376 ( .C ( clk ), .D ( new_AGEMA_signal_15875 ), .Q ( new_AGEMA_signal_15876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4424 ( .C ( clk ), .D ( new_AGEMA_signal_15923 ), .Q ( new_AGEMA_signal_15924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4432 ( .C ( clk ), .D ( new_AGEMA_signal_15931 ), .Q ( new_AGEMA_signal_15932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4440 ( .C ( clk ), .D ( new_AGEMA_signal_15939 ), .Q ( new_AGEMA_signal_15940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4448 ( .C ( clk ), .D ( new_AGEMA_signal_15947 ), .Q ( new_AGEMA_signal_15948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4552 ( .C ( clk ), .D ( new_AGEMA_signal_16051 ), .Q ( new_AGEMA_signal_16052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4560 ( .C ( clk ), .D ( new_AGEMA_signal_16059 ), .Q ( new_AGEMA_signal_16060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4568 ( .C ( clk ), .D ( new_AGEMA_signal_16067 ), .Q ( new_AGEMA_signal_16068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4576 ( .C ( clk ), .D ( new_AGEMA_signal_16075 ), .Q ( new_AGEMA_signal_16076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4584 ( .C ( clk ), .D ( new_AGEMA_signal_16083 ), .Q ( new_AGEMA_signal_16084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4592 ( .C ( clk ), .D ( new_AGEMA_signal_16091 ), .Q ( new_AGEMA_signal_16092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4600 ( .C ( clk ), .D ( new_AGEMA_signal_16099 ), .Q ( new_AGEMA_signal_16100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4608 ( .C ( clk ), .D ( new_AGEMA_signal_16107 ), .Q ( new_AGEMA_signal_16108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4928 ( .C ( clk ), .D ( new_AGEMA_signal_16427 ), .Q ( new_AGEMA_signal_16428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4938 ( .C ( clk ), .D ( new_AGEMA_signal_16437 ), .Q ( new_AGEMA_signal_16438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4948 ( .C ( clk ), .D ( new_AGEMA_signal_16447 ), .Q ( new_AGEMA_signal_16448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4958 ( .C ( clk ), .D ( new_AGEMA_signal_16457 ), .Q ( new_AGEMA_signal_16458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5128 ( .C ( clk ), .D ( new_AGEMA_signal_16627 ), .Q ( new_AGEMA_signal_16628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5138 ( .C ( clk ), .D ( new_AGEMA_signal_16637 ), .Q ( new_AGEMA_signal_16638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5148 ( .C ( clk ), .D ( new_AGEMA_signal_16647 ), .Q ( new_AGEMA_signal_16648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5158 ( .C ( clk ), .D ( new_AGEMA_signal_16657 ), .Q ( new_AGEMA_signal_16658 ) ) ;

    /* cells in depth 7 */
    buf_clk new_AGEMA_reg_buffer_2289 ( .C ( clk ), .D ( new_AGEMA_signal_13788 ), .Q ( new_AGEMA_signal_13789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2293 ( .C ( clk ), .D ( new_AGEMA_signal_13792 ), .Q ( new_AGEMA_signal_13793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2297 ( .C ( clk ), .D ( new_AGEMA_signal_13796 ), .Q ( new_AGEMA_signal_13797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2301 ( .C ( clk ), .D ( new_AGEMA_signal_13800 ), .Q ( new_AGEMA_signal_13801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2305 ( .C ( clk ), .D ( new_AGEMA_signal_13804 ), .Q ( new_AGEMA_signal_13805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2309 ( .C ( clk ), .D ( new_AGEMA_signal_13808 ), .Q ( new_AGEMA_signal_13809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2313 ( .C ( clk ), .D ( new_AGEMA_signal_13812 ), .Q ( new_AGEMA_signal_13813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2317 ( .C ( clk ), .D ( new_AGEMA_signal_13816 ), .Q ( new_AGEMA_signal_13817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2319 ( .C ( clk ), .D ( new_AGEMA_signal_13636 ), .Q ( new_AGEMA_signal_13819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2321 ( .C ( clk ), .D ( new_AGEMA_signal_13638 ), .Q ( new_AGEMA_signal_13821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2323 ( .C ( clk ), .D ( new_AGEMA_signal_13640 ), .Q ( new_AGEMA_signal_13823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2325 ( .C ( clk ), .D ( new_AGEMA_signal_13642 ), .Q ( new_AGEMA_signal_13825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2327 ( .C ( clk ), .D ( n1966 ), .Q ( new_AGEMA_signal_13827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2329 ( .C ( clk ), .D ( new_AGEMA_signal_2079 ), .Q ( new_AGEMA_signal_13829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2331 ( .C ( clk ), .D ( new_AGEMA_signal_2080 ), .Q ( new_AGEMA_signal_13831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2333 ( .C ( clk ), .D ( new_AGEMA_signal_2081 ), .Q ( new_AGEMA_signal_13833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2337 ( .C ( clk ), .D ( new_AGEMA_signal_13836 ), .Q ( new_AGEMA_signal_13837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2341 ( .C ( clk ), .D ( new_AGEMA_signal_13840 ), .Q ( new_AGEMA_signal_13841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2345 ( .C ( clk ), .D ( new_AGEMA_signal_13844 ), .Q ( new_AGEMA_signal_13845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2349 ( .C ( clk ), .D ( new_AGEMA_signal_13848 ), .Q ( new_AGEMA_signal_13849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2351 ( .C ( clk ), .D ( new_AGEMA_signal_13492 ), .Q ( new_AGEMA_signal_13851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2353 ( .C ( clk ), .D ( new_AGEMA_signal_13494 ), .Q ( new_AGEMA_signal_13853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2355 ( .C ( clk ), .D ( new_AGEMA_signal_13496 ), .Q ( new_AGEMA_signal_13855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2357 ( .C ( clk ), .D ( new_AGEMA_signal_13498 ), .Q ( new_AGEMA_signal_13857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2361 ( .C ( clk ), .D ( new_AGEMA_signal_13860 ), .Q ( new_AGEMA_signal_13861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2365 ( .C ( clk ), .D ( new_AGEMA_signal_13864 ), .Q ( new_AGEMA_signal_13865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2369 ( .C ( clk ), .D ( new_AGEMA_signal_13868 ), .Q ( new_AGEMA_signal_13869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2373 ( .C ( clk ), .D ( new_AGEMA_signal_13872 ), .Q ( new_AGEMA_signal_13873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2375 ( .C ( clk ), .D ( n1996 ), .Q ( new_AGEMA_signal_13875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2377 ( .C ( clk ), .D ( new_AGEMA_signal_2109 ), .Q ( new_AGEMA_signal_13877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2379 ( .C ( clk ), .D ( new_AGEMA_signal_2110 ), .Q ( new_AGEMA_signal_13879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2381 ( .C ( clk ), .D ( new_AGEMA_signal_2111 ), .Q ( new_AGEMA_signal_13881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2385 ( .C ( clk ), .D ( new_AGEMA_signal_13884 ), .Q ( new_AGEMA_signal_13885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2389 ( .C ( clk ), .D ( new_AGEMA_signal_13888 ), .Q ( new_AGEMA_signal_13889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2393 ( .C ( clk ), .D ( new_AGEMA_signal_13892 ), .Q ( new_AGEMA_signal_13893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2397 ( .C ( clk ), .D ( new_AGEMA_signal_13896 ), .Q ( new_AGEMA_signal_13897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2401 ( .C ( clk ), .D ( new_AGEMA_signal_13900 ), .Q ( new_AGEMA_signal_13901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2405 ( .C ( clk ), .D ( new_AGEMA_signal_13904 ), .Q ( new_AGEMA_signal_13905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2409 ( .C ( clk ), .D ( new_AGEMA_signal_13908 ), .Q ( new_AGEMA_signal_13909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2413 ( .C ( clk ), .D ( new_AGEMA_signal_13912 ), .Q ( new_AGEMA_signal_13913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2415 ( .C ( clk ), .D ( n2033 ), .Q ( new_AGEMA_signal_13915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2417 ( .C ( clk ), .D ( new_AGEMA_signal_2127 ), .Q ( new_AGEMA_signal_13917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2419 ( .C ( clk ), .D ( new_AGEMA_signal_2128 ), .Q ( new_AGEMA_signal_13919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2421 ( .C ( clk ), .D ( new_AGEMA_signal_2129 ), .Q ( new_AGEMA_signal_13921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2423 ( .C ( clk ), .D ( new_AGEMA_signal_13316 ), .Q ( new_AGEMA_signal_13923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2425 ( .C ( clk ), .D ( new_AGEMA_signal_13318 ), .Q ( new_AGEMA_signal_13925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2427 ( .C ( clk ), .D ( new_AGEMA_signal_13320 ), .Q ( new_AGEMA_signal_13927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2429 ( .C ( clk ), .D ( new_AGEMA_signal_13322 ), .Q ( new_AGEMA_signal_13929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2431 ( .C ( clk ), .D ( new_AGEMA_signal_13356 ), .Q ( new_AGEMA_signal_13931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2433 ( .C ( clk ), .D ( new_AGEMA_signal_13358 ), .Q ( new_AGEMA_signal_13933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2435 ( .C ( clk ), .D ( new_AGEMA_signal_13360 ), .Q ( new_AGEMA_signal_13935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2437 ( .C ( clk ), .D ( new_AGEMA_signal_13362 ), .Q ( new_AGEMA_signal_13937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2439 ( .C ( clk ), .D ( new_AGEMA_signal_13468 ), .Q ( new_AGEMA_signal_13939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2441 ( .C ( clk ), .D ( new_AGEMA_signal_13470 ), .Q ( new_AGEMA_signal_13941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2443 ( .C ( clk ), .D ( new_AGEMA_signal_13472 ), .Q ( new_AGEMA_signal_13943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2445 ( .C ( clk ), .D ( new_AGEMA_signal_13474 ), .Q ( new_AGEMA_signal_13945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2449 ( .C ( clk ), .D ( new_AGEMA_signal_13948 ), .Q ( new_AGEMA_signal_13949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2453 ( .C ( clk ), .D ( new_AGEMA_signal_13952 ), .Q ( new_AGEMA_signal_13953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2457 ( .C ( clk ), .D ( new_AGEMA_signal_13956 ), .Q ( new_AGEMA_signal_13957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2461 ( .C ( clk ), .D ( new_AGEMA_signal_13960 ), .Q ( new_AGEMA_signal_13961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2465 ( .C ( clk ), .D ( new_AGEMA_signal_13964 ), .Q ( new_AGEMA_signal_13965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2469 ( .C ( clk ), .D ( new_AGEMA_signal_13968 ), .Q ( new_AGEMA_signal_13969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2473 ( .C ( clk ), .D ( new_AGEMA_signal_13972 ), .Q ( new_AGEMA_signal_13973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2477 ( .C ( clk ), .D ( new_AGEMA_signal_13976 ), .Q ( new_AGEMA_signal_13977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2481 ( .C ( clk ), .D ( new_AGEMA_signal_13980 ), .Q ( new_AGEMA_signal_13981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2485 ( .C ( clk ), .D ( new_AGEMA_signal_13984 ), .Q ( new_AGEMA_signal_13985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2489 ( .C ( clk ), .D ( new_AGEMA_signal_13988 ), .Q ( new_AGEMA_signal_13989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2493 ( .C ( clk ), .D ( new_AGEMA_signal_13992 ), .Q ( new_AGEMA_signal_13993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2495 ( .C ( clk ), .D ( n2089 ), .Q ( new_AGEMA_signal_13995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2497 ( .C ( clk ), .D ( new_AGEMA_signal_2172 ), .Q ( new_AGEMA_signal_13997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2499 ( .C ( clk ), .D ( new_AGEMA_signal_2173 ), .Q ( new_AGEMA_signal_13999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2501 ( .C ( clk ), .D ( new_AGEMA_signal_2174 ), .Q ( new_AGEMA_signal_14001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2503 ( .C ( clk ), .D ( n2092 ), .Q ( new_AGEMA_signal_14003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2505 ( .C ( clk ), .D ( new_AGEMA_signal_2178 ), .Q ( new_AGEMA_signal_14005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2507 ( .C ( clk ), .D ( new_AGEMA_signal_2179 ), .Q ( new_AGEMA_signal_14007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2509 ( .C ( clk ), .D ( new_AGEMA_signal_2180 ), .Q ( new_AGEMA_signal_14009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2511 ( .C ( clk ), .D ( n2115 ), .Q ( new_AGEMA_signal_14011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2513 ( .C ( clk ), .D ( new_AGEMA_signal_1686 ), .Q ( new_AGEMA_signal_14013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2515 ( .C ( clk ), .D ( new_AGEMA_signal_1687 ), .Q ( new_AGEMA_signal_14015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2517 ( .C ( clk ), .D ( new_AGEMA_signal_1688 ), .Q ( new_AGEMA_signal_14017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2521 ( .C ( clk ), .D ( new_AGEMA_signal_14020 ), .Q ( new_AGEMA_signal_14021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2525 ( .C ( clk ), .D ( new_AGEMA_signal_14024 ), .Q ( new_AGEMA_signal_14025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2529 ( .C ( clk ), .D ( new_AGEMA_signal_14028 ), .Q ( new_AGEMA_signal_14029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2533 ( .C ( clk ), .D ( new_AGEMA_signal_14032 ), .Q ( new_AGEMA_signal_14033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2535 ( .C ( clk ), .D ( n2687 ), .Q ( new_AGEMA_signal_14035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2537 ( .C ( clk ), .D ( new_AGEMA_signal_2076 ), .Q ( new_AGEMA_signal_14037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2539 ( .C ( clk ), .D ( new_AGEMA_signal_2077 ), .Q ( new_AGEMA_signal_14039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2541 ( .C ( clk ), .D ( new_AGEMA_signal_2078 ), .Q ( new_AGEMA_signal_14041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2545 ( .C ( clk ), .D ( new_AGEMA_signal_14044 ), .Q ( new_AGEMA_signal_14045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2549 ( .C ( clk ), .D ( new_AGEMA_signal_14048 ), .Q ( new_AGEMA_signal_14049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2553 ( .C ( clk ), .D ( new_AGEMA_signal_14052 ), .Q ( new_AGEMA_signal_14053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2557 ( .C ( clk ), .D ( new_AGEMA_signal_14056 ), .Q ( new_AGEMA_signal_14057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2563 ( .C ( clk ), .D ( new_AGEMA_signal_14062 ), .Q ( new_AGEMA_signal_14063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2569 ( .C ( clk ), .D ( new_AGEMA_signal_14068 ), .Q ( new_AGEMA_signal_14069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2575 ( .C ( clk ), .D ( new_AGEMA_signal_14074 ), .Q ( new_AGEMA_signal_14075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2581 ( .C ( clk ), .D ( new_AGEMA_signal_14080 ), .Q ( new_AGEMA_signal_14081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2585 ( .C ( clk ), .D ( new_AGEMA_signal_14084 ), .Q ( new_AGEMA_signal_14085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2589 ( .C ( clk ), .D ( new_AGEMA_signal_14088 ), .Q ( new_AGEMA_signal_14089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2593 ( .C ( clk ), .D ( new_AGEMA_signal_14092 ), .Q ( new_AGEMA_signal_14093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2597 ( .C ( clk ), .D ( new_AGEMA_signal_14096 ), .Q ( new_AGEMA_signal_14097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2601 ( .C ( clk ), .D ( new_AGEMA_signal_14100 ), .Q ( new_AGEMA_signal_14101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2605 ( .C ( clk ), .D ( new_AGEMA_signal_14104 ), .Q ( new_AGEMA_signal_14105 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2609 ( .C ( clk ), .D ( new_AGEMA_signal_14108 ), .Q ( new_AGEMA_signal_14109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2613 ( .C ( clk ), .D ( new_AGEMA_signal_14112 ), .Q ( new_AGEMA_signal_14113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2615 ( .C ( clk ), .D ( n2193 ), .Q ( new_AGEMA_signal_14115 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2617 ( .C ( clk ), .D ( new_AGEMA_signal_2232 ), .Q ( new_AGEMA_signal_14117 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2619 ( .C ( clk ), .D ( new_AGEMA_signal_2233 ), .Q ( new_AGEMA_signal_14119 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2621 ( .C ( clk ), .D ( new_AGEMA_signal_2234 ), .Q ( new_AGEMA_signal_14121 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2623 ( .C ( clk ), .D ( n2202 ), .Q ( new_AGEMA_signal_14123 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2625 ( .C ( clk ), .D ( new_AGEMA_signal_2664 ), .Q ( new_AGEMA_signal_14125 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2627 ( .C ( clk ), .D ( new_AGEMA_signal_2665 ), .Q ( new_AGEMA_signal_14127 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2629 ( .C ( clk ), .D ( new_AGEMA_signal_2666 ), .Q ( new_AGEMA_signal_14129 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2631 ( .C ( clk ), .D ( n2228 ), .Q ( new_AGEMA_signal_14131 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2633 ( .C ( clk ), .D ( new_AGEMA_signal_1758 ), .Q ( new_AGEMA_signal_14133 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2635 ( .C ( clk ), .D ( new_AGEMA_signal_1759 ), .Q ( new_AGEMA_signal_14135 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2637 ( .C ( clk ), .D ( new_AGEMA_signal_1760 ), .Q ( new_AGEMA_signal_14137 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2639 ( .C ( clk ), .D ( n2235 ), .Q ( new_AGEMA_signal_14139 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2641 ( .C ( clk ), .D ( new_AGEMA_signal_2061 ), .Q ( new_AGEMA_signal_14141 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2643 ( .C ( clk ), .D ( new_AGEMA_signal_2062 ), .Q ( new_AGEMA_signal_14143 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2645 ( .C ( clk ), .D ( new_AGEMA_signal_2063 ), .Q ( new_AGEMA_signal_14145 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2649 ( .C ( clk ), .D ( new_AGEMA_signal_14148 ), .Q ( new_AGEMA_signal_14149 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2653 ( .C ( clk ), .D ( new_AGEMA_signal_14152 ), .Q ( new_AGEMA_signal_14153 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2657 ( .C ( clk ), .D ( new_AGEMA_signal_14156 ), .Q ( new_AGEMA_signal_14157 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2661 ( .C ( clk ), .D ( new_AGEMA_signal_14160 ), .Q ( new_AGEMA_signal_14161 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2667 ( .C ( clk ), .D ( new_AGEMA_signal_14166 ), .Q ( new_AGEMA_signal_14167 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2673 ( .C ( clk ), .D ( new_AGEMA_signal_14172 ), .Q ( new_AGEMA_signal_14173 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2679 ( .C ( clk ), .D ( new_AGEMA_signal_14178 ), .Q ( new_AGEMA_signal_14179 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2685 ( .C ( clk ), .D ( new_AGEMA_signal_14184 ), .Q ( new_AGEMA_signal_14185 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2689 ( .C ( clk ), .D ( new_AGEMA_signal_14188 ), .Q ( new_AGEMA_signal_14189 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2693 ( .C ( clk ), .D ( new_AGEMA_signal_14192 ), .Q ( new_AGEMA_signal_14193 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2697 ( .C ( clk ), .D ( new_AGEMA_signal_14196 ), .Q ( new_AGEMA_signal_14197 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2701 ( .C ( clk ), .D ( new_AGEMA_signal_14200 ), .Q ( new_AGEMA_signal_14201 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2703 ( .C ( clk ), .D ( n2752 ), .Q ( new_AGEMA_signal_14203 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2705 ( .C ( clk ), .D ( new_AGEMA_signal_2691 ), .Q ( new_AGEMA_signal_14205 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2707 ( .C ( clk ), .D ( new_AGEMA_signal_2692 ), .Q ( new_AGEMA_signal_14207 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2709 ( .C ( clk ), .D ( new_AGEMA_signal_2693 ), .Q ( new_AGEMA_signal_14209 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2711 ( .C ( clk ), .D ( new_AGEMA_signal_13576 ), .Q ( new_AGEMA_signal_14211 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2713 ( .C ( clk ), .D ( new_AGEMA_signal_13582 ), .Q ( new_AGEMA_signal_14213 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2715 ( .C ( clk ), .D ( new_AGEMA_signal_13588 ), .Q ( new_AGEMA_signal_14215 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2717 ( .C ( clk ), .D ( new_AGEMA_signal_13594 ), .Q ( new_AGEMA_signal_14217 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2719 ( .C ( clk ), .D ( n2293 ), .Q ( new_AGEMA_signal_14219 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2721 ( .C ( clk ), .D ( new_AGEMA_signal_2295 ), .Q ( new_AGEMA_signal_14221 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2723 ( .C ( clk ), .D ( new_AGEMA_signal_2296 ), .Q ( new_AGEMA_signal_14223 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2725 ( .C ( clk ), .D ( new_AGEMA_signal_2297 ), .Q ( new_AGEMA_signal_14225 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2729 ( .C ( clk ), .D ( new_AGEMA_signal_14228 ), .Q ( new_AGEMA_signal_14229 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2733 ( .C ( clk ), .D ( new_AGEMA_signal_14232 ), .Q ( new_AGEMA_signal_14233 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2737 ( .C ( clk ), .D ( new_AGEMA_signal_14236 ), .Q ( new_AGEMA_signal_14237 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2741 ( .C ( clk ), .D ( new_AGEMA_signal_14240 ), .Q ( new_AGEMA_signal_14241 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2743 ( .C ( clk ), .D ( n2357 ), .Q ( new_AGEMA_signal_14243 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2745 ( .C ( clk ), .D ( new_AGEMA_signal_2322 ), .Q ( new_AGEMA_signal_14245 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2747 ( .C ( clk ), .D ( new_AGEMA_signal_2323 ), .Q ( new_AGEMA_signal_14247 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2749 ( .C ( clk ), .D ( new_AGEMA_signal_2324 ), .Q ( new_AGEMA_signal_14249 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2751 ( .C ( clk ), .D ( n2386 ), .Q ( new_AGEMA_signal_14251 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2753 ( .C ( clk ), .D ( new_AGEMA_signal_2337 ), .Q ( new_AGEMA_signal_14253 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2755 ( .C ( clk ), .D ( new_AGEMA_signal_2338 ), .Q ( new_AGEMA_signal_14255 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2757 ( .C ( clk ), .D ( new_AGEMA_signal_2339 ), .Q ( new_AGEMA_signal_14257 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2761 ( .C ( clk ), .D ( new_AGEMA_signal_14260 ), .Q ( new_AGEMA_signal_14261 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2765 ( .C ( clk ), .D ( new_AGEMA_signal_14264 ), .Q ( new_AGEMA_signal_14265 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2769 ( .C ( clk ), .D ( new_AGEMA_signal_14268 ), .Q ( new_AGEMA_signal_14269 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2773 ( .C ( clk ), .D ( new_AGEMA_signal_14272 ), .Q ( new_AGEMA_signal_14273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2777 ( .C ( clk ), .D ( new_AGEMA_signal_14276 ), .Q ( new_AGEMA_signal_14277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2781 ( .C ( clk ), .D ( new_AGEMA_signal_14280 ), .Q ( new_AGEMA_signal_14281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2785 ( .C ( clk ), .D ( new_AGEMA_signal_14284 ), .Q ( new_AGEMA_signal_14285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2789 ( .C ( clk ), .D ( new_AGEMA_signal_14288 ), .Q ( new_AGEMA_signal_14289 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2793 ( .C ( clk ), .D ( new_AGEMA_signal_14292 ), .Q ( new_AGEMA_signal_14293 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2797 ( .C ( clk ), .D ( new_AGEMA_signal_14296 ), .Q ( new_AGEMA_signal_14297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2801 ( .C ( clk ), .D ( new_AGEMA_signal_14300 ), .Q ( new_AGEMA_signal_14301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2805 ( .C ( clk ), .D ( new_AGEMA_signal_14304 ), .Q ( new_AGEMA_signal_14305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2809 ( .C ( clk ), .D ( new_AGEMA_signal_14308 ), .Q ( new_AGEMA_signal_14309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2813 ( .C ( clk ), .D ( new_AGEMA_signal_14312 ), .Q ( new_AGEMA_signal_14313 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2817 ( .C ( clk ), .D ( new_AGEMA_signal_14316 ), .Q ( new_AGEMA_signal_14317 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2821 ( .C ( clk ), .D ( new_AGEMA_signal_14320 ), .Q ( new_AGEMA_signal_14321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2825 ( .C ( clk ), .D ( new_AGEMA_signal_14324 ), .Q ( new_AGEMA_signal_14325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2829 ( .C ( clk ), .D ( new_AGEMA_signal_14328 ), .Q ( new_AGEMA_signal_14329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2833 ( .C ( clk ), .D ( new_AGEMA_signal_14332 ), .Q ( new_AGEMA_signal_14333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2837 ( .C ( clk ), .D ( new_AGEMA_signal_14336 ), .Q ( new_AGEMA_signal_14337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2839 ( .C ( clk ), .D ( n2433 ), .Q ( new_AGEMA_signal_14339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2841 ( .C ( clk ), .D ( new_AGEMA_signal_2358 ), .Q ( new_AGEMA_signal_14341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2843 ( .C ( clk ), .D ( new_AGEMA_signal_2359 ), .Q ( new_AGEMA_signal_14343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2845 ( .C ( clk ), .D ( new_AGEMA_signal_2360 ), .Q ( new_AGEMA_signal_14345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2847 ( .C ( clk ), .D ( new_AGEMA_signal_13342 ), .Q ( new_AGEMA_signal_14347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2849 ( .C ( clk ), .D ( new_AGEMA_signal_13346 ), .Q ( new_AGEMA_signal_14349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2851 ( .C ( clk ), .D ( new_AGEMA_signal_13350 ), .Q ( new_AGEMA_signal_14351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2853 ( .C ( clk ), .D ( new_AGEMA_signal_13354 ), .Q ( new_AGEMA_signal_14353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2855 ( .C ( clk ), .D ( n2459 ), .Q ( new_AGEMA_signal_14355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2857 ( .C ( clk ), .D ( new_AGEMA_signal_2286 ), .Q ( new_AGEMA_signal_14357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2859 ( .C ( clk ), .D ( new_AGEMA_signal_2287 ), .Q ( new_AGEMA_signal_14359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2861 ( .C ( clk ), .D ( new_AGEMA_signal_2288 ), .Q ( new_AGEMA_signal_14361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2863 ( .C ( clk ), .D ( n2467 ), .Q ( new_AGEMA_signal_14363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2865 ( .C ( clk ), .D ( new_AGEMA_signal_1854 ), .Q ( new_AGEMA_signal_14365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2867 ( .C ( clk ), .D ( new_AGEMA_signal_1855 ), .Q ( new_AGEMA_signal_14367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2869 ( .C ( clk ), .D ( new_AGEMA_signal_1856 ), .Q ( new_AGEMA_signal_14369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2873 ( .C ( clk ), .D ( new_AGEMA_signal_14372 ), .Q ( new_AGEMA_signal_14373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2877 ( .C ( clk ), .D ( new_AGEMA_signal_14376 ), .Q ( new_AGEMA_signal_14377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2881 ( .C ( clk ), .D ( new_AGEMA_signal_14380 ), .Q ( new_AGEMA_signal_14381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2885 ( .C ( clk ), .D ( new_AGEMA_signal_14384 ), .Q ( new_AGEMA_signal_14385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2889 ( .C ( clk ), .D ( new_AGEMA_signal_14388 ), .Q ( new_AGEMA_signal_14389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2893 ( .C ( clk ), .D ( new_AGEMA_signal_14392 ), .Q ( new_AGEMA_signal_14393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2897 ( .C ( clk ), .D ( new_AGEMA_signal_14396 ), .Q ( new_AGEMA_signal_14397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2901 ( .C ( clk ), .D ( new_AGEMA_signal_14400 ), .Q ( new_AGEMA_signal_14401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2903 ( .C ( clk ), .D ( n2489 ), .Q ( new_AGEMA_signal_14403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2905 ( .C ( clk ), .D ( new_AGEMA_signal_1914 ), .Q ( new_AGEMA_signal_14405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2907 ( .C ( clk ), .D ( new_AGEMA_signal_1915 ), .Q ( new_AGEMA_signal_14407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2909 ( .C ( clk ), .D ( new_AGEMA_signal_1916 ), .Q ( new_AGEMA_signal_14409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2911 ( .C ( clk ), .D ( n2497 ), .Q ( new_AGEMA_signal_14411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2913 ( .C ( clk ), .D ( new_AGEMA_signal_1917 ), .Q ( new_AGEMA_signal_14413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2915 ( .C ( clk ), .D ( new_AGEMA_signal_1918 ), .Q ( new_AGEMA_signal_14415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2917 ( .C ( clk ), .D ( new_AGEMA_signal_1919 ), .Q ( new_AGEMA_signal_14417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2919 ( .C ( clk ), .D ( n2506 ), .Q ( new_AGEMA_signal_14419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2921 ( .C ( clk ), .D ( new_AGEMA_signal_2397 ), .Q ( new_AGEMA_signal_14421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2923 ( .C ( clk ), .D ( new_AGEMA_signal_2398 ), .Q ( new_AGEMA_signal_14423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2925 ( .C ( clk ), .D ( new_AGEMA_signal_2399 ), .Q ( new_AGEMA_signal_14425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2927 ( .C ( clk ), .D ( n2542 ), .Q ( new_AGEMA_signal_14427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2929 ( .C ( clk ), .D ( new_AGEMA_signal_2415 ), .Q ( new_AGEMA_signal_14429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2931 ( .C ( clk ), .D ( new_AGEMA_signal_2416 ), .Q ( new_AGEMA_signal_14431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2933 ( .C ( clk ), .D ( new_AGEMA_signal_2417 ), .Q ( new_AGEMA_signal_14433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2935 ( .C ( clk ), .D ( n2558 ), .Q ( new_AGEMA_signal_14435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2937 ( .C ( clk ), .D ( new_AGEMA_signal_2424 ), .Q ( new_AGEMA_signal_14437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2939 ( .C ( clk ), .D ( new_AGEMA_signal_2425 ), .Q ( new_AGEMA_signal_14439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2941 ( .C ( clk ), .D ( new_AGEMA_signal_2426 ), .Q ( new_AGEMA_signal_14441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2943 ( .C ( clk ), .D ( n2566 ), .Q ( new_AGEMA_signal_14443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2945 ( .C ( clk ), .D ( new_AGEMA_signal_2430 ), .Q ( new_AGEMA_signal_14445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2947 ( .C ( clk ), .D ( new_AGEMA_signal_2431 ), .Q ( new_AGEMA_signal_14447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2949 ( .C ( clk ), .D ( new_AGEMA_signal_2432 ), .Q ( new_AGEMA_signal_14449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2951 ( .C ( clk ), .D ( n2581 ), .Q ( new_AGEMA_signal_14451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2953 ( .C ( clk ), .D ( new_AGEMA_signal_1944 ), .Q ( new_AGEMA_signal_14453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2955 ( .C ( clk ), .D ( new_AGEMA_signal_1945 ), .Q ( new_AGEMA_signal_14455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2957 ( .C ( clk ), .D ( new_AGEMA_signal_1946 ), .Q ( new_AGEMA_signal_14457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2959 ( .C ( clk ), .D ( n2603 ), .Q ( new_AGEMA_signal_14459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2961 ( .C ( clk ), .D ( new_AGEMA_signal_2454 ), .Q ( new_AGEMA_signal_14461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2963 ( .C ( clk ), .D ( new_AGEMA_signal_2455 ), .Q ( new_AGEMA_signal_14463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2965 ( .C ( clk ), .D ( new_AGEMA_signal_2456 ), .Q ( new_AGEMA_signal_14465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2967 ( .C ( clk ), .D ( n2620 ), .Q ( new_AGEMA_signal_14467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2969 ( .C ( clk ), .D ( new_AGEMA_signal_2457 ), .Q ( new_AGEMA_signal_14469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2971 ( .C ( clk ), .D ( new_AGEMA_signal_2458 ), .Q ( new_AGEMA_signal_14471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2973 ( .C ( clk ), .D ( new_AGEMA_signal_2459 ), .Q ( new_AGEMA_signal_14473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2977 ( .C ( clk ), .D ( new_AGEMA_signal_14476 ), .Q ( new_AGEMA_signal_14477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2981 ( .C ( clk ), .D ( new_AGEMA_signal_14480 ), .Q ( new_AGEMA_signal_14481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2985 ( .C ( clk ), .D ( new_AGEMA_signal_14484 ), .Q ( new_AGEMA_signal_14485 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2989 ( .C ( clk ), .D ( new_AGEMA_signal_14488 ), .Q ( new_AGEMA_signal_14489 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2991 ( .C ( clk ), .D ( n2653 ), .Q ( new_AGEMA_signal_14491 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2993 ( .C ( clk ), .D ( new_AGEMA_signal_1983 ), .Q ( new_AGEMA_signal_14493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2995 ( .C ( clk ), .D ( new_AGEMA_signal_1984 ), .Q ( new_AGEMA_signal_14495 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2997 ( .C ( clk ), .D ( new_AGEMA_signal_1985 ), .Q ( new_AGEMA_signal_14497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2999 ( .C ( clk ), .D ( n2665 ), .Q ( new_AGEMA_signal_14499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3001 ( .C ( clk ), .D ( new_AGEMA_signal_2055 ), .Q ( new_AGEMA_signal_14501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3003 ( .C ( clk ), .D ( new_AGEMA_signal_2056 ), .Q ( new_AGEMA_signal_14503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3005 ( .C ( clk ), .D ( new_AGEMA_signal_2057 ), .Q ( new_AGEMA_signal_14505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3007 ( .C ( clk ), .D ( n2691 ), .Q ( new_AGEMA_signal_14507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3009 ( .C ( clk ), .D ( new_AGEMA_signal_1992 ), .Q ( new_AGEMA_signal_14509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3011 ( .C ( clk ), .D ( new_AGEMA_signal_1993 ), .Q ( new_AGEMA_signal_14511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3013 ( .C ( clk ), .D ( new_AGEMA_signal_1994 ), .Q ( new_AGEMA_signal_14513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3015 ( .C ( clk ), .D ( n2717 ), .Q ( new_AGEMA_signal_14515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3017 ( .C ( clk ), .D ( new_AGEMA_signal_2484 ), .Q ( new_AGEMA_signal_14517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3019 ( .C ( clk ), .D ( new_AGEMA_signal_2485 ), .Q ( new_AGEMA_signal_14519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3021 ( .C ( clk ), .D ( new_AGEMA_signal_2486 ), .Q ( new_AGEMA_signal_14521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3023 ( .C ( clk ), .D ( n2729 ), .Q ( new_AGEMA_signal_14523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3025 ( .C ( clk ), .D ( new_AGEMA_signal_2844 ), .Q ( new_AGEMA_signal_14525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3027 ( .C ( clk ), .D ( new_AGEMA_signal_2845 ), .Q ( new_AGEMA_signal_14527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3029 ( .C ( clk ), .D ( new_AGEMA_signal_2846 ), .Q ( new_AGEMA_signal_14529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3033 ( .C ( clk ), .D ( new_AGEMA_signal_14532 ), .Q ( new_AGEMA_signal_14533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3037 ( .C ( clk ), .D ( new_AGEMA_signal_14536 ), .Q ( new_AGEMA_signal_14537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3041 ( .C ( clk ), .D ( new_AGEMA_signal_14540 ), .Q ( new_AGEMA_signal_14541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3045 ( .C ( clk ), .D ( new_AGEMA_signal_14544 ), .Q ( new_AGEMA_signal_14545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3049 ( .C ( clk ), .D ( new_AGEMA_signal_14548 ), .Q ( new_AGEMA_signal_14549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3053 ( .C ( clk ), .D ( new_AGEMA_signal_14552 ), .Q ( new_AGEMA_signal_14553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3057 ( .C ( clk ), .D ( new_AGEMA_signal_14556 ), .Q ( new_AGEMA_signal_14557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3061 ( .C ( clk ), .D ( new_AGEMA_signal_14560 ), .Q ( new_AGEMA_signal_14561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3065 ( .C ( clk ), .D ( new_AGEMA_signal_14564 ), .Q ( new_AGEMA_signal_14565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3069 ( .C ( clk ), .D ( new_AGEMA_signal_14568 ), .Q ( new_AGEMA_signal_14569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3073 ( .C ( clk ), .D ( new_AGEMA_signal_14572 ), .Q ( new_AGEMA_signal_14573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3077 ( .C ( clk ), .D ( new_AGEMA_signal_14576 ), .Q ( new_AGEMA_signal_14577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3081 ( .C ( clk ), .D ( new_AGEMA_signal_14580 ), .Q ( new_AGEMA_signal_14581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3085 ( .C ( clk ), .D ( new_AGEMA_signal_14584 ), .Q ( new_AGEMA_signal_14585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3089 ( .C ( clk ), .D ( new_AGEMA_signal_14588 ), .Q ( new_AGEMA_signal_14589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3093 ( .C ( clk ), .D ( new_AGEMA_signal_14592 ), .Q ( new_AGEMA_signal_14593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3095 ( .C ( clk ), .D ( new_AGEMA_signal_13524 ), .Q ( new_AGEMA_signal_14595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3099 ( .C ( clk ), .D ( new_AGEMA_signal_13526 ), .Q ( new_AGEMA_signal_14599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3103 ( .C ( clk ), .D ( new_AGEMA_signal_13528 ), .Q ( new_AGEMA_signal_14603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3107 ( .C ( clk ), .D ( new_AGEMA_signal_13530 ), .Q ( new_AGEMA_signal_14607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3111 ( .C ( clk ), .D ( n1956 ), .Q ( new_AGEMA_signal_14611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3115 ( .C ( clk ), .D ( new_AGEMA_signal_2067 ), .Q ( new_AGEMA_signal_14615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3119 ( .C ( clk ), .D ( new_AGEMA_signal_2068 ), .Q ( new_AGEMA_signal_14619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3123 ( .C ( clk ), .D ( new_AGEMA_signal_2069 ), .Q ( new_AGEMA_signal_14623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3131 ( .C ( clk ), .D ( new_AGEMA_signal_14630 ), .Q ( new_AGEMA_signal_14631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3139 ( .C ( clk ), .D ( new_AGEMA_signal_14638 ), .Q ( new_AGEMA_signal_14639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3147 ( .C ( clk ), .D ( new_AGEMA_signal_14646 ), .Q ( new_AGEMA_signal_14647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3155 ( .C ( clk ), .D ( new_AGEMA_signal_14654 ), .Q ( new_AGEMA_signal_14655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3171 ( .C ( clk ), .D ( new_AGEMA_signal_14670 ), .Q ( new_AGEMA_signal_14671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3179 ( .C ( clk ), .D ( new_AGEMA_signal_14678 ), .Q ( new_AGEMA_signal_14679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3187 ( .C ( clk ), .D ( new_AGEMA_signal_14686 ), .Q ( new_AGEMA_signal_14687 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3195 ( .C ( clk ), .D ( new_AGEMA_signal_14694 ), .Q ( new_AGEMA_signal_14695 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3201 ( .C ( clk ), .D ( new_AGEMA_signal_14700 ), .Q ( new_AGEMA_signal_14701 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3207 ( .C ( clk ), .D ( new_AGEMA_signal_14706 ), .Q ( new_AGEMA_signal_14707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3213 ( .C ( clk ), .D ( new_AGEMA_signal_14712 ), .Q ( new_AGEMA_signal_14713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3219 ( .C ( clk ), .D ( new_AGEMA_signal_14718 ), .Q ( new_AGEMA_signal_14719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3223 ( .C ( clk ), .D ( n2023 ), .Q ( new_AGEMA_signal_14723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3227 ( .C ( clk ), .D ( new_AGEMA_signal_1614 ), .Q ( new_AGEMA_signal_14727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3231 ( .C ( clk ), .D ( new_AGEMA_signal_1615 ), .Q ( new_AGEMA_signal_14731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3235 ( .C ( clk ), .D ( new_AGEMA_signal_1616 ), .Q ( new_AGEMA_signal_14735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3241 ( .C ( clk ), .D ( new_AGEMA_signal_14740 ), .Q ( new_AGEMA_signal_14741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3247 ( .C ( clk ), .D ( new_AGEMA_signal_14746 ), .Q ( new_AGEMA_signal_14747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3253 ( .C ( clk ), .D ( new_AGEMA_signal_14752 ), .Q ( new_AGEMA_signal_14753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3259 ( .C ( clk ), .D ( new_AGEMA_signal_14758 ), .Q ( new_AGEMA_signal_14759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3273 ( .C ( clk ), .D ( new_AGEMA_signal_14772 ), .Q ( new_AGEMA_signal_14773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3279 ( .C ( clk ), .D ( new_AGEMA_signal_14778 ), .Q ( new_AGEMA_signal_14779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3285 ( .C ( clk ), .D ( new_AGEMA_signal_14784 ), .Q ( new_AGEMA_signal_14785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3291 ( .C ( clk ), .D ( new_AGEMA_signal_14790 ), .Q ( new_AGEMA_signal_14791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3297 ( .C ( clk ), .D ( new_AGEMA_signal_14796 ), .Q ( new_AGEMA_signal_14797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3303 ( .C ( clk ), .D ( new_AGEMA_signal_14802 ), .Q ( new_AGEMA_signal_14803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3309 ( .C ( clk ), .D ( new_AGEMA_signal_14808 ), .Q ( new_AGEMA_signal_14809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3315 ( .C ( clk ), .D ( new_AGEMA_signal_14814 ), .Q ( new_AGEMA_signal_14815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3327 ( .C ( clk ), .D ( n2094 ), .Q ( new_AGEMA_signal_14827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3331 ( .C ( clk ), .D ( new_AGEMA_signal_2181 ), .Q ( new_AGEMA_signal_14831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3335 ( .C ( clk ), .D ( new_AGEMA_signal_2182 ), .Q ( new_AGEMA_signal_14835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3339 ( .C ( clk ), .D ( new_AGEMA_signal_2183 ), .Q ( new_AGEMA_signal_14839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3345 ( .C ( clk ), .D ( new_AGEMA_signal_14844 ), .Q ( new_AGEMA_signal_14845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3351 ( .C ( clk ), .D ( new_AGEMA_signal_14850 ), .Q ( new_AGEMA_signal_14851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3357 ( .C ( clk ), .D ( new_AGEMA_signal_14856 ), .Q ( new_AGEMA_signal_14857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3363 ( .C ( clk ), .D ( new_AGEMA_signal_14862 ), .Q ( new_AGEMA_signal_14863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3369 ( .C ( clk ), .D ( new_AGEMA_signal_14868 ), .Q ( new_AGEMA_signal_14869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3375 ( .C ( clk ), .D ( new_AGEMA_signal_14874 ), .Q ( new_AGEMA_signal_14875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3381 ( .C ( clk ), .D ( new_AGEMA_signal_14880 ), .Q ( new_AGEMA_signal_14881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3387 ( .C ( clk ), .D ( new_AGEMA_signal_14886 ), .Q ( new_AGEMA_signal_14887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3401 ( .C ( clk ), .D ( new_AGEMA_signal_14900 ), .Q ( new_AGEMA_signal_14901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3407 ( .C ( clk ), .D ( new_AGEMA_signal_14906 ), .Q ( new_AGEMA_signal_14907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3413 ( .C ( clk ), .D ( new_AGEMA_signal_14912 ), .Q ( new_AGEMA_signal_14913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3419 ( .C ( clk ), .D ( new_AGEMA_signal_14918 ), .Q ( new_AGEMA_signal_14919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3431 ( .C ( clk ), .D ( n2181 ), .Q ( new_AGEMA_signal_14931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3435 ( .C ( clk ), .D ( new_AGEMA_signal_2223 ), .Q ( new_AGEMA_signal_14935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3439 ( .C ( clk ), .D ( new_AGEMA_signal_2224 ), .Q ( new_AGEMA_signal_14939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3443 ( .C ( clk ), .D ( new_AGEMA_signal_2225 ), .Q ( new_AGEMA_signal_14943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3447 ( .C ( clk ), .D ( n2195 ), .Q ( new_AGEMA_signal_14947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3451 ( .C ( clk ), .D ( new_AGEMA_signal_2229 ), .Q ( new_AGEMA_signal_14951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3455 ( .C ( clk ), .D ( new_AGEMA_signal_2230 ), .Q ( new_AGEMA_signal_14955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3459 ( .C ( clk ), .D ( new_AGEMA_signal_2231 ), .Q ( new_AGEMA_signal_14959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3475 ( .C ( clk ), .D ( new_AGEMA_signal_14974 ), .Q ( new_AGEMA_signal_14975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3483 ( .C ( clk ), .D ( new_AGEMA_signal_14982 ), .Q ( new_AGEMA_signal_14983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3491 ( .C ( clk ), .D ( new_AGEMA_signal_14990 ), .Q ( new_AGEMA_signal_14991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3499 ( .C ( clk ), .D ( new_AGEMA_signal_14998 ), .Q ( new_AGEMA_signal_14999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3505 ( .C ( clk ), .D ( new_AGEMA_signal_15004 ), .Q ( new_AGEMA_signal_15005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3511 ( .C ( clk ), .D ( new_AGEMA_signal_15010 ), .Q ( new_AGEMA_signal_15011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3517 ( .C ( clk ), .D ( new_AGEMA_signal_15016 ), .Q ( new_AGEMA_signal_15017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3523 ( .C ( clk ), .D ( new_AGEMA_signal_15022 ), .Q ( new_AGEMA_signal_15023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3527 ( .C ( clk ), .D ( n2237 ), .Q ( new_AGEMA_signal_15027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3531 ( .C ( clk ), .D ( new_AGEMA_signal_1761 ), .Q ( new_AGEMA_signal_15031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3535 ( .C ( clk ), .D ( new_AGEMA_signal_1762 ), .Q ( new_AGEMA_signal_15035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3539 ( .C ( clk ), .D ( new_AGEMA_signal_1763 ), .Q ( new_AGEMA_signal_15039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3543 ( .C ( clk ), .D ( n2248 ), .Q ( new_AGEMA_signal_15043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3547 ( .C ( clk ), .D ( new_AGEMA_signal_2256 ), .Q ( new_AGEMA_signal_15047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3551 ( .C ( clk ), .D ( new_AGEMA_signal_2257 ), .Q ( new_AGEMA_signal_15051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3555 ( .C ( clk ), .D ( new_AGEMA_signal_2258 ), .Q ( new_AGEMA_signal_15055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3575 ( .C ( clk ), .D ( n2294 ), .Q ( new_AGEMA_signal_15075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3579 ( .C ( clk ), .D ( new_AGEMA_signal_1806 ), .Q ( new_AGEMA_signal_15079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3583 ( .C ( clk ), .D ( new_AGEMA_signal_1807 ), .Q ( new_AGEMA_signal_15083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3587 ( .C ( clk ), .D ( new_AGEMA_signal_1808 ), .Q ( new_AGEMA_signal_15087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3591 ( .C ( clk ), .D ( n2323 ), .Q ( new_AGEMA_signal_15091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3595 ( .C ( clk ), .D ( new_AGEMA_signal_2301 ), .Q ( new_AGEMA_signal_15095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3599 ( .C ( clk ), .D ( new_AGEMA_signal_2302 ), .Q ( new_AGEMA_signal_15099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3603 ( .C ( clk ), .D ( new_AGEMA_signal_2303 ), .Q ( new_AGEMA_signal_15103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3617 ( .C ( clk ), .D ( new_AGEMA_signal_15116 ), .Q ( new_AGEMA_signal_15117 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3623 ( .C ( clk ), .D ( new_AGEMA_signal_15122 ), .Q ( new_AGEMA_signal_15123 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3629 ( .C ( clk ), .D ( new_AGEMA_signal_15128 ), .Q ( new_AGEMA_signal_15129 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3635 ( .C ( clk ), .D ( new_AGEMA_signal_15134 ), .Q ( new_AGEMA_signal_15135 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3639 ( .C ( clk ), .D ( n2360 ), .Q ( new_AGEMA_signal_15139 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3643 ( .C ( clk ), .D ( new_AGEMA_signal_2325 ), .Q ( new_AGEMA_signal_15143 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3647 ( .C ( clk ), .D ( new_AGEMA_signal_2326 ), .Q ( new_AGEMA_signal_15147 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3651 ( .C ( clk ), .D ( new_AGEMA_signal_2327 ), .Q ( new_AGEMA_signal_15151 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3663 ( .C ( clk ), .D ( n2394 ), .Q ( new_AGEMA_signal_15163 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3667 ( .C ( clk ), .D ( new_AGEMA_signal_1863 ), .Q ( new_AGEMA_signal_15167 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3671 ( .C ( clk ), .D ( new_AGEMA_signal_1864 ), .Q ( new_AGEMA_signal_15171 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3675 ( .C ( clk ), .D ( new_AGEMA_signal_1865 ), .Q ( new_AGEMA_signal_15175 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3679 ( .C ( clk ), .D ( n2406 ), .Q ( new_AGEMA_signal_15179 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3683 ( .C ( clk ), .D ( new_AGEMA_signal_2343 ), .Q ( new_AGEMA_signal_15183 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3687 ( .C ( clk ), .D ( new_AGEMA_signal_2344 ), .Q ( new_AGEMA_signal_15187 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3691 ( .C ( clk ), .D ( new_AGEMA_signal_2345 ), .Q ( new_AGEMA_signal_15191 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3695 ( .C ( clk ), .D ( new_AGEMA_signal_13124 ), .Q ( new_AGEMA_signal_15195 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3699 ( .C ( clk ), .D ( new_AGEMA_signal_13126 ), .Q ( new_AGEMA_signal_15199 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3703 ( .C ( clk ), .D ( new_AGEMA_signal_13128 ), .Q ( new_AGEMA_signal_15203 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3707 ( .C ( clk ), .D ( new_AGEMA_signal_13130 ), .Q ( new_AGEMA_signal_15207 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3719 ( .C ( clk ), .D ( new_AGEMA_signal_13132 ), .Q ( new_AGEMA_signal_15219 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3723 ( .C ( clk ), .D ( new_AGEMA_signal_13134 ), .Q ( new_AGEMA_signal_15223 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3727 ( .C ( clk ), .D ( new_AGEMA_signal_13136 ), .Q ( new_AGEMA_signal_15227 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3731 ( .C ( clk ), .D ( new_AGEMA_signal_13138 ), .Q ( new_AGEMA_signal_15231 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3745 ( .C ( clk ), .D ( new_AGEMA_signal_15244 ), .Q ( new_AGEMA_signal_15245 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3751 ( .C ( clk ), .D ( new_AGEMA_signal_15250 ), .Q ( new_AGEMA_signal_15251 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3757 ( .C ( clk ), .D ( new_AGEMA_signal_15256 ), .Q ( new_AGEMA_signal_15257 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3763 ( .C ( clk ), .D ( new_AGEMA_signal_15262 ), .Q ( new_AGEMA_signal_15263 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3769 ( .C ( clk ), .D ( new_AGEMA_signal_15268 ), .Q ( new_AGEMA_signal_15269 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3775 ( .C ( clk ), .D ( new_AGEMA_signal_15274 ), .Q ( new_AGEMA_signal_15275 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3781 ( .C ( clk ), .D ( new_AGEMA_signal_15280 ), .Q ( new_AGEMA_signal_15281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3787 ( .C ( clk ), .D ( new_AGEMA_signal_15286 ), .Q ( new_AGEMA_signal_15287 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3791 ( .C ( clk ), .D ( n2499 ), .Q ( new_AGEMA_signal_15291 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3795 ( .C ( clk ), .D ( new_AGEMA_signal_1923 ), .Q ( new_AGEMA_signal_15295 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3799 ( .C ( clk ), .D ( new_AGEMA_signal_1924 ), .Q ( new_AGEMA_signal_15299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3803 ( .C ( clk ), .D ( new_AGEMA_signal_1925 ), .Q ( new_AGEMA_signal_15303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3819 ( .C ( clk ), .D ( new_AGEMA_signal_15318 ), .Q ( new_AGEMA_signal_15319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3827 ( .C ( clk ), .D ( new_AGEMA_signal_15326 ), .Q ( new_AGEMA_signal_15327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3835 ( .C ( clk ), .D ( new_AGEMA_signal_15334 ), .Q ( new_AGEMA_signal_15335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3843 ( .C ( clk ), .D ( new_AGEMA_signal_15342 ), .Q ( new_AGEMA_signal_15343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3855 ( .C ( clk ), .D ( n2582 ), .Q ( new_AGEMA_signal_15355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3859 ( .C ( clk ), .D ( new_AGEMA_signal_2445 ), .Q ( new_AGEMA_signal_15359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3863 ( .C ( clk ), .D ( new_AGEMA_signal_2446 ), .Q ( new_AGEMA_signal_15363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3867 ( .C ( clk ), .D ( new_AGEMA_signal_2447 ), .Q ( new_AGEMA_signal_15367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3871 ( .C ( clk ), .D ( n2605 ), .Q ( new_AGEMA_signal_15371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3875 ( .C ( clk ), .D ( new_AGEMA_signal_2451 ), .Q ( new_AGEMA_signal_15375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3879 ( .C ( clk ), .D ( new_AGEMA_signal_2452 ), .Q ( new_AGEMA_signal_15379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3883 ( .C ( clk ), .D ( new_AGEMA_signal_2453 ), .Q ( new_AGEMA_signal_15383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3887 ( .C ( clk ), .D ( n2632 ), .Q ( new_AGEMA_signal_15387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3891 ( .C ( clk ), .D ( new_AGEMA_signal_1974 ), .Q ( new_AGEMA_signal_15391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3895 ( .C ( clk ), .D ( new_AGEMA_signal_1975 ), .Q ( new_AGEMA_signal_15395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3899 ( .C ( clk ), .D ( new_AGEMA_signal_1976 ), .Q ( new_AGEMA_signal_15399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3903 ( .C ( clk ), .D ( n2655 ), .Q ( new_AGEMA_signal_15403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3907 ( .C ( clk ), .D ( new_AGEMA_signal_2472 ), .Q ( new_AGEMA_signal_15407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3911 ( .C ( clk ), .D ( new_AGEMA_signal_2473 ), .Q ( new_AGEMA_signal_15411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3915 ( .C ( clk ), .D ( new_AGEMA_signal_2474 ), .Q ( new_AGEMA_signal_15415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3919 ( .C ( clk ), .D ( n2695 ), .Q ( new_AGEMA_signal_15419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3923 ( .C ( clk ), .D ( new_AGEMA_signal_2481 ), .Q ( new_AGEMA_signal_15423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3927 ( .C ( clk ), .D ( new_AGEMA_signal_2482 ), .Q ( new_AGEMA_signal_15427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3931 ( .C ( clk ), .D ( new_AGEMA_signal_2483 ), .Q ( new_AGEMA_signal_15431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3939 ( .C ( clk ), .D ( new_AGEMA_signal_15438 ), .Q ( new_AGEMA_signal_15439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3947 ( .C ( clk ), .D ( new_AGEMA_signal_15446 ), .Q ( new_AGEMA_signal_15447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3955 ( .C ( clk ), .D ( new_AGEMA_signal_15454 ), .Q ( new_AGEMA_signal_15455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3963 ( .C ( clk ), .D ( new_AGEMA_signal_15462 ), .Q ( new_AGEMA_signal_15463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3975 ( .C ( clk ), .D ( n2770 ), .Q ( new_AGEMA_signal_15475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3979 ( .C ( clk ), .D ( new_AGEMA_signal_2505 ), .Q ( new_AGEMA_signal_15479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3983 ( .C ( clk ), .D ( new_AGEMA_signal_2506 ), .Q ( new_AGEMA_signal_15483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3987 ( .C ( clk ), .D ( new_AGEMA_signal_2507 ), .Q ( new_AGEMA_signal_15487 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4001 ( .C ( clk ), .D ( new_AGEMA_signal_15500 ), .Q ( new_AGEMA_signal_15501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4007 ( .C ( clk ), .D ( new_AGEMA_signal_15506 ), .Q ( new_AGEMA_signal_15507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4013 ( .C ( clk ), .D ( new_AGEMA_signal_15512 ), .Q ( new_AGEMA_signal_15513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4019 ( .C ( clk ), .D ( new_AGEMA_signal_15518 ), .Q ( new_AGEMA_signal_15519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4033 ( .C ( clk ), .D ( new_AGEMA_signal_15532 ), .Q ( new_AGEMA_signal_15533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4041 ( .C ( clk ), .D ( new_AGEMA_signal_15540 ), .Q ( new_AGEMA_signal_15541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4049 ( .C ( clk ), .D ( new_AGEMA_signal_15548 ), .Q ( new_AGEMA_signal_15549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4057 ( .C ( clk ), .D ( new_AGEMA_signal_15556 ), .Q ( new_AGEMA_signal_15557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4089 ( .C ( clk ), .D ( new_AGEMA_signal_15588 ), .Q ( new_AGEMA_signal_15589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4097 ( .C ( clk ), .D ( new_AGEMA_signal_15596 ), .Q ( new_AGEMA_signal_15597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4105 ( .C ( clk ), .D ( new_AGEMA_signal_15604 ), .Q ( new_AGEMA_signal_15605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4113 ( .C ( clk ), .D ( new_AGEMA_signal_15612 ), .Q ( new_AGEMA_signal_15613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4127 ( .C ( clk ), .D ( n2050 ), .Q ( new_AGEMA_signal_15627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4133 ( .C ( clk ), .D ( new_AGEMA_signal_1629 ), .Q ( new_AGEMA_signal_15633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4139 ( .C ( clk ), .D ( new_AGEMA_signal_1630 ), .Q ( new_AGEMA_signal_15639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4145 ( .C ( clk ), .D ( new_AGEMA_signal_1631 ), .Q ( new_AGEMA_signal_15645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4169 ( .C ( clk ), .D ( new_AGEMA_signal_15668 ), .Q ( new_AGEMA_signal_15669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4177 ( .C ( clk ), .D ( new_AGEMA_signal_15676 ), .Q ( new_AGEMA_signal_15677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4185 ( .C ( clk ), .D ( new_AGEMA_signal_15684 ), .Q ( new_AGEMA_signal_15685 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4193 ( .C ( clk ), .D ( new_AGEMA_signal_15692 ), .Q ( new_AGEMA_signal_15693 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4215 ( .C ( clk ), .D ( n2183 ), .Q ( new_AGEMA_signal_15715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4221 ( .C ( clk ), .D ( new_AGEMA_signal_1374 ), .Q ( new_AGEMA_signal_15721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4227 ( .C ( clk ), .D ( new_AGEMA_signal_1375 ), .Q ( new_AGEMA_signal_15727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4233 ( .C ( clk ), .D ( new_AGEMA_signal_1376 ), .Q ( new_AGEMA_signal_15733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4239 ( .C ( clk ), .D ( n2196 ), .Q ( new_AGEMA_signal_15739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4245 ( .C ( clk ), .D ( new_AGEMA_signal_1743 ), .Q ( new_AGEMA_signal_15745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4251 ( .C ( clk ), .D ( new_AGEMA_signal_1744 ), .Q ( new_AGEMA_signal_15751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4257 ( .C ( clk ), .D ( new_AGEMA_signal_1745 ), .Q ( new_AGEMA_signal_15757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4263 ( .C ( clk ), .D ( n2238 ), .Q ( new_AGEMA_signal_15763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4269 ( .C ( clk ), .D ( new_AGEMA_signal_1764 ), .Q ( new_AGEMA_signal_15769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4275 ( .C ( clk ), .D ( new_AGEMA_signal_1765 ), .Q ( new_AGEMA_signal_15775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4281 ( .C ( clk ), .D ( new_AGEMA_signal_1766 ), .Q ( new_AGEMA_signal_15781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4287 ( .C ( clk ), .D ( n2249 ), .Q ( new_AGEMA_signal_15787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4293 ( .C ( clk ), .D ( new_AGEMA_signal_2262 ), .Q ( new_AGEMA_signal_15793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4299 ( .C ( clk ), .D ( new_AGEMA_signal_2263 ), .Q ( new_AGEMA_signal_15799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4305 ( .C ( clk ), .D ( new_AGEMA_signal_2264 ), .Q ( new_AGEMA_signal_15805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4311 ( .C ( clk ), .D ( n2273 ), .Q ( new_AGEMA_signal_15811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4317 ( .C ( clk ), .D ( new_AGEMA_signal_2688 ), .Q ( new_AGEMA_signal_15817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4323 ( .C ( clk ), .D ( new_AGEMA_signal_2689 ), .Q ( new_AGEMA_signal_15823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4329 ( .C ( clk ), .D ( new_AGEMA_signal_2690 ), .Q ( new_AGEMA_signal_15829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4353 ( .C ( clk ), .D ( new_AGEMA_signal_15852 ), .Q ( new_AGEMA_signal_15853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4361 ( .C ( clk ), .D ( new_AGEMA_signal_15860 ), .Q ( new_AGEMA_signal_15861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4369 ( .C ( clk ), .D ( new_AGEMA_signal_15868 ), .Q ( new_AGEMA_signal_15869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4377 ( .C ( clk ), .D ( new_AGEMA_signal_15876 ), .Q ( new_AGEMA_signal_15877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4399 ( .C ( clk ), .D ( n2349 ), .Q ( new_AGEMA_signal_15899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4405 ( .C ( clk ), .D ( new_AGEMA_signal_1836 ), .Q ( new_AGEMA_signal_15905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4411 ( .C ( clk ), .D ( new_AGEMA_signal_1837 ), .Q ( new_AGEMA_signal_15911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4417 ( .C ( clk ), .D ( new_AGEMA_signal_1838 ), .Q ( new_AGEMA_signal_15917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4425 ( .C ( clk ), .D ( new_AGEMA_signal_15924 ), .Q ( new_AGEMA_signal_15925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4433 ( .C ( clk ), .D ( new_AGEMA_signal_15932 ), .Q ( new_AGEMA_signal_15933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4441 ( .C ( clk ), .D ( new_AGEMA_signal_15940 ), .Q ( new_AGEMA_signal_15941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4449 ( .C ( clk ), .D ( new_AGEMA_signal_15948 ), .Q ( new_AGEMA_signal_15949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4463 ( .C ( clk ), .D ( n2396 ), .Q ( new_AGEMA_signal_15963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4469 ( .C ( clk ), .D ( new_AGEMA_signal_1869 ), .Q ( new_AGEMA_signal_15969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4475 ( .C ( clk ), .D ( new_AGEMA_signal_1870 ), .Q ( new_AGEMA_signal_15975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4481 ( .C ( clk ), .D ( new_AGEMA_signal_1871 ), .Q ( new_AGEMA_signal_15981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4503 ( .C ( clk ), .D ( n2439 ), .Q ( new_AGEMA_signal_16003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4509 ( .C ( clk ), .D ( new_AGEMA_signal_2367 ), .Q ( new_AGEMA_signal_16009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4515 ( .C ( clk ), .D ( new_AGEMA_signal_2368 ), .Q ( new_AGEMA_signal_16015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4521 ( .C ( clk ), .D ( new_AGEMA_signal_2369 ), .Q ( new_AGEMA_signal_16021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4527 ( .C ( clk ), .D ( n2470 ), .Q ( new_AGEMA_signal_16027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4533 ( .C ( clk ), .D ( new_AGEMA_signal_1899 ), .Q ( new_AGEMA_signal_16033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4539 ( .C ( clk ), .D ( new_AGEMA_signal_1900 ), .Q ( new_AGEMA_signal_16039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4545 ( .C ( clk ), .D ( new_AGEMA_signal_1901 ), .Q ( new_AGEMA_signal_16045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4553 ( .C ( clk ), .D ( new_AGEMA_signal_16052 ), .Q ( new_AGEMA_signal_16053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4561 ( .C ( clk ), .D ( new_AGEMA_signal_16060 ), .Q ( new_AGEMA_signal_16061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4569 ( .C ( clk ), .D ( new_AGEMA_signal_16068 ), .Q ( new_AGEMA_signal_16069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4577 ( .C ( clk ), .D ( new_AGEMA_signal_16076 ), .Q ( new_AGEMA_signal_16077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4585 ( .C ( clk ), .D ( new_AGEMA_signal_16084 ), .Q ( new_AGEMA_signal_16085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4593 ( .C ( clk ), .D ( new_AGEMA_signal_16092 ), .Q ( new_AGEMA_signal_16093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4601 ( .C ( clk ), .D ( new_AGEMA_signal_16100 ), .Q ( new_AGEMA_signal_16101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4609 ( .C ( clk ), .D ( new_AGEMA_signal_16108 ), .Q ( new_AGEMA_signal_16109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4615 ( .C ( clk ), .D ( n2585 ), .Q ( new_AGEMA_signal_16115 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4621 ( .C ( clk ), .D ( new_AGEMA_signal_2439 ), .Q ( new_AGEMA_signal_16121 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4627 ( .C ( clk ), .D ( new_AGEMA_signal_2440 ), .Q ( new_AGEMA_signal_16127 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4633 ( .C ( clk ), .D ( new_AGEMA_signal_2441 ), .Q ( new_AGEMA_signal_16133 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4639 ( .C ( clk ), .D ( n2607 ), .Q ( new_AGEMA_signal_16139 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4645 ( .C ( clk ), .D ( new_AGEMA_signal_1953 ), .Q ( new_AGEMA_signal_16145 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4651 ( .C ( clk ), .D ( new_AGEMA_signal_1954 ), .Q ( new_AGEMA_signal_16151 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4657 ( .C ( clk ), .D ( new_AGEMA_signal_1955 ), .Q ( new_AGEMA_signal_16157 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4775 ( .C ( clk ), .D ( n2013 ), .Q ( new_AGEMA_signal_16275 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4783 ( .C ( clk ), .D ( new_AGEMA_signal_2121 ), .Q ( new_AGEMA_signal_16283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4791 ( .C ( clk ), .D ( new_AGEMA_signal_2122 ), .Q ( new_AGEMA_signal_16291 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4799 ( .C ( clk ), .D ( new_AGEMA_signal_2123 ), .Q ( new_AGEMA_signal_16299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4807 ( .C ( clk ), .D ( n2028 ), .Q ( new_AGEMA_signal_16307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4815 ( .C ( clk ), .D ( new_AGEMA_signal_1329 ), .Q ( new_AGEMA_signal_16315 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4823 ( .C ( clk ), .D ( new_AGEMA_signal_1330 ), .Q ( new_AGEMA_signal_16323 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4831 ( .C ( clk ), .D ( new_AGEMA_signal_1331 ), .Q ( new_AGEMA_signal_16331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4839 ( .C ( clk ), .D ( n2051 ), .Q ( new_AGEMA_signal_16339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4847 ( .C ( clk ), .D ( new_AGEMA_signal_2139 ), .Q ( new_AGEMA_signal_16347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4855 ( .C ( clk ), .D ( new_AGEMA_signal_2140 ), .Q ( new_AGEMA_signal_16355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4863 ( .C ( clk ), .D ( new_AGEMA_signal_2141 ), .Q ( new_AGEMA_signal_16363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4871 ( .C ( clk ), .D ( n2069 ), .Q ( new_AGEMA_signal_16371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4879 ( .C ( clk ), .D ( new_AGEMA_signal_2154 ), .Q ( new_AGEMA_signal_16379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4887 ( .C ( clk ), .D ( new_AGEMA_signal_2155 ), .Q ( new_AGEMA_signal_16387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4895 ( .C ( clk ), .D ( new_AGEMA_signal_2156 ), .Q ( new_AGEMA_signal_16395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4929 ( .C ( clk ), .D ( new_AGEMA_signal_16428 ), .Q ( new_AGEMA_signal_16429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4939 ( .C ( clk ), .D ( new_AGEMA_signal_16438 ), .Q ( new_AGEMA_signal_16439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4949 ( .C ( clk ), .D ( new_AGEMA_signal_16448 ), .Q ( new_AGEMA_signal_16449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4959 ( .C ( clk ), .D ( new_AGEMA_signal_16458 ), .Q ( new_AGEMA_signal_16459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4967 ( .C ( clk ), .D ( n2144 ), .Q ( new_AGEMA_signal_16467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4975 ( .C ( clk ), .D ( new_AGEMA_signal_2205 ), .Q ( new_AGEMA_signal_16475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4983 ( .C ( clk ), .D ( new_AGEMA_signal_2206 ), .Q ( new_AGEMA_signal_16483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4991 ( .C ( clk ), .D ( new_AGEMA_signal_2207 ), .Q ( new_AGEMA_signal_16491 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4999 ( .C ( clk ), .D ( n2170 ), .Q ( new_AGEMA_signal_16499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5007 ( .C ( clk ), .D ( new_AGEMA_signal_2211 ), .Q ( new_AGEMA_signal_16507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5015 ( .C ( clk ), .D ( new_AGEMA_signal_2212 ), .Q ( new_AGEMA_signal_16515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5023 ( .C ( clk ), .D ( new_AGEMA_signal_2213 ), .Q ( new_AGEMA_signal_16523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5031 ( .C ( clk ), .D ( n2186 ), .Q ( new_AGEMA_signal_16531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5039 ( .C ( clk ), .D ( new_AGEMA_signal_1368 ), .Q ( new_AGEMA_signal_16539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5047 ( .C ( clk ), .D ( new_AGEMA_signal_1369 ), .Q ( new_AGEMA_signal_16547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5055 ( .C ( clk ), .D ( new_AGEMA_signal_1370 ), .Q ( new_AGEMA_signal_16555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5129 ( .C ( clk ), .D ( new_AGEMA_signal_16628 ), .Q ( new_AGEMA_signal_16629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5139 ( .C ( clk ), .D ( new_AGEMA_signal_16638 ), .Q ( new_AGEMA_signal_16639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5149 ( .C ( clk ), .D ( new_AGEMA_signal_16648 ), .Q ( new_AGEMA_signal_16649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5159 ( .C ( clk ), .D ( new_AGEMA_signal_16658 ), .Q ( new_AGEMA_signal_16659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5167 ( .C ( clk ), .D ( new_AGEMA_signal_13644 ), .Q ( new_AGEMA_signal_16667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5175 ( .C ( clk ), .D ( new_AGEMA_signal_13646 ), .Q ( new_AGEMA_signal_16675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5183 ( .C ( clk ), .D ( new_AGEMA_signal_13648 ), .Q ( new_AGEMA_signal_16683 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5191 ( .C ( clk ), .D ( new_AGEMA_signal_13650 ), .Q ( new_AGEMA_signal_16691 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5223 ( .C ( clk ), .D ( n2551 ), .Q ( new_AGEMA_signal_16723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5231 ( .C ( clk ), .D ( new_AGEMA_signal_2421 ), .Q ( new_AGEMA_signal_16731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5239 ( .C ( clk ), .D ( new_AGEMA_signal_2422 ), .Q ( new_AGEMA_signal_16739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5247 ( .C ( clk ), .D ( new_AGEMA_signal_2423 ), .Q ( new_AGEMA_signal_16747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5255 ( .C ( clk ), .D ( n2588 ), .Q ( new_AGEMA_signal_16755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5263 ( .C ( clk ), .D ( new_AGEMA_signal_2448 ), .Q ( new_AGEMA_signal_16763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5271 ( .C ( clk ), .D ( new_AGEMA_signal_2449 ), .Q ( new_AGEMA_signal_16771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5279 ( .C ( clk ), .D ( new_AGEMA_signal_2450 ), .Q ( new_AGEMA_signal_16779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5327 ( .C ( clk ), .D ( n2701 ), .Q ( new_AGEMA_signal_16827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5335 ( .C ( clk ), .D ( new_AGEMA_signal_1995 ), .Q ( new_AGEMA_signal_16835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5343 ( .C ( clk ), .D ( new_AGEMA_signal_1996 ), .Q ( new_AGEMA_signal_16843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5351 ( .C ( clk ), .D ( new_AGEMA_signal_1997 ), .Q ( new_AGEMA_signal_16851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5591 ( .C ( clk ), .D ( n2172 ), .Q ( new_AGEMA_signal_17091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5601 ( .C ( clk ), .D ( new_AGEMA_signal_2220 ), .Q ( new_AGEMA_signal_17101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5611 ( .C ( clk ), .D ( new_AGEMA_signal_2221 ), .Q ( new_AGEMA_signal_17111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5621 ( .C ( clk ), .D ( new_AGEMA_signal_2222 ), .Q ( new_AGEMA_signal_17121 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6375 ( .C ( clk ), .D ( n2150 ), .Q ( new_AGEMA_signal_17875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6389 ( .C ( clk ), .D ( new_AGEMA_signal_1707 ), .Q ( new_AGEMA_signal_17889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6403 ( .C ( clk ), .D ( new_AGEMA_signal_1708 ), .Q ( new_AGEMA_signal_17903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6417 ( .C ( clk ), .D ( new_AGEMA_signal_1709 ), .Q ( new_AGEMA_signal_17917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6463 ( .C ( clk ), .D ( n2369 ), .Q ( new_AGEMA_signal_17963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6477 ( .C ( clk ), .D ( new_AGEMA_signal_2736 ), .Q ( new_AGEMA_signal_17977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6491 ( .C ( clk ), .D ( new_AGEMA_signal_2737 ), .Q ( new_AGEMA_signal_17991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6505 ( .C ( clk ), .D ( new_AGEMA_signal_2738 ), .Q ( new_AGEMA_signal_18005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6607 ( .C ( clk ), .D ( n2152 ), .Q ( new_AGEMA_signal_18107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6623 ( .C ( clk ), .D ( new_AGEMA_signal_2208 ), .Q ( new_AGEMA_signal_18123 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6639 ( .C ( clk ), .D ( new_AGEMA_signal_2209 ), .Q ( new_AGEMA_signal_18139 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6655 ( .C ( clk ), .D ( new_AGEMA_signal_2210 ), .Q ( new_AGEMA_signal_18155 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6695 ( .C ( clk ), .D ( n2372 ), .Q ( new_AGEMA_signal_18195 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6711 ( .C ( clk ), .D ( new_AGEMA_signal_2328 ), .Q ( new_AGEMA_signal_18211 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6727 ( .C ( clk ), .D ( new_AGEMA_signal_2329 ), .Q ( new_AGEMA_signal_18227 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6743 ( .C ( clk ), .D ( new_AGEMA_signal_2330 ), .Q ( new_AGEMA_signal_18243 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6999 ( .C ( clk ), .D ( n2375 ), .Q ( new_AGEMA_signal_18499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7017 ( .C ( clk ), .D ( new_AGEMA_signal_1839 ), .Q ( new_AGEMA_signal_18517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7035 ( .C ( clk ), .D ( new_AGEMA_signal_1840 ), .Q ( new_AGEMA_signal_18535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7053 ( .C ( clk ), .D ( new_AGEMA_signal_1841 ), .Q ( new_AGEMA_signal_18553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7199 ( .C ( clk ), .D ( n2377 ), .Q ( new_AGEMA_signal_18699 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7219 ( .C ( clk ), .D ( new_AGEMA_signal_2331 ), .Q ( new_AGEMA_signal_18719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7239 ( .C ( clk ), .D ( new_AGEMA_signal_2332 ), .Q ( new_AGEMA_signal_18739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7259 ( .C ( clk ), .D ( new_AGEMA_signal_2333 ), .Q ( new_AGEMA_signal_18759 ) ) ;

    /* cells in depth 8 */
    nor_HPC1 #(.security_order(3), .pipeline(1)) U1968 ( .ina ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, new_AGEMA_signal_2043, n1924}), .inb ({new_AGEMA_signal_2048, new_AGEMA_signal_2047, new_AGEMA_signal_2046, n1923}), .clk ( clk ), .rnd ({Fresh[4519], Fresh[4518], Fresh[4517], Fresh[4516], Fresh[4515], Fresh[4514], Fresh[4513], Fresh[4512], Fresh[4511], Fresh[4510]}), .outt ({new_AGEMA_signal_2528, new_AGEMA_signal_2527, new_AGEMA_signal_2526, n1936}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U1982 ( .ina ({new_AGEMA_signal_13098, new_AGEMA_signal_13096, new_AGEMA_signal_13094, new_AGEMA_signal_13092}), .inb ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, new_AGEMA_signal_2049, n1927}), .clk ( clk ), .rnd ({Fresh[4529], Fresh[4528], Fresh[4527], Fresh[4526], Fresh[4525], Fresh[4524], Fresh[4523], Fresh[4522], Fresh[4521], Fresh[4520]}), .outt ({new_AGEMA_signal_2531, new_AGEMA_signal_2530, new_AGEMA_signal_2529, n1928}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U1994 ( .ina ({new_AGEMA_signal_13106, new_AGEMA_signal_13104, new_AGEMA_signal_13102, new_AGEMA_signal_13100}), .inb ({new_AGEMA_signal_2054, new_AGEMA_signal_2053, new_AGEMA_signal_2052, n1929}), .clk ( clk ), .rnd ({Fresh[4539], Fresh[4538], Fresh[4537], Fresh[4536], Fresh[4535], Fresh[4534], Fresh[4533], Fresh[4532], Fresh[4531], Fresh[4530]}), .outt ({new_AGEMA_signal_2534, new_AGEMA_signal_2533, new_AGEMA_signal_2532, n1931}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2012 ( .ina ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, new_AGEMA_signal_2055, n2665}), .inb ({new_AGEMA_signal_2060, new_AGEMA_signal_2059, new_AGEMA_signal_2058, n1938}), .clk ( clk ), .rnd ({Fresh[4549], Fresh[4548], Fresh[4547], Fresh[4546], Fresh[4545], Fresh[4544], Fresh[4543], Fresh[4542], Fresh[4541], Fresh[4540]}), .outt ({new_AGEMA_signal_2537, new_AGEMA_signal_2536, new_AGEMA_signal_2535, n1939}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2024 ( .ina ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, new_AGEMA_signal_2061, n2235}), .inb ({new_AGEMA_signal_1529, new_AGEMA_signal_1528, new_AGEMA_signal_1527, n1943}), .clk ( clk ), .rnd ({Fresh[4559], Fresh[4558], Fresh[4557], Fresh[4556], Fresh[4555], Fresh[4554], Fresh[4553], Fresh[4552], Fresh[4551], Fresh[4550]}), .outt ({new_AGEMA_signal_2540, new_AGEMA_signal_2539, new_AGEMA_signal_2538, n1948}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2032 ( .ina ({new_AGEMA_signal_1532, new_AGEMA_signal_1531, new_AGEMA_signal_1530, n1946}), .inb ({new_AGEMA_signal_2066, new_AGEMA_signal_2065, new_AGEMA_signal_2064, n1945}), .clk ( clk ), .rnd ({Fresh[4569], Fresh[4568], Fresh[4567], Fresh[4566], Fresh[4565], Fresh[4564], Fresh[4563], Fresh[4562], Fresh[4561], Fresh[4560]}), .outt ({new_AGEMA_signal_2543, new_AGEMA_signal_2542, new_AGEMA_signal_2541, n1947}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2041 ( .ina ({new_AGEMA_signal_13122, new_AGEMA_signal_13118, new_AGEMA_signal_13114, new_AGEMA_signal_13110}), .inb ({new_AGEMA_signal_2072, new_AGEMA_signal_2071, new_AGEMA_signal_2070, n1951}), .clk ( clk ), .rnd ({Fresh[4579], Fresh[4578], Fresh[4577], Fresh[4576], Fresh[4575], Fresh[4574], Fresh[4573], Fresh[4572], Fresh[4571], Fresh[4570]}), .outt ({new_AGEMA_signal_2546, new_AGEMA_signal_2545, new_AGEMA_signal_2544, n1954}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2049 ( .ina ({new_AGEMA_signal_13130, new_AGEMA_signal_13128, new_AGEMA_signal_13126, new_AGEMA_signal_13124}), .inb ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, new_AGEMA_signal_2073, n1952}), .clk ( clk ), .rnd ({Fresh[4589], Fresh[4588], Fresh[4587], Fresh[4586], Fresh[4585], Fresh[4584], Fresh[4583], Fresh[4582], Fresh[4581], Fresh[4580]}), .outt ({new_AGEMA_signal_2549, new_AGEMA_signal_2548, new_AGEMA_signal_2547, n1953}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2058 ( .ina ({new_AGEMA_signal_13138, new_AGEMA_signal_13136, new_AGEMA_signal_13134, new_AGEMA_signal_13132}), .inb ({new_AGEMA_signal_2078, new_AGEMA_signal_2077, new_AGEMA_signal_2076, n2687}), .clk ( clk ), .rnd ({Fresh[4599], Fresh[4598], Fresh[4597], Fresh[4596], Fresh[4595], Fresh[4594], Fresh[4593], Fresh[4592], Fresh[4591], Fresh[4590]}), .outt ({new_AGEMA_signal_2552, new_AGEMA_signal_2551, new_AGEMA_signal_2550, n2658}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2065 ( .ina ({new_AGEMA_signal_13146, new_AGEMA_signal_13144, new_AGEMA_signal_13142, new_AGEMA_signal_13140}), .inb ({new_AGEMA_signal_1547, new_AGEMA_signal_1546, new_AGEMA_signal_1545, n1963}), .clk ( clk ), .rnd ({Fresh[4609], Fresh[4608], Fresh[4607], Fresh[4606], Fresh[4605], Fresh[4604], Fresh[4603], Fresh[4602], Fresh[4601], Fresh[4600]}), .outt ({new_AGEMA_signal_2084, new_AGEMA_signal_2083, new_AGEMA_signal_2082, n1965}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2078 ( .ina ({new_AGEMA_signal_13154, new_AGEMA_signal_13152, new_AGEMA_signal_13150, new_AGEMA_signal_13148}), .inb ({new_AGEMA_signal_2558, new_AGEMA_signal_2557, new_AGEMA_signal_2556, n1968}), .clk ( clk ), .rnd ({Fresh[4619], Fresh[4618], Fresh[4617], Fresh[4616], Fresh[4615], Fresh[4614], Fresh[4613], Fresh[4612], Fresh[4611], Fresh[4610]}), .outt ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, new_AGEMA_signal_2889, n1970}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2084 ( .ina ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, new_AGEMA_signal_2091, n2684}), .inb ({new_AGEMA_signal_13162, new_AGEMA_signal_13160, new_AGEMA_signal_13158, new_AGEMA_signal_13156}), .clk ( clk ), .rnd ({Fresh[4629], Fresh[4628], Fresh[4627], Fresh[4626], Fresh[4625], Fresh[4624], Fresh[4623], Fresh[4622], Fresh[4621], Fresh[4620]}), .outt ({new_AGEMA_signal_2561, new_AGEMA_signal_2560, new_AGEMA_signal_2559, n1969}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2093 ( .ina ({new_AGEMA_signal_2096, new_AGEMA_signal_2095, new_AGEMA_signal_2094, n1972}), .inb ({new_AGEMA_signal_1565, new_AGEMA_signal_1564, new_AGEMA_signal_1563, n1971}), .clk ( clk ), .rnd ({Fresh[4639], Fresh[4638], Fresh[4637], Fresh[4636], Fresh[4635], Fresh[4634], Fresh[4633], Fresh[4632], Fresh[4631], Fresh[4630]}), .outt ({new_AGEMA_signal_2564, new_AGEMA_signal_2563, new_AGEMA_signal_2562, n1978}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2102 ( .ina ({new_AGEMA_signal_2099, new_AGEMA_signal_2098, new_AGEMA_signal_2097, n1974}), .inb ({new_AGEMA_signal_13170, new_AGEMA_signal_13168, new_AGEMA_signal_13166, new_AGEMA_signal_13164}), .clk ( clk ), .rnd ({Fresh[4649], Fresh[4648], Fresh[4647], Fresh[4646], Fresh[4645], Fresh[4644], Fresh[4643], Fresh[4642], Fresh[4641], Fresh[4640]}), .outt ({new_AGEMA_signal_2567, new_AGEMA_signal_2566, new_AGEMA_signal_2565, n1975}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2107 ( .ina ({new_AGEMA_signal_13178, new_AGEMA_signal_13176, new_AGEMA_signal_13174, new_AGEMA_signal_13172}), .inb ({new_AGEMA_signal_2102, new_AGEMA_signal_2101, new_AGEMA_signal_2100, n1979}), .clk ( clk ), .rnd ({Fresh[4659], Fresh[4658], Fresh[4657], Fresh[4656], Fresh[4655], Fresh[4654], Fresh[4653], Fresh[4652], Fresh[4651], Fresh[4650]}), .outt ({new_AGEMA_signal_2570, new_AGEMA_signal_2569, new_AGEMA_signal_2568, n1980}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2114 ( .ina ({new_AGEMA_signal_1574, new_AGEMA_signal_1573, new_AGEMA_signal_1572, n1985}), .inb ({new_AGEMA_signal_13186, new_AGEMA_signal_13184, new_AGEMA_signal_13182, new_AGEMA_signal_13180}), .clk ( clk ), .rnd ({Fresh[4669], Fresh[4668], Fresh[4667], Fresh[4666], Fresh[4665], Fresh[4664], Fresh[4663], Fresh[4662], Fresh[4661], Fresh[4660]}), .outt ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, new_AGEMA_signal_2103, n1986}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2124 ( .ina ({new_AGEMA_signal_2108, new_AGEMA_signal_2107, new_AGEMA_signal_2106, n1994}), .inb ({new_AGEMA_signal_13194, new_AGEMA_signal_13192, new_AGEMA_signal_13190, new_AGEMA_signal_13188}), .clk ( clk ), .rnd ({Fresh[4679], Fresh[4678], Fresh[4677], Fresh[4676], Fresh[4675], Fresh[4674], Fresh[4673], Fresh[4672], Fresh[4671], Fresh[4670]}), .outt ({new_AGEMA_signal_2576, new_AGEMA_signal_2575, new_AGEMA_signal_2574, n1997}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2137 ( .ina ({new_AGEMA_signal_13202, new_AGEMA_signal_13200, new_AGEMA_signal_13198, new_AGEMA_signal_13196}), .inb ({new_AGEMA_signal_2114, new_AGEMA_signal_2113, new_AGEMA_signal_2112, n2137}), .clk ( clk ), .rnd ({Fresh[4689], Fresh[4688], Fresh[4687], Fresh[4686], Fresh[4685], Fresh[4684], Fresh[4683], Fresh[4682], Fresh[4681], Fresh[4680]}), .outt ({new_AGEMA_signal_2579, new_AGEMA_signal_2578, new_AGEMA_signal_2577, n2012}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2145 ( .ina ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, new_AGEMA_signal_2115, n2006}), .inb ({new_AGEMA_signal_2120, new_AGEMA_signal_2119, new_AGEMA_signal_2118, n2005}), .clk ( clk ), .rnd ({Fresh[4699], Fresh[4698], Fresh[4697], Fresh[4696], Fresh[4695], Fresh[4694], Fresh[4693], Fresh[4692], Fresh[4691], Fresh[4690]}), .outt ({new_AGEMA_signal_2582, new_AGEMA_signal_2581, new_AGEMA_signal_2580, n2007}) ) ;
    mux2_HPC1 #(.security_order(3), .pipeline(1)) U2161 ( .ins ({new_AGEMA_signal_13210, new_AGEMA_signal_13208, new_AGEMA_signal_13206, new_AGEMA_signal_13204}), .inb ({new_AGEMA_signal_1613, new_AGEMA_signal_1612, new_AGEMA_signal_1611, n2020}), .ina ({new_AGEMA_signal_13226, new_AGEMA_signal_13222, new_AGEMA_signal_13218, new_AGEMA_signal_13214}), .clk ( clk ), .rnd ({Fresh[4709], Fresh[4708], Fresh[4707], Fresh[4706], Fresh[4705], Fresh[4704], Fresh[4703], Fresh[4702], Fresh[4701], Fresh[4700]}), .outt ({new_AGEMA_signal_2126, new_AGEMA_signal_2125, new_AGEMA_signal_2124, n2021}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2176 ( .ina ({new_AGEMA_signal_13234, new_AGEMA_signal_13232, new_AGEMA_signal_13230, new_AGEMA_signal_13228}), .inb ({new_AGEMA_signal_2132, new_AGEMA_signal_2131, new_AGEMA_signal_2130, n2031}), .clk ( clk ), .rnd ({Fresh[4719], Fresh[4718], Fresh[4717], Fresh[4716], Fresh[4715], Fresh[4714], Fresh[4713], Fresh[4712], Fresh[4711], Fresh[4710]}), .outt ({new_AGEMA_signal_2588, new_AGEMA_signal_2587, new_AGEMA_signal_2586, n2032}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2185 ( .ina ({new_AGEMA_signal_13242, new_AGEMA_signal_13240, new_AGEMA_signal_13238, new_AGEMA_signal_13236}), .inb ({new_AGEMA_signal_2135, new_AGEMA_signal_2134, new_AGEMA_signal_2133, n2040}), .clk ( clk ), .rnd ({Fresh[4729], Fresh[4728], Fresh[4727], Fresh[4726], Fresh[4725], Fresh[4724], Fresh[4723], Fresh[4722], Fresh[4721], Fresh[4720]}), .outt ({new_AGEMA_signal_2591, new_AGEMA_signal_2590, new_AGEMA_signal_2589, n2041}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2189 ( .ina ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, new_AGEMA_signal_2055, n2665}), .inb ({new_AGEMA_signal_13250, new_AGEMA_signal_13248, new_AGEMA_signal_13246, new_AGEMA_signal_13244}), .clk ( clk ), .rnd ({Fresh[4739], Fresh[4738], Fresh[4737], Fresh[4736], Fresh[4735], Fresh[4734], Fresh[4733], Fresh[4732], Fresh[4731], Fresh[4730]}), .outt ({new_AGEMA_signal_2594, new_AGEMA_signal_2593, new_AGEMA_signal_2592, n2043}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2194 ( .ina ({new_AGEMA_signal_13258, new_AGEMA_signal_13256, new_AGEMA_signal_13254, new_AGEMA_signal_13252}), .inb ({new_AGEMA_signal_2138, new_AGEMA_signal_2137, new_AGEMA_signal_2136, n2045}), .clk ( clk ), .rnd ({Fresh[4749], Fresh[4748], Fresh[4747], Fresh[4746], Fresh[4745], Fresh[4744], Fresh[4743], Fresh[4742], Fresh[4741], Fresh[4740]}), .outt ({new_AGEMA_signal_2597, new_AGEMA_signal_2596, new_AGEMA_signal_2595, n2046}) ) ;
    mux2_HPC1 #(.security_order(3), .pipeline(1)) U2204 ( .ins ({new_AGEMA_signal_13210, new_AGEMA_signal_13208, new_AGEMA_signal_13206, new_AGEMA_signal_13204}), .inb ({new_AGEMA_signal_2144, new_AGEMA_signal_2143, new_AGEMA_signal_2142, n2056}), .ina ({new_AGEMA_signal_13266, new_AGEMA_signal_13264, new_AGEMA_signal_13262, new_AGEMA_signal_13260}), .clk ( clk ), .rnd ({Fresh[4759], Fresh[4758], Fresh[4757], Fresh[4756], Fresh[4755], Fresh[4754], Fresh[4753], Fresh[4752], Fresh[4751], Fresh[4750]}), .outt ({new_AGEMA_signal_2600, new_AGEMA_signal_2599, new_AGEMA_signal_2598, n2058}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2210 ( .ina ({new_AGEMA_signal_13274, new_AGEMA_signal_13272, new_AGEMA_signal_13270, new_AGEMA_signal_13268}), .inb ({new_AGEMA_signal_2147, new_AGEMA_signal_2146, new_AGEMA_signal_2145, n2060}), .clk ( clk ), .rnd ({Fresh[4769], Fresh[4768], Fresh[4767], Fresh[4766], Fresh[4765], Fresh[4764], Fresh[4763], Fresh[4762], Fresh[4761], Fresh[4760]}), .outt ({new_AGEMA_signal_2603, new_AGEMA_signal_2602, new_AGEMA_signal_2601, n2063}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2218 ( .ina ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, new_AGEMA_signal_2148, n2066}), .inb ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, new_AGEMA_signal_2151, n2065}), .clk ( clk ), .rnd ({Fresh[4779], Fresh[4778], Fresh[4777], Fresh[4776], Fresh[4775], Fresh[4774], Fresh[4773], Fresh[4772], Fresh[4771], Fresh[4770]}), .outt ({new_AGEMA_signal_2606, new_AGEMA_signal_2605, new_AGEMA_signal_2604, n2652}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2227 ( .ina ({new_AGEMA_signal_13282, new_AGEMA_signal_13280, new_AGEMA_signal_13278, new_AGEMA_signal_13276}), .inb ({new_AGEMA_signal_2159, new_AGEMA_signal_2158, new_AGEMA_signal_2157, n2074}), .clk ( clk ), .rnd ({Fresh[4789], Fresh[4788], Fresh[4787], Fresh[4786], Fresh[4785], Fresh[4784], Fresh[4783], Fresh[4782], Fresh[4781], Fresh[4780]}), .outt ({new_AGEMA_signal_2609, new_AGEMA_signal_2608, new_AGEMA_signal_2607, n2076}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2236 ( .ina ({new_AGEMA_signal_13298, new_AGEMA_signal_13294, new_AGEMA_signal_13290, new_AGEMA_signal_13286}), .inb ({new_AGEMA_signal_2162, new_AGEMA_signal_2161, new_AGEMA_signal_2160, n2082}), .clk ( clk ), .rnd ({Fresh[4799], Fresh[4798], Fresh[4797], Fresh[4796], Fresh[4795], Fresh[4794], Fresh[4793], Fresh[4792], Fresh[4791], Fresh[4790]}), .outt ({new_AGEMA_signal_2612, new_AGEMA_signal_2611, new_AGEMA_signal_2610, n2105}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2241 ( .ina ({new_AGEMA_signal_13306, new_AGEMA_signal_13304, new_AGEMA_signal_13302, new_AGEMA_signal_13300}), .inb ({new_AGEMA_signal_2165, new_AGEMA_signal_2164, new_AGEMA_signal_2163, n2084}), .clk ( clk ), .rnd ({Fresh[4809], Fresh[4808], Fresh[4807], Fresh[4806], Fresh[4805], Fresh[4804], Fresh[4803], Fresh[4802], Fresh[4801], Fresh[4800]}), .outt ({new_AGEMA_signal_2615, new_AGEMA_signal_2614, new_AGEMA_signal_2613, n2099}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2243 ( .ina ({new_AGEMA_signal_2168, new_AGEMA_signal_2167, new_AGEMA_signal_2166, n2085}), .inb ({new_AGEMA_signal_13314, new_AGEMA_signal_13312, new_AGEMA_signal_13310, new_AGEMA_signal_13308}), .clk ( clk ), .rnd ({Fresh[4819], Fresh[4818], Fresh[4817], Fresh[4816], Fresh[4815], Fresh[4814], Fresh[4813], Fresh[4812], Fresh[4811], Fresh[4810]}), .outt ({new_AGEMA_signal_2618, new_AGEMA_signal_2617, new_AGEMA_signal_2616, n2091}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(1)) U2246 ( .ina ({new_AGEMA_signal_13322, new_AGEMA_signal_13320, new_AGEMA_signal_13318, new_AGEMA_signal_13316}), .inb ({new_AGEMA_signal_2171, new_AGEMA_signal_2170, new_AGEMA_signal_2169, n2131}), .clk ( clk ), .rnd ({Fresh[4829], Fresh[4828], Fresh[4827], Fresh[4826], Fresh[4825], Fresh[4824], Fresh[4823], Fresh[4822], Fresh[4821], Fresh[4820]}), .outt ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, new_AGEMA_signal_2619, n2090}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2253 ( .ina ({new_AGEMA_signal_13330, new_AGEMA_signal_13328, new_AGEMA_signal_13326, new_AGEMA_signal_13324}), .inb ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, new_AGEMA_signal_2175, n2330}), .clk ( clk ), .rnd ({Fresh[4839], Fresh[4838], Fresh[4837], Fresh[4836], Fresh[4835], Fresh[4834], Fresh[4833], Fresh[4832], Fresh[4831], Fresh[4830]}), .outt ({new_AGEMA_signal_2624, new_AGEMA_signal_2623, new_AGEMA_signal_2622, n2093}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2262 ( .ina ({new_AGEMA_signal_13338, new_AGEMA_signal_13336, new_AGEMA_signal_13334, new_AGEMA_signal_13332}), .inb ({new_AGEMA_signal_2186, new_AGEMA_signal_2185, new_AGEMA_signal_2184, n2160}), .clk ( clk ), .rnd ({Fresh[4849], Fresh[4848], Fresh[4847], Fresh[4846], Fresh[4845], Fresh[4844], Fresh[4843], Fresh[4842], Fresh[4841], Fresh[4840]}), .outt ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, new_AGEMA_signal_2625, n2102}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2266 ( .ina ({new_AGEMA_signal_1685, new_AGEMA_signal_1684, new_AGEMA_signal_1683, n2504}), .inb ({new_AGEMA_signal_13354, new_AGEMA_signal_13350, new_AGEMA_signal_13346, new_AGEMA_signal_13342}), .clk ( clk ), .rnd ({Fresh[4859], Fresh[4858], Fresh[4857], Fresh[4856], Fresh[4855], Fresh[4854], Fresh[4853], Fresh[4852], Fresh[4851], Fresh[4850]}), .outt ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, new_AGEMA_signal_2187, n2106}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2272 ( .ina ({new_AGEMA_signal_13362, new_AGEMA_signal_13360, new_AGEMA_signal_13358, new_AGEMA_signal_13356}), .inb ({new_AGEMA_signal_2630, new_AGEMA_signal_2629, new_AGEMA_signal_2628, n2114}), .clk ( clk ), .rnd ({Fresh[4869], Fresh[4868], Fresh[4867], Fresh[4866], Fresh[4865], Fresh[4864], Fresh[4863], Fresh[4862], Fresh[4861], Fresh[4860]}), .outt ({new_AGEMA_signal_2936, new_AGEMA_signal_2935, new_AGEMA_signal_2934, n2116}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2282 ( .ina ({new_AGEMA_signal_2192, new_AGEMA_signal_2191, new_AGEMA_signal_2190, n2291}), .inb ({new_AGEMA_signal_1694, new_AGEMA_signal_1693, new_AGEMA_signal_1692, n2119}), .clk ( clk ), .rnd ({Fresh[4879], Fresh[4878], Fresh[4877], Fresh[4876], Fresh[4875], Fresh[4874], Fresh[4873], Fresh[4872], Fresh[4871], Fresh[4870]}), .outt ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, new_AGEMA_signal_2631, n2120}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2293 ( .ina ({new_AGEMA_signal_1703, new_AGEMA_signal_1702, new_AGEMA_signal_1701, n2130}), .inb ({new_AGEMA_signal_1706, new_AGEMA_signal_1705, new_AGEMA_signal_1704, n2129}), .clk ( clk ), .rnd ({Fresh[4889], Fresh[4888], Fresh[4887], Fresh[4886], Fresh[4885], Fresh[4884], Fresh[4883], Fresh[4882], Fresh[4881], Fresh[4880]}), .outt ({new_AGEMA_signal_2195, new_AGEMA_signal_2194, new_AGEMA_signal_2193, n2155}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2296 ( .ina ({new_AGEMA_signal_13370, new_AGEMA_signal_13368, new_AGEMA_signal_13366, new_AGEMA_signal_13364}), .inb ({new_AGEMA_signal_2171, new_AGEMA_signal_2170, new_AGEMA_signal_2169, n2131}), .clk ( clk ), .rnd ({Fresh[4899], Fresh[4898], Fresh[4897], Fresh[4896], Fresh[4895], Fresh[4894], Fresh[4893], Fresh[4892], Fresh[4891], Fresh[4890]}), .outt ({new_AGEMA_signal_2636, new_AGEMA_signal_2635, new_AGEMA_signal_2634, n2543}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2299 ( .ina ({new_AGEMA_signal_1712, new_AGEMA_signal_1711, new_AGEMA_signal_1710, n2133}), .inb ({new_AGEMA_signal_13378, new_AGEMA_signal_13376, new_AGEMA_signal_13374, new_AGEMA_signal_13372}), .clk ( clk ), .rnd ({Fresh[4909], Fresh[4908], Fresh[4907], Fresh[4906], Fresh[4905], Fresh[4904], Fresh[4903], Fresh[4902], Fresh[4901], Fresh[4900]}), .outt ({new_AGEMA_signal_2198, new_AGEMA_signal_2197, new_AGEMA_signal_2196, n2134}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2303 ( .ina ({new_AGEMA_signal_2114, new_AGEMA_signal_2113, new_AGEMA_signal_2112, n2137}), .inb ({new_AGEMA_signal_2201, new_AGEMA_signal_2200, new_AGEMA_signal_2199, n2136}), .clk ( clk ), .rnd ({Fresh[4919], Fresh[4918], Fresh[4917], Fresh[4916], Fresh[4915], Fresh[4914], Fresh[4913], Fresh[4912], Fresh[4911], Fresh[4910]}), .outt ({new_AGEMA_signal_2642, new_AGEMA_signal_2641, new_AGEMA_signal_2640, n2143}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2308 ( .ina ({new_AGEMA_signal_2204, new_AGEMA_signal_2203, new_AGEMA_signal_2202, n2139}), .inb ({new_AGEMA_signal_13394, new_AGEMA_signal_13390, new_AGEMA_signal_13386, new_AGEMA_signal_13382}), .clk ( clk ), .rnd ({Fresh[4929], Fresh[4928], Fresh[4927], Fresh[4926], Fresh[4925], Fresh[4924], Fresh[4923], Fresh[4922], Fresh[4921], Fresh[4920]}), .outt ({new_AGEMA_signal_2645, new_AGEMA_signal_2644, new_AGEMA_signal_2643, n2140}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2324 ( .ina ({new_AGEMA_signal_2216, new_AGEMA_signal_2215, new_AGEMA_signal_2214, n2157}), .inb ({new_AGEMA_signal_13402, new_AGEMA_signal_13400, new_AGEMA_signal_13398, new_AGEMA_signal_13396}), .clk ( clk ), .rnd ({Fresh[4939], Fresh[4938], Fresh[4937], Fresh[4936], Fresh[4935], Fresh[4934], Fresh[4933], Fresh[4932], Fresh[4931], Fresh[4930]}), .outt ({new_AGEMA_signal_2648, new_AGEMA_signal_2647, new_AGEMA_signal_2646, n2159}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2326 ( .ina ({new_AGEMA_signal_2186, new_AGEMA_signal_2185, new_AGEMA_signal_2184, n2160}), .inb ({new_AGEMA_signal_13410, new_AGEMA_signal_13408, new_AGEMA_signal_13406, new_AGEMA_signal_13404}), .clk ( clk ), .rnd ({Fresh[4949], Fresh[4948], Fresh[4947], Fresh[4946], Fresh[4945], Fresh[4944], Fresh[4943], Fresh[4942], Fresh[4941], Fresh[4940]}), .outt ({new_AGEMA_signal_2651, new_AGEMA_signal_2650, new_AGEMA_signal_2649, n2161}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2330 ( .ina ({new_AGEMA_signal_13122, new_AGEMA_signal_13118, new_AGEMA_signal_13114, new_AGEMA_signal_13110}), .inb ({new_AGEMA_signal_1727, new_AGEMA_signal_1726, new_AGEMA_signal_1725, n2163}), .clk ( clk ), .rnd ({Fresh[4959], Fresh[4958], Fresh[4957], Fresh[4956], Fresh[4955], Fresh[4954], Fresh[4953], Fresh[4952], Fresh[4951], Fresh[4950]}), .outt ({new_AGEMA_signal_2219, new_AGEMA_signal_2218, new_AGEMA_signal_2217, n2164}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2345 ( .ina ({new_AGEMA_signal_13418, new_AGEMA_signal_13416, new_AGEMA_signal_13414, new_AGEMA_signal_13412}), .inb ({new_AGEMA_signal_2228, new_AGEMA_signal_2227, new_AGEMA_signal_2226, n2177}), .clk ( clk ), .rnd ({Fresh[4969], Fresh[4968], Fresh[4967], Fresh[4966], Fresh[4965], Fresh[4964], Fresh[4963], Fresh[4962], Fresh[4961], Fresh[4960]}), .outt ({new_AGEMA_signal_2657, new_AGEMA_signal_2656, new_AGEMA_signal_2655, n2179}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2359 ( .ina ({new_AGEMA_signal_13434, new_AGEMA_signal_13430, new_AGEMA_signal_13426, new_AGEMA_signal_13422}), .inb ({new_AGEMA_signal_2237, new_AGEMA_signal_2236, new_AGEMA_signal_2235, n2191}), .clk ( clk ), .rnd ({Fresh[4979], Fresh[4978], Fresh[4977], Fresh[4976], Fresh[4975], Fresh[4974], Fresh[4973], Fresh[4972], Fresh[4971], Fresh[4970]}), .outt ({new_AGEMA_signal_2660, new_AGEMA_signal_2659, new_AGEMA_signal_2658, n2192}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2370 ( .ina ({new_AGEMA_signal_2240, new_AGEMA_signal_2239, new_AGEMA_signal_2238, n2201}), .inb ({new_AGEMA_signal_2663, new_AGEMA_signal_2662, new_AGEMA_signal_2661, n2200}), .clk ( clk ), .rnd ({Fresh[4989], Fresh[4988], Fresh[4987], Fresh[4986], Fresh[4985], Fresh[4984], Fresh[4983], Fresh[4982], Fresh[4981], Fresh[4980]}), .outt ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, new_AGEMA_signal_2955, n2203}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2382 ( .ina ({new_AGEMA_signal_2246, new_AGEMA_signal_2245, new_AGEMA_signal_2244, n2217}), .inb ({new_AGEMA_signal_1748, new_AGEMA_signal_1747, new_AGEMA_signal_1746, n2216}), .clk ( clk ), .rnd ({Fresh[4999], Fresh[4998], Fresh[4997], Fresh[4996], Fresh[4995], Fresh[4994], Fresh[4993], Fresh[4992], Fresh[4991], Fresh[4990]}), .outt ({new_AGEMA_signal_2669, new_AGEMA_signal_2668, new_AGEMA_signal_2667, n2224}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2388 ( .ina ({new_AGEMA_signal_2249, new_AGEMA_signal_2248, new_AGEMA_signal_2247, n2222}), .inb ({new_AGEMA_signal_2252, new_AGEMA_signal_2251, new_AGEMA_signal_2250, n2221}), .clk ( clk ), .rnd ({Fresh[5009], Fresh[5008], Fresh[5007], Fresh[5006], Fresh[5005], Fresh[5004], Fresh[5003], Fresh[5002], Fresh[5001], Fresh[5000]}), .outt ({new_AGEMA_signal_2672, new_AGEMA_signal_2671, new_AGEMA_signal_2670, n2223}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2392 ( .ina ({new_AGEMA_signal_1685, new_AGEMA_signal_1684, new_AGEMA_signal_1683, n2504}), .inb ({new_AGEMA_signal_1757, new_AGEMA_signal_1756, new_AGEMA_signal_1755, n2226}), .clk ( clk ), .rnd ({Fresh[5019], Fresh[5018], Fresh[5017], Fresh[5016], Fresh[5015], Fresh[5014], Fresh[5013], Fresh[5012], Fresh[5011], Fresh[5010]}), .outt ({new_AGEMA_signal_2255, new_AGEMA_signal_2254, new_AGEMA_signal_2253, n2229}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2399 ( .ina ({new_AGEMA_signal_13130, new_AGEMA_signal_13128, new_AGEMA_signal_13126, new_AGEMA_signal_13124}), .inb ({new_AGEMA_signal_2678, new_AGEMA_signal_2677, new_AGEMA_signal_2676, n2233}), .clk ( clk ), .rnd ({Fresh[5029], Fresh[5028], Fresh[5027], Fresh[5026], Fresh[5025], Fresh[5024], Fresh[5023], Fresh[5022], Fresh[5021], Fresh[5020]}), .outt ({new_AGEMA_signal_2966, new_AGEMA_signal_2965, new_AGEMA_signal_2964, n2234}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2410 ( .ina ({new_AGEMA_signal_13138, new_AGEMA_signal_13136, new_AGEMA_signal_13134, new_AGEMA_signal_13132}), .inb ({new_AGEMA_signal_2261, new_AGEMA_signal_2260, new_AGEMA_signal_2259, n2244}), .clk ( clk ), .rnd ({Fresh[5039], Fresh[5038], Fresh[5037], Fresh[5036], Fresh[5035], Fresh[5034], Fresh[5033], Fresh[5032], Fresh[5031], Fresh[5030]}), .outt ({new_AGEMA_signal_2681, new_AGEMA_signal_2680, new_AGEMA_signal_2679, n2246}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2418 ( .ina ({new_AGEMA_signal_13442, new_AGEMA_signal_13440, new_AGEMA_signal_13438, new_AGEMA_signal_13436}), .inb ({new_AGEMA_signal_2267, new_AGEMA_signal_2266, new_AGEMA_signal_2265, n2253}), .clk ( clk ), .rnd ({Fresh[5049], Fresh[5048], Fresh[5047], Fresh[5046], Fresh[5045], Fresh[5044], Fresh[5043], Fresh[5042], Fresh[5041], Fresh[5040]}), .outt ({new_AGEMA_signal_2684, new_AGEMA_signal_2683, new_AGEMA_signal_2682, n2254}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2425 ( .ina ({new_AGEMA_signal_13450, new_AGEMA_signal_13448, new_AGEMA_signal_13446, new_AGEMA_signal_13444}), .inb ({new_AGEMA_signal_2270, new_AGEMA_signal_2269, new_AGEMA_signal_2268, n2260}), .clk ( clk ), .rnd ({Fresh[5059], Fresh[5058], Fresh[5057], Fresh[5056], Fresh[5055], Fresh[5054], Fresh[5053], Fresh[5052], Fresh[5051], Fresh[5050]}), .outt ({new_AGEMA_signal_2687, new_AGEMA_signal_2686, new_AGEMA_signal_2685, n2263}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2434 ( .ina ({new_AGEMA_signal_13458, new_AGEMA_signal_13456, new_AGEMA_signal_13454, new_AGEMA_signal_13452}), .inb ({new_AGEMA_signal_1787, new_AGEMA_signal_1786, new_AGEMA_signal_1785, n2265}), .clk ( clk ), .rnd ({Fresh[5069], Fresh[5068], Fresh[5067], Fresh[5066], Fresh[5065], Fresh[5064], Fresh[5063], Fresh[5062], Fresh[5061], Fresh[5060]}), .outt ({new_AGEMA_signal_2273, new_AGEMA_signal_2272, new_AGEMA_signal_2271, n2267}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2438 ( .ina ({new_AGEMA_signal_13130, new_AGEMA_signal_13128, new_AGEMA_signal_13126, new_AGEMA_signal_13124}), .inb ({new_AGEMA_signal_1790, new_AGEMA_signal_1789, new_AGEMA_signal_1788, n2269}), .clk ( clk ), .rnd ({Fresh[5079], Fresh[5078], Fresh[5077], Fresh[5076], Fresh[5075], Fresh[5074], Fresh[5073], Fresh[5072], Fresh[5071], Fresh[5070]}), .outt ({new_AGEMA_signal_2276, new_AGEMA_signal_2275, new_AGEMA_signal_2274, n2270}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2445 ( .ina ({new_AGEMA_signal_13466, new_AGEMA_signal_13464, new_AGEMA_signal_13462, new_AGEMA_signal_13460}), .inb ({new_AGEMA_signal_1796, new_AGEMA_signal_1795, new_AGEMA_signal_1794, n2277}), .clk ( clk ), .rnd ({Fresh[5089], Fresh[5088], Fresh[5087], Fresh[5086], Fresh[5085], Fresh[5084], Fresh[5083], Fresh[5082], Fresh[5081], Fresh[5080]}), .outt ({new_AGEMA_signal_2279, new_AGEMA_signal_2278, new_AGEMA_signal_2277, n2279}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2450 ( .ina ({new_AGEMA_signal_13226, new_AGEMA_signal_13222, new_AGEMA_signal_13218, new_AGEMA_signal_13214}), .inb ({new_AGEMA_signal_1799, new_AGEMA_signal_1798, new_AGEMA_signal_1797, n2282}), .clk ( clk ), .rnd ({Fresh[5099], Fresh[5098], Fresh[5097], Fresh[5096], Fresh[5095], Fresh[5094], Fresh[5093], Fresh[5092], Fresh[5091], Fresh[5090]}), .outt ({new_AGEMA_signal_2282, new_AGEMA_signal_2281, new_AGEMA_signal_2280, n2283}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2453 ( .ina ({new_AGEMA_signal_13306, new_AGEMA_signal_13304, new_AGEMA_signal_13302, new_AGEMA_signal_13300}), .inb ({new_AGEMA_signal_2285, new_AGEMA_signal_2284, new_AGEMA_signal_2283, n2284}), .clk ( clk ), .rnd ({Fresh[5109], Fresh[5108], Fresh[5107], Fresh[5106], Fresh[5105], Fresh[5104], Fresh[5103], Fresh[5102], Fresh[5101], Fresh[5100]}), .outt ({new_AGEMA_signal_2702, new_AGEMA_signal_2701, new_AGEMA_signal_2700, n2285}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2457 ( .ina ({new_AGEMA_signal_13122, new_AGEMA_signal_13118, new_AGEMA_signal_13114, new_AGEMA_signal_13110}), .inb ({new_AGEMA_signal_2288, new_AGEMA_signal_2287, new_AGEMA_signal_2286, n2459}), .clk ( clk ), .rnd ({Fresh[5119], Fresh[5118], Fresh[5117], Fresh[5116], Fresh[5115], Fresh[5114], Fresh[5113], Fresh[5112], Fresh[5111], Fresh[5110]}), .outt ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, new_AGEMA_signal_2703, n2686}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2460 ( .ina ({new_AGEMA_signal_13138, new_AGEMA_signal_13136, new_AGEMA_signal_13134, new_AGEMA_signal_13132}), .inb ({new_AGEMA_signal_2291, new_AGEMA_signal_2290, new_AGEMA_signal_2289, n2288}), .clk ( clk ), .rnd ({Fresh[5129], Fresh[5128], Fresh[5127], Fresh[5126], Fresh[5125], Fresh[5124], Fresh[5123], Fresh[5122], Fresh[5121], Fresh[5120]}), .outt ({new_AGEMA_signal_2708, new_AGEMA_signal_2707, new_AGEMA_signal_2706, n2289}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2463 ( .ina ({new_AGEMA_signal_2294, new_AGEMA_signal_2293, new_AGEMA_signal_2292, n2458}), .inb ({new_AGEMA_signal_13474, new_AGEMA_signal_13472, new_AGEMA_signal_13470, new_AGEMA_signal_13468}), .clk ( clk ), .rnd ({Fresh[5139], Fresh[5138], Fresh[5137], Fresh[5136], Fresh[5135], Fresh[5134], Fresh[5133], Fresh[5132], Fresh[5131], Fresh[5130]}), .outt ({new_AGEMA_signal_2711, new_AGEMA_signal_2710, new_AGEMA_signal_2709, n2297}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2465 ( .ina ({new_AGEMA_signal_13482, new_AGEMA_signal_13480, new_AGEMA_signal_13478, new_AGEMA_signal_13476}), .inb ({new_AGEMA_signal_2192, new_AGEMA_signal_2191, new_AGEMA_signal_2190, n2291}), .clk ( clk ), .rnd ({Fresh[5149], Fresh[5148], Fresh[5147], Fresh[5146], Fresh[5145], Fresh[5144], Fresh[5143], Fresh[5142], Fresh[5141], Fresh[5140]}), .outt ({new_AGEMA_signal_2714, new_AGEMA_signal_2713, new_AGEMA_signal_2712, n2292}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2473 ( .ina ({new_AGEMA_signal_13490, new_AGEMA_signal_13488, new_AGEMA_signal_13486, new_AGEMA_signal_13484}), .inb ({new_AGEMA_signal_2300, new_AGEMA_signal_2299, new_AGEMA_signal_2298, n2300}), .clk ( clk ), .rnd ({Fresh[5159], Fresh[5158], Fresh[5157], Fresh[5156], Fresh[5155], Fresh[5154], Fresh[5153], Fresh[5152], Fresh[5151], Fresh[5150]}), .outt ({new_AGEMA_signal_2717, new_AGEMA_signal_2716, new_AGEMA_signal_2715, n2301}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2483 ( .ina ({new_AGEMA_signal_13498, new_AGEMA_signal_13496, new_AGEMA_signal_13494, new_AGEMA_signal_13492}), .inb ({new_AGEMA_signal_2306, new_AGEMA_signal_2305, new_AGEMA_signal_2304, n2314}), .clk ( clk ), .rnd ({Fresh[5169], Fresh[5168], Fresh[5167], Fresh[5166], Fresh[5165], Fresh[5164], Fresh[5163], Fresh[5162], Fresh[5161], Fresh[5160]}), .outt ({new_AGEMA_signal_2720, new_AGEMA_signal_2719, new_AGEMA_signal_2718, n2321}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2487 ( .ina ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, new_AGEMA_signal_1407, n2319}), .inb ({new_AGEMA_signal_13506, new_AGEMA_signal_13504, new_AGEMA_signal_13502, new_AGEMA_signal_13500}), .clk ( clk ), .rnd ({Fresh[5179], Fresh[5178], Fresh[5177], Fresh[5176], Fresh[5175], Fresh[5174], Fresh[5173], Fresh[5172], Fresh[5171], Fresh[5170]}), .outt ({new_AGEMA_signal_1817, new_AGEMA_signal_1816, new_AGEMA_signal_1815, n2320}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2493 ( .ina ({new_AGEMA_signal_1820, new_AGEMA_signal_1819, new_AGEMA_signal_1818, n2326}), .inb ({new_AGEMA_signal_13514, new_AGEMA_signal_13512, new_AGEMA_signal_13510, new_AGEMA_signal_13508}), .clk ( clk ), .rnd ({Fresh[5189], Fresh[5188], Fresh[5187], Fresh[5186], Fresh[5185], Fresh[5184], Fresh[5183], Fresh[5182], Fresh[5181], Fresh[5180]}), .outt ({new_AGEMA_signal_2309, new_AGEMA_signal_2308, new_AGEMA_signal_2307, n2334}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2497 ( .ina ({new_AGEMA_signal_2312, new_AGEMA_signal_2311, new_AGEMA_signal_2310, n2329}), .inb ({new_AGEMA_signal_13226, new_AGEMA_signal_13222, new_AGEMA_signal_13218, new_AGEMA_signal_13214}), .clk ( clk ), .rnd ({Fresh[5199], Fresh[5198], Fresh[5197], Fresh[5196], Fresh[5195], Fresh[5194], Fresh[5193], Fresh[5192], Fresh[5191], Fresh[5190]}), .outt ({new_AGEMA_signal_2723, new_AGEMA_signal_2722, new_AGEMA_signal_2721, n2332}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2498 ( .ina ({new_AGEMA_signal_13522, new_AGEMA_signal_13520, new_AGEMA_signal_13518, new_AGEMA_signal_13516}), .inb ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, new_AGEMA_signal_2175, n2330}), .clk ( clk ), .rnd ({Fresh[5209], Fresh[5208], Fresh[5207], Fresh[5206], Fresh[5205], Fresh[5204], Fresh[5203], Fresh[5202], Fresh[5201], Fresh[5200]}), .outt ({new_AGEMA_signal_2726, new_AGEMA_signal_2725, new_AGEMA_signal_2724, n2331}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2502 ( .ina ({new_AGEMA_signal_13530, new_AGEMA_signal_13528, new_AGEMA_signal_13526, new_AGEMA_signal_13524}), .inb ({new_AGEMA_signal_2729, new_AGEMA_signal_2728, new_AGEMA_signal_2727, n2335}), .clk ( clk ), .rnd ({Fresh[5219], Fresh[5218], Fresh[5217], Fresh[5216], Fresh[5215], Fresh[5214], Fresh[5213], Fresh[5212], Fresh[5211], Fresh[5210]}), .outt ({new_AGEMA_signal_2996, new_AGEMA_signal_2995, new_AGEMA_signal_2994, n2336}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2508 ( .ina ({new_AGEMA_signal_2315, new_AGEMA_signal_2314, new_AGEMA_signal_2313, n2341}), .inb ({new_AGEMA_signal_1832, new_AGEMA_signal_1831, new_AGEMA_signal_1830, n2340}), .clk ( clk ), .rnd ({Fresh[5229], Fresh[5228], Fresh[5227], Fresh[5226], Fresh[5225], Fresh[5224], Fresh[5223], Fresh[5222], Fresh[5221], Fresh[5220]}), .outt ({new_AGEMA_signal_2732, new_AGEMA_signal_2731, new_AGEMA_signal_2730, n2342}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2519 ( .ina ({new_AGEMA_signal_1844, new_AGEMA_signal_1843, new_AGEMA_signal_1842, n2352}), .inb ({new_AGEMA_signal_13538, new_AGEMA_signal_13536, new_AGEMA_signal_13534, new_AGEMA_signal_13532}), .clk ( clk ), .rnd ({Fresh[5239], Fresh[5238], Fresh[5237], Fresh[5236], Fresh[5235], Fresh[5234], Fresh[5233], Fresh[5232], Fresh[5231], Fresh[5230]}), .outt ({new_AGEMA_signal_2318, new_AGEMA_signal_2317, new_AGEMA_signal_2316, n2367}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2523 ( .ina ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, new_AGEMA_signal_2319, n2354}), .inb ({new_AGEMA_signal_13546, new_AGEMA_signal_13544, new_AGEMA_signal_13542, new_AGEMA_signal_13540}), .clk ( clk ), .rnd ({Fresh[5249], Fresh[5248], Fresh[5247], Fresh[5246], Fresh[5245], Fresh[5244], Fresh[5243], Fresh[5242], Fresh[5241], Fresh[5240]}), .outt ({new_AGEMA_signal_2735, new_AGEMA_signal_2734, new_AGEMA_signal_2733, n2358}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2547 ( .ina ({new_AGEMA_signal_1859, new_AGEMA_signal_1858, new_AGEMA_signal_1857, n2385}), .inb ({new_AGEMA_signal_1862, new_AGEMA_signal_1861, new_AGEMA_signal_1860, n2384}), .clk ( clk ), .rnd ({Fresh[5259], Fresh[5258], Fresh[5257], Fresh[5256], Fresh[5255], Fresh[5254], Fresh[5253], Fresh[5252], Fresh[5251], Fresh[5250]}), .outt ({new_AGEMA_signal_2336, new_AGEMA_signal_2335, new_AGEMA_signal_2334, n2387}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2555 ( .ina ({new_AGEMA_signal_1868, new_AGEMA_signal_1867, new_AGEMA_signal_1866, n2391}), .inb ({new_AGEMA_signal_2342, new_AGEMA_signal_2341, new_AGEMA_signal_2340, n2390}), .clk ( clk ), .rnd ({Fresh[5269], Fresh[5268], Fresh[5267], Fresh[5266], Fresh[5265], Fresh[5264], Fresh[5263], Fresh[5262], Fresh[5261], Fresh[5260]}), .outt ({new_AGEMA_signal_2744, new_AGEMA_signal_2743, new_AGEMA_signal_2742, n2392}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2566 ( .ina ({new_AGEMA_signal_1874, new_AGEMA_signal_1873, new_AGEMA_signal_1872, n2403}), .inb ({new_AGEMA_signal_13554, new_AGEMA_signal_13552, new_AGEMA_signal_13550, new_AGEMA_signal_13548}), .clk ( clk ), .rnd ({Fresh[5279], Fresh[5278], Fresh[5277], Fresh[5276], Fresh[5275], Fresh[5274], Fresh[5273], Fresh[5272], Fresh[5271], Fresh[5270]}), .outt ({new_AGEMA_signal_2348, new_AGEMA_signal_2347, new_AGEMA_signal_2346, n2404}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2570 ( .ina ({new_AGEMA_signal_13274, new_AGEMA_signal_13272, new_AGEMA_signal_13270, new_AGEMA_signal_13268}), .inb ({new_AGEMA_signal_2351, new_AGEMA_signal_2350, new_AGEMA_signal_2349, n2408}), .clk ( clk ), .rnd ({Fresh[5289], Fresh[5288], Fresh[5287], Fresh[5286], Fresh[5285], Fresh[5284], Fresh[5283], Fresh[5282], Fresh[5281], Fresh[5280]}), .outt ({new_AGEMA_signal_2750, new_AGEMA_signal_2749, new_AGEMA_signal_2748, n2409}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2575 ( .ina ({new_AGEMA_signal_2354, new_AGEMA_signal_2353, new_AGEMA_signal_2352, n2574}), .inb ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, new_AGEMA_signal_1875, n2413}), .clk ( clk ), .rnd ({Fresh[5299], Fresh[5298], Fresh[5297], Fresh[5296], Fresh[5295], Fresh[5294], Fresh[5293], Fresh[5292], Fresh[5291], Fresh[5290]}), .outt ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, new_AGEMA_signal_2751, n2414}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2578 ( .ina ({new_AGEMA_signal_13562, new_AGEMA_signal_13560, new_AGEMA_signal_13558, new_AGEMA_signal_13556}), .inb ({new_AGEMA_signal_1880, new_AGEMA_signal_1879, new_AGEMA_signal_1878, n2416}), .clk ( clk ), .rnd ({Fresh[5309], Fresh[5308], Fresh[5307], Fresh[5306], Fresh[5305], Fresh[5304], Fresh[5303], Fresh[5302], Fresh[5301], Fresh[5300]}), .outt ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, new_AGEMA_signal_2355, n2418}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2589 ( .ina ({new_AGEMA_signal_2363, new_AGEMA_signal_2362, new_AGEMA_signal_2361, n2689}), .inb ({new_AGEMA_signal_13570, new_AGEMA_signal_13568, new_AGEMA_signal_13566, new_AGEMA_signal_13564}), .clk ( clk ), .rnd ({Fresh[5319], Fresh[5318], Fresh[5317], Fresh[5316], Fresh[5315], Fresh[5314], Fresh[5313], Fresh[5312], Fresh[5311], Fresh[5310]}), .outt ({new_AGEMA_signal_2759, new_AGEMA_signal_2758, new_AGEMA_signal_2757, n2432}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2592 ( .ina ({new_AGEMA_signal_13594, new_AGEMA_signal_13588, new_AGEMA_signal_13582, new_AGEMA_signal_13576}), .inb ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, new_AGEMA_signal_1887, n2434}), .clk ( clk ), .rnd ({Fresh[5329], Fresh[5328], Fresh[5327], Fresh[5326], Fresh[5325], Fresh[5324], Fresh[5323], Fresh[5322], Fresh[5321], Fresh[5320]}), .outt ({new_AGEMA_signal_2366, new_AGEMA_signal_2365, new_AGEMA_signal_2364, n2435}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2601 ( .ina ({new_AGEMA_signal_2372, new_AGEMA_signal_2371, new_AGEMA_signal_2370, n2445}), .inb ({new_AGEMA_signal_2375, new_AGEMA_signal_2374, new_AGEMA_signal_2373, n2444}), .clk ( clk ), .rnd ({Fresh[5339], Fresh[5338], Fresh[5337], Fresh[5336], Fresh[5335], Fresh[5334], Fresh[5333], Fresh[5332], Fresh[5331], Fresh[5330]}), .outt ({new_AGEMA_signal_2762, new_AGEMA_signal_2761, new_AGEMA_signal_2760, n2449}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2603 ( .ina ({new_AGEMA_signal_13498, new_AGEMA_signal_13496, new_AGEMA_signal_13494, new_AGEMA_signal_13492}), .inb ({new_AGEMA_signal_2378, new_AGEMA_signal_2377, new_AGEMA_signal_2376, n2447}), .clk ( clk ), .rnd ({Fresh[5349], Fresh[5348], Fresh[5347], Fresh[5346], Fresh[5345], Fresh[5344], Fresh[5343], Fresh[5342], Fresh[5341], Fresh[5340]}), .outt ({new_AGEMA_signal_2765, new_AGEMA_signal_2764, new_AGEMA_signal_2763, n2448}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2609 ( .ina ({new_AGEMA_signal_2381, new_AGEMA_signal_2380, new_AGEMA_signal_2379, n2454}), .inb ({new_AGEMA_signal_13602, new_AGEMA_signal_13600, new_AGEMA_signal_13598, new_AGEMA_signal_13596}), .clk ( clk ), .rnd ({Fresh[5359], Fresh[5358], Fresh[5357], Fresh[5356], Fresh[5355], Fresh[5354], Fresh[5353], Fresh[5352], Fresh[5351], Fresh[5350]}), .outt ({new_AGEMA_signal_2768, new_AGEMA_signal_2767, new_AGEMA_signal_2766, n2455}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2612 ( .ina ({new_AGEMA_signal_2078, new_AGEMA_signal_2077, new_AGEMA_signal_2076, n2687}), .inb ({new_AGEMA_signal_2294, new_AGEMA_signal_2293, new_AGEMA_signal_2292, n2458}), .clk ( clk ), .rnd ({Fresh[5369], Fresh[5368], Fresh[5367], Fresh[5366], Fresh[5365], Fresh[5364], Fresh[5363], Fresh[5362], Fresh[5361], Fresh[5360]}), .outt ({new_AGEMA_signal_2771, new_AGEMA_signal_2770, new_AGEMA_signal_2769, n2460}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2618 ( .ina ({new_AGEMA_signal_13482, new_AGEMA_signal_13480, new_AGEMA_signal_13478, new_AGEMA_signal_13476}), .inb ({new_AGEMA_signal_1898, new_AGEMA_signal_1897, new_AGEMA_signal_1896, n2465}), .clk ( clk ), .rnd ({Fresh[5379], Fresh[5378], Fresh[5377], Fresh[5376], Fresh[5375], Fresh[5374], Fresh[5373], Fresh[5372], Fresh[5371], Fresh[5370]}), .outt ({new_AGEMA_signal_2384, new_AGEMA_signal_2383, new_AGEMA_signal_2382, n2466}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2629 ( .ina ({new_AGEMA_signal_1904, new_AGEMA_signal_1903, new_AGEMA_signal_1902, n2476}), .inb ({new_AGEMA_signal_13610, new_AGEMA_signal_13608, new_AGEMA_signal_13606, new_AGEMA_signal_13604}), .clk ( clk ), .rnd ({Fresh[5389], Fresh[5388], Fresh[5387], Fresh[5386], Fresh[5385], Fresh[5384], Fresh[5383], Fresh[5382], Fresh[5381], Fresh[5380]}), .outt ({new_AGEMA_signal_2387, new_AGEMA_signal_2386, new_AGEMA_signal_2385, n2477}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2634 ( .ina ({new_AGEMA_signal_13266, new_AGEMA_signal_13264, new_AGEMA_signal_13262, new_AGEMA_signal_13260}), .inb ({new_AGEMA_signal_2390, new_AGEMA_signal_2389, new_AGEMA_signal_2388, n2481}), .clk ( clk ), .rnd ({Fresh[5399], Fresh[5398], Fresh[5397], Fresh[5396], Fresh[5395], Fresh[5394], Fresh[5393], Fresh[5392], Fresh[5391], Fresh[5390]}), .outt ({new_AGEMA_signal_2780, new_AGEMA_signal_2779, new_AGEMA_signal_2778, n2482}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2640 ( .ina ({new_AGEMA_signal_13618, new_AGEMA_signal_13616, new_AGEMA_signal_13614, new_AGEMA_signal_13612}), .inb ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, new_AGEMA_signal_1911, n2486}), .clk ( clk ), .rnd ({Fresh[5409], Fresh[5408], Fresh[5407], Fresh[5406], Fresh[5405], Fresh[5404], Fresh[5403], Fresh[5402], Fresh[5401], Fresh[5400]}), .outt ({new_AGEMA_signal_2393, new_AGEMA_signal_2392, new_AGEMA_signal_2391, n2490}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2648 ( .ina ({new_AGEMA_signal_1922, new_AGEMA_signal_1921, new_AGEMA_signal_1920, n2495}), .inb ({new_AGEMA_signal_2396, new_AGEMA_signal_2395, new_AGEMA_signal_2394, n2494}), .clk ( clk ), .rnd ({Fresh[5419], Fresh[5418], Fresh[5417], Fresh[5416], Fresh[5415], Fresh[5414], Fresh[5413], Fresh[5412], Fresh[5411], Fresh[5410]}), .outt ({new_AGEMA_signal_2786, new_AGEMA_signal_2785, new_AGEMA_signal_2784, n2496}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2654 ( .ina ({new_AGEMA_signal_1685, new_AGEMA_signal_1684, new_AGEMA_signal_1683, n2504}), .inb ({new_AGEMA_signal_2789, new_AGEMA_signal_2788, new_AGEMA_signal_2787, n2503}), .clk ( clk ), .rnd ({Fresh[5429], Fresh[5428], Fresh[5427], Fresh[5426], Fresh[5425], Fresh[5424], Fresh[5423], Fresh[5422], Fresh[5421], Fresh[5420]}), .outt ({new_AGEMA_signal_3047, new_AGEMA_signal_3046, new_AGEMA_signal_3045, n2507}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2664 ( .ina ({new_AGEMA_signal_2402, new_AGEMA_signal_2401, new_AGEMA_signal_2400, n2518}), .inb ({new_AGEMA_signal_2792, new_AGEMA_signal_2791, new_AGEMA_signal_2790, n2517}), .clk ( clk ), .rnd ({Fresh[5439], Fresh[5438], Fresh[5437], Fresh[5436], Fresh[5435], Fresh[5434], Fresh[5433], Fresh[5432], Fresh[5431], Fresh[5430]}), .outt ({new_AGEMA_signal_3050, new_AGEMA_signal_3049, new_AGEMA_signal_3048, n2525}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2669 ( .ina ({new_AGEMA_signal_2405, new_AGEMA_signal_2404, new_AGEMA_signal_2403, n2523}), .inb ({new_AGEMA_signal_2408, new_AGEMA_signal_2407, new_AGEMA_signal_2406, n2522}), .clk ( clk ), .rnd ({Fresh[5449], Fresh[5448], Fresh[5447], Fresh[5446], Fresh[5445], Fresh[5444], Fresh[5443], Fresh[5442], Fresh[5441], Fresh[5440]}), .outt ({new_AGEMA_signal_2795, new_AGEMA_signal_2794, new_AGEMA_signal_2793, n2524}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2676 ( .ina ({new_AGEMA_signal_2411, new_AGEMA_signal_2410, new_AGEMA_signal_2409, n2532}), .inb ({new_AGEMA_signal_13634, new_AGEMA_signal_13630, new_AGEMA_signal_13626, new_AGEMA_signal_13622}), .clk ( clk ), .rnd ({Fresh[5459], Fresh[5458], Fresh[5457], Fresh[5456], Fresh[5455], Fresh[5454], Fresh[5453], Fresh[5452], Fresh[5451], Fresh[5450]}), .outt ({new_AGEMA_signal_2798, new_AGEMA_signal_2797, new_AGEMA_signal_2796, n2537}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2678 ( .ina ({new_AGEMA_signal_13274, new_AGEMA_signal_13272, new_AGEMA_signal_13270, new_AGEMA_signal_13268}), .inb ({new_AGEMA_signal_2414, new_AGEMA_signal_2413, new_AGEMA_signal_2412, n2534}), .clk ( clk ), .rnd ({Fresh[5469], Fresh[5468], Fresh[5467], Fresh[5466], Fresh[5465], Fresh[5464], Fresh[5463], Fresh[5462], Fresh[5461], Fresh[5460]}), .outt ({new_AGEMA_signal_2801, new_AGEMA_signal_2800, new_AGEMA_signal_2799, n2536}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2684 ( .ina ({new_AGEMA_signal_13642, new_AGEMA_signal_13640, new_AGEMA_signal_13638, new_AGEMA_signal_13636}), .inb ({new_AGEMA_signal_1934, new_AGEMA_signal_1933, new_AGEMA_signal_1932, n2546}), .clk ( clk ), .rnd ({Fresh[5479], Fresh[5478], Fresh[5477], Fresh[5476], Fresh[5475], Fresh[5474], Fresh[5473], Fresh[5472], Fresh[5471], Fresh[5470]}), .outt ({new_AGEMA_signal_2420, new_AGEMA_signal_2419, new_AGEMA_signal_2418, n2547}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2693 ( .ina ({new_AGEMA_signal_13650, new_AGEMA_signal_13648, new_AGEMA_signal_13646, new_AGEMA_signal_13644}), .inb ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, new_AGEMA_signal_2427, n2556}), .clk ( clk ), .rnd ({Fresh[5489], Fresh[5488], Fresh[5487], Fresh[5486], Fresh[5485], Fresh[5484], Fresh[5483], Fresh[5482], Fresh[5481], Fresh[5480]}), .outt ({new_AGEMA_signal_2804, new_AGEMA_signal_2803, new_AGEMA_signal_2802, n2557}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2699 ( .ina ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, new_AGEMA_signal_2433, n2715}), .inb ({new_AGEMA_signal_13658, new_AGEMA_signal_13656, new_AGEMA_signal_13654, new_AGEMA_signal_13652}), .clk ( clk ), .rnd ({Fresh[5499], Fresh[5498], Fresh[5497], Fresh[5496], Fresh[5495], Fresh[5494], Fresh[5493], Fresh[5492], Fresh[5491], Fresh[5490]}), .outt ({new_AGEMA_signal_2807, new_AGEMA_signal_2806, new_AGEMA_signal_2805, n2565}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2704 ( .ina ({new_AGEMA_signal_2354, new_AGEMA_signal_2353, new_AGEMA_signal_2352, n2574}), .inb ({new_AGEMA_signal_2438, new_AGEMA_signal_2437, new_AGEMA_signal_2436, n2573}), .clk ( clk ), .rnd ({Fresh[5509], Fresh[5508], Fresh[5507], Fresh[5506], Fresh[5505], Fresh[5504], Fresh[5503], Fresh[5502], Fresh[5501], Fresh[5500]}), .outt ({new_AGEMA_signal_2810, new_AGEMA_signal_2809, new_AGEMA_signal_2808, n2591}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2709 ( .ina ({new_AGEMA_signal_2444, new_AGEMA_signal_2443, new_AGEMA_signal_2442, n2579}), .inb ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, new_AGEMA_signal_1947, n2578}), .clk ( clk ), .rnd ({Fresh[5519], Fresh[5518], Fresh[5517], Fresh[5516], Fresh[5515], Fresh[5514], Fresh[5513], Fresh[5512], Fresh[5511], Fresh[5510]}), .outt ({new_AGEMA_signal_2813, new_AGEMA_signal_2812, new_AGEMA_signal_2811, n2580}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2727 ( .ina ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, new_AGEMA_signal_1470, n2601}), .inb ({new_AGEMA_signal_13674, new_AGEMA_signal_13670, new_AGEMA_signal_13666, new_AGEMA_signal_13662}), .clk ( clk ), .rnd ({Fresh[5529], Fresh[5528], Fresh[5527], Fresh[5526], Fresh[5525], Fresh[5524], Fresh[5523], Fresh[5522], Fresh[5521], Fresh[5520]}), .outt ({new_AGEMA_signal_1964, new_AGEMA_signal_1963, new_AGEMA_signal_1962, n2602}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2738 ( .ina ({new_AGEMA_signal_2462, new_AGEMA_signal_2461, new_AGEMA_signal_2460, n2618}), .inb ({new_AGEMA_signal_13682, new_AGEMA_signal_13680, new_AGEMA_signal_13678, new_AGEMA_signal_13676}), .clk ( clk ), .rnd ({Fresh[5539], Fresh[5538], Fresh[5537], Fresh[5536], Fresh[5535], Fresh[5534], Fresh[5533], Fresh[5532], Fresh[5531], Fresh[5530]}), .outt ({new_AGEMA_signal_2819, new_AGEMA_signal_2818, new_AGEMA_signal_2817, n2619}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2744 ( .ina ({new_AGEMA_signal_13314, new_AGEMA_signal_13312, new_AGEMA_signal_13310, new_AGEMA_signal_13308}), .inb ({new_AGEMA_signal_2465, new_AGEMA_signal_2464, new_AGEMA_signal_2463, n2626}), .clk ( clk ), .rnd ({Fresh[5549], Fresh[5548], Fresh[5547], Fresh[5546], Fresh[5545], Fresh[5544], Fresh[5543], Fresh[5542], Fresh[5541], Fresh[5540]}), .outt ({new_AGEMA_signal_2822, new_AGEMA_signal_2821, new_AGEMA_signal_2820, n2628}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2753 ( .ina ({new_AGEMA_signal_2468, new_AGEMA_signal_2467, new_AGEMA_signal_2466, n2644}), .inb ({new_AGEMA_signal_13370, new_AGEMA_signal_13368, new_AGEMA_signal_13366, new_AGEMA_signal_13364}), .clk ( clk ), .rnd ({Fresh[5559], Fresh[5558], Fresh[5557], Fresh[5556], Fresh[5555], Fresh[5554], Fresh[5553], Fresh[5552], Fresh[5551], Fresh[5550]}), .outt ({new_AGEMA_signal_2825, new_AGEMA_signal_2824, new_AGEMA_signal_2823, n2649}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2755 ( .ina ({new_AGEMA_signal_13690, new_AGEMA_signal_13688, new_AGEMA_signal_13686, new_AGEMA_signal_13684}), .inb ({new_AGEMA_signal_1982, new_AGEMA_signal_1981, new_AGEMA_signal_1980, n2646}), .clk ( clk ), .rnd ({Fresh[5569], Fresh[5568], Fresh[5567], Fresh[5566], Fresh[5565], Fresh[5564], Fresh[5563], Fresh[5562], Fresh[5561], Fresh[5560]}), .outt ({new_AGEMA_signal_2471, new_AGEMA_signal_2470, new_AGEMA_signal_2469, n2648}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2765 ( .ina ({new_AGEMA_signal_13138, new_AGEMA_signal_13136, new_AGEMA_signal_13134, new_AGEMA_signal_13132}), .inb ({new_AGEMA_signal_2477, new_AGEMA_signal_2476, new_AGEMA_signal_2475, n2663}), .clk ( clk ), .rnd ({Fresh[5579], Fresh[5578], Fresh[5577], Fresh[5576], Fresh[5575], Fresh[5574], Fresh[5573], Fresh[5572], Fresh[5571], Fresh[5570]}), .outt ({new_AGEMA_signal_2828, new_AGEMA_signal_2827, new_AGEMA_signal_2826, n2664}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2771 ( .ina ({new_AGEMA_signal_1988, new_AGEMA_signal_1987, new_AGEMA_signal_1986, n2675}), .inb ({new_AGEMA_signal_13698, new_AGEMA_signal_13696, new_AGEMA_signal_13694, new_AGEMA_signal_13692}), .clk ( clk ), .rnd ({Fresh[5589], Fresh[5588], Fresh[5587], Fresh[5586], Fresh[5585], Fresh[5584], Fresh[5583], Fresh[5582], Fresh[5581], Fresh[5580]}), .outt ({new_AGEMA_signal_2831, new_AGEMA_signal_2830, new_AGEMA_signal_2829, n2681}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2773 ( .ina ({new_AGEMA_signal_13402, new_AGEMA_signal_13400, new_AGEMA_signal_13398, new_AGEMA_signal_13396}), .inb ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, new_AGEMA_signal_1989, n2678}), .clk ( clk ), .rnd ({Fresh[5599], Fresh[5598], Fresh[5597], Fresh[5596], Fresh[5595], Fresh[5594], Fresh[5593], Fresh[5592], Fresh[5591], Fresh[5590]}), .outt ({new_AGEMA_signal_2480, new_AGEMA_signal_2479, new_AGEMA_signal_2478, n2680}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2776 ( .ina ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, new_AGEMA_signal_2091, n2684}), .inb ({new_AGEMA_signal_13706, new_AGEMA_signal_13704, new_AGEMA_signal_13702, new_AGEMA_signal_13700}), .clk ( clk ), .rnd ({Fresh[5609], Fresh[5608], Fresh[5607], Fresh[5606], Fresh[5605], Fresh[5604], Fresh[5603], Fresh[5602], Fresh[5601], Fresh[5600]}), .outt ({new_AGEMA_signal_2834, new_AGEMA_signal_2833, new_AGEMA_signal_2832, n2685}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2778 ( .ina ({new_AGEMA_signal_2078, new_AGEMA_signal_2077, new_AGEMA_signal_2076, n2687}), .inb ({new_AGEMA_signal_13642, new_AGEMA_signal_13640, new_AGEMA_signal_13638, new_AGEMA_signal_13636}), .clk ( clk ), .rnd ({Fresh[5619], Fresh[5618], Fresh[5617], Fresh[5616], Fresh[5615], Fresh[5614], Fresh[5613], Fresh[5612], Fresh[5611], Fresh[5610]}), .outt ({new_AGEMA_signal_2837, new_AGEMA_signal_2836, new_AGEMA_signal_2835, n2698}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2779 ( .ina ({new_AGEMA_signal_2363, new_AGEMA_signal_2362, new_AGEMA_signal_2361, n2689}), .inb ({new_AGEMA_signal_13650, new_AGEMA_signal_13648, new_AGEMA_signal_13646, new_AGEMA_signal_13644}), .clk ( clk ), .rnd ({Fresh[5629], Fresh[5628], Fresh[5627], Fresh[5626], Fresh[5625], Fresh[5624], Fresh[5623], Fresh[5622], Fresh[5621], Fresh[5620]}), .outt ({new_AGEMA_signal_2840, new_AGEMA_signal_2839, new_AGEMA_signal_2838, n2692}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2793 ( .ina ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, new_AGEMA_signal_2433, n2715}), .inb ({new_AGEMA_signal_13714, new_AGEMA_signal_13712, new_AGEMA_signal_13710, new_AGEMA_signal_13708}), .clk ( clk ), .rnd ({Fresh[5639], Fresh[5638], Fresh[5637], Fresh[5636], Fresh[5635], Fresh[5634], Fresh[5633], Fresh[5632], Fresh[5631], Fresh[5630]}), .outt ({new_AGEMA_signal_2843, new_AGEMA_signal_2842, new_AGEMA_signal_2841, n2716}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2800 ( .ina ({new_AGEMA_signal_2006, new_AGEMA_signal_2005, new_AGEMA_signal_2004, n2727}), .inb ({new_AGEMA_signal_13722, new_AGEMA_signal_13720, new_AGEMA_signal_13718, new_AGEMA_signal_13716}), .clk ( clk ), .rnd ({Fresh[5649], Fresh[5648], Fresh[5647], Fresh[5646], Fresh[5645], Fresh[5644], Fresh[5643], Fresh[5642], Fresh[5641], Fresh[5640]}), .outt ({new_AGEMA_signal_2489, new_AGEMA_signal_2488, new_AGEMA_signal_2487, n2728}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2804 ( .ina ({new_AGEMA_signal_13730, new_AGEMA_signal_13728, new_AGEMA_signal_13726, new_AGEMA_signal_13724}), .inb ({new_AGEMA_signal_2492, new_AGEMA_signal_2491, new_AGEMA_signal_2490, n2733}), .clk ( clk ), .rnd ({Fresh[5659], Fresh[5658], Fresh[5657], Fresh[5656], Fresh[5655], Fresh[5654], Fresh[5653], Fresh[5652], Fresh[5651], Fresh[5650]}), .outt ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, new_AGEMA_signal_2847, n2735}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2808 ( .ina ({new_AGEMA_signal_13186, new_AGEMA_signal_13184, new_AGEMA_signal_13182, new_AGEMA_signal_13180}), .inb ({new_AGEMA_signal_2495, new_AGEMA_signal_2494, new_AGEMA_signal_2493, n2740}), .clk ( clk ), .rnd ({Fresh[5669], Fresh[5668], Fresh[5667], Fresh[5666], Fresh[5665], Fresh[5664], Fresh[5663], Fresh[5662], Fresh[5661], Fresh[5660]}), .outt ({new_AGEMA_signal_2852, new_AGEMA_signal_2851, new_AGEMA_signal_2850, n2743}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2813 ( .ina ({new_AGEMA_signal_13746, new_AGEMA_signal_13742, new_AGEMA_signal_13738, new_AGEMA_signal_13734}), .inb ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, new_AGEMA_signal_2013, n2749}), .clk ( clk ), .rnd ({Fresh[5679], Fresh[5678], Fresh[5677], Fresh[5676], Fresh[5675], Fresh[5674], Fresh[5673], Fresh[5672], Fresh[5671], Fresh[5670]}), .outt ({new_AGEMA_signal_2498, new_AGEMA_signal_2497, new_AGEMA_signal_2496, n2751}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2817 ( .ina ({new_AGEMA_signal_2501, new_AGEMA_signal_2500, new_AGEMA_signal_2499, n2757}), .inb ({new_AGEMA_signal_2018, new_AGEMA_signal_2017, new_AGEMA_signal_2016, n2756}), .clk ( clk ), .rnd ({Fresh[5689], Fresh[5688], Fresh[5687], Fresh[5686], Fresh[5685], Fresh[5684], Fresh[5683], Fresh[5682], Fresh[5681], Fresh[5680]}), .outt ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, new_AGEMA_signal_2853, n2758}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2820 ( .ina ({new_AGEMA_signal_13754, new_AGEMA_signal_13752, new_AGEMA_signal_13750, new_AGEMA_signal_13748}), .inb ({new_AGEMA_signal_2504, new_AGEMA_signal_2503, new_AGEMA_signal_2502, n2762}), .clk ( clk ), .rnd ({Fresh[5699], Fresh[5698], Fresh[5697], Fresh[5696], Fresh[5695], Fresh[5694], Fresh[5693], Fresh[5692], Fresh[5691], Fresh[5690]}), .outt ({new_AGEMA_signal_2858, new_AGEMA_signal_2857, new_AGEMA_signal_2856, n2764}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2827 ( .ina ({new_AGEMA_signal_2510, new_AGEMA_signal_2509, new_AGEMA_signal_2508, n2776}), .inb ({new_AGEMA_signal_2513, new_AGEMA_signal_2512, new_AGEMA_signal_2511, n2775}), .clk ( clk ), .rnd ({Fresh[5709], Fresh[5708], Fresh[5707], Fresh[5706], Fresh[5705], Fresh[5704], Fresh[5703], Fresh[5702], Fresh[5701], Fresh[5700]}), .outt ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, new_AGEMA_signal_2859, n2800}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2831 ( .ina ({new_AGEMA_signal_13762, new_AGEMA_signal_13760, new_AGEMA_signal_13758, new_AGEMA_signal_13756}), .inb ({new_AGEMA_signal_2024, new_AGEMA_signal_2023, new_AGEMA_signal_2022, n2783}), .clk ( clk ), .rnd ({Fresh[5719], Fresh[5718], Fresh[5717], Fresh[5716], Fresh[5715], Fresh[5714], Fresh[5713], Fresh[5712], Fresh[5711], Fresh[5710]}), .outt ({new_AGEMA_signal_2516, new_AGEMA_signal_2515, new_AGEMA_signal_2514, n2788}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2837 ( .ina ({new_AGEMA_signal_13778, new_AGEMA_signal_13774, new_AGEMA_signal_13770, new_AGEMA_signal_13766}), .inb ({new_AGEMA_signal_2519, new_AGEMA_signal_2518, new_AGEMA_signal_2517, n2795}), .clk ( clk ), .rnd ({Fresh[5729], Fresh[5728], Fresh[5727], Fresh[5726], Fresh[5725], Fresh[5724], Fresh[5723], Fresh[5722], Fresh[5721], Fresh[5720]}), .outt ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, new_AGEMA_signal_2865, n2797}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2846 ( .ina ({new_AGEMA_signal_2522, new_AGEMA_signal_2521, new_AGEMA_signal_2520, n2814}), .inb ({new_AGEMA_signal_13210, new_AGEMA_signal_13208, new_AGEMA_signal_13206, new_AGEMA_signal_13204}), .clk ( clk ), .rnd ({Fresh[5739], Fresh[5738], Fresh[5737], Fresh[5736], Fresh[5735], Fresh[5734], Fresh[5733], Fresh[5732], Fresh[5731], Fresh[5730]}), .outt ({new_AGEMA_signal_2870, new_AGEMA_signal_2869, new_AGEMA_signal_2868, n2822}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2849 ( .ina ({new_AGEMA_signal_13786, new_AGEMA_signal_13784, new_AGEMA_signal_13782, new_AGEMA_signal_13780}), .inb ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, new_AGEMA_signal_2037, n2819}), .clk ( clk ), .rnd ({Fresh[5749], Fresh[5748], Fresh[5747], Fresh[5746], Fresh[5745], Fresh[5744], Fresh[5743], Fresh[5742], Fresh[5741], Fresh[5740]}), .outt ({new_AGEMA_signal_2525, new_AGEMA_signal_2524, new_AGEMA_signal_2523, n2821}) ) ;
    buf_clk new_AGEMA_reg_buffer_2290 ( .C ( clk ), .D ( new_AGEMA_signal_13789 ), .Q ( new_AGEMA_signal_13790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2294 ( .C ( clk ), .D ( new_AGEMA_signal_13793 ), .Q ( new_AGEMA_signal_13794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2298 ( .C ( clk ), .D ( new_AGEMA_signal_13797 ), .Q ( new_AGEMA_signal_13798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2302 ( .C ( clk ), .D ( new_AGEMA_signal_13801 ), .Q ( new_AGEMA_signal_13802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2306 ( .C ( clk ), .D ( new_AGEMA_signal_13805 ), .Q ( new_AGEMA_signal_13806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2310 ( .C ( clk ), .D ( new_AGEMA_signal_13809 ), .Q ( new_AGEMA_signal_13810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2314 ( .C ( clk ), .D ( new_AGEMA_signal_13813 ), .Q ( new_AGEMA_signal_13814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2318 ( .C ( clk ), .D ( new_AGEMA_signal_13817 ), .Q ( new_AGEMA_signal_13818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2320 ( .C ( clk ), .D ( new_AGEMA_signal_13819 ), .Q ( new_AGEMA_signal_13820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2322 ( .C ( clk ), .D ( new_AGEMA_signal_13821 ), .Q ( new_AGEMA_signal_13822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2324 ( .C ( clk ), .D ( new_AGEMA_signal_13823 ), .Q ( new_AGEMA_signal_13824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2326 ( .C ( clk ), .D ( new_AGEMA_signal_13825 ), .Q ( new_AGEMA_signal_13826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2328 ( .C ( clk ), .D ( new_AGEMA_signal_13827 ), .Q ( new_AGEMA_signal_13828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2330 ( .C ( clk ), .D ( new_AGEMA_signal_13829 ), .Q ( new_AGEMA_signal_13830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2332 ( .C ( clk ), .D ( new_AGEMA_signal_13831 ), .Q ( new_AGEMA_signal_13832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2334 ( .C ( clk ), .D ( new_AGEMA_signal_13833 ), .Q ( new_AGEMA_signal_13834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2338 ( .C ( clk ), .D ( new_AGEMA_signal_13837 ), .Q ( new_AGEMA_signal_13838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2342 ( .C ( clk ), .D ( new_AGEMA_signal_13841 ), .Q ( new_AGEMA_signal_13842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2346 ( .C ( clk ), .D ( new_AGEMA_signal_13845 ), .Q ( new_AGEMA_signal_13846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2350 ( .C ( clk ), .D ( new_AGEMA_signal_13849 ), .Q ( new_AGEMA_signal_13850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2352 ( .C ( clk ), .D ( new_AGEMA_signal_13851 ), .Q ( new_AGEMA_signal_13852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2354 ( .C ( clk ), .D ( new_AGEMA_signal_13853 ), .Q ( new_AGEMA_signal_13854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2356 ( .C ( clk ), .D ( new_AGEMA_signal_13855 ), .Q ( new_AGEMA_signal_13856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2358 ( .C ( clk ), .D ( new_AGEMA_signal_13857 ), .Q ( new_AGEMA_signal_13858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2362 ( .C ( clk ), .D ( new_AGEMA_signal_13861 ), .Q ( new_AGEMA_signal_13862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2366 ( .C ( clk ), .D ( new_AGEMA_signal_13865 ), .Q ( new_AGEMA_signal_13866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2370 ( .C ( clk ), .D ( new_AGEMA_signal_13869 ), .Q ( new_AGEMA_signal_13870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2374 ( .C ( clk ), .D ( new_AGEMA_signal_13873 ), .Q ( new_AGEMA_signal_13874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2376 ( .C ( clk ), .D ( new_AGEMA_signal_13875 ), .Q ( new_AGEMA_signal_13876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2378 ( .C ( clk ), .D ( new_AGEMA_signal_13877 ), .Q ( new_AGEMA_signal_13878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2380 ( .C ( clk ), .D ( new_AGEMA_signal_13879 ), .Q ( new_AGEMA_signal_13880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2382 ( .C ( clk ), .D ( new_AGEMA_signal_13881 ), .Q ( new_AGEMA_signal_13882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2386 ( .C ( clk ), .D ( new_AGEMA_signal_13885 ), .Q ( new_AGEMA_signal_13886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2390 ( .C ( clk ), .D ( new_AGEMA_signal_13889 ), .Q ( new_AGEMA_signal_13890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2394 ( .C ( clk ), .D ( new_AGEMA_signal_13893 ), .Q ( new_AGEMA_signal_13894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2398 ( .C ( clk ), .D ( new_AGEMA_signal_13897 ), .Q ( new_AGEMA_signal_13898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2402 ( .C ( clk ), .D ( new_AGEMA_signal_13901 ), .Q ( new_AGEMA_signal_13902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2406 ( .C ( clk ), .D ( new_AGEMA_signal_13905 ), .Q ( new_AGEMA_signal_13906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2410 ( .C ( clk ), .D ( new_AGEMA_signal_13909 ), .Q ( new_AGEMA_signal_13910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2414 ( .C ( clk ), .D ( new_AGEMA_signal_13913 ), .Q ( new_AGEMA_signal_13914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2416 ( .C ( clk ), .D ( new_AGEMA_signal_13915 ), .Q ( new_AGEMA_signal_13916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2418 ( .C ( clk ), .D ( new_AGEMA_signal_13917 ), .Q ( new_AGEMA_signal_13918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2420 ( .C ( clk ), .D ( new_AGEMA_signal_13919 ), .Q ( new_AGEMA_signal_13920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2422 ( .C ( clk ), .D ( new_AGEMA_signal_13921 ), .Q ( new_AGEMA_signal_13922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2424 ( .C ( clk ), .D ( new_AGEMA_signal_13923 ), .Q ( new_AGEMA_signal_13924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2426 ( .C ( clk ), .D ( new_AGEMA_signal_13925 ), .Q ( new_AGEMA_signal_13926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2428 ( .C ( clk ), .D ( new_AGEMA_signal_13927 ), .Q ( new_AGEMA_signal_13928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2430 ( .C ( clk ), .D ( new_AGEMA_signal_13929 ), .Q ( new_AGEMA_signal_13930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2432 ( .C ( clk ), .D ( new_AGEMA_signal_13931 ), .Q ( new_AGEMA_signal_13932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2434 ( .C ( clk ), .D ( new_AGEMA_signal_13933 ), .Q ( new_AGEMA_signal_13934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2436 ( .C ( clk ), .D ( new_AGEMA_signal_13935 ), .Q ( new_AGEMA_signal_13936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2438 ( .C ( clk ), .D ( new_AGEMA_signal_13937 ), .Q ( new_AGEMA_signal_13938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2440 ( .C ( clk ), .D ( new_AGEMA_signal_13939 ), .Q ( new_AGEMA_signal_13940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2442 ( .C ( clk ), .D ( new_AGEMA_signal_13941 ), .Q ( new_AGEMA_signal_13942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2444 ( .C ( clk ), .D ( new_AGEMA_signal_13943 ), .Q ( new_AGEMA_signal_13944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2446 ( .C ( clk ), .D ( new_AGEMA_signal_13945 ), .Q ( new_AGEMA_signal_13946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2450 ( .C ( clk ), .D ( new_AGEMA_signal_13949 ), .Q ( new_AGEMA_signal_13950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2454 ( .C ( clk ), .D ( new_AGEMA_signal_13953 ), .Q ( new_AGEMA_signal_13954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2458 ( .C ( clk ), .D ( new_AGEMA_signal_13957 ), .Q ( new_AGEMA_signal_13958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2462 ( .C ( clk ), .D ( new_AGEMA_signal_13961 ), .Q ( new_AGEMA_signal_13962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2466 ( .C ( clk ), .D ( new_AGEMA_signal_13965 ), .Q ( new_AGEMA_signal_13966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2470 ( .C ( clk ), .D ( new_AGEMA_signal_13969 ), .Q ( new_AGEMA_signal_13970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2474 ( .C ( clk ), .D ( new_AGEMA_signal_13973 ), .Q ( new_AGEMA_signal_13974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2478 ( .C ( clk ), .D ( new_AGEMA_signal_13977 ), .Q ( new_AGEMA_signal_13978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2482 ( .C ( clk ), .D ( new_AGEMA_signal_13981 ), .Q ( new_AGEMA_signal_13982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2486 ( .C ( clk ), .D ( new_AGEMA_signal_13985 ), .Q ( new_AGEMA_signal_13986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2490 ( .C ( clk ), .D ( new_AGEMA_signal_13989 ), .Q ( new_AGEMA_signal_13990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2494 ( .C ( clk ), .D ( new_AGEMA_signal_13993 ), .Q ( new_AGEMA_signal_13994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2496 ( .C ( clk ), .D ( new_AGEMA_signal_13995 ), .Q ( new_AGEMA_signal_13996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2498 ( .C ( clk ), .D ( new_AGEMA_signal_13997 ), .Q ( new_AGEMA_signal_13998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2500 ( .C ( clk ), .D ( new_AGEMA_signal_13999 ), .Q ( new_AGEMA_signal_14000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2502 ( .C ( clk ), .D ( new_AGEMA_signal_14001 ), .Q ( new_AGEMA_signal_14002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2504 ( .C ( clk ), .D ( new_AGEMA_signal_14003 ), .Q ( new_AGEMA_signal_14004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2506 ( .C ( clk ), .D ( new_AGEMA_signal_14005 ), .Q ( new_AGEMA_signal_14006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2508 ( .C ( clk ), .D ( new_AGEMA_signal_14007 ), .Q ( new_AGEMA_signal_14008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2510 ( .C ( clk ), .D ( new_AGEMA_signal_14009 ), .Q ( new_AGEMA_signal_14010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2512 ( .C ( clk ), .D ( new_AGEMA_signal_14011 ), .Q ( new_AGEMA_signal_14012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2514 ( .C ( clk ), .D ( new_AGEMA_signal_14013 ), .Q ( new_AGEMA_signal_14014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2516 ( .C ( clk ), .D ( new_AGEMA_signal_14015 ), .Q ( new_AGEMA_signal_14016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2518 ( .C ( clk ), .D ( new_AGEMA_signal_14017 ), .Q ( new_AGEMA_signal_14018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2522 ( .C ( clk ), .D ( new_AGEMA_signal_14021 ), .Q ( new_AGEMA_signal_14022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2526 ( .C ( clk ), .D ( new_AGEMA_signal_14025 ), .Q ( new_AGEMA_signal_14026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2530 ( .C ( clk ), .D ( new_AGEMA_signal_14029 ), .Q ( new_AGEMA_signal_14030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2534 ( .C ( clk ), .D ( new_AGEMA_signal_14033 ), .Q ( new_AGEMA_signal_14034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2536 ( .C ( clk ), .D ( new_AGEMA_signal_14035 ), .Q ( new_AGEMA_signal_14036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2538 ( .C ( clk ), .D ( new_AGEMA_signal_14037 ), .Q ( new_AGEMA_signal_14038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2540 ( .C ( clk ), .D ( new_AGEMA_signal_14039 ), .Q ( new_AGEMA_signal_14040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2542 ( .C ( clk ), .D ( new_AGEMA_signal_14041 ), .Q ( new_AGEMA_signal_14042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2546 ( .C ( clk ), .D ( new_AGEMA_signal_14045 ), .Q ( new_AGEMA_signal_14046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2550 ( .C ( clk ), .D ( new_AGEMA_signal_14049 ), .Q ( new_AGEMA_signal_14050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2554 ( .C ( clk ), .D ( new_AGEMA_signal_14053 ), .Q ( new_AGEMA_signal_14054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2558 ( .C ( clk ), .D ( new_AGEMA_signal_14057 ), .Q ( new_AGEMA_signal_14058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2564 ( .C ( clk ), .D ( new_AGEMA_signal_14063 ), .Q ( new_AGEMA_signal_14064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2570 ( .C ( clk ), .D ( new_AGEMA_signal_14069 ), .Q ( new_AGEMA_signal_14070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2576 ( .C ( clk ), .D ( new_AGEMA_signal_14075 ), .Q ( new_AGEMA_signal_14076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2582 ( .C ( clk ), .D ( new_AGEMA_signal_14081 ), .Q ( new_AGEMA_signal_14082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2586 ( .C ( clk ), .D ( new_AGEMA_signal_14085 ), .Q ( new_AGEMA_signal_14086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2590 ( .C ( clk ), .D ( new_AGEMA_signal_14089 ), .Q ( new_AGEMA_signal_14090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2594 ( .C ( clk ), .D ( new_AGEMA_signal_14093 ), .Q ( new_AGEMA_signal_14094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2598 ( .C ( clk ), .D ( new_AGEMA_signal_14097 ), .Q ( new_AGEMA_signal_14098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2602 ( .C ( clk ), .D ( new_AGEMA_signal_14101 ), .Q ( new_AGEMA_signal_14102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2606 ( .C ( clk ), .D ( new_AGEMA_signal_14105 ), .Q ( new_AGEMA_signal_14106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2610 ( .C ( clk ), .D ( new_AGEMA_signal_14109 ), .Q ( new_AGEMA_signal_14110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2614 ( .C ( clk ), .D ( new_AGEMA_signal_14113 ), .Q ( new_AGEMA_signal_14114 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2616 ( .C ( clk ), .D ( new_AGEMA_signal_14115 ), .Q ( new_AGEMA_signal_14116 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2618 ( .C ( clk ), .D ( new_AGEMA_signal_14117 ), .Q ( new_AGEMA_signal_14118 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2620 ( .C ( clk ), .D ( new_AGEMA_signal_14119 ), .Q ( new_AGEMA_signal_14120 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2622 ( .C ( clk ), .D ( new_AGEMA_signal_14121 ), .Q ( new_AGEMA_signal_14122 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2624 ( .C ( clk ), .D ( new_AGEMA_signal_14123 ), .Q ( new_AGEMA_signal_14124 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2626 ( .C ( clk ), .D ( new_AGEMA_signal_14125 ), .Q ( new_AGEMA_signal_14126 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2628 ( .C ( clk ), .D ( new_AGEMA_signal_14127 ), .Q ( new_AGEMA_signal_14128 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2630 ( .C ( clk ), .D ( new_AGEMA_signal_14129 ), .Q ( new_AGEMA_signal_14130 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2632 ( .C ( clk ), .D ( new_AGEMA_signal_14131 ), .Q ( new_AGEMA_signal_14132 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2634 ( .C ( clk ), .D ( new_AGEMA_signal_14133 ), .Q ( new_AGEMA_signal_14134 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2636 ( .C ( clk ), .D ( new_AGEMA_signal_14135 ), .Q ( new_AGEMA_signal_14136 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2638 ( .C ( clk ), .D ( new_AGEMA_signal_14137 ), .Q ( new_AGEMA_signal_14138 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2640 ( .C ( clk ), .D ( new_AGEMA_signal_14139 ), .Q ( new_AGEMA_signal_14140 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2642 ( .C ( clk ), .D ( new_AGEMA_signal_14141 ), .Q ( new_AGEMA_signal_14142 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2644 ( .C ( clk ), .D ( new_AGEMA_signal_14143 ), .Q ( new_AGEMA_signal_14144 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2646 ( .C ( clk ), .D ( new_AGEMA_signal_14145 ), .Q ( new_AGEMA_signal_14146 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2650 ( .C ( clk ), .D ( new_AGEMA_signal_14149 ), .Q ( new_AGEMA_signal_14150 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2654 ( .C ( clk ), .D ( new_AGEMA_signal_14153 ), .Q ( new_AGEMA_signal_14154 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2658 ( .C ( clk ), .D ( new_AGEMA_signal_14157 ), .Q ( new_AGEMA_signal_14158 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2662 ( .C ( clk ), .D ( new_AGEMA_signal_14161 ), .Q ( new_AGEMA_signal_14162 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2668 ( .C ( clk ), .D ( new_AGEMA_signal_14167 ), .Q ( new_AGEMA_signal_14168 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2674 ( .C ( clk ), .D ( new_AGEMA_signal_14173 ), .Q ( new_AGEMA_signal_14174 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2680 ( .C ( clk ), .D ( new_AGEMA_signal_14179 ), .Q ( new_AGEMA_signal_14180 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2686 ( .C ( clk ), .D ( new_AGEMA_signal_14185 ), .Q ( new_AGEMA_signal_14186 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2690 ( .C ( clk ), .D ( new_AGEMA_signal_14189 ), .Q ( new_AGEMA_signal_14190 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2694 ( .C ( clk ), .D ( new_AGEMA_signal_14193 ), .Q ( new_AGEMA_signal_14194 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2698 ( .C ( clk ), .D ( new_AGEMA_signal_14197 ), .Q ( new_AGEMA_signal_14198 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2702 ( .C ( clk ), .D ( new_AGEMA_signal_14201 ), .Q ( new_AGEMA_signal_14202 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2704 ( .C ( clk ), .D ( new_AGEMA_signal_14203 ), .Q ( new_AGEMA_signal_14204 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2706 ( .C ( clk ), .D ( new_AGEMA_signal_14205 ), .Q ( new_AGEMA_signal_14206 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2708 ( .C ( clk ), .D ( new_AGEMA_signal_14207 ), .Q ( new_AGEMA_signal_14208 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2710 ( .C ( clk ), .D ( new_AGEMA_signal_14209 ), .Q ( new_AGEMA_signal_14210 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2712 ( .C ( clk ), .D ( new_AGEMA_signal_14211 ), .Q ( new_AGEMA_signal_14212 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2714 ( .C ( clk ), .D ( new_AGEMA_signal_14213 ), .Q ( new_AGEMA_signal_14214 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2716 ( .C ( clk ), .D ( new_AGEMA_signal_14215 ), .Q ( new_AGEMA_signal_14216 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2718 ( .C ( clk ), .D ( new_AGEMA_signal_14217 ), .Q ( new_AGEMA_signal_14218 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2720 ( .C ( clk ), .D ( new_AGEMA_signal_14219 ), .Q ( new_AGEMA_signal_14220 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2722 ( .C ( clk ), .D ( new_AGEMA_signal_14221 ), .Q ( new_AGEMA_signal_14222 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2724 ( .C ( clk ), .D ( new_AGEMA_signal_14223 ), .Q ( new_AGEMA_signal_14224 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2726 ( .C ( clk ), .D ( new_AGEMA_signal_14225 ), .Q ( new_AGEMA_signal_14226 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2730 ( .C ( clk ), .D ( new_AGEMA_signal_14229 ), .Q ( new_AGEMA_signal_14230 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2734 ( .C ( clk ), .D ( new_AGEMA_signal_14233 ), .Q ( new_AGEMA_signal_14234 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2738 ( .C ( clk ), .D ( new_AGEMA_signal_14237 ), .Q ( new_AGEMA_signal_14238 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2742 ( .C ( clk ), .D ( new_AGEMA_signal_14241 ), .Q ( new_AGEMA_signal_14242 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2744 ( .C ( clk ), .D ( new_AGEMA_signal_14243 ), .Q ( new_AGEMA_signal_14244 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2746 ( .C ( clk ), .D ( new_AGEMA_signal_14245 ), .Q ( new_AGEMA_signal_14246 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2748 ( .C ( clk ), .D ( new_AGEMA_signal_14247 ), .Q ( new_AGEMA_signal_14248 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2750 ( .C ( clk ), .D ( new_AGEMA_signal_14249 ), .Q ( new_AGEMA_signal_14250 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2752 ( .C ( clk ), .D ( new_AGEMA_signal_14251 ), .Q ( new_AGEMA_signal_14252 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2754 ( .C ( clk ), .D ( new_AGEMA_signal_14253 ), .Q ( new_AGEMA_signal_14254 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2756 ( .C ( clk ), .D ( new_AGEMA_signal_14255 ), .Q ( new_AGEMA_signal_14256 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2758 ( .C ( clk ), .D ( new_AGEMA_signal_14257 ), .Q ( new_AGEMA_signal_14258 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2762 ( .C ( clk ), .D ( new_AGEMA_signal_14261 ), .Q ( new_AGEMA_signal_14262 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2766 ( .C ( clk ), .D ( new_AGEMA_signal_14265 ), .Q ( new_AGEMA_signal_14266 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2770 ( .C ( clk ), .D ( new_AGEMA_signal_14269 ), .Q ( new_AGEMA_signal_14270 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2774 ( .C ( clk ), .D ( new_AGEMA_signal_14273 ), .Q ( new_AGEMA_signal_14274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2778 ( .C ( clk ), .D ( new_AGEMA_signal_14277 ), .Q ( new_AGEMA_signal_14278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2782 ( .C ( clk ), .D ( new_AGEMA_signal_14281 ), .Q ( new_AGEMA_signal_14282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2786 ( .C ( clk ), .D ( new_AGEMA_signal_14285 ), .Q ( new_AGEMA_signal_14286 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2790 ( .C ( clk ), .D ( new_AGEMA_signal_14289 ), .Q ( new_AGEMA_signal_14290 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2794 ( .C ( clk ), .D ( new_AGEMA_signal_14293 ), .Q ( new_AGEMA_signal_14294 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2798 ( .C ( clk ), .D ( new_AGEMA_signal_14297 ), .Q ( new_AGEMA_signal_14298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2802 ( .C ( clk ), .D ( new_AGEMA_signal_14301 ), .Q ( new_AGEMA_signal_14302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2806 ( .C ( clk ), .D ( new_AGEMA_signal_14305 ), .Q ( new_AGEMA_signal_14306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2810 ( .C ( clk ), .D ( new_AGEMA_signal_14309 ), .Q ( new_AGEMA_signal_14310 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2814 ( .C ( clk ), .D ( new_AGEMA_signal_14313 ), .Q ( new_AGEMA_signal_14314 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2818 ( .C ( clk ), .D ( new_AGEMA_signal_14317 ), .Q ( new_AGEMA_signal_14318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2822 ( .C ( clk ), .D ( new_AGEMA_signal_14321 ), .Q ( new_AGEMA_signal_14322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2826 ( .C ( clk ), .D ( new_AGEMA_signal_14325 ), .Q ( new_AGEMA_signal_14326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2830 ( .C ( clk ), .D ( new_AGEMA_signal_14329 ), .Q ( new_AGEMA_signal_14330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2834 ( .C ( clk ), .D ( new_AGEMA_signal_14333 ), .Q ( new_AGEMA_signal_14334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2838 ( .C ( clk ), .D ( new_AGEMA_signal_14337 ), .Q ( new_AGEMA_signal_14338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2840 ( .C ( clk ), .D ( new_AGEMA_signal_14339 ), .Q ( new_AGEMA_signal_14340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2842 ( .C ( clk ), .D ( new_AGEMA_signal_14341 ), .Q ( new_AGEMA_signal_14342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2844 ( .C ( clk ), .D ( new_AGEMA_signal_14343 ), .Q ( new_AGEMA_signal_14344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2846 ( .C ( clk ), .D ( new_AGEMA_signal_14345 ), .Q ( new_AGEMA_signal_14346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2848 ( .C ( clk ), .D ( new_AGEMA_signal_14347 ), .Q ( new_AGEMA_signal_14348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2850 ( .C ( clk ), .D ( new_AGEMA_signal_14349 ), .Q ( new_AGEMA_signal_14350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2852 ( .C ( clk ), .D ( new_AGEMA_signal_14351 ), .Q ( new_AGEMA_signal_14352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2854 ( .C ( clk ), .D ( new_AGEMA_signal_14353 ), .Q ( new_AGEMA_signal_14354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2856 ( .C ( clk ), .D ( new_AGEMA_signal_14355 ), .Q ( new_AGEMA_signal_14356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2858 ( .C ( clk ), .D ( new_AGEMA_signal_14357 ), .Q ( new_AGEMA_signal_14358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2860 ( .C ( clk ), .D ( new_AGEMA_signal_14359 ), .Q ( new_AGEMA_signal_14360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2862 ( .C ( clk ), .D ( new_AGEMA_signal_14361 ), .Q ( new_AGEMA_signal_14362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2864 ( .C ( clk ), .D ( new_AGEMA_signal_14363 ), .Q ( new_AGEMA_signal_14364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2866 ( .C ( clk ), .D ( new_AGEMA_signal_14365 ), .Q ( new_AGEMA_signal_14366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2868 ( .C ( clk ), .D ( new_AGEMA_signal_14367 ), .Q ( new_AGEMA_signal_14368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2870 ( .C ( clk ), .D ( new_AGEMA_signal_14369 ), .Q ( new_AGEMA_signal_14370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2874 ( .C ( clk ), .D ( new_AGEMA_signal_14373 ), .Q ( new_AGEMA_signal_14374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2878 ( .C ( clk ), .D ( new_AGEMA_signal_14377 ), .Q ( new_AGEMA_signal_14378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2882 ( .C ( clk ), .D ( new_AGEMA_signal_14381 ), .Q ( new_AGEMA_signal_14382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2886 ( .C ( clk ), .D ( new_AGEMA_signal_14385 ), .Q ( new_AGEMA_signal_14386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2890 ( .C ( clk ), .D ( new_AGEMA_signal_14389 ), .Q ( new_AGEMA_signal_14390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2894 ( .C ( clk ), .D ( new_AGEMA_signal_14393 ), .Q ( new_AGEMA_signal_14394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2898 ( .C ( clk ), .D ( new_AGEMA_signal_14397 ), .Q ( new_AGEMA_signal_14398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2902 ( .C ( clk ), .D ( new_AGEMA_signal_14401 ), .Q ( new_AGEMA_signal_14402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2904 ( .C ( clk ), .D ( new_AGEMA_signal_14403 ), .Q ( new_AGEMA_signal_14404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2906 ( .C ( clk ), .D ( new_AGEMA_signal_14405 ), .Q ( new_AGEMA_signal_14406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2908 ( .C ( clk ), .D ( new_AGEMA_signal_14407 ), .Q ( new_AGEMA_signal_14408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2910 ( .C ( clk ), .D ( new_AGEMA_signal_14409 ), .Q ( new_AGEMA_signal_14410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2912 ( .C ( clk ), .D ( new_AGEMA_signal_14411 ), .Q ( new_AGEMA_signal_14412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2914 ( .C ( clk ), .D ( new_AGEMA_signal_14413 ), .Q ( new_AGEMA_signal_14414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2916 ( .C ( clk ), .D ( new_AGEMA_signal_14415 ), .Q ( new_AGEMA_signal_14416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2918 ( .C ( clk ), .D ( new_AGEMA_signal_14417 ), .Q ( new_AGEMA_signal_14418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2920 ( .C ( clk ), .D ( new_AGEMA_signal_14419 ), .Q ( new_AGEMA_signal_14420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2922 ( .C ( clk ), .D ( new_AGEMA_signal_14421 ), .Q ( new_AGEMA_signal_14422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2924 ( .C ( clk ), .D ( new_AGEMA_signal_14423 ), .Q ( new_AGEMA_signal_14424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2926 ( .C ( clk ), .D ( new_AGEMA_signal_14425 ), .Q ( new_AGEMA_signal_14426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2928 ( .C ( clk ), .D ( new_AGEMA_signal_14427 ), .Q ( new_AGEMA_signal_14428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2930 ( .C ( clk ), .D ( new_AGEMA_signal_14429 ), .Q ( new_AGEMA_signal_14430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2932 ( .C ( clk ), .D ( new_AGEMA_signal_14431 ), .Q ( new_AGEMA_signal_14432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2934 ( .C ( clk ), .D ( new_AGEMA_signal_14433 ), .Q ( new_AGEMA_signal_14434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2936 ( .C ( clk ), .D ( new_AGEMA_signal_14435 ), .Q ( new_AGEMA_signal_14436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2938 ( .C ( clk ), .D ( new_AGEMA_signal_14437 ), .Q ( new_AGEMA_signal_14438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2940 ( .C ( clk ), .D ( new_AGEMA_signal_14439 ), .Q ( new_AGEMA_signal_14440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2942 ( .C ( clk ), .D ( new_AGEMA_signal_14441 ), .Q ( new_AGEMA_signal_14442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2944 ( .C ( clk ), .D ( new_AGEMA_signal_14443 ), .Q ( new_AGEMA_signal_14444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2946 ( .C ( clk ), .D ( new_AGEMA_signal_14445 ), .Q ( new_AGEMA_signal_14446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2948 ( .C ( clk ), .D ( new_AGEMA_signal_14447 ), .Q ( new_AGEMA_signal_14448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2950 ( .C ( clk ), .D ( new_AGEMA_signal_14449 ), .Q ( new_AGEMA_signal_14450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2952 ( .C ( clk ), .D ( new_AGEMA_signal_14451 ), .Q ( new_AGEMA_signal_14452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2954 ( .C ( clk ), .D ( new_AGEMA_signal_14453 ), .Q ( new_AGEMA_signal_14454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2956 ( .C ( clk ), .D ( new_AGEMA_signal_14455 ), .Q ( new_AGEMA_signal_14456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2958 ( .C ( clk ), .D ( new_AGEMA_signal_14457 ), .Q ( new_AGEMA_signal_14458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2960 ( .C ( clk ), .D ( new_AGEMA_signal_14459 ), .Q ( new_AGEMA_signal_14460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2962 ( .C ( clk ), .D ( new_AGEMA_signal_14461 ), .Q ( new_AGEMA_signal_14462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2964 ( .C ( clk ), .D ( new_AGEMA_signal_14463 ), .Q ( new_AGEMA_signal_14464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2966 ( .C ( clk ), .D ( new_AGEMA_signal_14465 ), .Q ( new_AGEMA_signal_14466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2968 ( .C ( clk ), .D ( new_AGEMA_signal_14467 ), .Q ( new_AGEMA_signal_14468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2970 ( .C ( clk ), .D ( new_AGEMA_signal_14469 ), .Q ( new_AGEMA_signal_14470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2972 ( .C ( clk ), .D ( new_AGEMA_signal_14471 ), .Q ( new_AGEMA_signal_14472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2974 ( .C ( clk ), .D ( new_AGEMA_signal_14473 ), .Q ( new_AGEMA_signal_14474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2978 ( .C ( clk ), .D ( new_AGEMA_signal_14477 ), .Q ( new_AGEMA_signal_14478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2982 ( .C ( clk ), .D ( new_AGEMA_signal_14481 ), .Q ( new_AGEMA_signal_14482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2986 ( .C ( clk ), .D ( new_AGEMA_signal_14485 ), .Q ( new_AGEMA_signal_14486 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2990 ( .C ( clk ), .D ( new_AGEMA_signal_14489 ), .Q ( new_AGEMA_signal_14490 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2992 ( .C ( clk ), .D ( new_AGEMA_signal_14491 ), .Q ( new_AGEMA_signal_14492 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2994 ( .C ( clk ), .D ( new_AGEMA_signal_14493 ), .Q ( new_AGEMA_signal_14494 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2996 ( .C ( clk ), .D ( new_AGEMA_signal_14495 ), .Q ( new_AGEMA_signal_14496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2998 ( .C ( clk ), .D ( new_AGEMA_signal_14497 ), .Q ( new_AGEMA_signal_14498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3000 ( .C ( clk ), .D ( new_AGEMA_signal_14499 ), .Q ( new_AGEMA_signal_14500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3002 ( .C ( clk ), .D ( new_AGEMA_signal_14501 ), .Q ( new_AGEMA_signal_14502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3004 ( .C ( clk ), .D ( new_AGEMA_signal_14503 ), .Q ( new_AGEMA_signal_14504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3006 ( .C ( clk ), .D ( new_AGEMA_signal_14505 ), .Q ( new_AGEMA_signal_14506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3008 ( .C ( clk ), .D ( new_AGEMA_signal_14507 ), .Q ( new_AGEMA_signal_14508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3010 ( .C ( clk ), .D ( new_AGEMA_signal_14509 ), .Q ( new_AGEMA_signal_14510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3012 ( .C ( clk ), .D ( new_AGEMA_signal_14511 ), .Q ( new_AGEMA_signal_14512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3014 ( .C ( clk ), .D ( new_AGEMA_signal_14513 ), .Q ( new_AGEMA_signal_14514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3016 ( .C ( clk ), .D ( new_AGEMA_signal_14515 ), .Q ( new_AGEMA_signal_14516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3018 ( .C ( clk ), .D ( new_AGEMA_signal_14517 ), .Q ( new_AGEMA_signal_14518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3020 ( .C ( clk ), .D ( new_AGEMA_signal_14519 ), .Q ( new_AGEMA_signal_14520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3022 ( .C ( clk ), .D ( new_AGEMA_signal_14521 ), .Q ( new_AGEMA_signal_14522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3024 ( .C ( clk ), .D ( new_AGEMA_signal_14523 ), .Q ( new_AGEMA_signal_14524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3026 ( .C ( clk ), .D ( new_AGEMA_signal_14525 ), .Q ( new_AGEMA_signal_14526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3028 ( .C ( clk ), .D ( new_AGEMA_signal_14527 ), .Q ( new_AGEMA_signal_14528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3030 ( .C ( clk ), .D ( new_AGEMA_signal_14529 ), .Q ( new_AGEMA_signal_14530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3034 ( .C ( clk ), .D ( new_AGEMA_signal_14533 ), .Q ( new_AGEMA_signal_14534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3038 ( .C ( clk ), .D ( new_AGEMA_signal_14537 ), .Q ( new_AGEMA_signal_14538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3042 ( .C ( clk ), .D ( new_AGEMA_signal_14541 ), .Q ( new_AGEMA_signal_14542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3046 ( .C ( clk ), .D ( new_AGEMA_signal_14545 ), .Q ( new_AGEMA_signal_14546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3050 ( .C ( clk ), .D ( new_AGEMA_signal_14549 ), .Q ( new_AGEMA_signal_14550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3054 ( .C ( clk ), .D ( new_AGEMA_signal_14553 ), .Q ( new_AGEMA_signal_14554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3058 ( .C ( clk ), .D ( new_AGEMA_signal_14557 ), .Q ( new_AGEMA_signal_14558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3062 ( .C ( clk ), .D ( new_AGEMA_signal_14561 ), .Q ( new_AGEMA_signal_14562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3066 ( .C ( clk ), .D ( new_AGEMA_signal_14565 ), .Q ( new_AGEMA_signal_14566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3070 ( .C ( clk ), .D ( new_AGEMA_signal_14569 ), .Q ( new_AGEMA_signal_14570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3074 ( .C ( clk ), .D ( new_AGEMA_signal_14573 ), .Q ( new_AGEMA_signal_14574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3078 ( .C ( clk ), .D ( new_AGEMA_signal_14577 ), .Q ( new_AGEMA_signal_14578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3082 ( .C ( clk ), .D ( new_AGEMA_signal_14581 ), .Q ( new_AGEMA_signal_14582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3086 ( .C ( clk ), .D ( new_AGEMA_signal_14585 ), .Q ( new_AGEMA_signal_14586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3090 ( .C ( clk ), .D ( new_AGEMA_signal_14589 ), .Q ( new_AGEMA_signal_14590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3094 ( .C ( clk ), .D ( new_AGEMA_signal_14593 ), .Q ( new_AGEMA_signal_14594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3096 ( .C ( clk ), .D ( new_AGEMA_signal_14595 ), .Q ( new_AGEMA_signal_14596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3100 ( .C ( clk ), .D ( new_AGEMA_signal_14599 ), .Q ( new_AGEMA_signal_14600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3104 ( .C ( clk ), .D ( new_AGEMA_signal_14603 ), .Q ( new_AGEMA_signal_14604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3108 ( .C ( clk ), .D ( new_AGEMA_signal_14607 ), .Q ( new_AGEMA_signal_14608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3112 ( .C ( clk ), .D ( new_AGEMA_signal_14611 ), .Q ( new_AGEMA_signal_14612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3116 ( .C ( clk ), .D ( new_AGEMA_signal_14615 ), .Q ( new_AGEMA_signal_14616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3120 ( .C ( clk ), .D ( new_AGEMA_signal_14619 ), .Q ( new_AGEMA_signal_14620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3124 ( .C ( clk ), .D ( new_AGEMA_signal_14623 ), .Q ( new_AGEMA_signal_14624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3132 ( .C ( clk ), .D ( new_AGEMA_signal_14631 ), .Q ( new_AGEMA_signal_14632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3140 ( .C ( clk ), .D ( new_AGEMA_signal_14639 ), .Q ( new_AGEMA_signal_14640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3148 ( .C ( clk ), .D ( new_AGEMA_signal_14647 ), .Q ( new_AGEMA_signal_14648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3156 ( .C ( clk ), .D ( new_AGEMA_signal_14655 ), .Q ( new_AGEMA_signal_14656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3172 ( .C ( clk ), .D ( new_AGEMA_signal_14671 ), .Q ( new_AGEMA_signal_14672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3180 ( .C ( clk ), .D ( new_AGEMA_signal_14679 ), .Q ( new_AGEMA_signal_14680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3188 ( .C ( clk ), .D ( new_AGEMA_signal_14687 ), .Q ( new_AGEMA_signal_14688 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3196 ( .C ( clk ), .D ( new_AGEMA_signal_14695 ), .Q ( new_AGEMA_signal_14696 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3202 ( .C ( clk ), .D ( new_AGEMA_signal_14701 ), .Q ( new_AGEMA_signal_14702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3208 ( .C ( clk ), .D ( new_AGEMA_signal_14707 ), .Q ( new_AGEMA_signal_14708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3214 ( .C ( clk ), .D ( new_AGEMA_signal_14713 ), .Q ( new_AGEMA_signal_14714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3220 ( .C ( clk ), .D ( new_AGEMA_signal_14719 ), .Q ( new_AGEMA_signal_14720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3224 ( .C ( clk ), .D ( new_AGEMA_signal_14723 ), .Q ( new_AGEMA_signal_14724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3228 ( .C ( clk ), .D ( new_AGEMA_signal_14727 ), .Q ( new_AGEMA_signal_14728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3232 ( .C ( clk ), .D ( new_AGEMA_signal_14731 ), .Q ( new_AGEMA_signal_14732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3236 ( .C ( clk ), .D ( new_AGEMA_signal_14735 ), .Q ( new_AGEMA_signal_14736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3242 ( .C ( clk ), .D ( new_AGEMA_signal_14741 ), .Q ( new_AGEMA_signal_14742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3248 ( .C ( clk ), .D ( new_AGEMA_signal_14747 ), .Q ( new_AGEMA_signal_14748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3254 ( .C ( clk ), .D ( new_AGEMA_signal_14753 ), .Q ( new_AGEMA_signal_14754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3260 ( .C ( clk ), .D ( new_AGEMA_signal_14759 ), .Q ( new_AGEMA_signal_14760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3274 ( .C ( clk ), .D ( new_AGEMA_signal_14773 ), .Q ( new_AGEMA_signal_14774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3280 ( .C ( clk ), .D ( new_AGEMA_signal_14779 ), .Q ( new_AGEMA_signal_14780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3286 ( .C ( clk ), .D ( new_AGEMA_signal_14785 ), .Q ( new_AGEMA_signal_14786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3292 ( .C ( clk ), .D ( new_AGEMA_signal_14791 ), .Q ( new_AGEMA_signal_14792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3298 ( .C ( clk ), .D ( new_AGEMA_signal_14797 ), .Q ( new_AGEMA_signal_14798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3304 ( .C ( clk ), .D ( new_AGEMA_signal_14803 ), .Q ( new_AGEMA_signal_14804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3310 ( .C ( clk ), .D ( new_AGEMA_signal_14809 ), .Q ( new_AGEMA_signal_14810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3316 ( .C ( clk ), .D ( new_AGEMA_signal_14815 ), .Q ( new_AGEMA_signal_14816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3328 ( .C ( clk ), .D ( new_AGEMA_signal_14827 ), .Q ( new_AGEMA_signal_14828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3332 ( .C ( clk ), .D ( new_AGEMA_signal_14831 ), .Q ( new_AGEMA_signal_14832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3336 ( .C ( clk ), .D ( new_AGEMA_signal_14835 ), .Q ( new_AGEMA_signal_14836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3340 ( .C ( clk ), .D ( new_AGEMA_signal_14839 ), .Q ( new_AGEMA_signal_14840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3346 ( .C ( clk ), .D ( new_AGEMA_signal_14845 ), .Q ( new_AGEMA_signal_14846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3352 ( .C ( clk ), .D ( new_AGEMA_signal_14851 ), .Q ( new_AGEMA_signal_14852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3358 ( .C ( clk ), .D ( new_AGEMA_signal_14857 ), .Q ( new_AGEMA_signal_14858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3364 ( .C ( clk ), .D ( new_AGEMA_signal_14863 ), .Q ( new_AGEMA_signal_14864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3370 ( .C ( clk ), .D ( new_AGEMA_signal_14869 ), .Q ( new_AGEMA_signal_14870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3376 ( .C ( clk ), .D ( new_AGEMA_signal_14875 ), .Q ( new_AGEMA_signal_14876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3382 ( .C ( clk ), .D ( new_AGEMA_signal_14881 ), .Q ( new_AGEMA_signal_14882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3388 ( .C ( clk ), .D ( new_AGEMA_signal_14887 ), .Q ( new_AGEMA_signal_14888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3402 ( .C ( clk ), .D ( new_AGEMA_signal_14901 ), .Q ( new_AGEMA_signal_14902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3408 ( .C ( clk ), .D ( new_AGEMA_signal_14907 ), .Q ( new_AGEMA_signal_14908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3414 ( .C ( clk ), .D ( new_AGEMA_signal_14913 ), .Q ( new_AGEMA_signal_14914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3420 ( .C ( clk ), .D ( new_AGEMA_signal_14919 ), .Q ( new_AGEMA_signal_14920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3432 ( .C ( clk ), .D ( new_AGEMA_signal_14931 ), .Q ( new_AGEMA_signal_14932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3436 ( .C ( clk ), .D ( new_AGEMA_signal_14935 ), .Q ( new_AGEMA_signal_14936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3440 ( .C ( clk ), .D ( new_AGEMA_signal_14939 ), .Q ( new_AGEMA_signal_14940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3444 ( .C ( clk ), .D ( new_AGEMA_signal_14943 ), .Q ( new_AGEMA_signal_14944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3448 ( .C ( clk ), .D ( new_AGEMA_signal_14947 ), .Q ( new_AGEMA_signal_14948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3452 ( .C ( clk ), .D ( new_AGEMA_signal_14951 ), .Q ( new_AGEMA_signal_14952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3456 ( .C ( clk ), .D ( new_AGEMA_signal_14955 ), .Q ( new_AGEMA_signal_14956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3460 ( .C ( clk ), .D ( new_AGEMA_signal_14959 ), .Q ( new_AGEMA_signal_14960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3476 ( .C ( clk ), .D ( new_AGEMA_signal_14975 ), .Q ( new_AGEMA_signal_14976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3484 ( .C ( clk ), .D ( new_AGEMA_signal_14983 ), .Q ( new_AGEMA_signal_14984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3492 ( .C ( clk ), .D ( new_AGEMA_signal_14991 ), .Q ( new_AGEMA_signal_14992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3500 ( .C ( clk ), .D ( new_AGEMA_signal_14999 ), .Q ( new_AGEMA_signal_15000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3506 ( .C ( clk ), .D ( new_AGEMA_signal_15005 ), .Q ( new_AGEMA_signal_15006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3512 ( .C ( clk ), .D ( new_AGEMA_signal_15011 ), .Q ( new_AGEMA_signal_15012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3518 ( .C ( clk ), .D ( new_AGEMA_signal_15017 ), .Q ( new_AGEMA_signal_15018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3524 ( .C ( clk ), .D ( new_AGEMA_signal_15023 ), .Q ( new_AGEMA_signal_15024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3528 ( .C ( clk ), .D ( new_AGEMA_signal_15027 ), .Q ( new_AGEMA_signal_15028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3532 ( .C ( clk ), .D ( new_AGEMA_signal_15031 ), .Q ( new_AGEMA_signal_15032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3536 ( .C ( clk ), .D ( new_AGEMA_signal_15035 ), .Q ( new_AGEMA_signal_15036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3540 ( .C ( clk ), .D ( new_AGEMA_signal_15039 ), .Q ( new_AGEMA_signal_15040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3544 ( .C ( clk ), .D ( new_AGEMA_signal_15043 ), .Q ( new_AGEMA_signal_15044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3548 ( .C ( clk ), .D ( new_AGEMA_signal_15047 ), .Q ( new_AGEMA_signal_15048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3552 ( .C ( clk ), .D ( new_AGEMA_signal_15051 ), .Q ( new_AGEMA_signal_15052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3556 ( .C ( clk ), .D ( new_AGEMA_signal_15055 ), .Q ( new_AGEMA_signal_15056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3576 ( .C ( clk ), .D ( new_AGEMA_signal_15075 ), .Q ( new_AGEMA_signal_15076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3580 ( .C ( clk ), .D ( new_AGEMA_signal_15079 ), .Q ( new_AGEMA_signal_15080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3584 ( .C ( clk ), .D ( new_AGEMA_signal_15083 ), .Q ( new_AGEMA_signal_15084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3588 ( .C ( clk ), .D ( new_AGEMA_signal_15087 ), .Q ( new_AGEMA_signal_15088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3592 ( .C ( clk ), .D ( new_AGEMA_signal_15091 ), .Q ( new_AGEMA_signal_15092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3596 ( .C ( clk ), .D ( new_AGEMA_signal_15095 ), .Q ( new_AGEMA_signal_15096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3600 ( .C ( clk ), .D ( new_AGEMA_signal_15099 ), .Q ( new_AGEMA_signal_15100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3604 ( .C ( clk ), .D ( new_AGEMA_signal_15103 ), .Q ( new_AGEMA_signal_15104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3618 ( .C ( clk ), .D ( new_AGEMA_signal_15117 ), .Q ( new_AGEMA_signal_15118 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3624 ( .C ( clk ), .D ( new_AGEMA_signal_15123 ), .Q ( new_AGEMA_signal_15124 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3630 ( .C ( clk ), .D ( new_AGEMA_signal_15129 ), .Q ( new_AGEMA_signal_15130 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3636 ( .C ( clk ), .D ( new_AGEMA_signal_15135 ), .Q ( new_AGEMA_signal_15136 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3640 ( .C ( clk ), .D ( new_AGEMA_signal_15139 ), .Q ( new_AGEMA_signal_15140 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3644 ( .C ( clk ), .D ( new_AGEMA_signal_15143 ), .Q ( new_AGEMA_signal_15144 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3648 ( .C ( clk ), .D ( new_AGEMA_signal_15147 ), .Q ( new_AGEMA_signal_15148 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3652 ( .C ( clk ), .D ( new_AGEMA_signal_15151 ), .Q ( new_AGEMA_signal_15152 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3664 ( .C ( clk ), .D ( new_AGEMA_signal_15163 ), .Q ( new_AGEMA_signal_15164 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3668 ( .C ( clk ), .D ( new_AGEMA_signal_15167 ), .Q ( new_AGEMA_signal_15168 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3672 ( .C ( clk ), .D ( new_AGEMA_signal_15171 ), .Q ( new_AGEMA_signal_15172 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3676 ( .C ( clk ), .D ( new_AGEMA_signal_15175 ), .Q ( new_AGEMA_signal_15176 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3680 ( .C ( clk ), .D ( new_AGEMA_signal_15179 ), .Q ( new_AGEMA_signal_15180 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3684 ( .C ( clk ), .D ( new_AGEMA_signal_15183 ), .Q ( new_AGEMA_signal_15184 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3688 ( .C ( clk ), .D ( new_AGEMA_signal_15187 ), .Q ( new_AGEMA_signal_15188 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3692 ( .C ( clk ), .D ( new_AGEMA_signal_15191 ), .Q ( new_AGEMA_signal_15192 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3696 ( .C ( clk ), .D ( new_AGEMA_signal_15195 ), .Q ( new_AGEMA_signal_15196 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3700 ( .C ( clk ), .D ( new_AGEMA_signal_15199 ), .Q ( new_AGEMA_signal_15200 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3704 ( .C ( clk ), .D ( new_AGEMA_signal_15203 ), .Q ( new_AGEMA_signal_15204 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3708 ( .C ( clk ), .D ( new_AGEMA_signal_15207 ), .Q ( new_AGEMA_signal_15208 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3720 ( .C ( clk ), .D ( new_AGEMA_signal_15219 ), .Q ( new_AGEMA_signal_15220 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3724 ( .C ( clk ), .D ( new_AGEMA_signal_15223 ), .Q ( new_AGEMA_signal_15224 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3728 ( .C ( clk ), .D ( new_AGEMA_signal_15227 ), .Q ( new_AGEMA_signal_15228 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3732 ( .C ( clk ), .D ( new_AGEMA_signal_15231 ), .Q ( new_AGEMA_signal_15232 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3746 ( .C ( clk ), .D ( new_AGEMA_signal_15245 ), .Q ( new_AGEMA_signal_15246 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3752 ( .C ( clk ), .D ( new_AGEMA_signal_15251 ), .Q ( new_AGEMA_signal_15252 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3758 ( .C ( clk ), .D ( new_AGEMA_signal_15257 ), .Q ( new_AGEMA_signal_15258 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3764 ( .C ( clk ), .D ( new_AGEMA_signal_15263 ), .Q ( new_AGEMA_signal_15264 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3770 ( .C ( clk ), .D ( new_AGEMA_signal_15269 ), .Q ( new_AGEMA_signal_15270 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3776 ( .C ( clk ), .D ( new_AGEMA_signal_15275 ), .Q ( new_AGEMA_signal_15276 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3782 ( .C ( clk ), .D ( new_AGEMA_signal_15281 ), .Q ( new_AGEMA_signal_15282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3788 ( .C ( clk ), .D ( new_AGEMA_signal_15287 ), .Q ( new_AGEMA_signal_15288 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3792 ( .C ( clk ), .D ( new_AGEMA_signal_15291 ), .Q ( new_AGEMA_signal_15292 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3796 ( .C ( clk ), .D ( new_AGEMA_signal_15295 ), .Q ( new_AGEMA_signal_15296 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3800 ( .C ( clk ), .D ( new_AGEMA_signal_15299 ), .Q ( new_AGEMA_signal_15300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3804 ( .C ( clk ), .D ( new_AGEMA_signal_15303 ), .Q ( new_AGEMA_signal_15304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3820 ( .C ( clk ), .D ( new_AGEMA_signal_15319 ), .Q ( new_AGEMA_signal_15320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3828 ( .C ( clk ), .D ( new_AGEMA_signal_15327 ), .Q ( new_AGEMA_signal_15328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3836 ( .C ( clk ), .D ( new_AGEMA_signal_15335 ), .Q ( new_AGEMA_signal_15336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3844 ( .C ( clk ), .D ( new_AGEMA_signal_15343 ), .Q ( new_AGEMA_signal_15344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3856 ( .C ( clk ), .D ( new_AGEMA_signal_15355 ), .Q ( new_AGEMA_signal_15356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3860 ( .C ( clk ), .D ( new_AGEMA_signal_15359 ), .Q ( new_AGEMA_signal_15360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3864 ( .C ( clk ), .D ( new_AGEMA_signal_15363 ), .Q ( new_AGEMA_signal_15364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3868 ( .C ( clk ), .D ( new_AGEMA_signal_15367 ), .Q ( new_AGEMA_signal_15368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3872 ( .C ( clk ), .D ( new_AGEMA_signal_15371 ), .Q ( new_AGEMA_signal_15372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3876 ( .C ( clk ), .D ( new_AGEMA_signal_15375 ), .Q ( new_AGEMA_signal_15376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3880 ( .C ( clk ), .D ( new_AGEMA_signal_15379 ), .Q ( new_AGEMA_signal_15380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3884 ( .C ( clk ), .D ( new_AGEMA_signal_15383 ), .Q ( new_AGEMA_signal_15384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3888 ( .C ( clk ), .D ( new_AGEMA_signal_15387 ), .Q ( new_AGEMA_signal_15388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3892 ( .C ( clk ), .D ( new_AGEMA_signal_15391 ), .Q ( new_AGEMA_signal_15392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3896 ( .C ( clk ), .D ( new_AGEMA_signal_15395 ), .Q ( new_AGEMA_signal_15396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3900 ( .C ( clk ), .D ( new_AGEMA_signal_15399 ), .Q ( new_AGEMA_signal_15400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3904 ( .C ( clk ), .D ( new_AGEMA_signal_15403 ), .Q ( new_AGEMA_signal_15404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3908 ( .C ( clk ), .D ( new_AGEMA_signal_15407 ), .Q ( new_AGEMA_signal_15408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3912 ( .C ( clk ), .D ( new_AGEMA_signal_15411 ), .Q ( new_AGEMA_signal_15412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3916 ( .C ( clk ), .D ( new_AGEMA_signal_15415 ), .Q ( new_AGEMA_signal_15416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3920 ( .C ( clk ), .D ( new_AGEMA_signal_15419 ), .Q ( new_AGEMA_signal_15420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3924 ( .C ( clk ), .D ( new_AGEMA_signal_15423 ), .Q ( new_AGEMA_signal_15424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3928 ( .C ( clk ), .D ( new_AGEMA_signal_15427 ), .Q ( new_AGEMA_signal_15428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3932 ( .C ( clk ), .D ( new_AGEMA_signal_15431 ), .Q ( new_AGEMA_signal_15432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3940 ( .C ( clk ), .D ( new_AGEMA_signal_15439 ), .Q ( new_AGEMA_signal_15440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3948 ( .C ( clk ), .D ( new_AGEMA_signal_15447 ), .Q ( new_AGEMA_signal_15448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3956 ( .C ( clk ), .D ( new_AGEMA_signal_15455 ), .Q ( new_AGEMA_signal_15456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3964 ( .C ( clk ), .D ( new_AGEMA_signal_15463 ), .Q ( new_AGEMA_signal_15464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3976 ( .C ( clk ), .D ( new_AGEMA_signal_15475 ), .Q ( new_AGEMA_signal_15476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3980 ( .C ( clk ), .D ( new_AGEMA_signal_15479 ), .Q ( new_AGEMA_signal_15480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3984 ( .C ( clk ), .D ( new_AGEMA_signal_15483 ), .Q ( new_AGEMA_signal_15484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3988 ( .C ( clk ), .D ( new_AGEMA_signal_15487 ), .Q ( new_AGEMA_signal_15488 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4002 ( .C ( clk ), .D ( new_AGEMA_signal_15501 ), .Q ( new_AGEMA_signal_15502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4008 ( .C ( clk ), .D ( new_AGEMA_signal_15507 ), .Q ( new_AGEMA_signal_15508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4014 ( .C ( clk ), .D ( new_AGEMA_signal_15513 ), .Q ( new_AGEMA_signal_15514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4020 ( .C ( clk ), .D ( new_AGEMA_signal_15519 ), .Q ( new_AGEMA_signal_15520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4034 ( .C ( clk ), .D ( new_AGEMA_signal_15533 ), .Q ( new_AGEMA_signal_15534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4042 ( .C ( clk ), .D ( new_AGEMA_signal_15541 ), .Q ( new_AGEMA_signal_15542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4050 ( .C ( clk ), .D ( new_AGEMA_signal_15549 ), .Q ( new_AGEMA_signal_15550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4058 ( .C ( clk ), .D ( new_AGEMA_signal_15557 ), .Q ( new_AGEMA_signal_15558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4090 ( .C ( clk ), .D ( new_AGEMA_signal_15589 ), .Q ( new_AGEMA_signal_15590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4098 ( .C ( clk ), .D ( new_AGEMA_signal_15597 ), .Q ( new_AGEMA_signal_15598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4106 ( .C ( clk ), .D ( new_AGEMA_signal_15605 ), .Q ( new_AGEMA_signal_15606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4114 ( .C ( clk ), .D ( new_AGEMA_signal_15613 ), .Q ( new_AGEMA_signal_15614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4128 ( .C ( clk ), .D ( new_AGEMA_signal_15627 ), .Q ( new_AGEMA_signal_15628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4134 ( .C ( clk ), .D ( new_AGEMA_signal_15633 ), .Q ( new_AGEMA_signal_15634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4140 ( .C ( clk ), .D ( new_AGEMA_signal_15639 ), .Q ( new_AGEMA_signal_15640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4146 ( .C ( clk ), .D ( new_AGEMA_signal_15645 ), .Q ( new_AGEMA_signal_15646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4170 ( .C ( clk ), .D ( new_AGEMA_signal_15669 ), .Q ( new_AGEMA_signal_15670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4178 ( .C ( clk ), .D ( new_AGEMA_signal_15677 ), .Q ( new_AGEMA_signal_15678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4186 ( .C ( clk ), .D ( new_AGEMA_signal_15685 ), .Q ( new_AGEMA_signal_15686 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4194 ( .C ( clk ), .D ( new_AGEMA_signal_15693 ), .Q ( new_AGEMA_signal_15694 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4216 ( .C ( clk ), .D ( new_AGEMA_signal_15715 ), .Q ( new_AGEMA_signal_15716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4222 ( .C ( clk ), .D ( new_AGEMA_signal_15721 ), .Q ( new_AGEMA_signal_15722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4228 ( .C ( clk ), .D ( new_AGEMA_signal_15727 ), .Q ( new_AGEMA_signal_15728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4234 ( .C ( clk ), .D ( new_AGEMA_signal_15733 ), .Q ( new_AGEMA_signal_15734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4240 ( .C ( clk ), .D ( new_AGEMA_signal_15739 ), .Q ( new_AGEMA_signal_15740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4246 ( .C ( clk ), .D ( new_AGEMA_signal_15745 ), .Q ( new_AGEMA_signal_15746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4252 ( .C ( clk ), .D ( new_AGEMA_signal_15751 ), .Q ( new_AGEMA_signal_15752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4258 ( .C ( clk ), .D ( new_AGEMA_signal_15757 ), .Q ( new_AGEMA_signal_15758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4264 ( .C ( clk ), .D ( new_AGEMA_signal_15763 ), .Q ( new_AGEMA_signal_15764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4270 ( .C ( clk ), .D ( new_AGEMA_signal_15769 ), .Q ( new_AGEMA_signal_15770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4276 ( .C ( clk ), .D ( new_AGEMA_signal_15775 ), .Q ( new_AGEMA_signal_15776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4282 ( .C ( clk ), .D ( new_AGEMA_signal_15781 ), .Q ( new_AGEMA_signal_15782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4288 ( .C ( clk ), .D ( new_AGEMA_signal_15787 ), .Q ( new_AGEMA_signal_15788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4294 ( .C ( clk ), .D ( new_AGEMA_signal_15793 ), .Q ( new_AGEMA_signal_15794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4300 ( .C ( clk ), .D ( new_AGEMA_signal_15799 ), .Q ( new_AGEMA_signal_15800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4306 ( .C ( clk ), .D ( new_AGEMA_signal_15805 ), .Q ( new_AGEMA_signal_15806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4312 ( .C ( clk ), .D ( new_AGEMA_signal_15811 ), .Q ( new_AGEMA_signal_15812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4318 ( .C ( clk ), .D ( new_AGEMA_signal_15817 ), .Q ( new_AGEMA_signal_15818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4324 ( .C ( clk ), .D ( new_AGEMA_signal_15823 ), .Q ( new_AGEMA_signal_15824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4330 ( .C ( clk ), .D ( new_AGEMA_signal_15829 ), .Q ( new_AGEMA_signal_15830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4354 ( .C ( clk ), .D ( new_AGEMA_signal_15853 ), .Q ( new_AGEMA_signal_15854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4362 ( .C ( clk ), .D ( new_AGEMA_signal_15861 ), .Q ( new_AGEMA_signal_15862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4370 ( .C ( clk ), .D ( new_AGEMA_signal_15869 ), .Q ( new_AGEMA_signal_15870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4378 ( .C ( clk ), .D ( new_AGEMA_signal_15877 ), .Q ( new_AGEMA_signal_15878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4400 ( .C ( clk ), .D ( new_AGEMA_signal_15899 ), .Q ( new_AGEMA_signal_15900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4406 ( .C ( clk ), .D ( new_AGEMA_signal_15905 ), .Q ( new_AGEMA_signal_15906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4412 ( .C ( clk ), .D ( new_AGEMA_signal_15911 ), .Q ( new_AGEMA_signal_15912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4418 ( .C ( clk ), .D ( new_AGEMA_signal_15917 ), .Q ( new_AGEMA_signal_15918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4426 ( .C ( clk ), .D ( new_AGEMA_signal_15925 ), .Q ( new_AGEMA_signal_15926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4434 ( .C ( clk ), .D ( new_AGEMA_signal_15933 ), .Q ( new_AGEMA_signal_15934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4442 ( .C ( clk ), .D ( new_AGEMA_signal_15941 ), .Q ( new_AGEMA_signal_15942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4450 ( .C ( clk ), .D ( new_AGEMA_signal_15949 ), .Q ( new_AGEMA_signal_15950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4464 ( .C ( clk ), .D ( new_AGEMA_signal_15963 ), .Q ( new_AGEMA_signal_15964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4470 ( .C ( clk ), .D ( new_AGEMA_signal_15969 ), .Q ( new_AGEMA_signal_15970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4476 ( .C ( clk ), .D ( new_AGEMA_signal_15975 ), .Q ( new_AGEMA_signal_15976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4482 ( .C ( clk ), .D ( new_AGEMA_signal_15981 ), .Q ( new_AGEMA_signal_15982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4504 ( .C ( clk ), .D ( new_AGEMA_signal_16003 ), .Q ( new_AGEMA_signal_16004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4510 ( .C ( clk ), .D ( new_AGEMA_signal_16009 ), .Q ( new_AGEMA_signal_16010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4516 ( .C ( clk ), .D ( new_AGEMA_signal_16015 ), .Q ( new_AGEMA_signal_16016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4522 ( .C ( clk ), .D ( new_AGEMA_signal_16021 ), .Q ( new_AGEMA_signal_16022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4528 ( .C ( clk ), .D ( new_AGEMA_signal_16027 ), .Q ( new_AGEMA_signal_16028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4534 ( .C ( clk ), .D ( new_AGEMA_signal_16033 ), .Q ( new_AGEMA_signal_16034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4540 ( .C ( clk ), .D ( new_AGEMA_signal_16039 ), .Q ( new_AGEMA_signal_16040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4546 ( .C ( clk ), .D ( new_AGEMA_signal_16045 ), .Q ( new_AGEMA_signal_16046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4554 ( .C ( clk ), .D ( new_AGEMA_signal_16053 ), .Q ( new_AGEMA_signal_16054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4562 ( .C ( clk ), .D ( new_AGEMA_signal_16061 ), .Q ( new_AGEMA_signal_16062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4570 ( .C ( clk ), .D ( new_AGEMA_signal_16069 ), .Q ( new_AGEMA_signal_16070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4578 ( .C ( clk ), .D ( new_AGEMA_signal_16077 ), .Q ( new_AGEMA_signal_16078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4586 ( .C ( clk ), .D ( new_AGEMA_signal_16085 ), .Q ( new_AGEMA_signal_16086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4594 ( .C ( clk ), .D ( new_AGEMA_signal_16093 ), .Q ( new_AGEMA_signal_16094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4602 ( .C ( clk ), .D ( new_AGEMA_signal_16101 ), .Q ( new_AGEMA_signal_16102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4610 ( .C ( clk ), .D ( new_AGEMA_signal_16109 ), .Q ( new_AGEMA_signal_16110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4616 ( .C ( clk ), .D ( new_AGEMA_signal_16115 ), .Q ( new_AGEMA_signal_16116 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4622 ( .C ( clk ), .D ( new_AGEMA_signal_16121 ), .Q ( new_AGEMA_signal_16122 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4628 ( .C ( clk ), .D ( new_AGEMA_signal_16127 ), .Q ( new_AGEMA_signal_16128 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4634 ( .C ( clk ), .D ( new_AGEMA_signal_16133 ), .Q ( new_AGEMA_signal_16134 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4640 ( .C ( clk ), .D ( new_AGEMA_signal_16139 ), .Q ( new_AGEMA_signal_16140 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4646 ( .C ( clk ), .D ( new_AGEMA_signal_16145 ), .Q ( new_AGEMA_signal_16146 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4652 ( .C ( clk ), .D ( new_AGEMA_signal_16151 ), .Q ( new_AGEMA_signal_16152 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4658 ( .C ( clk ), .D ( new_AGEMA_signal_16157 ), .Q ( new_AGEMA_signal_16158 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4776 ( .C ( clk ), .D ( new_AGEMA_signal_16275 ), .Q ( new_AGEMA_signal_16276 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4784 ( .C ( clk ), .D ( new_AGEMA_signal_16283 ), .Q ( new_AGEMA_signal_16284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4792 ( .C ( clk ), .D ( new_AGEMA_signal_16291 ), .Q ( new_AGEMA_signal_16292 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4800 ( .C ( clk ), .D ( new_AGEMA_signal_16299 ), .Q ( new_AGEMA_signal_16300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4808 ( .C ( clk ), .D ( new_AGEMA_signal_16307 ), .Q ( new_AGEMA_signal_16308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4816 ( .C ( clk ), .D ( new_AGEMA_signal_16315 ), .Q ( new_AGEMA_signal_16316 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4824 ( .C ( clk ), .D ( new_AGEMA_signal_16323 ), .Q ( new_AGEMA_signal_16324 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4832 ( .C ( clk ), .D ( new_AGEMA_signal_16331 ), .Q ( new_AGEMA_signal_16332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4840 ( .C ( clk ), .D ( new_AGEMA_signal_16339 ), .Q ( new_AGEMA_signal_16340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4848 ( .C ( clk ), .D ( new_AGEMA_signal_16347 ), .Q ( new_AGEMA_signal_16348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4856 ( .C ( clk ), .D ( new_AGEMA_signal_16355 ), .Q ( new_AGEMA_signal_16356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4864 ( .C ( clk ), .D ( new_AGEMA_signal_16363 ), .Q ( new_AGEMA_signal_16364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4872 ( .C ( clk ), .D ( new_AGEMA_signal_16371 ), .Q ( new_AGEMA_signal_16372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4880 ( .C ( clk ), .D ( new_AGEMA_signal_16379 ), .Q ( new_AGEMA_signal_16380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4888 ( .C ( clk ), .D ( new_AGEMA_signal_16387 ), .Q ( new_AGEMA_signal_16388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4896 ( .C ( clk ), .D ( new_AGEMA_signal_16395 ), .Q ( new_AGEMA_signal_16396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4930 ( .C ( clk ), .D ( new_AGEMA_signal_16429 ), .Q ( new_AGEMA_signal_16430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4940 ( .C ( clk ), .D ( new_AGEMA_signal_16439 ), .Q ( new_AGEMA_signal_16440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4950 ( .C ( clk ), .D ( new_AGEMA_signal_16449 ), .Q ( new_AGEMA_signal_16450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4960 ( .C ( clk ), .D ( new_AGEMA_signal_16459 ), .Q ( new_AGEMA_signal_16460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4968 ( .C ( clk ), .D ( new_AGEMA_signal_16467 ), .Q ( new_AGEMA_signal_16468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4976 ( .C ( clk ), .D ( new_AGEMA_signal_16475 ), .Q ( new_AGEMA_signal_16476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4984 ( .C ( clk ), .D ( new_AGEMA_signal_16483 ), .Q ( new_AGEMA_signal_16484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4992 ( .C ( clk ), .D ( new_AGEMA_signal_16491 ), .Q ( new_AGEMA_signal_16492 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5000 ( .C ( clk ), .D ( new_AGEMA_signal_16499 ), .Q ( new_AGEMA_signal_16500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5008 ( .C ( clk ), .D ( new_AGEMA_signal_16507 ), .Q ( new_AGEMA_signal_16508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5016 ( .C ( clk ), .D ( new_AGEMA_signal_16515 ), .Q ( new_AGEMA_signal_16516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5024 ( .C ( clk ), .D ( new_AGEMA_signal_16523 ), .Q ( new_AGEMA_signal_16524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5032 ( .C ( clk ), .D ( new_AGEMA_signal_16531 ), .Q ( new_AGEMA_signal_16532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5040 ( .C ( clk ), .D ( new_AGEMA_signal_16539 ), .Q ( new_AGEMA_signal_16540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5048 ( .C ( clk ), .D ( new_AGEMA_signal_16547 ), .Q ( new_AGEMA_signal_16548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5056 ( .C ( clk ), .D ( new_AGEMA_signal_16555 ), .Q ( new_AGEMA_signal_16556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5130 ( .C ( clk ), .D ( new_AGEMA_signal_16629 ), .Q ( new_AGEMA_signal_16630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5140 ( .C ( clk ), .D ( new_AGEMA_signal_16639 ), .Q ( new_AGEMA_signal_16640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5150 ( .C ( clk ), .D ( new_AGEMA_signal_16649 ), .Q ( new_AGEMA_signal_16650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5160 ( .C ( clk ), .D ( new_AGEMA_signal_16659 ), .Q ( new_AGEMA_signal_16660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5168 ( .C ( clk ), .D ( new_AGEMA_signal_16667 ), .Q ( new_AGEMA_signal_16668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5176 ( .C ( clk ), .D ( new_AGEMA_signal_16675 ), .Q ( new_AGEMA_signal_16676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5184 ( .C ( clk ), .D ( new_AGEMA_signal_16683 ), .Q ( new_AGEMA_signal_16684 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5192 ( .C ( clk ), .D ( new_AGEMA_signal_16691 ), .Q ( new_AGEMA_signal_16692 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5224 ( .C ( clk ), .D ( new_AGEMA_signal_16723 ), .Q ( new_AGEMA_signal_16724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5232 ( .C ( clk ), .D ( new_AGEMA_signal_16731 ), .Q ( new_AGEMA_signal_16732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5240 ( .C ( clk ), .D ( new_AGEMA_signal_16739 ), .Q ( new_AGEMA_signal_16740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5248 ( .C ( clk ), .D ( new_AGEMA_signal_16747 ), .Q ( new_AGEMA_signal_16748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5256 ( .C ( clk ), .D ( new_AGEMA_signal_16755 ), .Q ( new_AGEMA_signal_16756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5264 ( .C ( clk ), .D ( new_AGEMA_signal_16763 ), .Q ( new_AGEMA_signal_16764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5272 ( .C ( clk ), .D ( new_AGEMA_signal_16771 ), .Q ( new_AGEMA_signal_16772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5280 ( .C ( clk ), .D ( new_AGEMA_signal_16779 ), .Q ( new_AGEMA_signal_16780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5328 ( .C ( clk ), .D ( new_AGEMA_signal_16827 ), .Q ( new_AGEMA_signal_16828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5336 ( .C ( clk ), .D ( new_AGEMA_signal_16835 ), .Q ( new_AGEMA_signal_16836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5344 ( .C ( clk ), .D ( new_AGEMA_signal_16843 ), .Q ( new_AGEMA_signal_16844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5352 ( .C ( clk ), .D ( new_AGEMA_signal_16851 ), .Q ( new_AGEMA_signal_16852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5592 ( .C ( clk ), .D ( new_AGEMA_signal_17091 ), .Q ( new_AGEMA_signal_17092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5602 ( .C ( clk ), .D ( new_AGEMA_signal_17101 ), .Q ( new_AGEMA_signal_17102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5612 ( .C ( clk ), .D ( new_AGEMA_signal_17111 ), .Q ( new_AGEMA_signal_17112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5622 ( .C ( clk ), .D ( new_AGEMA_signal_17121 ), .Q ( new_AGEMA_signal_17122 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6376 ( .C ( clk ), .D ( new_AGEMA_signal_17875 ), .Q ( new_AGEMA_signal_17876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6390 ( .C ( clk ), .D ( new_AGEMA_signal_17889 ), .Q ( new_AGEMA_signal_17890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6404 ( .C ( clk ), .D ( new_AGEMA_signal_17903 ), .Q ( new_AGEMA_signal_17904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6418 ( .C ( clk ), .D ( new_AGEMA_signal_17917 ), .Q ( new_AGEMA_signal_17918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6464 ( .C ( clk ), .D ( new_AGEMA_signal_17963 ), .Q ( new_AGEMA_signal_17964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6478 ( .C ( clk ), .D ( new_AGEMA_signal_17977 ), .Q ( new_AGEMA_signal_17978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6492 ( .C ( clk ), .D ( new_AGEMA_signal_17991 ), .Q ( new_AGEMA_signal_17992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6506 ( .C ( clk ), .D ( new_AGEMA_signal_18005 ), .Q ( new_AGEMA_signal_18006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6608 ( .C ( clk ), .D ( new_AGEMA_signal_18107 ), .Q ( new_AGEMA_signal_18108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6624 ( .C ( clk ), .D ( new_AGEMA_signal_18123 ), .Q ( new_AGEMA_signal_18124 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6640 ( .C ( clk ), .D ( new_AGEMA_signal_18139 ), .Q ( new_AGEMA_signal_18140 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6656 ( .C ( clk ), .D ( new_AGEMA_signal_18155 ), .Q ( new_AGEMA_signal_18156 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6696 ( .C ( clk ), .D ( new_AGEMA_signal_18195 ), .Q ( new_AGEMA_signal_18196 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6712 ( .C ( clk ), .D ( new_AGEMA_signal_18211 ), .Q ( new_AGEMA_signal_18212 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6728 ( .C ( clk ), .D ( new_AGEMA_signal_18227 ), .Q ( new_AGEMA_signal_18228 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6744 ( .C ( clk ), .D ( new_AGEMA_signal_18243 ), .Q ( new_AGEMA_signal_18244 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7000 ( .C ( clk ), .D ( new_AGEMA_signal_18499 ), .Q ( new_AGEMA_signal_18500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7018 ( .C ( clk ), .D ( new_AGEMA_signal_18517 ), .Q ( new_AGEMA_signal_18518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7036 ( .C ( clk ), .D ( new_AGEMA_signal_18535 ), .Q ( new_AGEMA_signal_18536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7054 ( .C ( clk ), .D ( new_AGEMA_signal_18553 ), .Q ( new_AGEMA_signal_18554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7200 ( .C ( clk ), .D ( new_AGEMA_signal_18699 ), .Q ( new_AGEMA_signal_18700 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7220 ( .C ( clk ), .D ( new_AGEMA_signal_18719 ), .Q ( new_AGEMA_signal_18720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7240 ( .C ( clk ), .D ( new_AGEMA_signal_18739 ), .Q ( new_AGEMA_signal_18740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7260 ( .C ( clk ), .D ( new_AGEMA_signal_18759 ), .Q ( new_AGEMA_signal_18760 ) ) ;

    /* cells in depth 9 */
    buf_clk new_AGEMA_reg_buffer_3097 ( .C ( clk ), .D ( new_AGEMA_signal_14596 ), .Q ( new_AGEMA_signal_14597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3101 ( .C ( clk ), .D ( new_AGEMA_signal_14600 ), .Q ( new_AGEMA_signal_14601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3105 ( .C ( clk ), .D ( new_AGEMA_signal_14604 ), .Q ( new_AGEMA_signal_14605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3109 ( .C ( clk ), .D ( new_AGEMA_signal_14608 ), .Q ( new_AGEMA_signal_14609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3113 ( .C ( clk ), .D ( new_AGEMA_signal_14612 ), .Q ( new_AGEMA_signal_14613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3117 ( .C ( clk ), .D ( new_AGEMA_signal_14616 ), .Q ( new_AGEMA_signal_14617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3121 ( .C ( clk ), .D ( new_AGEMA_signal_14620 ), .Q ( new_AGEMA_signal_14621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3125 ( .C ( clk ), .D ( new_AGEMA_signal_14624 ), .Q ( new_AGEMA_signal_14625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3133 ( .C ( clk ), .D ( new_AGEMA_signal_14632 ), .Q ( new_AGEMA_signal_14633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3141 ( .C ( clk ), .D ( new_AGEMA_signal_14640 ), .Q ( new_AGEMA_signal_14641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3149 ( .C ( clk ), .D ( new_AGEMA_signal_14648 ), .Q ( new_AGEMA_signal_14649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3157 ( .C ( clk ), .D ( new_AGEMA_signal_14656 ), .Q ( new_AGEMA_signal_14657 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3159 ( .C ( clk ), .D ( n1978 ), .Q ( new_AGEMA_signal_14659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3161 ( .C ( clk ), .D ( new_AGEMA_signal_2562 ), .Q ( new_AGEMA_signal_14661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3163 ( .C ( clk ), .D ( new_AGEMA_signal_2563 ), .Q ( new_AGEMA_signal_14663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3165 ( .C ( clk ), .D ( new_AGEMA_signal_2564 ), .Q ( new_AGEMA_signal_14665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3173 ( .C ( clk ), .D ( new_AGEMA_signal_14672 ), .Q ( new_AGEMA_signal_14673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3181 ( .C ( clk ), .D ( new_AGEMA_signal_14680 ), .Q ( new_AGEMA_signal_14681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3189 ( .C ( clk ), .D ( new_AGEMA_signal_14688 ), .Q ( new_AGEMA_signal_14689 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3197 ( .C ( clk ), .D ( new_AGEMA_signal_14696 ), .Q ( new_AGEMA_signal_14697 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3203 ( .C ( clk ), .D ( new_AGEMA_signal_14702 ), .Q ( new_AGEMA_signal_14703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3209 ( .C ( clk ), .D ( new_AGEMA_signal_14708 ), .Q ( new_AGEMA_signal_14709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3215 ( .C ( clk ), .D ( new_AGEMA_signal_14714 ), .Q ( new_AGEMA_signal_14715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3221 ( .C ( clk ), .D ( new_AGEMA_signal_14720 ), .Q ( new_AGEMA_signal_14721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3225 ( .C ( clk ), .D ( new_AGEMA_signal_14724 ), .Q ( new_AGEMA_signal_14725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3229 ( .C ( clk ), .D ( new_AGEMA_signal_14728 ), .Q ( new_AGEMA_signal_14729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3233 ( .C ( clk ), .D ( new_AGEMA_signal_14732 ), .Q ( new_AGEMA_signal_14733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3237 ( .C ( clk ), .D ( new_AGEMA_signal_14736 ), .Q ( new_AGEMA_signal_14737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3243 ( .C ( clk ), .D ( new_AGEMA_signal_14742 ), .Q ( new_AGEMA_signal_14743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3249 ( .C ( clk ), .D ( new_AGEMA_signal_14748 ), .Q ( new_AGEMA_signal_14749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3255 ( .C ( clk ), .D ( new_AGEMA_signal_14754 ), .Q ( new_AGEMA_signal_14755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3261 ( .C ( clk ), .D ( new_AGEMA_signal_14760 ), .Q ( new_AGEMA_signal_14761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3263 ( .C ( clk ), .D ( new_AGEMA_signal_14374 ), .Q ( new_AGEMA_signal_14763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3265 ( .C ( clk ), .D ( new_AGEMA_signal_14378 ), .Q ( new_AGEMA_signal_14765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3267 ( .C ( clk ), .D ( new_AGEMA_signal_14382 ), .Q ( new_AGEMA_signal_14767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3269 ( .C ( clk ), .D ( new_AGEMA_signal_14386 ), .Q ( new_AGEMA_signal_14769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3275 ( .C ( clk ), .D ( new_AGEMA_signal_14774 ), .Q ( new_AGEMA_signal_14775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3281 ( .C ( clk ), .D ( new_AGEMA_signal_14780 ), .Q ( new_AGEMA_signal_14781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3287 ( .C ( clk ), .D ( new_AGEMA_signal_14786 ), .Q ( new_AGEMA_signal_14787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3293 ( .C ( clk ), .D ( new_AGEMA_signal_14792 ), .Q ( new_AGEMA_signal_14793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3299 ( .C ( clk ), .D ( new_AGEMA_signal_14798 ), .Q ( new_AGEMA_signal_14799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3305 ( .C ( clk ), .D ( new_AGEMA_signal_14804 ), .Q ( new_AGEMA_signal_14805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3311 ( .C ( clk ), .D ( new_AGEMA_signal_14810 ), .Q ( new_AGEMA_signal_14811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3317 ( .C ( clk ), .D ( new_AGEMA_signal_14816 ), .Q ( new_AGEMA_signal_14817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3319 ( .C ( clk ), .D ( n2091 ), .Q ( new_AGEMA_signal_14819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3321 ( .C ( clk ), .D ( new_AGEMA_signal_2616 ), .Q ( new_AGEMA_signal_14821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3323 ( .C ( clk ), .D ( new_AGEMA_signal_2617 ), .Q ( new_AGEMA_signal_14823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3325 ( .C ( clk ), .D ( new_AGEMA_signal_2618 ), .Q ( new_AGEMA_signal_14825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3329 ( .C ( clk ), .D ( new_AGEMA_signal_14828 ), .Q ( new_AGEMA_signal_14829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3333 ( .C ( clk ), .D ( new_AGEMA_signal_14832 ), .Q ( new_AGEMA_signal_14833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3337 ( .C ( clk ), .D ( new_AGEMA_signal_14836 ), .Q ( new_AGEMA_signal_14837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3341 ( .C ( clk ), .D ( new_AGEMA_signal_14840 ), .Q ( new_AGEMA_signal_14841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3347 ( .C ( clk ), .D ( new_AGEMA_signal_14846 ), .Q ( new_AGEMA_signal_14847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3353 ( .C ( clk ), .D ( new_AGEMA_signal_14852 ), .Q ( new_AGEMA_signal_14853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3359 ( .C ( clk ), .D ( new_AGEMA_signal_14858 ), .Q ( new_AGEMA_signal_14859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3365 ( .C ( clk ), .D ( new_AGEMA_signal_14864 ), .Q ( new_AGEMA_signal_14865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3371 ( .C ( clk ), .D ( new_AGEMA_signal_14870 ), .Q ( new_AGEMA_signal_14871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3377 ( .C ( clk ), .D ( new_AGEMA_signal_14876 ), .Q ( new_AGEMA_signal_14877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3383 ( .C ( clk ), .D ( new_AGEMA_signal_14882 ), .Q ( new_AGEMA_signal_14883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3389 ( .C ( clk ), .D ( new_AGEMA_signal_14888 ), .Q ( new_AGEMA_signal_14889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3391 ( .C ( clk ), .D ( n2543 ), .Q ( new_AGEMA_signal_14891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3393 ( .C ( clk ), .D ( new_AGEMA_signal_2634 ), .Q ( new_AGEMA_signal_14893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3395 ( .C ( clk ), .D ( new_AGEMA_signal_2635 ), .Q ( new_AGEMA_signal_14895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3397 ( .C ( clk ), .D ( new_AGEMA_signal_2636 ), .Q ( new_AGEMA_signal_14897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3403 ( .C ( clk ), .D ( new_AGEMA_signal_14902 ), .Q ( new_AGEMA_signal_14903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3409 ( .C ( clk ), .D ( new_AGEMA_signal_14908 ), .Q ( new_AGEMA_signal_14909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3415 ( .C ( clk ), .D ( new_AGEMA_signal_14914 ), .Q ( new_AGEMA_signal_14915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3421 ( .C ( clk ), .D ( new_AGEMA_signal_14920 ), .Q ( new_AGEMA_signal_14921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3423 ( .C ( clk ), .D ( n2159 ), .Q ( new_AGEMA_signal_14923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3425 ( .C ( clk ), .D ( new_AGEMA_signal_2646 ), .Q ( new_AGEMA_signal_14925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3427 ( .C ( clk ), .D ( new_AGEMA_signal_2647 ), .Q ( new_AGEMA_signal_14927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3429 ( .C ( clk ), .D ( new_AGEMA_signal_2648 ), .Q ( new_AGEMA_signal_14929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3433 ( .C ( clk ), .D ( new_AGEMA_signal_14932 ), .Q ( new_AGEMA_signal_14933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3437 ( .C ( clk ), .D ( new_AGEMA_signal_14936 ), .Q ( new_AGEMA_signal_14937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3441 ( .C ( clk ), .D ( new_AGEMA_signal_14940 ), .Q ( new_AGEMA_signal_14941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3445 ( .C ( clk ), .D ( new_AGEMA_signal_14944 ), .Q ( new_AGEMA_signal_14945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3449 ( .C ( clk ), .D ( new_AGEMA_signal_14948 ), .Q ( new_AGEMA_signal_14949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3453 ( .C ( clk ), .D ( new_AGEMA_signal_14952 ), .Q ( new_AGEMA_signal_14953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3457 ( .C ( clk ), .D ( new_AGEMA_signal_14956 ), .Q ( new_AGEMA_signal_14957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3461 ( .C ( clk ), .D ( new_AGEMA_signal_14960 ), .Q ( new_AGEMA_signal_14961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3463 ( .C ( clk ), .D ( new_AGEMA_signal_14348 ), .Q ( new_AGEMA_signal_14963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3465 ( .C ( clk ), .D ( new_AGEMA_signal_14350 ), .Q ( new_AGEMA_signal_14965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3467 ( .C ( clk ), .D ( new_AGEMA_signal_14352 ), .Q ( new_AGEMA_signal_14967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3469 ( .C ( clk ), .D ( new_AGEMA_signal_14354 ), .Q ( new_AGEMA_signal_14969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3477 ( .C ( clk ), .D ( new_AGEMA_signal_14976 ), .Q ( new_AGEMA_signal_14977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3485 ( .C ( clk ), .D ( new_AGEMA_signal_14984 ), .Q ( new_AGEMA_signal_14985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3493 ( .C ( clk ), .D ( new_AGEMA_signal_14992 ), .Q ( new_AGEMA_signal_14993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3501 ( .C ( clk ), .D ( new_AGEMA_signal_15000 ), .Q ( new_AGEMA_signal_15001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3507 ( .C ( clk ), .D ( new_AGEMA_signal_15006 ), .Q ( new_AGEMA_signal_15007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3513 ( .C ( clk ), .D ( new_AGEMA_signal_15012 ), .Q ( new_AGEMA_signal_15013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3519 ( .C ( clk ), .D ( new_AGEMA_signal_15018 ), .Q ( new_AGEMA_signal_15019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3525 ( .C ( clk ), .D ( new_AGEMA_signal_15024 ), .Q ( new_AGEMA_signal_15025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3529 ( .C ( clk ), .D ( new_AGEMA_signal_15028 ), .Q ( new_AGEMA_signal_15029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3533 ( .C ( clk ), .D ( new_AGEMA_signal_15032 ), .Q ( new_AGEMA_signal_15033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3537 ( .C ( clk ), .D ( new_AGEMA_signal_15036 ), .Q ( new_AGEMA_signal_15037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3541 ( .C ( clk ), .D ( new_AGEMA_signal_15040 ), .Q ( new_AGEMA_signal_15041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3545 ( .C ( clk ), .D ( new_AGEMA_signal_15044 ), .Q ( new_AGEMA_signal_15045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3549 ( .C ( clk ), .D ( new_AGEMA_signal_15048 ), .Q ( new_AGEMA_signal_15049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3553 ( .C ( clk ), .D ( new_AGEMA_signal_15052 ), .Q ( new_AGEMA_signal_15053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3557 ( .C ( clk ), .D ( new_AGEMA_signal_15056 ), .Q ( new_AGEMA_signal_15057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3559 ( .C ( clk ), .D ( n2270 ), .Q ( new_AGEMA_signal_15059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3561 ( .C ( clk ), .D ( new_AGEMA_signal_2274 ), .Q ( new_AGEMA_signal_15061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3563 ( .C ( clk ), .D ( new_AGEMA_signal_2275 ), .Q ( new_AGEMA_signal_15063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3565 ( .C ( clk ), .D ( new_AGEMA_signal_2276 ), .Q ( new_AGEMA_signal_15065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3567 ( .C ( clk ), .D ( n2285 ), .Q ( new_AGEMA_signal_15067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3569 ( .C ( clk ), .D ( new_AGEMA_signal_2700 ), .Q ( new_AGEMA_signal_15069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3571 ( .C ( clk ), .D ( new_AGEMA_signal_2701 ), .Q ( new_AGEMA_signal_15071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3573 ( .C ( clk ), .D ( new_AGEMA_signal_2702 ), .Q ( new_AGEMA_signal_15073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3577 ( .C ( clk ), .D ( new_AGEMA_signal_15076 ), .Q ( new_AGEMA_signal_15077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3581 ( .C ( clk ), .D ( new_AGEMA_signal_15080 ), .Q ( new_AGEMA_signal_15081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3585 ( .C ( clk ), .D ( new_AGEMA_signal_15084 ), .Q ( new_AGEMA_signal_15085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3589 ( .C ( clk ), .D ( new_AGEMA_signal_15088 ), .Q ( new_AGEMA_signal_15089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3593 ( .C ( clk ), .D ( new_AGEMA_signal_15092 ), .Q ( new_AGEMA_signal_15093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3597 ( .C ( clk ), .D ( new_AGEMA_signal_15096 ), .Q ( new_AGEMA_signal_15097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3601 ( .C ( clk ), .D ( new_AGEMA_signal_15100 ), .Q ( new_AGEMA_signal_15101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3605 ( .C ( clk ), .D ( new_AGEMA_signal_15104 ), .Q ( new_AGEMA_signal_15105 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3607 ( .C ( clk ), .D ( n2334 ), .Q ( new_AGEMA_signal_15107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3609 ( .C ( clk ), .D ( new_AGEMA_signal_2307 ), .Q ( new_AGEMA_signal_15109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3611 ( .C ( clk ), .D ( new_AGEMA_signal_2308 ), .Q ( new_AGEMA_signal_15111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3613 ( .C ( clk ), .D ( new_AGEMA_signal_2309 ), .Q ( new_AGEMA_signal_15113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3619 ( .C ( clk ), .D ( new_AGEMA_signal_15118 ), .Q ( new_AGEMA_signal_15119 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3625 ( .C ( clk ), .D ( new_AGEMA_signal_15124 ), .Q ( new_AGEMA_signal_15125 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3631 ( .C ( clk ), .D ( new_AGEMA_signal_15130 ), .Q ( new_AGEMA_signal_15131 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3637 ( .C ( clk ), .D ( new_AGEMA_signal_15136 ), .Q ( new_AGEMA_signal_15137 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3641 ( .C ( clk ), .D ( new_AGEMA_signal_15140 ), .Q ( new_AGEMA_signal_15141 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3645 ( .C ( clk ), .D ( new_AGEMA_signal_15144 ), .Q ( new_AGEMA_signal_15145 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3649 ( .C ( clk ), .D ( new_AGEMA_signal_15148 ), .Q ( new_AGEMA_signal_15149 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3653 ( .C ( clk ), .D ( new_AGEMA_signal_15152 ), .Q ( new_AGEMA_signal_15153 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3655 ( .C ( clk ), .D ( new_AGEMA_signal_14364 ), .Q ( new_AGEMA_signal_15155 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3657 ( .C ( clk ), .D ( new_AGEMA_signal_14366 ), .Q ( new_AGEMA_signal_15157 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3659 ( .C ( clk ), .D ( new_AGEMA_signal_14368 ), .Q ( new_AGEMA_signal_15159 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3661 ( .C ( clk ), .D ( new_AGEMA_signal_14370 ), .Q ( new_AGEMA_signal_15161 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3665 ( .C ( clk ), .D ( new_AGEMA_signal_15164 ), .Q ( new_AGEMA_signal_15165 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3669 ( .C ( clk ), .D ( new_AGEMA_signal_15168 ), .Q ( new_AGEMA_signal_15169 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3673 ( .C ( clk ), .D ( new_AGEMA_signal_15172 ), .Q ( new_AGEMA_signal_15173 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3677 ( .C ( clk ), .D ( new_AGEMA_signal_15176 ), .Q ( new_AGEMA_signal_15177 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3681 ( .C ( clk ), .D ( new_AGEMA_signal_15180 ), .Q ( new_AGEMA_signal_15181 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3685 ( .C ( clk ), .D ( new_AGEMA_signal_15184 ), .Q ( new_AGEMA_signal_15185 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3689 ( .C ( clk ), .D ( new_AGEMA_signal_15188 ), .Q ( new_AGEMA_signal_15189 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3693 ( .C ( clk ), .D ( new_AGEMA_signal_15192 ), .Q ( new_AGEMA_signal_15193 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3697 ( .C ( clk ), .D ( new_AGEMA_signal_15196 ), .Q ( new_AGEMA_signal_15197 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3701 ( .C ( clk ), .D ( new_AGEMA_signal_15200 ), .Q ( new_AGEMA_signal_15201 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3705 ( .C ( clk ), .D ( new_AGEMA_signal_15204 ), .Q ( new_AGEMA_signal_15205 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3709 ( .C ( clk ), .D ( new_AGEMA_signal_15208 ), .Q ( new_AGEMA_signal_15209 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3711 ( .C ( clk ), .D ( n2435 ), .Q ( new_AGEMA_signal_15211 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3713 ( .C ( clk ), .D ( new_AGEMA_signal_2364 ), .Q ( new_AGEMA_signal_15213 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3715 ( .C ( clk ), .D ( new_AGEMA_signal_2365 ), .Q ( new_AGEMA_signal_15215 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3717 ( .C ( clk ), .D ( new_AGEMA_signal_2366 ), .Q ( new_AGEMA_signal_15217 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3721 ( .C ( clk ), .D ( new_AGEMA_signal_15220 ), .Q ( new_AGEMA_signal_15221 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3725 ( .C ( clk ), .D ( new_AGEMA_signal_15224 ), .Q ( new_AGEMA_signal_15225 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3729 ( .C ( clk ), .D ( new_AGEMA_signal_15228 ), .Q ( new_AGEMA_signal_15229 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3733 ( .C ( clk ), .D ( new_AGEMA_signal_15232 ), .Q ( new_AGEMA_signal_15233 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3735 ( .C ( clk ), .D ( new_AGEMA_signal_14212 ), .Q ( new_AGEMA_signal_15235 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3737 ( .C ( clk ), .D ( new_AGEMA_signal_14214 ), .Q ( new_AGEMA_signal_15237 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3739 ( .C ( clk ), .D ( new_AGEMA_signal_14216 ), .Q ( new_AGEMA_signal_15239 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3741 ( .C ( clk ), .D ( new_AGEMA_signal_14218 ), .Q ( new_AGEMA_signal_15241 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3747 ( .C ( clk ), .D ( new_AGEMA_signal_15246 ), .Q ( new_AGEMA_signal_15247 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3753 ( .C ( clk ), .D ( new_AGEMA_signal_15252 ), .Q ( new_AGEMA_signal_15253 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3759 ( .C ( clk ), .D ( new_AGEMA_signal_15258 ), .Q ( new_AGEMA_signal_15259 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3765 ( .C ( clk ), .D ( new_AGEMA_signal_15264 ), .Q ( new_AGEMA_signal_15265 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3771 ( .C ( clk ), .D ( new_AGEMA_signal_15270 ), .Q ( new_AGEMA_signal_15271 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3777 ( .C ( clk ), .D ( new_AGEMA_signal_15276 ), .Q ( new_AGEMA_signal_15277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3783 ( .C ( clk ), .D ( new_AGEMA_signal_15282 ), .Q ( new_AGEMA_signal_15283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3789 ( .C ( clk ), .D ( new_AGEMA_signal_15288 ), .Q ( new_AGEMA_signal_15289 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3793 ( .C ( clk ), .D ( new_AGEMA_signal_15292 ), .Q ( new_AGEMA_signal_15293 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3797 ( .C ( clk ), .D ( new_AGEMA_signal_15296 ), .Q ( new_AGEMA_signal_15297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3801 ( .C ( clk ), .D ( new_AGEMA_signal_15300 ), .Q ( new_AGEMA_signal_15301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3805 ( .C ( clk ), .D ( new_AGEMA_signal_15304 ), .Q ( new_AGEMA_signal_15305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3807 ( .C ( clk ), .D ( new_AGEMA_signal_14168 ), .Q ( new_AGEMA_signal_15307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3809 ( .C ( clk ), .D ( new_AGEMA_signal_14174 ), .Q ( new_AGEMA_signal_15309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3811 ( .C ( clk ), .D ( new_AGEMA_signal_14180 ), .Q ( new_AGEMA_signal_15311 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3813 ( .C ( clk ), .D ( new_AGEMA_signal_14186 ), .Q ( new_AGEMA_signal_15313 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3821 ( .C ( clk ), .D ( new_AGEMA_signal_15320 ), .Q ( new_AGEMA_signal_15321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3829 ( .C ( clk ), .D ( new_AGEMA_signal_15328 ), .Q ( new_AGEMA_signal_15329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3837 ( .C ( clk ), .D ( new_AGEMA_signal_15336 ), .Q ( new_AGEMA_signal_15337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3845 ( .C ( clk ), .D ( new_AGEMA_signal_15344 ), .Q ( new_AGEMA_signal_15345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3847 ( .C ( clk ), .D ( n2547 ), .Q ( new_AGEMA_signal_15347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3849 ( .C ( clk ), .D ( new_AGEMA_signal_2418 ), .Q ( new_AGEMA_signal_15349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3851 ( .C ( clk ), .D ( new_AGEMA_signal_2419 ), .Q ( new_AGEMA_signal_15351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3853 ( .C ( clk ), .D ( new_AGEMA_signal_2420 ), .Q ( new_AGEMA_signal_15353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3857 ( .C ( clk ), .D ( new_AGEMA_signal_15356 ), .Q ( new_AGEMA_signal_15357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3861 ( .C ( clk ), .D ( new_AGEMA_signal_15360 ), .Q ( new_AGEMA_signal_15361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3865 ( .C ( clk ), .D ( new_AGEMA_signal_15364 ), .Q ( new_AGEMA_signal_15365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3869 ( .C ( clk ), .D ( new_AGEMA_signal_15368 ), .Q ( new_AGEMA_signal_15369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3873 ( .C ( clk ), .D ( new_AGEMA_signal_15372 ), .Q ( new_AGEMA_signal_15373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3877 ( .C ( clk ), .D ( new_AGEMA_signal_15376 ), .Q ( new_AGEMA_signal_15377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3881 ( .C ( clk ), .D ( new_AGEMA_signal_15380 ), .Q ( new_AGEMA_signal_15381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3885 ( .C ( clk ), .D ( new_AGEMA_signal_15384 ), .Q ( new_AGEMA_signal_15385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3889 ( .C ( clk ), .D ( new_AGEMA_signal_15388 ), .Q ( new_AGEMA_signal_15389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3893 ( .C ( clk ), .D ( new_AGEMA_signal_15392 ), .Q ( new_AGEMA_signal_15393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3897 ( .C ( clk ), .D ( new_AGEMA_signal_15396 ), .Q ( new_AGEMA_signal_15397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3901 ( .C ( clk ), .D ( new_AGEMA_signal_15400 ), .Q ( new_AGEMA_signal_15401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3905 ( .C ( clk ), .D ( new_AGEMA_signal_15404 ), .Q ( new_AGEMA_signal_15405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3909 ( .C ( clk ), .D ( new_AGEMA_signal_15408 ), .Q ( new_AGEMA_signal_15409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3913 ( .C ( clk ), .D ( new_AGEMA_signal_15412 ), .Q ( new_AGEMA_signal_15413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3917 ( .C ( clk ), .D ( new_AGEMA_signal_15416 ), .Q ( new_AGEMA_signal_15417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3921 ( .C ( clk ), .D ( new_AGEMA_signal_15420 ), .Q ( new_AGEMA_signal_15421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3925 ( .C ( clk ), .D ( new_AGEMA_signal_15424 ), .Q ( new_AGEMA_signal_15425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3929 ( .C ( clk ), .D ( new_AGEMA_signal_15428 ), .Q ( new_AGEMA_signal_15429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3933 ( .C ( clk ), .D ( new_AGEMA_signal_15432 ), .Q ( new_AGEMA_signal_15433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3941 ( .C ( clk ), .D ( new_AGEMA_signal_15440 ), .Q ( new_AGEMA_signal_15441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3949 ( .C ( clk ), .D ( new_AGEMA_signal_15448 ), .Q ( new_AGEMA_signal_15449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3957 ( .C ( clk ), .D ( new_AGEMA_signal_15456 ), .Q ( new_AGEMA_signal_15457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3965 ( .C ( clk ), .D ( new_AGEMA_signal_15464 ), .Q ( new_AGEMA_signal_15465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3967 ( .C ( clk ), .D ( n2758 ), .Q ( new_AGEMA_signal_15467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3969 ( .C ( clk ), .D ( new_AGEMA_signal_2853 ), .Q ( new_AGEMA_signal_15469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3971 ( .C ( clk ), .D ( new_AGEMA_signal_2854 ), .Q ( new_AGEMA_signal_15471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3973 ( .C ( clk ), .D ( new_AGEMA_signal_2855 ), .Q ( new_AGEMA_signal_15473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3977 ( .C ( clk ), .D ( new_AGEMA_signal_15476 ), .Q ( new_AGEMA_signal_15477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3981 ( .C ( clk ), .D ( new_AGEMA_signal_15480 ), .Q ( new_AGEMA_signal_15481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3985 ( .C ( clk ), .D ( new_AGEMA_signal_15484 ), .Q ( new_AGEMA_signal_15485 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3989 ( .C ( clk ), .D ( new_AGEMA_signal_15488 ), .Q ( new_AGEMA_signal_15489 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3991 ( .C ( clk ), .D ( n2797 ), .Q ( new_AGEMA_signal_15491 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3993 ( .C ( clk ), .D ( new_AGEMA_signal_2865 ), .Q ( new_AGEMA_signal_15493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3995 ( .C ( clk ), .D ( new_AGEMA_signal_2866 ), .Q ( new_AGEMA_signal_15495 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3997 ( .C ( clk ), .D ( new_AGEMA_signal_2867 ), .Q ( new_AGEMA_signal_15497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4003 ( .C ( clk ), .D ( new_AGEMA_signal_15502 ), .Q ( new_AGEMA_signal_15503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4009 ( .C ( clk ), .D ( new_AGEMA_signal_15508 ), .Q ( new_AGEMA_signal_15509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4015 ( .C ( clk ), .D ( new_AGEMA_signal_15514 ), .Q ( new_AGEMA_signal_15515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4021 ( .C ( clk ), .D ( new_AGEMA_signal_15520 ), .Q ( new_AGEMA_signal_15521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4035 ( .C ( clk ), .D ( new_AGEMA_signal_15534 ), .Q ( new_AGEMA_signal_15535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4043 ( .C ( clk ), .D ( new_AGEMA_signal_15542 ), .Q ( new_AGEMA_signal_15543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4051 ( .C ( clk ), .D ( new_AGEMA_signal_15550 ), .Q ( new_AGEMA_signal_15551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4059 ( .C ( clk ), .D ( new_AGEMA_signal_15558 ), .Q ( new_AGEMA_signal_15559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4071 ( .C ( clk ), .D ( n2012 ), .Q ( new_AGEMA_signal_15571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4075 ( .C ( clk ), .D ( new_AGEMA_signal_2577 ), .Q ( new_AGEMA_signal_15575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4079 ( .C ( clk ), .D ( new_AGEMA_signal_2578 ), .Q ( new_AGEMA_signal_15579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4083 ( .C ( clk ), .D ( new_AGEMA_signal_2579 ), .Q ( new_AGEMA_signal_15583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4091 ( .C ( clk ), .D ( new_AGEMA_signal_15590 ), .Q ( new_AGEMA_signal_15591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4099 ( .C ( clk ), .D ( new_AGEMA_signal_15598 ), .Q ( new_AGEMA_signal_15599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4107 ( .C ( clk ), .D ( new_AGEMA_signal_15606 ), .Q ( new_AGEMA_signal_15607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4115 ( .C ( clk ), .D ( new_AGEMA_signal_15614 ), .Q ( new_AGEMA_signal_15615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4129 ( .C ( clk ), .D ( new_AGEMA_signal_15628 ), .Q ( new_AGEMA_signal_15629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4135 ( .C ( clk ), .D ( new_AGEMA_signal_15634 ), .Q ( new_AGEMA_signal_15635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4141 ( .C ( clk ), .D ( new_AGEMA_signal_15640 ), .Q ( new_AGEMA_signal_15641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4147 ( .C ( clk ), .D ( new_AGEMA_signal_15646 ), .Q ( new_AGEMA_signal_15647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4151 ( .C ( clk ), .D ( n2652 ), .Q ( new_AGEMA_signal_15651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4155 ( .C ( clk ), .D ( new_AGEMA_signal_2604 ), .Q ( new_AGEMA_signal_15655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4159 ( .C ( clk ), .D ( new_AGEMA_signal_2605 ), .Q ( new_AGEMA_signal_15659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4163 ( .C ( clk ), .D ( new_AGEMA_signal_2606 ), .Q ( new_AGEMA_signal_15663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4171 ( .C ( clk ), .D ( new_AGEMA_signal_15670 ), .Q ( new_AGEMA_signal_15671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4179 ( .C ( clk ), .D ( new_AGEMA_signal_15678 ), .Q ( new_AGEMA_signal_15679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4187 ( .C ( clk ), .D ( new_AGEMA_signal_15686 ), .Q ( new_AGEMA_signal_15687 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4195 ( .C ( clk ), .D ( new_AGEMA_signal_15694 ), .Q ( new_AGEMA_signal_15695 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4199 ( .C ( clk ), .D ( n2143 ), .Q ( new_AGEMA_signal_15699 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4203 ( .C ( clk ), .D ( new_AGEMA_signal_2640 ), .Q ( new_AGEMA_signal_15703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4207 ( .C ( clk ), .D ( new_AGEMA_signal_2641 ), .Q ( new_AGEMA_signal_15707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4211 ( .C ( clk ), .D ( new_AGEMA_signal_2642 ), .Q ( new_AGEMA_signal_15711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4217 ( .C ( clk ), .D ( new_AGEMA_signal_15716 ), .Q ( new_AGEMA_signal_15717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4223 ( .C ( clk ), .D ( new_AGEMA_signal_15722 ), .Q ( new_AGEMA_signal_15723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4229 ( .C ( clk ), .D ( new_AGEMA_signal_15728 ), .Q ( new_AGEMA_signal_15729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4235 ( .C ( clk ), .D ( new_AGEMA_signal_15734 ), .Q ( new_AGEMA_signal_15735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4241 ( .C ( clk ), .D ( new_AGEMA_signal_15740 ), .Q ( new_AGEMA_signal_15741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4247 ( .C ( clk ), .D ( new_AGEMA_signal_15746 ), .Q ( new_AGEMA_signal_15747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4253 ( .C ( clk ), .D ( new_AGEMA_signal_15752 ), .Q ( new_AGEMA_signal_15753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4259 ( .C ( clk ), .D ( new_AGEMA_signal_15758 ), .Q ( new_AGEMA_signal_15759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4265 ( .C ( clk ), .D ( new_AGEMA_signal_15764 ), .Q ( new_AGEMA_signal_15765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4271 ( .C ( clk ), .D ( new_AGEMA_signal_15770 ), .Q ( new_AGEMA_signal_15771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4277 ( .C ( clk ), .D ( new_AGEMA_signal_15776 ), .Q ( new_AGEMA_signal_15777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4283 ( .C ( clk ), .D ( new_AGEMA_signal_15782 ), .Q ( new_AGEMA_signal_15783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4289 ( .C ( clk ), .D ( new_AGEMA_signal_15788 ), .Q ( new_AGEMA_signal_15789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4295 ( .C ( clk ), .D ( new_AGEMA_signal_15794 ), .Q ( new_AGEMA_signal_15795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4301 ( .C ( clk ), .D ( new_AGEMA_signal_15800 ), .Q ( new_AGEMA_signal_15801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4307 ( .C ( clk ), .D ( new_AGEMA_signal_15806 ), .Q ( new_AGEMA_signal_15807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4313 ( .C ( clk ), .D ( new_AGEMA_signal_15812 ), .Q ( new_AGEMA_signal_15813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4319 ( .C ( clk ), .D ( new_AGEMA_signal_15818 ), .Q ( new_AGEMA_signal_15819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4325 ( .C ( clk ), .D ( new_AGEMA_signal_15824 ), .Q ( new_AGEMA_signal_15825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4331 ( .C ( clk ), .D ( new_AGEMA_signal_15830 ), .Q ( new_AGEMA_signal_15831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4335 ( .C ( clk ), .D ( n2297 ), .Q ( new_AGEMA_signal_15835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4339 ( .C ( clk ), .D ( new_AGEMA_signal_2709 ), .Q ( new_AGEMA_signal_15839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4343 ( .C ( clk ), .D ( new_AGEMA_signal_2710 ), .Q ( new_AGEMA_signal_15843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4347 ( .C ( clk ), .D ( new_AGEMA_signal_2711 ), .Q ( new_AGEMA_signal_15847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4355 ( .C ( clk ), .D ( new_AGEMA_signal_15854 ), .Q ( new_AGEMA_signal_15855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4363 ( .C ( clk ), .D ( new_AGEMA_signal_15862 ), .Q ( new_AGEMA_signal_15863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4371 ( .C ( clk ), .D ( new_AGEMA_signal_15870 ), .Q ( new_AGEMA_signal_15871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4379 ( .C ( clk ), .D ( new_AGEMA_signal_15878 ), .Q ( new_AGEMA_signal_15879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4383 ( .C ( clk ), .D ( n2336 ), .Q ( new_AGEMA_signal_15883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4387 ( .C ( clk ), .D ( new_AGEMA_signal_2994 ), .Q ( new_AGEMA_signal_15887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4391 ( .C ( clk ), .D ( new_AGEMA_signal_2995 ), .Q ( new_AGEMA_signal_15891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4395 ( .C ( clk ), .D ( new_AGEMA_signal_2996 ), .Q ( new_AGEMA_signal_15895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4401 ( .C ( clk ), .D ( new_AGEMA_signal_15900 ), .Q ( new_AGEMA_signal_15901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4407 ( .C ( clk ), .D ( new_AGEMA_signal_15906 ), .Q ( new_AGEMA_signal_15907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4413 ( .C ( clk ), .D ( new_AGEMA_signal_15912 ), .Q ( new_AGEMA_signal_15913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4419 ( .C ( clk ), .D ( new_AGEMA_signal_15918 ), .Q ( new_AGEMA_signal_15919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4427 ( .C ( clk ), .D ( new_AGEMA_signal_15926 ), .Q ( new_AGEMA_signal_15927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4435 ( .C ( clk ), .D ( new_AGEMA_signal_15934 ), .Q ( new_AGEMA_signal_15935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4443 ( .C ( clk ), .D ( new_AGEMA_signal_15942 ), .Q ( new_AGEMA_signal_15943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4451 ( .C ( clk ), .D ( new_AGEMA_signal_15950 ), .Q ( new_AGEMA_signal_15951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4465 ( .C ( clk ), .D ( new_AGEMA_signal_15964 ), .Q ( new_AGEMA_signal_15965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4471 ( .C ( clk ), .D ( new_AGEMA_signal_15970 ), .Q ( new_AGEMA_signal_15971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4477 ( .C ( clk ), .D ( new_AGEMA_signal_15976 ), .Q ( new_AGEMA_signal_15977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4483 ( .C ( clk ), .D ( new_AGEMA_signal_15982 ), .Q ( new_AGEMA_signal_15983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4505 ( .C ( clk ), .D ( new_AGEMA_signal_16004 ), .Q ( new_AGEMA_signal_16005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4511 ( .C ( clk ), .D ( new_AGEMA_signal_16010 ), .Q ( new_AGEMA_signal_16011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4517 ( .C ( clk ), .D ( new_AGEMA_signal_16016 ), .Q ( new_AGEMA_signal_16017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4523 ( .C ( clk ), .D ( new_AGEMA_signal_16022 ), .Q ( new_AGEMA_signal_16023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4529 ( .C ( clk ), .D ( new_AGEMA_signal_16028 ), .Q ( new_AGEMA_signal_16029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4535 ( .C ( clk ), .D ( new_AGEMA_signal_16034 ), .Q ( new_AGEMA_signal_16035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4541 ( .C ( clk ), .D ( new_AGEMA_signal_16040 ), .Q ( new_AGEMA_signal_16041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4547 ( .C ( clk ), .D ( new_AGEMA_signal_16046 ), .Q ( new_AGEMA_signal_16047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4555 ( .C ( clk ), .D ( new_AGEMA_signal_16054 ), .Q ( new_AGEMA_signal_16055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4563 ( .C ( clk ), .D ( new_AGEMA_signal_16062 ), .Q ( new_AGEMA_signal_16063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4571 ( .C ( clk ), .D ( new_AGEMA_signal_16070 ), .Q ( new_AGEMA_signal_16071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4579 ( .C ( clk ), .D ( new_AGEMA_signal_16078 ), .Q ( new_AGEMA_signal_16079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4587 ( .C ( clk ), .D ( new_AGEMA_signal_16086 ), .Q ( new_AGEMA_signal_16087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4595 ( .C ( clk ), .D ( new_AGEMA_signal_16094 ), .Q ( new_AGEMA_signal_16095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4603 ( .C ( clk ), .D ( new_AGEMA_signal_16102 ), .Q ( new_AGEMA_signal_16103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4611 ( .C ( clk ), .D ( new_AGEMA_signal_16110 ), .Q ( new_AGEMA_signal_16111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4617 ( .C ( clk ), .D ( new_AGEMA_signal_16116 ), .Q ( new_AGEMA_signal_16117 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4623 ( .C ( clk ), .D ( new_AGEMA_signal_16122 ), .Q ( new_AGEMA_signal_16123 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4629 ( .C ( clk ), .D ( new_AGEMA_signal_16128 ), .Q ( new_AGEMA_signal_16129 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4635 ( .C ( clk ), .D ( new_AGEMA_signal_16134 ), .Q ( new_AGEMA_signal_16135 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4641 ( .C ( clk ), .D ( new_AGEMA_signal_16140 ), .Q ( new_AGEMA_signal_16141 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4647 ( .C ( clk ), .D ( new_AGEMA_signal_16146 ), .Q ( new_AGEMA_signal_16147 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4653 ( .C ( clk ), .D ( new_AGEMA_signal_16152 ), .Q ( new_AGEMA_signal_16153 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4659 ( .C ( clk ), .D ( new_AGEMA_signal_16158 ), .Q ( new_AGEMA_signal_16159 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4671 ( .C ( clk ), .D ( n2658 ), .Q ( new_AGEMA_signal_16171 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4675 ( .C ( clk ), .D ( new_AGEMA_signal_2550 ), .Q ( new_AGEMA_signal_16175 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4679 ( .C ( clk ), .D ( new_AGEMA_signal_2551 ), .Q ( new_AGEMA_signal_16179 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4683 ( .C ( clk ), .D ( new_AGEMA_signal_2552 ), .Q ( new_AGEMA_signal_16183 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4687 ( .C ( clk ), .D ( n2698 ), .Q ( new_AGEMA_signal_16187 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4691 ( .C ( clk ), .D ( new_AGEMA_signal_2835 ), .Q ( new_AGEMA_signal_16191 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4695 ( .C ( clk ), .D ( new_AGEMA_signal_2836 ), .Q ( new_AGEMA_signal_16195 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4699 ( .C ( clk ), .D ( new_AGEMA_signal_2837 ), .Q ( new_AGEMA_signal_16199 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4703 ( .C ( clk ), .D ( n2800 ), .Q ( new_AGEMA_signal_16203 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4707 ( .C ( clk ), .D ( new_AGEMA_signal_2859 ), .Q ( new_AGEMA_signal_16207 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4711 ( .C ( clk ), .D ( new_AGEMA_signal_2860 ), .Q ( new_AGEMA_signal_16211 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4715 ( .C ( clk ), .D ( new_AGEMA_signal_2861 ), .Q ( new_AGEMA_signal_16215 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4727 ( .C ( clk ), .D ( n1936 ), .Q ( new_AGEMA_signal_16227 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4733 ( .C ( clk ), .D ( new_AGEMA_signal_2526 ), .Q ( new_AGEMA_signal_16233 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4739 ( .C ( clk ), .D ( new_AGEMA_signal_2527 ), .Q ( new_AGEMA_signal_16239 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4745 ( .C ( clk ), .D ( new_AGEMA_signal_2528 ), .Q ( new_AGEMA_signal_16245 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4777 ( .C ( clk ), .D ( new_AGEMA_signal_16276 ), .Q ( new_AGEMA_signal_16277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4785 ( .C ( clk ), .D ( new_AGEMA_signal_16284 ), .Q ( new_AGEMA_signal_16285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4793 ( .C ( clk ), .D ( new_AGEMA_signal_16292 ), .Q ( new_AGEMA_signal_16293 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4801 ( .C ( clk ), .D ( new_AGEMA_signal_16300 ), .Q ( new_AGEMA_signal_16301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4809 ( .C ( clk ), .D ( new_AGEMA_signal_16308 ), .Q ( new_AGEMA_signal_16309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4817 ( .C ( clk ), .D ( new_AGEMA_signal_16316 ), .Q ( new_AGEMA_signal_16317 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4825 ( .C ( clk ), .D ( new_AGEMA_signal_16324 ), .Q ( new_AGEMA_signal_16325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4833 ( .C ( clk ), .D ( new_AGEMA_signal_16332 ), .Q ( new_AGEMA_signal_16333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4841 ( .C ( clk ), .D ( new_AGEMA_signal_16340 ), .Q ( new_AGEMA_signal_16341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4849 ( .C ( clk ), .D ( new_AGEMA_signal_16348 ), .Q ( new_AGEMA_signal_16349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4857 ( .C ( clk ), .D ( new_AGEMA_signal_16356 ), .Q ( new_AGEMA_signal_16357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4865 ( .C ( clk ), .D ( new_AGEMA_signal_16364 ), .Q ( new_AGEMA_signal_16365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4873 ( .C ( clk ), .D ( new_AGEMA_signal_16372 ), .Q ( new_AGEMA_signal_16373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4881 ( .C ( clk ), .D ( new_AGEMA_signal_16380 ), .Q ( new_AGEMA_signal_16381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4889 ( .C ( clk ), .D ( new_AGEMA_signal_16388 ), .Q ( new_AGEMA_signal_16389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4897 ( .C ( clk ), .D ( new_AGEMA_signal_16396 ), .Q ( new_AGEMA_signal_16397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4903 ( .C ( clk ), .D ( n2099 ), .Q ( new_AGEMA_signal_16403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4909 ( .C ( clk ), .D ( new_AGEMA_signal_2613 ), .Q ( new_AGEMA_signal_16409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4915 ( .C ( clk ), .D ( new_AGEMA_signal_2614 ), .Q ( new_AGEMA_signal_16415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4921 ( .C ( clk ), .D ( new_AGEMA_signal_2615 ), .Q ( new_AGEMA_signal_16421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4931 ( .C ( clk ), .D ( new_AGEMA_signal_16430 ), .Q ( new_AGEMA_signal_16431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4941 ( .C ( clk ), .D ( new_AGEMA_signal_16440 ), .Q ( new_AGEMA_signal_16441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4951 ( .C ( clk ), .D ( new_AGEMA_signal_16450 ), .Q ( new_AGEMA_signal_16451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4961 ( .C ( clk ), .D ( new_AGEMA_signal_16460 ), .Q ( new_AGEMA_signal_16461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4969 ( .C ( clk ), .D ( new_AGEMA_signal_16468 ), .Q ( new_AGEMA_signal_16469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4977 ( .C ( clk ), .D ( new_AGEMA_signal_16476 ), .Q ( new_AGEMA_signal_16477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4985 ( .C ( clk ), .D ( new_AGEMA_signal_16484 ), .Q ( new_AGEMA_signal_16485 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4993 ( .C ( clk ), .D ( new_AGEMA_signal_16492 ), .Q ( new_AGEMA_signal_16493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5001 ( .C ( clk ), .D ( new_AGEMA_signal_16500 ), .Q ( new_AGEMA_signal_16501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5009 ( .C ( clk ), .D ( new_AGEMA_signal_16508 ), .Q ( new_AGEMA_signal_16509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5017 ( .C ( clk ), .D ( new_AGEMA_signal_16516 ), .Q ( new_AGEMA_signal_16517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5025 ( .C ( clk ), .D ( new_AGEMA_signal_16524 ), .Q ( new_AGEMA_signal_16525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5033 ( .C ( clk ), .D ( new_AGEMA_signal_16532 ), .Q ( new_AGEMA_signal_16533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5041 ( .C ( clk ), .D ( new_AGEMA_signal_16540 ), .Q ( new_AGEMA_signal_16541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5049 ( .C ( clk ), .D ( new_AGEMA_signal_16548 ), .Q ( new_AGEMA_signal_16549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5057 ( .C ( clk ), .D ( new_AGEMA_signal_16556 ), .Q ( new_AGEMA_signal_16557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5087 ( .C ( clk ), .D ( n2301 ), .Q ( new_AGEMA_signal_16587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5093 ( .C ( clk ), .D ( new_AGEMA_signal_2715 ), .Q ( new_AGEMA_signal_16593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5099 ( .C ( clk ), .D ( new_AGEMA_signal_2716 ), .Q ( new_AGEMA_signal_16599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5105 ( .C ( clk ), .D ( new_AGEMA_signal_2717 ), .Q ( new_AGEMA_signal_16605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5131 ( .C ( clk ), .D ( new_AGEMA_signal_16630 ), .Q ( new_AGEMA_signal_16631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5141 ( .C ( clk ), .D ( new_AGEMA_signal_16640 ), .Q ( new_AGEMA_signal_16641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5151 ( .C ( clk ), .D ( new_AGEMA_signal_16650 ), .Q ( new_AGEMA_signal_16651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5161 ( .C ( clk ), .D ( new_AGEMA_signal_16660 ), .Q ( new_AGEMA_signal_16661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5169 ( .C ( clk ), .D ( new_AGEMA_signal_16668 ), .Q ( new_AGEMA_signal_16669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5177 ( .C ( clk ), .D ( new_AGEMA_signal_16676 ), .Q ( new_AGEMA_signal_16677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5185 ( .C ( clk ), .D ( new_AGEMA_signal_16684 ), .Q ( new_AGEMA_signal_16685 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5193 ( .C ( clk ), .D ( new_AGEMA_signal_16692 ), .Q ( new_AGEMA_signal_16693 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5225 ( .C ( clk ), .D ( new_AGEMA_signal_16724 ), .Q ( new_AGEMA_signal_16725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5233 ( .C ( clk ), .D ( new_AGEMA_signal_16732 ), .Q ( new_AGEMA_signal_16733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5241 ( .C ( clk ), .D ( new_AGEMA_signal_16740 ), .Q ( new_AGEMA_signal_16741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5249 ( .C ( clk ), .D ( new_AGEMA_signal_16748 ), .Q ( new_AGEMA_signal_16749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5257 ( .C ( clk ), .D ( new_AGEMA_signal_16756 ), .Q ( new_AGEMA_signal_16757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5265 ( .C ( clk ), .D ( new_AGEMA_signal_16764 ), .Q ( new_AGEMA_signal_16765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5273 ( .C ( clk ), .D ( new_AGEMA_signal_16772 ), .Q ( new_AGEMA_signal_16773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5281 ( .C ( clk ), .D ( new_AGEMA_signal_16780 ), .Q ( new_AGEMA_signal_16781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5287 ( .C ( clk ), .D ( new_AGEMA_signal_14102 ), .Q ( new_AGEMA_signal_16787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5293 ( .C ( clk ), .D ( new_AGEMA_signal_14106 ), .Q ( new_AGEMA_signal_16793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5299 ( .C ( clk ), .D ( new_AGEMA_signal_14110 ), .Q ( new_AGEMA_signal_16799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5305 ( .C ( clk ), .D ( new_AGEMA_signal_14114 ), .Q ( new_AGEMA_signal_16805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5329 ( .C ( clk ), .D ( new_AGEMA_signal_16828 ), .Q ( new_AGEMA_signal_16829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5337 ( .C ( clk ), .D ( new_AGEMA_signal_16836 ), .Q ( new_AGEMA_signal_16837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5345 ( .C ( clk ), .D ( new_AGEMA_signal_16844 ), .Q ( new_AGEMA_signal_16845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5353 ( .C ( clk ), .D ( new_AGEMA_signal_16852 ), .Q ( new_AGEMA_signal_16853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5455 ( .C ( clk ), .D ( new_AGEMA_signal_14550 ), .Q ( new_AGEMA_signal_16955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5463 ( .C ( clk ), .D ( new_AGEMA_signal_14554 ), .Q ( new_AGEMA_signal_16963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5471 ( .C ( clk ), .D ( new_AGEMA_signal_14558 ), .Q ( new_AGEMA_signal_16971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5479 ( .C ( clk ), .D ( new_AGEMA_signal_14562 ), .Q ( new_AGEMA_signal_16979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5527 ( .C ( clk ), .D ( n2102 ), .Q ( new_AGEMA_signal_17027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5535 ( .C ( clk ), .D ( new_AGEMA_signal_2625 ), .Q ( new_AGEMA_signal_17035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5543 ( .C ( clk ), .D ( new_AGEMA_signal_2626 ), .Q ( new_AGEMA_signal_17043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5551 ( .C ( clk ), .D ( new_AGEMA_signal_2627 ), .Q ( new_AGEMA_signal_17051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5559 ( .C ( clk ), .D ( new_AGEMA_signal_13940 ), .Q ( new_AGEMA_signal_17059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5567 ( .C ( clk ), .D ( new_AGEMA_signal_13942 ), .Q ( new_AGEMA_signal_17067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5575 ( .C ( clk ), .D ( new_AGEMA_signal_13944 ), .Q ( new_AGEMA_signal_17075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5583 ( .C ( clk ), .D ( new_AGEMA_signal_13946 ), .Q ( new_AGEMA_signal_17083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5593 ( .C ( clk ), .D ( new_AGEMA_signal_17092 ), .Q ( new_AGEMA_signal_17093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5603 ( .C ( clk ), .D ( new_AGEMA_signal_17102 ), .Q ( new_AGEMA_signal_17103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5613 ( .C ( clk ), .D ( new_AGEMA_signal_17112 ), .Q ( new_AGEMA_signal_17113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5623 ( .C ( clk ), .D ( new_AGEMA_signal_17122 ), .Q ( new_AGEMA_signal_17123 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5631 ( .C ( clk ), .D ( new_AGEMA_signal_14310 ), .Q ( new_AGEMA_signal_17131 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5639 ( .C ( clk ), .D ( new_AGEMA_signal_14314 ), .Q ( new_AGEMA_signal_17139 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5647 ( .C ( clk ), .D ( new_AGEMA_signal_14318 ), .Q ( new_AGEMA_signal_17147 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5655 ( .C ( clk ), .D ( new_AGEMA_signal_14322 ), .Q ( new_AGEMA_signal_17155 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5727 ( .C ( clk ), .D ( n2367 ), .Q ( new_AGEMA_signal_17227 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5735 ( .C ( clk ), .D ( new_AGEMA_signal_2316 ), .Q ( new_AGEMA_signal_17235 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5743 ( .C ( clk ), .D ( new_AGEMA_signal_2317 ), .Q ( new_AGEMA_signal_17243 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5751 ( .C ( clk ), .D ( new_AGEMA_signal_2318 ), .Q ( new_AGEMA_signal_17251 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5791 ( .C ( clk ), .D ( n2591 ), .Q ( new_AGEMA_signal_17291 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5799 ( .C ( clk ), .D ( new_AGEMA_signal_2808 ), .Q ( new_AGEMA_signal_17299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5807 ( .C ( clk ), .D ( new_AGEMA_signal_2809 ), .Q ( new_AGEMA_signal_17307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5815 ( .C ( clk ), .D ( new_AGEMA_signal_2810 ), .Q ( new_AGEMA_signal_17315 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5967 ( .C ( clk ), .D ( n2105 ), .Q ( new_AGEMA_signal_17467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5977 ( .C ( clk ), .D ( new_AGEMA_signal_2610 ), .Q ( new_AGEMA_signal_17477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5987 ( .C ( clk ), .D ( new_AGEMA_signal_2611 ), .Q ( new_AGEMA_signal_17487 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5997 ( .C ( clk ), .D ( new_AGEMA_signal_2612 ), .Q ( new_AGEMA_signal_17497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6327 ( .C ( clk ), .D ( n2106 ), .Q ( new_AGEMA_signal_17827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6339 ( .C ( clk ), .D ( new_AGEMA_signal_2187 ), .Q ( new_AGEMA_signal_17839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6351 ( .C ( clk ), .D ( new_AGEMA_signal_2188 ), .Q ( new_AGEMA_signal_17851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6363 ( .C ( clk ), .D ( new_AGEMA_signal_2189 ), .Q ( new_AGEMA_signal_17863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6377 ( .C ( clk ), .D ( new_AGEMA_signal_17876 ), .Q ( new_AGEMA_signal_17877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6391 ( .C ( clk ), .D ( new_AGEMA_signal_17890 ), .Q ( new_AGEMA_signal_17891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6405 ( .C ( clk ), .D ( new_AGEMA_signal_17904 ), .Q ( new_AGEMA_signal_17905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6419 ( .C ( clk ), .D ( new_AGEMA_signal_17918 ), .Q ( new_AGEMA_signal_17919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6465 ( .C ( clk ), .D ( new_AGEMA_signal_17964 ), .Q ( new_AGEMA_signal_17965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6479 ( .C ( clk ), .D ( new_AGEMA_signal_17978 ), .Q ( new_AGEMA_signal_17979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6493 ( .C ( clk ), .D ( new_AGEMA_signal_17992 ), .Q ( new_AGEMA_signal_17993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6507 ( .C ( clk ), .D ( new_AGEMA_signal_18006 ), .Q ( new_AGEMA_signal_18007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6609 ( .C ( clk ), .D ( new_AGEMA_signal_18108 ), .Q ( new_AGEMA_signal_18109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6625 ( .C ( clk ), .D ( new_AGEMA_signal_18124 ), .Q ( new_AGEMA_signal_18125 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6641 ( .C ( clk ), .D ( new_AGEMA_signal_18140 ), .Q ( new_AGEMA_signal_18141 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6657 ( .C ( clk ), .D ( new_AGEMA_signal_18156 ), .Q ( new_AGEMA_signal_18157 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6697 ( .C ( clk ), .D ( new_AGEMA_signal_18196 ), .Q ( new_AGEMA_signal_18197 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6713 ( .C ( clk ), .D ( new_AGEMA_signal_18212 ), .Q ( new_AGEMA_signal_18213 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6729 ( .C ( clk ), .D ( new_AGEMA_signal_18228 ), .Q ( new_AGEMA_signal_18229 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6745 ( .C ( clk ), .D ( new_AGEMA_signal_18244 ), .Q ( new_AGEMA_signal_18245 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6895 ( .C ( clk ), .D ( n2155 ), .Q ( new_AGEMA_signal_18395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6911 ( .C ( clk ), .D ( new_AGEMA_signal_2193 ), .Q ( new_AGEMA_signal_18411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6927 ( .C ( clk ), .D ( new_AGEMA_signal_2194 ), .Q ( new_AGEMA_signal_18427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6943 ( .C ( clk ), .D ( new_AGEMA_signal_2195 ), .Q ( new_AGEMA_signal_18443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7001 ( .C ( clk ), .D ( new_AGEMA_signal_18500 ), .Q ( new_AGEMA_signal_18501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7019 ( .C ( clk ), .D ( new_AGEMA_signal_18518 ), .Q ( new_AGEMA_signal_18519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7037 ( .C ( clk ), .D ( new_AGEMA_signal_18536 ), .Q ( new_AGEMA_signal_18537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7055 ( .C ( clk ), .D ( new_AGEMA_signal_18554 ), .Q ( new_AGEMA_signal_18555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7201 ( .C ( clk ), .D ( new_AGEMA_signal_18700 ), .Q ( new_AGEMA_signal_18701 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7221 ( .C ( clk ), .D ( new_AGEMA_signal_18720 ), .Q ( new_AGEMA_signal_18721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7241 ( .C ( clk ), .D ( new_AGEMA_signal_18740 ), .Q ( new_AGEMA_signal_18741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7261 ( .C ( clk ), .D ( new_AGEMA_signal_18760 ), .Q ( new_AGEMA_signal_18761 ) ) ;

    /* cells in depth 10 */
    nor_HPC1 #(.security_order(3), .pipeline(1)) U1983 ( .ina ({new_AGEMA_signal_13802, new_AGEMA_signal_13798, new_AGEMA_signal_13794, new_AGEMA_signal_13790}), .inb ({new_AGEMA_signal_2531, new_AGEMA_signal_2530, new_AGEMA_signal_2529, n1928}), .clk ( clk ), .rnd ({Fresh[5759], Fresh[5758], Fresh[5757], Fresh[5756], Fresh[5755], Fresh[5754], Fresh[5753], Fresh[5752], Fresh[5751], Fresh[5750]}), .outt ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, new_AGEMA_signal_2871, n1934}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U1998 ( .ina ({new_AGEMA_signal_2534, new_AGEMA_signal_2533, new_AGEMA_signal_2532, n1931}), .inb ({new_AGEMA_signal_13818, new_AGEMA_signal_13814, new_AGEMA_signal_13810, new_AGEMA_signal_13806}), .clk ( clk ), .rnd ({Fresh[5769], Fresh[5768], Fresh[5767], Fresh[5766], Fresh[5765], Fresh[5764], Fresh[5763], Fresh[5762], Fresh[5761], Fresh[5760]}), .outt ({new_AGEMA_signal_2876, new_AGEMA_signal_2875, new_AGEMA_signal_2874, n1932}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2015 ( .ina ({new_AGEMA_signal_2537, new_AGEMA_signal_2536, new_AGEMA_signal_2535, n1939}), .inb ({new_AGEMA_signal_13826, new_AGEMA_signal_13824, new_AGEMA_signal_13822, new_AGEMA_signal_13820}), .clk ( clk ), .rnd ({Fresh[5779], Fresh[5778], Fresh[5777], Fresh[5776], Fresh[5775], Fresh[5774], Fresh[5773], Fresh[5772], Fresh[5771], Fresh[5770]}), .outt ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, new_AGEMA_signal_2877, n1940}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2033 ( .ina ({new_AGEMA_signal_2540, new_AGEMA_signal_2539, new_AGEMA_signal_2538, n1948}), .inb ({new_AGEMA_signal_2543, new_AGEMA_signal_2542, new_AGEMA_signal_2541, n1947}), .clk ( clk ), .rnd ({Fresh[5789], Fresh[5788], Fresh[5787], Fresh[5786], Fresh[5785], Fresh[5784], Fresh[5783], Fresh[5782], Fresh[5781], Fresh[5780]}), .outt ({new_AGEMA_signal_2882, new_AGEMA_signal_2881, new_AGEMA_signal_2880, n1961}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2050 ( .ina ({new_AGEMA_signal_2546, new_AGEMA_signal_2545, new_AGEMA_signal_2544, n1954}), .inb ({new_AGEMA_signal_2549, new_AGEMA_signal_2548, new_AGEMA_signal_2547, n1953}), .clk ( clk ), .rnd ({Fresh[5799], Fresh[5798], Fresh[5797], Fresh[5796], Fresh[5795], Fresh[5794], Fresh[5793], Fresh[5792], Fresh[5791], Fresh[5790]}), .outt ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, new_AGEMA_signal_2883, n1955}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2066 ( .ina ({new_AGEMA_signal_13834, new_AGEMA_signal_13832, new_AGEMA_signal_13830, new_AGEMA_signal_13828}), .inb ({new_AGEMA_signal_2084, new_AGEMA_signal_2083, new_AGEMA_signal_2082, n1965}), .clk ( clk ), .rnd ({Fresh[5809], Fresh[5808], Fresh[5807], Fresh[5806], Fresh[5805], Fresh[5804], Fresh[5803], Fresh[5802], Fresh[5801], Fresh[5800]}), .outt ({new_AGEMA_signal_2555, new_AGEMA_signal_2554, new_AGEMA_signal_2553, n1967}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2085 ( .ina ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, new_AGEMA_signal_2889, n1970}), .inb ({new_AGEMA_signal_2561, new_AGEMA_signal_2560, new_AGEMA_signal_2559, n1969}), .clk ( clk ), .rnd ({Fresh[5819], Fresh[5818], Fresh[5817], Fresh[5816], Fresh[5815], Fresh[5814], Fresh[5813], Fresh[5812], Fresh[5811], Fresh[5810]}), .outt ({new_AGEMA_signal_3125, new_AGEMA_signal_3124, new_AGEMA_signal_3123, n1984}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2103 ( .ina ({new_AGEMA_signal_13850, new_AGEMA_signal_13846, new_AGEMA_signal_13842, new_AGEMA_signal_13838}), .inb ({new_AGEMA_signal_2567, new_AGEMA_signal_2566, new_AGEMA_signal_2565, n1975}), .clk ( clk ), .rnd ({Fresh[5829], Fresh[5828], Fresh[5827], Fresh[5826], Fresh[5825], Fresh[5824], Fresh[5823], Fresh[5822], Fresh[5821], Fresh[5820]}), .outt ({new_AGEMA_signal_2894, new_AGEMA_signal_2893, new_AGEMA_signal_2892, n1977}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2108 ( .ina ({new_AGEMA_signal_13858, new_AGEMA_signal_13856, new_AGEMA_signal_13854, new_AGEMA_signal_13852}), .inb ({new_AGEMA_signal_2570, new_AGEMA_signal_2569, new_AGEMA_signal_2568, n1980}), .clk ( clk ), .rnd ({Fresh[5839], Fresh[5838], Fresh[5837], Fresh[5836], Fresh[5835], Fresh[5834], Fresh[5833], Fresh[5832], Fresh[5831], Fresh[5830]}), .outt ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, new_AGEMA_signal_2895, n1981}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2115 ( .ina ({new_AGEMA_signal_13874, new_AGEMA_signal_13870, new_AGEMA_signal_13866, new_AGEMA_signal_13862}), .inb ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, new_AGEMA_signal_2103, n1986}), .clk ( clk ), .rnd ({Fresh[5849], Fresh[5848], Fresh[5847], Fresh[5846], Fresh[5845], Fresh[5844], Fresh[5843], Fresh[5842], Fresh[5841], Fresh[5840]}), .outt ({new_AGEMA_signal_2573, new_AGEMA_signal_2572, new_AGEMA_signal_2571, n1987}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2127 ( .ina ({new_AGEMA_signal_2576, new_AGEMA_signal_2575, new_AGEMA_signal_2574, n1997}), .inb ({new_AGEMA_signal_13882, new_AGEMA_signal_13880, new_AGEMA_signal_13878, new_AGEMA_signal_13876}), .clk ( clk ), .rnd ({Fresh[5859], Fresh[5858], Fresh[5857], Fresh[5856], Fresh[5855], Fresh[5854], Fresh[5853], Fresh[5852], Fresh[5851], Fresh[5850]}), .outt ({new_AGEMA_signal_2900, new_AGEMA_signal_2899, new_AGEMA_signal_2898, n1998}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2146 ( .ina ({new_AGEMA_signal_13898, new_AGEMA_signal_13894, new_AGEMA_signal_13890, new_AGEMA_signal_13886}), .inb ({new_AGEMA_signal_2582, new_AGEMA_signal_2581, new_AGEMA_signal_2580, n2007}), .clk ( clk ), .rnd ({Fresh[5869], Fresh[5868], Fresh[5867], Fresh[5866], Fresh[5865], Fresh[5864], Fresh[5863], Fresh[5862], Fresh[5861], Fresh[5860]}), .outt ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, new_AGEMA_signal_2901, n2010}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2162 ( .ina ({new_AGEMA_signal_13914, new_AGEMA_signal_13910, new_AGEMA_signal_13906, new_AGEMA_signal_13902}), .inb ({new_AGEMA_signal_2126, new_AGEMA_signal_2125, new_AGEMA_signal_2124, n2021}), .clk ( clk ), .rnd ({Fresh[5879], Fresh[5878], Fresh[5877], Fresh[5876], Fresh[5875], Fresh[5874], Fresh[5873], Fresh[5872], Fresh[5871], Fresh[5870]}), .outt ({new_AGEMA_signal_2585, new_AGEMA_signal_2584, new_AGEMA_signal_2583, n2024}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2177 ( .ina ({new_AGEMA_signal_13922, new_AGEMA_signal_13920, new_AGEMA_signal_13918, new_AGEMA_signal_13916}), .inb ({new_AGEMA_signal_2588, new_AGEMA_signal_2587, new_AGEMA_signal_2586, n2032}), .clk ( clk ), .rnd ({Fresh[5889], Fresh[5888], Fresh[5887], Fresh[5886], Fresh[5885], Fresh[5884], Fresh[5883], Fresh[5882], Fresh[5881], Fresh[5880]}), .outt ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, new_AGEMA_signal_2907, n2035}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2186 ( .ina ({new_AGEMA_signal_2591, new_AGEMA_signal_2590, new_AGEMA_signal_2589, n2041}), .inb ({new_AGEMA_signal_13930, new_AGEMA_signal_13928, new_AGEMA_signal_13926, new_AGEMA_signal_13924}), .clk ( clk ), .rnd ({Fresh[5899], Fresh[5898], Fresh[5897], Fresh[5896], Fresh[5895], Fresh[5894], Fresh[5893], Fresh[5892], Fresh[5891], Fresh[5890]}), .outt ({new_AGEMA_signal_2912, new_AGEMA_signal_2911, new_AGEMA_signal_2910, n2054}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2190 ( .ina ({new_AGEMA_signal_13938, new_AGEMA_signal_13936, new_AGEMA_signal_13934, new_AGEMA_signal_13932}), .inb ({new_AGEMA_signal_2594, new_AGEMA_signal_2593, new_AGEMA_signal_2592, n2043}), .clk ( clk ), .rnd ({Fresh[5909], Fresh[5908], Fresh[5907], Fresh[5906], Fresh[5905], Fresh[5904], Fresh[5903], Fresh[5902], Fresh[5901], Fresh[5900]}), .outt ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, new_AGEMA_signal_2913, n2048}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2195 ( .ina ({new_AGEMA_signal_2597, new_AGEMA_signal_2596, new_AGEMA_signal_2595, n2046}), .inb ({new_AGEMA_signal_13946, new_AGEMA_signal_13944, new_AGEMA_signal_13942, new_AGEMA_signal_13940}), .clk ( clk ), .rnd ({Fresh[5919], Fresh[5918], Fresh[5917], Fresh[5916], Fresh[5915], Fresh[5914], Fresh[5913], Fresh[5912], Fresh[5911], Fresh[5910]}), .outt ({new_AGEMA_signal_2918, new_AGEMA_signal_2917, new_AGEMA_signal_2916, n2047}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2206 ( .ina ({new_AGEMA_signal_2600, new_AGEMA_signal_2599, new_AGEMA_signal_2598, n2058}), .inb ({new_AGEMA_signal_13962, new_AGEMA_signal_13958, new_AGEMA_signal_13954, new_AGEMA_signal_13950}), .clk ( clk ), .rnd ({Fresh[5929], Fresh[5928], Fresh[5927], Fresh[5926], Fresh[5925], Fresh[5924], Fresh[5923], Fresh[5922], Fresh[5921], Fresh[5920]}), .outt ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, new_AGEMA_signal_2919, n2059}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2213 ( .ina ({new_AGEMA_signal_2603, new_AGEMA_signal_2602, new_AGEMA_signal_2601, n2063}), .inb ({new_AGEMA_signal_13978, new_AGEMA_signal_13974, new_AGEMA_signal_13970, new_AGEMA_signal_13966}), .clk ( clk ), .rnd ({Fresh[5939], Fresh[5938], Fresh[5937], Fresh[5936], Fresh[5935], Fresh[5934], Fresh[5933], Fresh[5932], Fresh[5931], Fresh[5930]}), .outt ({new_AGEMA_signal_2924, new_AGEMA_signal_2923, new_AGEMA_signal_2922, n2064}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2229 ( .ina ({new_AGEMA_signal_2609, new_AGEMA_signal_2608, new_AGEMA_signal_2607, n2076}), .inb ({new_AGEMA_signal_13994, new_AGEMA_signal_13990, new_AGEMA_signal_13986, new_AGEMA_signal_13982}), .clk ( clk ), .rnd ({Fresh[5949], Fresh[5948], Fresh[5947], Fresh[5946], Fresh[5945], Fresh[5944], Fresh[5943], Fresh[5942], Fresh[5941], Fresh[5940]}), .outt ({new_AGEMA_signal_2927, new_AGEMA_signal_2926, new_AGEMA_signal_2925, n2077}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2249 ( .ina ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, new_AGEMA_signal_2619, n2090}), .inb ({new_AGEMA_signal_14002, new_AGEMA_signal_14000, new_AGEMA_signal_13998, new_AGEMA_signal_13996}), .clk ( clk ), .rnd ({Fresh[5959], Fresh[5958], Fresh[5957], Fresh[5956], Fresh[5955], Fresh[5954], Fresh[5953], Fresh[5952], Fresh[5951], Fresh[5950]}), .outt ({new_AGEMA_signal_2930, new_AGEMA_signal_2929, new_AGEMA_signal_2928, n2158}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2255 ( .ina ({new_AGEMA_signal_2624, new_AGEMA_signal_2623, new_AGEMA_signal_2622, n2093}), .inb ({new_AGEMA_signal_14010, new_AGEMA_signal_14008, new_AGEMA_signal_14006, new_AGEMA_signal_14004}), .clk ( clk ), .rnd ({Fresh[5969], Fresh[5968], Fresh[5967], Fresh[5966], Fresh[5965], Fresh[5964], Fresh[5963], Fresh[5962], Fresh[5961], Fresh[5960]}), .outt ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, new_AGEMA_signal_2931, n2095}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2274 ( .ina ({new_AGEMA_signal_2936, new_AGEMA_signal_2935, new_AGEMA_signal_2934, n2116}), .inb ({new_AGEMA_signal_14018, new_AGEMA_signal_14016, new_AGEMA_signal_14014, new_AGEMA_signal_14012}), .clk ( clk ), .rnd ({Fresh[5979], Fresh[5978], Fresh[5977], Fresh[5976], Fresh[5975], Fresh[5974], Fresh[5973], Fresh[5972], Fresh[5971], Fresh[5970]}), .outt ({new_AGEMA_signal_3161, new_AGEMA_signal_3160, new_AGEMA_signal_3159, n2117}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2283 ( .ina ({new_AGEMA_signal_14034, new_AGEMA_signal_14030, new_AGEMA_signal_14026, new_AGEMA_signal_14022}), .inb ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, new_AGEMA_signal_2631, n2120}), .clk ( clk ), .rnd ({Fresh[5989], Fresh[5988], Fresh[5987], Fresh[5986], Fresh[5985], Fresh[5984], Fresh[5983], Fresh[5982], Fresh[5981], Fresh[5980]}), .outt ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, new_AGEMA_signal_2937, n2123}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2300 ( .ina ({new_AGEMA_signal_14042, new_AGEMA_signal_14040, new_AGEMA_signal_14038, new_AGEMA_signal_14036}), .inb ({new_AGEMA_signal_2198, new_AGEMA_signal_2197, new_AGEMA_signal_2196, n2134}), .clk ( clk ), .rnd ({Fresh[5999], Fresh[5998], Fresh[5997], Fresh[5996], Fresh[5995], Fresh[5994], Fresh[5993], Fresh[5992], Fresh[5991], Fresh[5990]}), .outt ({new_AGEMA_signal_2639, new_AGEMA_signal_2638, new_AGEMA_signal_2637, n2135}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2309 ( .ina ({new_AGEMA_signal_14058, new_AGEMA_signal_14054, new_AGEMA_signal_14050, new_AGEMA_signal_14046}), .inb ({new_AGEMA_signal_2645, new_AGEMA_signal_2644, new_AGEMA_signal_2643, n2140}), .clk ( clk ), .rnd ({Fresh[6009], Fresh[6008], Fresh[6007], Fresh[6006], Fresh[6005], Fresh[6004], Fresh[6003], Fresh[6002], Fresh[6001], Fresh[6000]}), .outt ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, new_AGEMA_signal_2943, n2141}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2327 ( .ina ({new_AGEMA_signal_14082, new_AGEMA_signal_14076, new_AGEMA_signal_14070, new_AGEMA_signal_14064}), .inb ({new_AGEMA_signal_2651, new_AGEMA_signal_2650, new_AGEMA_signal_2649, n2161}), .clk ( clk ), .rnd ({Fresh[6019], Fresh[6018], Fresh[6017], Fresh[6016], Fresh[6015], Fresh[6014], Fresh[6013], Fresh[6012], Fresh[6011], Fresh[6010]}), .outt ({new_AGEMA_signal_2948, new_AGEMA_signal_2947, new_AGEMA_signal_2946, n2166}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2331 ( .ina ({new_AGEMA_signal_14098, new_AGEMA_signal_14094, new_AGEMA_signal_14090, new_AGEMA_signal_14086}), .inb ({new_AGEMA_signal_2219, new_AGEMA_signal_2218, new_AGEMA_signal_2217, n2164}), .clk ( clk ), .rnd ({Fresh[6029], Fresh[6028], Fresh[6027], Fresh[6026], Fresh[6025], Fresh[6024], Fresh[6023], Fresh[6022], Fresh[6021], Fresh[6020]}), .outt ({new_AGEMA_signal_2654, new_AGEMA_signal_2653, new_AGEMA_signal_2652, n2165}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2346 ( .ina ({new_AGEMA_signal_2657, new_AGEMA_signal_2656, new_AGEMA_signal_2655, n2179}), .inb ({new_AGEMA_signal_14114, new_AGEMA_signal_14110, new_AGEMA_signal_14106, new_AGEMA_signal_14102}), .clk ( clk ), .rnd ({Fresh[6039], Fresh[6038], Fresh[6037], Fresh[6036], Fresh[6035], Fresh[6034], Fresh[6033], Fresh[6032], Fresh[6031], Fresh[6030]}), .outt ({new_AGEMA_signal_2951, new_AGEMA_signal_2950, new_AGEMA_signal_2949, n2180}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2360 ( .ina ({new_AGEMA_signal_14122, new_AGEMA_signal_14120, new_AGEMA_signal_14118, new_AGEMA_signal_14116}), .inb ({new_AGEMA_signal_2660, new_AGEMA_signal_2659, new_AGEMA_signal_2658, n2192}), .clk ( clk ), .rnd ({Fresh[6049], Fresh[6048], Fresh[6047], Fresh[6046], Fresh[6045], Fresh[6044], Fresh[6043], Fresh[6042], Fresh[6041], Fresh[6040]}), .outt ({new_AGEMA_signal_2954, new_AGEMA_signal_2953, new_AGEMA_signal_2952, n2194}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2372 ( .ina ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, new_AGEMA_signal_2955, n2203}), .inb ({new_AGEMA_signal_14130, new_AGEMA_signal_14128, new_AGEMA_signal_14126, new_AGEMA_signal_14124}), .clk ( clk ), .rnd ({Fresh[6059], Fresh[6058], Fresh[6057], Fresh[6056], Fresh[6055], Fresh[6054], Fresh[6053], Fresh[6052], Fresh[6051], Fresh[6050]}), .outt ({new_AGEMA_signal_3182, new_AGEMA_signal_3181, new_AGEMA_signal_3180, n2204}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2389 ( .ina ({new_AGEMA_signal_2669, new_AGEMA_signal_2668, new_AGEMA_signal_2667, n2224}), .inb ({new_AGEMA_signal_2672, new_AGEMA_signal_2671, new_AGEMA_signal_2670, n2223}), .clk ( clk ), .rnd ({Fresh[6069], Fresh[6068], Fresh[6067], Fresh[6066], Fresh[6065], Fresh[6064], Fresh[6063], Fresh[6062], Fresh[6061], Fresh[6060]}), .outt ({new_AGEMA_signal_2960, new_AGEMA_signal_2959, new_AGEMA_signal_2958, n2225}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2394 ( .ina ({new_AGEMA_signal_2255, new_AGEMA_signal_2254, new_AGEMA_signal_2253, n2229}), .inb ({new_AGEMA_signal_14138, new_AGEMA_signal_14136, new_AGEMA_signal_14134, new_AGEMA_signal_14132}), .clk ( clk ), .rnd ({Fresh[6079], Fresh[6078], Fresh[6077], Fresh[6076], Fresh[6075], Fresh[6074], Fresh[6073], Fresh[6072], Fresh[6071], Fresh[6070]}), .outt ({new_AGEMA_signal_2675, new_AGEMA_signal_2674, new_AGEMA_signal_2673, n2230}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2400 ( .ina ({new_AGEMA_signal_14146, new_AGEMA_signal_14144, new_AGEMA_signal_14142, new_AGEMA_signal_14140}), .inb ({new_AGEMA_signal_2966, new_AGEMA_signal_2965, new_AGEMA_signal_2964, n2234}), .clk ( clk ), .rnd ({Fresh[6089], Fresh[6088], Fresh[6087], Fresh[6086], Fresh[6085], Fresh[6084], Fresh[6083], Fresh[6082], Fresh[6081], Fresh[6080]}), .outt ({new_AGEMA_signal_3188, new_AGEMA_signal_3187, new_AGEMA_signal_3186, n2236}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2412 ( .ina ({new_AGEMA_signal_2681, new_AGEMA_signal_2680, new_AGEMA_signal_2679, n2246}), .inb ({new_AGEMA_signal_14162, new_AGEMA_signal_14158, new_AGEMA_signal_14154, new_AGEMA_signal_14150}), .clk ( clk ), .rnd ({Fresh[6099], Fresh[6098], Fresh[6097], Fresh[6096], Fresh[6095], Fresh[6094], Fresh[6093], Fresh[6092], Fresh[6091], Fresh[6090]}), .outt ({new_AGEMA_signal_2969, new_AGEMA_signal_2968, new_AGEMA_signal_2967, n2247}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2419 ( .ina ({new_AGEMA_signal_2684, new_AGEMA_signal_2683, new_AGEMA_signal_2682, n2254}), .inb ({new_AGEMA_signal_14186, new_AGEMA_signal_14180, new_AGEMA_signal_14174, new_AGEMA_signal_14168}), .clk ( clk ), .rnd ({Fresh[6109], Fresh[6108], Fresh[6107], Fresh[6106], Fresh[6105], Fresh[6104], Fresh[6103], Fresh[6102], Fresh[6101], Fresh[6100]}), .outt ({new_AGEMA_signal_2972, new_AGEMA_signal_2971, new_AGEMA_signal_2970, n2255}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2427 ( .ina ({new_AGEMA_signal_2687, new_AGEMA_signal_2686, new_AGEMA_signal_2685, n2263}), .inb ({new_AGEMA_signal_14202, new_AGEMA_signal_14198, new_AGEMA_signal_14194, new_AGEMA_signal_14190}), .clk ( clk ), .rnd ({Fresh[6119], Fresh[6118], Fresh[6117], Fresh[6116], Fresh[6115], Fresh[6114], Fresh[6113], Fresh[6112], Fresh[6111], Fresh[6110]}), .outt ({new_AGEMA_signal_2975, new_AGEMA_signal_2974, new_AGEMA_signal_2973, n2264}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2435 ( .ina ({new_AGEMA_signal_14210, new_AGEMA_signal_14208, new_AGEMA_signal_14206, new_AGEMA_signal_14204}), .inb ({new_AGEMA_signal_2273, new_AGEMA_signal_2272, new_AGEMA_signal_2271, n2267}), .clk ( clk ), .rnd ({Fresh[6129], Fresh[6128], Fresh[6127], Fresh[6126], Fresh[6125], Fresh[6124], Fresh[6123], Fresh[6122], Fresh[6121], Fresh[6120]}), .outt ({new_AGEMA_signal_2978, new_AGEMA_signal_2977, new_AGEMA_signal_2976, n2271}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2446 ( .ina ({new_AGEMA_signal_13874, new_AGEMA_signal_13870, new_AGEMA_signal_13866, new_AGEMA_signal_13862}), .inb ({new_AGEMA_signal_2279, new_AGEMA_signal_2278, new_AGEMA_signal_2277, n2279}), .clk ( clk ), .rnd ({Fresh[6139], Fresh[6138], Fresh[6137], Fresh[6136], Fresh[6135], Fresh[6134], Fresh[6133], Fresh[6132], Fresh[6131], Fresh[6130]}), .outt ({new_AGEMA_signal_2696, new_AGEMA_signal_2695, new_AGEMA_signal_2694, n2280}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2451 ( .ina ({new_AGEMA_signal_14218, new_AGEMA_signal_14216, new_AGEMA_signal_14214, new_AGEMA_signal_14212}), .inb ({new_AGEMA_signal_2282, new_AGEMA_signal_2281, new_AGEMA_signal_2280, n2283}), .clk ( clk ), .rnd ({Fresh[6149], Fresh[6148], Fresh[6147], Fresh[6146], Fresh[6145], Fresh[6144], Fresh[6143], Fresh[6142], Fresh[6141], Fresh[6140]}), .outt ({new_AGEMA_signal_2699, new_AGEMA_signal_2698, new_AGEMA_signal_2697, n2286}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2461 ( .ina ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, new_AGEMA_signal_2703, n2686}), .inb ({new_AGEMA_signal_2708, new_AGEMA_signal_2707, new_AGEMA_signal_2706, n2289}), .clk ( clk ), .rnd ({Fresh[6159], Fresh[6158], Fresh[6157], Fresh[6156], Fresh[6155], Fresh[6154], Fresh[6153], Fresh[6152], Fresh[6151], Fresh[6150]}), .outt ({new_AGEMA_signal_2984, new_AGEMA_signal_2983, new_AGEMA_signal_2982, n2304}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2466 ( .ina ({new_AGEMA_signal_14226, new_AGEMA_signal_14224, new_AGEMA_signal_14222, new_AGEMA_signal_14220}), .inb ({new_AGEMA_signal_2714, new_AGEMA_signal_2713, new_AGEMA_signal_2712, n2292}), .clk ( clk ), .rnd ({Fresh[6169], Fresh[6168], Fresh[6167], Fresh[6166], Fresh[6165], Fresh[6164], Fresh[6163], Fresh[6162], Fresh[6161], Fresh[6160]}), .outt ({new_AGEMA_signal_2987, new_AGEMA_signal_2986, new_AGEMA_signal_2985, n2295}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2488 ( .ina ({new_AGEMA_signal_2720, new_AGEMA_signal_2719, new_AGEMA_signal_2718, n2321}), .inb ({new_AGEMA_signal_1817, new_AGEMA_signal_1816, new_AGEMA_signal_1815, n2320}), .clk ( clk ), .rnd ({Fresh[6179], Fresh[6178], Fresh[6177], Fresh[6176], Fresh[6175], Fresh[6174], Fresh[6173], Fresh[6172], Fresh[6171], Fresh[6170]}), .outt ({new_AGEMA_signal_2990, new_AGEMA_signal_2989, new_AGEMA_signal_2988, n2322}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2499 ( .ina ({new_AGEMA_signal_2723, new_AGEMA_signal_2722, new_AGEMA_signal_2721, n2332}), .inb ({new_AGEMA_signal_2726, new_AGEMA_signal_2725, new_AGEMA_signal_2724, n2331}), .clk ( clk ), .rnd ({Fresh[6189], Fresh[6188], Fresh[6187], Fresh[6186], Fresh[6185], Fresh[6184], Fresh[6183], Fresh[6182], Fresh[6181], Fresh[6180]}), .outt ({new_AGEMA_signal_2993, new_AGEMA_signal_2992, new_AGEMA_signal_2991, n2333}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2509 ( .ina ({new_AGEMA_signal_14242, new_AGEMA_signal_14238, new_AGEMA_signal_14234, new_AGEMA_signal_14230}), .inb ({new_AGEMA_signal_2732, new_AGEMA_signal_2731, new_AGEMA_signal_2730, n2342}), .clk ( clk ), .rnd ({Fresh[6199], Fresh[6198], Fresh[6197], Fresh[6196], Fresh[6195], Fresh[6194], Fresh[6193], Fresh[6192], Fresh[6191], Fresh[6190]}), .outt ({new_AGEMA_signal_2999, new_AGEMA_signal_2998, new_AGEMA_signal_2997, n2345}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2526 ( .ina ({new_AGEMA_signal_2735, new_AGEMA_signal_2734, new_AGEMA_signal_2733, n2358}), .inb ({new_AGEMA_signal_14250, new_AGEMA_signal_14248, new_AGEMA_signal_14246, new_AGEMA_signal_14244}), .clk ( clk ), .rnd ({Fresh[6209], Fresh[6208], Fresh[6207], Fresh[6206], Fresh[6205], Fresh[6204], Fresh[6203], Fresh[6202], Fresh[6201], Fresh[6200]}), .outt ({new_AGEMA_signal_3002, new_AGEMA_signal_3001, new_AGEMA_signal_3000, n2361}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2549 ( .ina ({new_AGEMA_signal_2336, new_AGEMA_signal_2335, new_AGEMA_signal_2334, n2387}), .inb ({new_AGEMA_signal_14258, new_AGEMA_signal_14256, new_AGEMA_signal_14254, new_AGEMA_signal_14252}), .clk ( clk ), .rnd ({Fresh[6219], Fresh[6218], Fresh[6217], Fresh[6216], Fresh[6215], Fresh[6214], Fresh[6213], Fresh[6212], Fresh[6211], Fresh[6210]}), .outt ({new_AGEMA_signal_2741, new_AGEMA_signal_2740, new_AGEMA_signal_2739, n2388}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2556 ( .ina ({new_AGEMA_signal_14274, new_AGEMA_signal_14270, new_AGEMA_signal_14266, new_AGEMA_signal_14262}), .inb ({new_AGEMA_signal_2744, new_AGEMA_signal_2743, new_AGEMA_signal_2742, n2392}), .clk ( clk ), .rnd ({Fresh[6229], Fresh[6228], Fresh[6227], Fresh[6226], Fresh[6225], Fresh[6224], Fresh[6223], Fresh[6222], Fresh[6221], Fresh[6220]}), .outt ({new_AGEMA_signal_3008, new_AGEMA_signal_3007, new_AGEMA_signal_3006, n2393}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2567 ( .ina ({new_AGEMA_signal_14290, new_AGEMA_signal_14286, new_AGEMA_signal_14282, new_AGEMA_signal_14278}), .inb ({new_AGEMA_signal_2348, new_AGEMA_signal_2347, new_AGEMA_signal_2346, n2404}), .clk ( clk ), .rnd ({Fresh[6239], Fresh[6238], Fresh[6237], Fresh[6236], Fresh[6235], Fresh[6234], Fresh[6233], Fresh[6232], Fresh[6231], Fresh[6230]}), .outt ({new_AGEMA_signal_2747, new_AGEMA_signal_2746, new_AGEMA_signal_2745, n2405}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2571 ( .ina ({new_AGEMA_signal_2750, new_AGEMA_signal_2749, new_AGEMA_signal_2748, n2409}), .inb ({new_AGEMA_signal_14306, new_AGEMA_signal_14302, new_AGEMA_signal_14298, new_AGEMA_signal_14294}), .clk ( clk ), .rnd ({Fresh[6249], Fresh[6248], Fresh[6247], Fresh[6246], Fresh[6245], Fresh[6244], Fresh[6243], Fresh[6242], Fresh[6241], Fresh[6240]}), .outt ({new_AGEMA_signal_3014, new_AGEMA_signal_3013, new_AGEMA_signal_3012, n2410}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2576 ( .ina ({new_AGEMA_signal_14322, new_AGEMA_signal_14318, new_AGEMA_signal_14314, new_AGEMA_signal_14310}), .inb ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, new_AGEMA_signal_2751, n2414}), .clk ( clk ), .rnd ({Fresh[6259], Fresh[6258], Fresh[6257], Fresh[6256], Fresh[6255], Fresh[6254], Fresh[6253], Fresh[6252], Fresh[6251], Fresh[6250]}), .outt ({new_AGEMA_signal_3017, new_AGEMA_signal_3016, new_AGEMA_signal_3015, n2421}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2579 ( .ina ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, new_AGEMA_signal_2355, n2418}), .inb ({new_AGEMA_signal_14338, new_AGEMA_signal_14334, new_AGEMA_signal_14330, new_AGEMA_signal_14326}), .clk ( clk ), .rnd ({Fresh[6269], Fresh[6268], Fresh[6267], Fresh[6266], Fresh[6265], Fresh[6264], Fresh[6263], Fresh[6262], Fresh[6261], Fresh[6260]}), .outt ({new_AGEMA_signal_2756, new_AGEMA_signal_2755, new_AGEMA_signal_2754, n2419}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2590 ( .ina ({new_AGEMA_signal_14346, new_AGEMA_signal_14344, new_AGEMA_signal_14342, new_AGEMA_signal_14340}), .inb ({new_AGEMA_signal_2759, new_AGEMA_signal_2758, new_AGEMA_signal_2757, n2432}), .clk ( clk ), .rnd ({Fresh[6279], Fresh[6278], Fresh[6277], Fresh[6276], Fresh[6275], Fresh[6274], Fresh[6273], Fresh[6272], Fresh[6271], Fresh[6270]}), .outt ({new_AGEMA_signal_3023, new_AGEMA_signal_3022, new_AGEMA_signal_3021, n2436}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2604 ( .ina ({new_AGEMA_signal_2762, new_AGEMA_signal_2761, new_AGEMA_signal_2760, n2449}), .inb ({new_AGEMA_signal_2765, new_AGEMA_signal_2764, new_AGEMA_signal_2763, n2448}), .clk ( clk ), .rnd ({Fresh[6289], Fresh[6288], Fresh[6287], Fresh[6286], Fresh[6285], Fresh[6284], Fresh[6283], Fresh[6282], Fresh[6281], Fresh[6280]}), .outt ({new_AGEMA_signal_3026, new_AGEMA_signal_3025, new_AGEMA_signal_3024, n2450}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2610 ( .ina ({new_AGEMA_signal_14354, new_AGEMA_signal_14352, new_AGEMA_signal_14350, new_AGEMA_signal_14348}), .inb ({new_AGEMA_signal_2768, new_AGEMA_signal_2767, new_AGEMA_signal_2766, n2455}), .clk ( clk ), .rnd ({Fresh[6299], Fresh[6298], Fresh[6297], Fresh[6296], Fresh[6295], Fresh[6294], Fresh[6293], Fresh[6292], Fresh[6291], Fresh[6290]}), .outt ({new_AGEMA_signal_3029, new_AGEMA_signal_3028, new_AGEMA_signal_3027, n2456}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2613 ( .ina ({new_AGEMA_signal_2771, new_AGEMA_signal_2770, new_AGEMA_signal_2769, n2460}), .inb ({new_AGEMA_signal_14362, new_AGEMA_signal_14360, new_AGEMA_signal_14358, new_AGEMA_signal_14356}), .clk ( clk ), .rnd ({Fresh[6309], Fresh[6308], Fresh[6307], Fresh[6306], Fresh[6305], Fresh[6304], Fresh[6303], Fresh[6302], Fresh[6301], Fresh[6300]}), .outt ({new_AGEMA_signal_3032, new_AGEMA_signal_3031, new_AGEMA_signal_3030, n2461}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2619 ( .ina ({new_AGEMA_signal_14370, new_AGEMA_signal_14368, new_AGEMA_signal_14366, new_AGEMA_signal_14364}), .inb ({new_AGEMA_signal_2384, new_AGEMA_signal_2383, new_AGEMA_signal_2382, n2466}), .clk ( clk ), .rnd ({Fresh[6319], Fresh[6318], Fresh[6317], Fresh[6316], Fresh[6315], Fresh[6314], Fresh[6313], Fresh[6312], Fresh[6311], Fresh[6310]}), .outt ({new_AGEMA_signal_2774, new_AGEMA_signal_2773, new_AGEMA_signal_2772, n2469}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2630 ( .ina ({new_AGEMA_signal_14386, new_AGEMA_signal_14382, new_AGEMA_signal_14378, new_AGEMA_signal_14374}), .inb ({new_AGEMA_signal_2387, new_AGEMA_signal_2386, new_AGEMA_signal_2385, n2477}), .clk ( clk ), .rnd ({Fresh[6329], Fresh[6328], Fresh[6327], Fresh[6326], Fresh[6325], Fresh[6324], Fresh[6323], Fresh[6322], Fresh[6321], Fresh[6320]}), .outt ({new_AGEMA_signal_2777, new_AGEMA_signal_2776, new_AGEMA_signal_2775, n2478}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2635 ( .ina ({new_AGEMA_signal_14402, new_AGEMA_signal_14398, new_AGEMA_signal_14394, new_AGEMA_signal_14390}), .inb ({new_AGEMA_signal_2780, new_AGEMA_signal_2779, new_AGEMA_signal_2778, n2482}), .clk ( clk ), .rnd ({Fresh[6339], Fresh[6338], Fresh[6337], Fresh[6336], Fresh[6335], Fresh[6334], Fresh[6333], Fresh[6332], Fresh[6331], Fresh[6330]}), .outt ({new_AGEMA_signal_3038, new_AGEMA_signal_3037, new_AGEMA_signal_3036, n2484}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2643 ( .ina ({new_AGEMA_signal_2393, new_AGEMA_signal_2392, new_AGEMA_signal_2391, n2490}), .inb ({new_AGEMA_signal_14410, new_AGEMA_signal_14408, new_AGEMA_signal_14406, new_AGEMA_signal_14404}), .clk ( clk ), .rnd ({Fresh[6349], Fresh[6348], Fresh[6347], Fresh[6346], Fresh[6345], Fresh[6344], Fresh[6343], Fresh[6342], Fresh[6341], Fresh[6340]}), .outt ({new_AGEMA_signal_2783, new_AGEMA_signal_2782, new_AGEMA_signal_2781, n2491}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2649 ( .ina ({new_AGEMA_signal_14418, new_AGEMA_signal_14416, new_AGEMA_signal_14414, new_AGEMA_signal_14412}), .inb ({new_AGEMA_signal_2786, new_AGEMA_signal_2785, new_AGEMA_signal_2784, n2496}), .clk ( clk ), .rnd ({Fresh[6359], Fresh[6358], Fresh[6357], Fresh[6356], Fresh[6355], Fresh[6354], Fresh[6353], Fresh[6352], Fresh[6351], Fresh[6350]}), .outt ({new_AGEMA_signal_3044, new_AGEMA_signal_3043, new_AGEMA_signal_3042, n2500}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2656 ( .ina ({new_AGEMA_signal_3047, new_AGEMA_signal_3046, new_AGEMA_signal_3045, n2507}), .inb ({new_AGEMA_signal_14426, new_AGEMA_signal_14424, new_AGEMA_signal_14422, new_AGEMA_signal_14420}), .clk ( clk ), .rnd ({Fresh[6369], Fresh[6368], Fresh[6367], Fresh[6366], Fresh[6365], Fresh[6364], Fresh[6363], Fresh[6362], Fresh[6361], Fresh[6360]}), .outt ({new_AGEMA_signal_3242, new_AGEMA_signal_3241, new_AGEMA_signal_3240, n2508}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2670 ( .ina ({new_AGEMA_signal_3050, new_AGEMA_signal_3049, new_AGEMA_signal_3048, n2525}), .inb ({new_AGEMA_signal_2795, new_AGEMA_signal_2794, new_AGEMA_signal_2793, n2524}), .clk ( clk ), .rnd ({Fresh[6379], Fresh[6378], Fresh[6377], Fresh[6376], Fresh[6375], Fresh[6374], Fresh[6373], Fresh[6372], Fresh[6371], Fresh[6370]}), .outt ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, new_AGEMA_signal_3243, n2526}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2679 ( .ina ({new_AGEMA_signal_2798, new_AGEMA_signal_2797, new_AGEMA_signal_2796, n2537}), .inb ({new_AGEMA_signal_2801, new_AGEMA_signal_2800, new_AGEMA_signal_2799, n2536}), .clk ( clk ), .rnd ({Fresh[6389], Fresh[6388], Fresh[6387], Fresh[6386], Fresh[6385], Fresh[6384], Fresh[6383], Fresh[6382], Fresh[6381], Fresh[6380]}), .outt ({new_AGEMA_signal_3053, new_AGEMA_signal_3052, new_AGEMA_signal_3051, n2539}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2682 ( .ina ({new_AGEMA_signal_2636, new_AGEMA_signal_2635, new_AGEMA_signal_2634, n2543}), .inb ({new_AGEMA_signal_14434, new_AGEMA_signal_14432, new_AGEMA_signal_14430, new_AGEMA_signal_14428}), .clk ( clk ), .rnd ({Fresh[6399], Fresh[6398], Fresh[6397], Fresh[6396], Fresh[6395], Fresh[6394], Fresh[6393], Fresh[6392], Fresh[6391], Fresh[6390]}), .outt ({new_AGEMA_signal_3056, new_AGEMA_signal_3055, new_AGEMA_signal_3054, n2548}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2694 ( .ina ({new_AGEMA_signal_14442, new_AGEMA_signal_14440, new_AGEMA_signal_14438, new_AGEMA_signal_14436}), .inb ({new_AGEMA_signal_2804, new_AGEMA_signal_2803, new_AGEMA_signal_2802, n2557}), .clk ( clk ), .rnd ({Fresh[6409], Fresh[6408], Fresh[6407], Fresh[6406], Fresh[6405], Fresh[6404], Fresh[6403], Fresh[6402], Fresh[6401], Fresh[6400]}), .outt ({new_AGEMA_signal_3059, new_AGEMA_signal_3058, new_AGEMA_signal_3057, n2568}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2700 ( .ina ({new_AGEMA_signal_14450, new_AGEMA_signal_14448, new_AGEMA_signal_14446, new_AGEMA_signal_14444}), .inb ({new_AGEMA_signal_2807, new_AGEMA_signal_2806, new_AGEMA_signal_2805, n2565}), .clk ( clk ), .rnd ({Fresh[6419], Fresh[6418], Fresh[6417], Fresh[6416], Fresh[6415], Fresh[6414], Fresh[6413], Fresh[6412], Fresh[6411], Fresh[6410]}), .outt ({new_AGEMA_signal_3062, new_AGEMA_signal_3061, new_AGEMA_signal_3060, n2567}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2710 ( .ina ({new_AGEMA_signal_14458, new_AGEMA_signal_14456, new_AGEMA_signal_14454, new_AGEMA_signal_14452}), .inb ({new_AGEMA_signal_2813, new_AGEMA_signal_2812, new_AGEMA_signal_2811, n2580}), .clk ( clk ), .rnd ({Fresh[6429], Fresh[6428], Fresh[6427], Fresh[6426], Fresh[6425], Fresh[6424], Fresh[6423], Fresh[6422], Fresh[6421], Fresh[6420]}), .outt ({new_AGEMA_signal_3065, new_AGEMA_signal_3064, new_AGEMA_signal_3063, n2583}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2728 ( .ina ({new_AGEMA_signal_14466, new_AGEMA_signal_14464, new_AGEMA_signal_14462, new_AGEMA_signal_14460}), .inb ({new_AGEMA_signal_1964, new_AGEMA_signal_1963, new_AGEMA_signal_1962, n2602}), .clk ( clk ), .rnd ({Fresh[6439], Fresh[6438], Fresh[6437], Fresh[6436], Fresh[6435], Fresh[6434], Fresh[6433], Fresh[6432], Fresh[6431], Fresh[6430]}), .outt ({new_AGEMA_signal_2816, new_AGEMA_signal_2815, new_AGEMA_signal_2814, n2604}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2739 ( .ina ({new_AGEMA_signal_14474, new_AGEMA_signal_14472, new_AGEMA_signal_14470, new_AGEMA_signal_14468}), .inb ({new_AGEMA_signal_2819, new_AGEMA_signal_2818, new_AGEMA_signal_2817, n2619}), .clk ( clk ), .rnd ({Fresh[6449], Fresh[6448], Fresh[6447], Fresh[6446], Fresh[6445], Fresh[6444], Fresh[6443], Fresh[6442], Fresh[6441], Fresh[6440]}), .outt ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, new_AGEMA_signal_3069, n2621}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2745 ( .ina ({new_AGEMA_signal_14490, new_AGEMA_signal_14486, new_AGEMA_signal_14482, new_AGEMA_signal_14478}), .inb ({new_AGEMA_signal_2822, new_AGEMA_signal_2821, new_AGEMA_signal_2820, n2628}), .clk ( clk ), .rnd ({Fresh[6459], Fresh[6458], Fresh[6457], Fresh[6456], Fresh[6455], Fresh[6454], Fresh[6453], Fresh[6452], Fresh[6451], Fresh[6450]}), .outt ({new_AGEMA_signal_3074, new_AGEMA_signal_3073, new_AGEMA_signal_3072, n2633}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2756 ( .ina ({new_AGEMA_signal_2825, new_AGEMA_signal_2824, new_AGEMA_signal_2823, n2649}), .inb ({new_AGEMA_signal_2471, new_AGEMA_signal_2470, new_AGEMA_signal_2469, n2648}), .clk ( clk ), .rnd ({Fresh[6469], Fresh[6468], Fresh[6467], Fresh[6466], Fresh[6465], Fresh[6464], Fresh[6463], Fresh[6462], Fresh[6461], Fresh[6460]}), .outt ({new_AGEMA_signal_3077, new_AGEMA_signal_3076, new_AGEMA_signal_3075, n2660}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2759 ( .ina ({new_AGEMA_signal_14498, new_AGEMA_signal_14496, new_AGEMA_signal_14494, new_AGEMA_signal_14492}), .inb ({new_AGEMA_signal_2606, new_AGEMA_signal_2605, new_AGEMA_signal_2604, n2652}), .clk ( clk ), .rnd ({Fresh[6479], Fresh[6478], Fresh[6477], Fresh[6476], Fresh[6475], Fresh[6474], Fresh[6473], Fresh[6472], Fresh[6471], Fresh[6470]}), .outt ({new_AGEMA_signal_3080, new_AGEMA_signal_3079, new_AGEMA_signal_3078, n2656}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2766 ( .ina ({new_AGEMA_signal_14506, new_AGEMA_signal_14504, new_AGEMA_signal_14502, new_AGEMA_signal_14500}), .inb ({new_AGEMA_signal_2828, new_AGEMA_signal_2827, new_AGEMA_signal_2826, n2664}), .clk ( clk ), .rnd ({Fresh[6489], Fresh[6488], Fresh[6487], Fresh[6486], Fresh[6485], Fresh[6484], Fresh[6483], Fresh[6482], Fresh[6481], Fresh[6480]}), .outt ({new_AGEMA_signal_3083, new_AGEMA_signal_3082, new_AGEMA_signal_3081, n2666}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2774 ( .ina ({new_AGEMA_signal_2831, new_AGEMA_signal_2830, new_AGEMA_signal_2829, n2681}), .inb ({new_AGEMA_signal_2480, new_AGEMA_signal_2479, new_AGEMA_signal_2478, n2680}), .clk ( clk ), .rnd ({Fresh[6499], Fresh[6498], Fresh[6497], Fresh[6496], Fresh[6495], Fresh[6494], Fresh[6493], Fresh[6492], Fresh[6491], Fresh[6490]}), .outt ({new_AGEMA_signal_3086, new_AGEMA_signal_3085, new_AGEMA_signal_3084, n2706}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2777 ( .ina ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, new_AGEMA_signal_2703, n2686}), .inb ({new_AGEMA_signal_2834, new_AGEMA_signal_2833, new_AGEMA_signal_2832, n2685}), .clk ( clk ), .rnd ({Fresh[6509], Fresh[6508], Fresh[6507], Fresh[6506], Fresh[6505], Fresh[6504], Fresh[6503], Fresh[6502], Fresh[6501], Fresh[6500]}), .outt ({new_AGEMA_signal_3089, new_AGEMA_signal_3088, new_AGEMA_signal_3087, n2704}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2781 ( .ina ({new_AGEMA_signal_2840, new_AGEMA_signal_2839, new_AGEMA_signal_2838, n2692}), .inb ({new_AGEMA_signal_14514, new_AGEMA_signal_14512, new_AGEMA_signal_14510, new_AGEMA_signal_14508}), .clk ( clk ), .rnd ({Fresh[6519], Fresh[6518], Fresh[6517], Fresh[6516], Fresh[6515], Fresh[6514], Fresh[6513], Fresh[6512], Fresh[6511], Fresh[6510]}), .outt ({new_AGEMA_signal_3092, new_AGEMA_signal_3091, new_AGEMA_signal_3090, n2696}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2794 ( .ina ({new_AGEMA_signal_14522, new_AGEMA_signal_14520, new_AGEMA_signal_14518, new_AGEMA_signal_14516}), .inb ({new_AGEMA_signal_2843, new_AGEMA_signal_2842, new_AGEMA_signal_2841, n2716}), .clk ( clk ), .rnd ({Fresh[6529], Fresh[6528], Fresh[6527], Fresh[6526], Fresh[6525], Fresh[6524], Fresh[6523], Fresh[6522], Fresh[6521], Fresh[6520]}), .outt ({new_AGEMA_signal_3095, new_AGEMA_signal_3094, new_AGEMA_signal_3093, n2718}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2801 ( .ina ({new_AGEMA_signal_14530, new_AGEMA_signal_14528, new_AGEMA_signal_14526, new_AGEMA_signal_14524}), .inb ({new_AGEMA_signal_2489, new_AGEMA_signal_2488, new_AGEMA_signal_2487, n2728}), .clk ( clk ), .rnd ({Fresh[6539], Fresh[6538], Fresh[6537], Fresh[6536], Fresh[6535], Fresh[6534], Fresh[6533], Fresh[6532], Fresh[6531], Fresh[6530]}), .outt ({new_AGEMA_signal_3098, new_AGEMA_signal_3097, new_AGEMA_signal_3096, n2730}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2805 ( .ina ({new_AGEMA_signal_14546, new_AGEMA_signal_14542, new_AGEMA_signal_14538, new_AGEMA_signal_14534}), .inb ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, new_AGEMA_signal_2847, n2735}), .clk ( clk ), .rnd ({Fresh[6549], Fresh[6548], Fresh[6547], Fresh[6546], Fresh[6545], Fresh[6544], Fresh[6543], Fresh[6542], Fresh[6541], Fresh[6540]}), .outt ({new_AGEMA_signal_3101, new_AGEMA_signal_3100, new_AGEMA_signal_3099, n2745}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2809 ( .ina ({new_AGEMA_signal_2852, new_AGEMA_signal_2851, new_AGEMA_signal_2850, n2743}), .inb ({new_AGEMA_signal_14562, new_AGEMA_signal_14558, new_AGEMA_signal_14554, new_AGEMA_signal_14550}), .clk ( clk ), .rnd ({Fresh[6559], Fresh[6558], Fresh[6557], Fresh[6556], Fresh[6555], Fresh[6554], Fresh[6553], Fresh[6552], Fresh[6551], Fresh[6550]}), .outt ({new_AGEMA_signal_3104, new_AGEMA_signal_3103, new_AGEMA_signal_3102, n2744}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2814 ( .ina ({new_AGEMA_signal_14210, new_AGEMA_signal_14208, new_AGEMA_signal_14206, new_AGEMA_signal_14204}), .inb ({new_AGEMA_signal_2498, new_AGEMA_signal_2497, new_AGEMA_signal_2496, n2751}), .clk ( clk ), .rnd ({Fresh[6569], Fresh[6568], Fresh[6567], Fresh[6566], Fresh[6565], Fresh[6564], Fresh[6563], Fresh[6562], Fresh[6561], Fresh[6560]}), .outt ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, new_AGEMA_signal_3105, n2759}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2821 ( .ina ({new_AGEMA_signal_14578, new_AGEMA_signal_14574, new_AGEMA_signal_14570, new_AGEMA_signal_14566}), .inb ({new_AGEMA_signal_2858, new_AGEMA_signal_2857, new_AGEMA_signal_2856, n2764}), .clk ( clk ), .rnd ({Fresh[6579], Fresh[6578], Fresh[6577], Fresh[6576], Fresh[6575], Fresh[6574], Fresh[6573], Fresh[6572], Fresh[6571], Fresh[6570]}), .outt ({new_AGEMA_signal_3110, new_AGEMA_signal_3109, new_AGEMA_signal_3108, n2771}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2833 ( .ina ({new_AGEMA_signal_2516, new_AGEMA_signal_2515, new_AGEMA_signal_2514, n2788}), .inb ({new_AGEMA_signal_14594, new_AGEMA_signal_14590, new_AGEMA_signal_14586, new_AGEMA_signal_14582}), .clk ( clk ), .rnd ({Fresh[6589], Fresh[6588], Fresh[6587], Fresh[6586], Fresh[6585], Fresh[6584], Fresh[6583], Fresh[6582], Fresh[6581], Fresh[6580]}), .outt ({new_AGEMA_signal_2864, new_AGEMA_signal_2863, new_AGEMA_signal_2862, n2798}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2850 ( .ina ({new_AGEMA_signal_2870, new_AGEMA_signal_2869, new_AGEMA_signal_2868, n2822}), .inb ({new_AGEMA_signal_2525, new_AGEMA_signal_2524, new_AGEMA_signal_2523, n2821}), .clk ( clk ), .rnd ({Fresh[6599], Fresh[6598], Fresh[6597], Fresh[6596], Fresh[6595], Fresh[6594], Fresh[6593], Fresh[6592], Fresh[6591], Fresh[6590]}), .outt ({new_AGEMA_signal_3116, new_AGEMA_signal_3115, new_AGEMA_signal_3114, n2826}) ) ;
    buf_clk new_AGEMA_reg_buffer_3098 ( .C ( clk ), .D ( new_AGEMA_signal_14597 ), .Q ( new_AGEMA_signal_14598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3102 ( .C ( clk ), .D ( new_AGEMA_signal_14601 ), .Q ( new_AGEMA_signal_14602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3106 ( .C ( clk ), .D ( new_AGEMA_signal_14605 ), .Q ( new_AGEMA_signal_14606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3110 ( .C ( clk ), .D ( new_AGEMA_signal_14609 ), .Q ( new_AGEMA_signal_14610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3114 ( .C ( clk ), .D ( new_AGEMA_signal_14613 ), .Q ( new_AGEMA_signal_14614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3118 ( .C ( clk ), .D ( new_AGEMA_signal_14617 ), .Q ( new_AGEMA_signal_14618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3122 ( .C ( clk ), .D ( new_AGEMA_signal_14621 ), .Q ( new_AGEMA_signal_14622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3126 ( .C ( clk ), .D ( new_AGEMA_signal_14625 ), .Q ( new_AGEMA_signal_14626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3134 ( .C ( clk ), .D ( new_AGEMA_signal_14633 ), .Q ( new_AGEMA_signal_14634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3142 ( .C ( clk ), .D ( new_AGEMA_signal_14641 ), .Q ( new_AGEMA_signal_14642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3150 ( .C ( clk ), .D ( new_AGEMA_signal_14649 ), .Q ( new_AGEMA_signal_14650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3158 ( .C ( clk ), .D ( new_AGEMA_signal_14657 ), .Q ( new_AGEMA_signal_14658 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3160 ( .C ( clk ), .D ( new_AGEMA_signal_14659 ), .Q ( new_AGEMA_signal_14660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3162 ( .C ( clk ), .D ( new_AGEMA_signal_14661 ), .Q ( new_AGEMA_signal_14662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3164 ( .C ( clk ), .D ( new_AGEMA_signal_14663 ), .Q ( new_AGEMA_signal_14664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3166 ( .C ( clk ), .D ( new_AGEMA_signal_14665 ), .Q ( new_AGEMA_signal_14666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3174 ( .C ( clk ), .D ( new_AGEMA_signal_14673 ), .Q ( new_AGEMA_signal_14674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3182 ( .C ( clk ), .D ( new_AGEMA_signal_14681 ), .Q ( new_AGEMA_signal_14682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3190 ( .C ( clk ), .D ( new_AGEMA_signal_14689 ), .Q ( new_AGEMA_signal_14690 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3198 ( .C ( clk ), .D ( new_AGEMA_signal_14697 ), .Q ( new_AGEMA_signal_14698 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3204 ( .C ( clk ), .D ( new_AGEMA_signal_14703 ), .Q ( new_AGEMA_signal_14704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3210 ( .C ( clk ), .D ( new_AGEMA_signal_14709 ), .Q ( new_AGEMA_signal_14710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3216 ( .C ( clk ), .D ( new_AGEMA_signal_14715 ), .Q ( new_AGEMA_signal_14716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3222 ( .C ( clk ), .D ( new_AGEMA_signal_14721 ), .Q ( new_AGEMA_signal_14722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3226 ( .C ( clk ), .D ( new_AGEMA_signal_14725 ), .Q ( new_AGEMA_signal_14726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3230 ( .C ( clk ), .D ( new_AGEMA_signal_14729 ), .Q ( new_AGEMA_signal_14730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3234 ( .C ( clk ), .D ( new_AGEMA_signal_14733 ), .Q ( new_AGEMA_signal_14734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3238 ( .C ( clk ), .D ( new_AGEMA_signal_14737 ), .Q ( new_AGEMA_signal_14738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3244 ( .C ( clk ), .D ( new_AGEMA_signal_14743 ), .Q ( new_AGEMA_signal_14744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3250 ( .C ( clk ), .D ( new_AGEMA_signal_14749 ), .Q ( new_AGEMA_signal_14750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3256 ( .C ( clk ), .D ( new_AGEMA_signal_14755 ), .Q ( new_AGEMA_signal_14756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3262 ( .C ( clk ), .D ( new_AGEMA_signal_14761 ), .Q ( new_AGEMA_signal_14762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3264 ( .C ( clk ), .D ( new_AGEMA_signal_14763 ), .Q ( new_AGEMA_signal_14764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3266 ( .C ( clk ), .D ( new_AGEMA_signal_14765 ), .Q ( new_AGEMA_signal_14766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3268 ( .C ( clk ), .D ( new_AGEMA_signal_14767 ), .Q ( new_AGEMA_signal_14768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3270 ( .C ( clk ), .D ( new_AGEMA_signal_14769 ), .Q ( new_AGEMA_signal_14770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3276 ( .C ( clk ), .D ( new_AGEMA_signal_14775 ), .Q ( new_AGEMA_signal_14776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3282 ( .C ( clk ), .D ( new_AGEMA_signal_14781 ), .Q ( new_AGEMA_signal_14782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3288 ( .C ( clk ), .D ( new_AGEMA_signal_14787 ), .Q ( new_AGEMA_signal_14788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3294 ( .C ( clk ), .D ( new_AGEMA_signal_14793 ), .Q ( new_AGEMA_signal_14794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3300 ( .C ( clk ), .D ( new_AGEMA_signal_14799 ), .Q ( new_AGEMA_signal_14800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3306 ( .C ( clk ), .D ( new_AGEMA_signal_14805 ), .Q ( new_AGEMA_signal_14806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3312 ( .C ( clk ), .D ( new_AGEMA_signal_14811 ), .Q ( new_AGEMA_signal_14812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3318 ( .C ( clk ), .D ( new_AGEMA_signal_14817 ), .Q ( new_AGEMA_signal_14818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3320 ( .C ( clk ), .D ( new_AGEMA_signal_14819 ), .Q ( new_AGEMA_signal_14820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3322 ( .C ( clk ), .D ( new_AGEMA_signal_14821 ), .Q ( new_AGEMA_signal_14822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3324 ( .C ( clk ), .D ( new_AGEMA_signal_14823 ), .Q ( new_AGEMA_signal_14824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3326 ( .C ( clk ), .D ( new_AGEMA_signal_14825 ), .Q ( new_AGEMA_signal_14826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3330 ( .C ( clk ), .D ( new_AGEMA_signal_14829 ), .Q ( new_AGEMA_signal_14830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3334 ( .C ( clk ), .D ( new_AGEMA_signal_14833 ), .Q ( new_AGEMA_signal_14834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3338 ( .C ( clk ), .D ( new_AGEMA_signal_14837 ), .Q ( new_AGEMA_signal_14838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3342 ( .C ( clk ), .D ( new_AGEMA_signal_14841 ), .Q ( new_AGEMA_signal_14842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3348 ( .C ( clk ), .D ( new_AGEMA_signal_14847 ), .Q ( new_AGEMA_signal_14848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3354 ( .C ( clk ), .D ( new_AGEMA_signal_14853 ), .Q ( new_AGEMA_signal_14854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3360 ( .C ( clk ), .D ( new_AGEMA_signal_14859 ), .Q ( new_AGEMA_signal_14860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3366 ( .C ( clk ), .D ( new_AGEMA_signal_14865 ), .Q ( new_AGEMA_signal_14866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3372 ( .C ( clk ), .D ( new_AGEMA_signal_14871 ), .Q ( new_AGEMA_signal_14872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3378 ( .C ( clk ), .D ( new_AGEMA_signal_14877 ), .Q ( new_AGEMA_signal_14878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3384 ( .C ( clk ), .D ( new_AGEMA_signal_14883 ), .Q ( new_AGEMA_signal_14884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3390 ( .C ( clk ), .D ( new_AGEMA_signal_14889 ), .Q ( new_AGEMA_signal_14890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3392 ( .C ( clk ), .D ( new_AGEMA_signal_14891 ), .Q ( new_AGEMA_signal_14892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3394 ( .C ( clk ), .D ( new_AGEMA_signal_14893 ), .Q ( new_AGEMA_signal_14894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3396 ( .C ( clk ), .D ( new_AGEMA_signal_14895 ), .Q ( new_AGEMA_signal_14896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3398 ( .C ( clk ), .D ( new_AGEMA_signal_14897 ), .Q ( new_AGEMA_signal_14898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3404 ( .C ( clk ), .D ( new_AGEMA_signal_14903 ), .Q ( new_AGEMA_signal_14904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3410 ( .C ( clk ), .D ( new_AGEMA_signal_14909 ), .Q ( new_AGEMA_signal_14910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3416 ( .C ( clk ), .D ( new_AGEMA_signal_14915 ), .Q ( new_AGEMA_signal_14916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3422 ( .C ( clk ), .D ( new_AGEMA_signal_14921 ), .Q ( new_AGEMA_signal_14922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3424 ( .C ( clk ), .D ( new_AGEMA_signal_14923 ), .Q ( new_AGEMA_signal_14924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3426 ( .C ( clk ), .D ( new_AGEMA_signal_14925 ), .Q ( new_AGEMA_signal_14926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3428 ( .C ( clk ), .D ( new_AGEMA_signal_14927 ), .Q ( new_AGEMA_signal_14928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3430 ( .C ( clk ), .D ( new_AGEMA_signal_14929 ), .Q ( new_AGEMA_signal_14930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3434 ( .C ( clk ), .D ( new_AGEMA_signal_14933 ), .Q ( new_AGEMA_signal_14934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3438 ( .C ( clk ), .D ( new_AGEMA_signal_14937 ), .Q ( new_AGEMA_signal_14938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3442 ( .C ( clk ), .D ( new_AGEMA_signal_14941 ), .Q ( new_AGEMA_signal_14942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3446 ( .C ( clk ), .D ( new_AGEMA_signal_14945 ), .Q ( new_AGEMA_signal_14946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3450 ( .C ( clk ), .D ( new_AGEMA_signal_14949 ), .Q ( new_AGEMA_signal_14950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3454 ( .C ( clk ), .D ( new_AGEMA_signal_14953 ), .Q ( new_AGEMA_signal_14954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3458 ( .C ( clk ), .D ( new_AGEMA_signal_14957 ), .Q ( new_AGEMA_signal_14958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3462 ( .C ( clk ), .D ( new_AGEMA_signal_14961 ), .Q ( new_AGEMA_signal_14962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3464 ( .C ( clk ), .D ( new_AGEMA_signal_14963 ), .Q ( new_AGEMA_signal_14964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3466 ( .C ( clk ), .D ( new_AGEMA_signal_14965 ), .Q ( new_AGEMA_signal_14966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3468 ( .C ( clk ), .D ( new_AGEMA_signal_14967 ), .Q ( new_AGEMA_signal_14968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3470 ( .C ( clk ), .D ( new_AGEMA_signal_14969 ), .Q ( new_AGEMA_signal_14970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3478 ( .C ( clk ), .D ( new_AGEMA_signal_14977 ), .Q ( new_AGEMA_signal_14978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3486 ( .C ( clk ), .D ( new_AGEMA_signal_14985 ), .Q ( new_AGEMA_signal_14986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3494 ( .C ( clk ), .D ( new_AGEMA_signal_14993 ), .Q ( new_AGEMA_signal_14994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3502 ( .C ( clk ), .D ( new_AGEMA_signal_15001 ), .Q ( new_AGEMA_signal_15002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3508 ( .C ( clk ), .D ( new_AGEMA_signal_15007 ), .Q ( new_AGEMA_signal_15008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3514 ( .C ( clk ), .D ( new_AGEMA_signal_15013 ), .Q ( new_AGEMA_signal_15014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3520 ( .C ( clk ), .D ( new_AGEMA_signal_15019 ), .Q ( new_AGEMA_signal_15020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3526 ( .C ( clk ), .D ( new_AGEMA_signal_15025 ), .Q ( new_AGEMA_signal_15026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3530 ( .C ( clk ), .D ( new_AGEMA_signal_15029 ), .Q ( new_AGEMA_signal_15030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3534 ( .C ( clk ), .D ( new_AGEMA_signal_15033 ), .Q ( new_AGEMA_signal_15034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3538 ( .C ( clk ), .D ( new_AGEMA_signal_15037 ), .Q ( new_AGEMA_signal_15038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3542 ( .C ( clk ), .D ( new_AGEMA_signal_15041 ), .Q ( new_AGEMA_signal_15042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3546 ( .C ( clk ), .D ( new_AGEMA_signal_15045 ), .Q ( new_AGEMA_signal_15046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3550 ( .C ( clk ), .D ( new_AGEMA_signal_15049 ), .Q ( new_AGEMA_signal_15050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3554 ( .C ( clk ), .D ( new_AGEMA_signal_15053 ), .Q ( new_AGEMA_signal_15054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3558 ( .C ( clk ), .D ( new_AGEMA_signal_15057 ), .Q ( new_AGEMA_signal_15058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3560 ( .C ( clk ), .D ( new_AGEMA_signal_15059 ), .Q ( new_AGEMA_signal_15060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3562 ( .C ( clk ), .D ( new_AGEMA_signal_15061 ), .Q ( new_AGEMA_signal_15062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3564 ( .C ( clk ), .D ( new_AGEMA_signal_15063 ), .Q ( new_AGEMA_signal_15064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3566 ( .C ( clk ), .D ( new_AGEMA_signal_15065 ), .Q ( new_AGEMA_signal_15066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3568 ( .C ( clk ), .D ( new_AGEMA_signal_15067 ), .Q ( new_AGEMA_signal_15068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3570 ( .C ( clk ), .D ( new_AGEMA_signal_15069 ), .Q ( new_AGEMA_signal_15070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3572 ( .C ( clk ), .D ( new_AGEMA_signal_15071 ), .Q ( new_AGEMA_signal_15072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3574 ( .C ( clk ), .D ( new_AGEMA_signal_15073 ), .Q ( new_AGEMA_signal_15074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3578 ( .C ( clk ), .D ( new_AGEMA_signal_15077 ), .Q ( new_AGEMA_signal_15078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3582 ( .C ( clk ), .D ( new_AGEMA_signal_15081 ), .Q ( new_AGEMA_signal_15082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3586 ( .C ( clk ), .D ( new_AGEMA_signal_15085 ), .Q ( new_AGEMA_signal_15086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3590 ( .C ( clk ), .D ( new_AGEMA_signal_15089 ), .Q ( new_AGEMA_signal_15090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3594 ( .C ( clk ), .D ( new_AGEMA_signal_15093 ), .Q ( new_AGEMA_signal_15094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3598 ( .C ( clk ), .D ( new_AGEMA_signal_15097 ), .Q ( new_AGEMA_signal_15098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3602 ( .C ( clk ), .D ( new_AGEMA_signal_15101 ), .Q ( new_AGEMA_signal_15102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3606 ( .C ( clk ), .D ( new_AGEMA_signal_15105 ), .Q ( new_AGEMA_signal_15106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3608 ( .C ( clk ), .D ( new_AGEMA_signal_15107 ), .Q ( new_AGEMA_signal_15108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3610 ( .C ( clk ), .D ( new_AGEMA_signal_15109 ), .Q ( new_AGEMA_signal_15110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3612 ( .C ( clk ), .D ( new_AGEMA_signal_15111 ), .Q ( new_AGEMA_signal_15112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3614 ( .C ( clk ), .D ( new_AGEMA_signal_15113 ), .Q ( new_AGEMA_signal_15114 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3620 ( .C ( clk ), .D ( new_AGEMA_signal_15119 ), .Q ( new_AGEMA_signal_15120 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3626 ( .C ( clk ), .D ( new_AGEMA_signal_15125 ), .Q ( new_AGEMA_signal_15126 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3632 ( .C ( clk ), .D ( new_AGEMA_signal_15131 ), .Q ( new_AGEMA_signal_15132 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3638 ( .C ( clk ), .D ( new_AGEMA_signal_15137 ), .Q ( new_AGEMA_signal_15138 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3642 ( .C ( clk ), .D ( new_AGEMA_signal_15141 ), .Q ( new_AGEMA_signal_15142 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3646 ( .C ( clk ), .D ( new_AGEMA_signal_15145 ), .Q ( new_AGEMA_signal_15146 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3650 ( .C ( clk ), .D ( new_AGEMA_signal_15149 ), .Q ( new_AGEMA_signal_15150 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3654 ( .C ( clk ), .D ( new_AGEMA_signal_15153 ), .Q ( new_AGEMA_signal_15154 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3656 ( .C ( clk ), .D ( new_AGEMA_signal_15155 ), .Q ( new_AGEMA_signal_15156 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3658 ( .C ( clk ), .D ( new_AGEMA_signal_15157 ), .Q ( new_AGEMA_signal_15158 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3660 ( .C ( clk ), .D ( new_AGEMA_signal_15159 ), .Q ( new_AGEMA_signal_15160 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3662 ( .C ( clk ), .D ( new_AGEMA_signal_15161 ), .Q ( new_AGEMA_signal_15162 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3666 ( .C ( clk ), .D ( new_AGEMA_signal_15165 ), .Q ( new_AGEMA_signal_15166 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3670 ( .C ( clk ), .D ( new_AGEMA_signal_15169 ), .Q ( new_AGEMA_signal_15170 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3674 ( .C ( clk ), .D ( new_AGEMA_signal_15173 ), .Q ( new_AGEMA_signal_15174 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3678 ( .C ( clk ), .D ( new_AGEMA_signal_15177 ), .Q ( new_AGEMA_signal_15178 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3682 ( .C ( clk ), .D ( new_AGEMA_signal_15181 ), .Q ( new_AGEMA_signal_15182 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3686 ( .C ( clk ), .D ( new_AGEMA_signal_15185 ), .Q ( new_AGEMA_signal_15186 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3690 ( .C ( clk ), .D ( new_AGEMA_signal_15189 ), .Q ( new_AGEMA_signal_15190 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3694 ( .C ( clk ), .D ( new_AGEMA_signal_15193 ), .Q ( new_AGEMA_signal_15194 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3698 ( .C ( clk ), .D ( new_AGEMA_signal_15197 ), .Q ( new_AGEMA_signal_15198 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3702 ( .C ( clk ), .D ( new_AGEMA_signal_15201 ), .Q ( new_AGEMA_signal_15202 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3706 ( .C ( clk ), .D ( new_AGEMA_signal_15205 ), .Q ( new_AGEMA_signal_15206 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3710 ( .C ( clk ), .D ( new_AGEMA_signal_15209 ), .Q ( new_AGEMA_signal_15210 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3712 ( .C ( clk ), .D ( new_AGEMA_signal_15211 ), .Q ( new_AGEMA_signal_15212 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3714 ( .C ( clk ), .D ( new_AGEMA_signal_15213 ), .Q ( new_AGEMA_signal_15214 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3716 ( .C ( clk ), .D ( new_AGEMA_signal_15215 ), .Q ( new_AGEMA_signal_15216 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3718 ( .C ( clk ), .D ( new_AGEMA_signal_15217 ), .Q ( new_AGEMA_signal_15218 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3722 ( .C ( clk ), .D ( new_AGEMA_signal_15221 ), .Q ( new_AGEMA_signal_15222 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3726 ( .C ( clk ), .D ( new_AGEMA_signal_15225 ), .Q ( new_AGEMA_signal_15226 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3730 ( .C ( clk ), .D ( new_AGEMA_signal_15229 ), .Q ( new_AGEMA_signal_15230 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3734 ( .C ( clk ), .D ( new_AGEMA_signal_15233 ), .Q ( new_AGEMA_signal_15234 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3736 ( .C ( clk ), .D ( new_AGEMA_signal_15235 ), .Q ( new_AGEMA_signal_15236 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3738 ( .C ( clk ), .D ( new_AGEMA_signal_15237 ), .Q ( new_AGEMA_signal_15238 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3740 ( .C ( clk ), .D ( new_AGEMA_signal_15239 ), .Q ( new_AGEMA_signal_15240 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3742 ( .C ( clk ), .D ( new_AGEMA_signal_15241 ), .Q ( new_AGEMA_signal_15242 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3748 ( .C ( clk ), .D ( new_AGEMA_signal_15247 ), .Q ( new_AGEMA_signal_15248 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3754 ( .C ( clk ), .D ( new_AGEMA_signal_15253 ), .Q ( new_AGEMA_signal_15254 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3760 ( .C ( clk ), .D ( new_AGEMA_signal_15259 ), .Q ( new_AGEMA_signal_15260 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3766 ( .C ( clk ), .D ( new_AGEMA_signal_15265 ), .Q ( new_AGEMA_signal_15266 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3772 ( .C ( clk ), .D ( new_AGEMA_signal_15271 ), .Q ( new_AGEMA_signal_15272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3778 ( .C ( clk ), .D ( new_AGEMA_signal_15277 ), .Q ( new_AGEMA_signal_15278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3784 ( .C ( clk ), .D ( new_AGEMA_signal_15283 ), .Q ( new_AGEMA_signal_15284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3790 ( .C ( clk ), .D ( new_AGEMA_signal_15289 ), .Q ( new_AGEMA_signal_15290 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3794 ( .C ( clk ), .D ( new_AGEMA_signal_15293 ), .Q ( new_AGEMA_signal_15294 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3798 ( .C ( clk ), .D ( new_AGEMA_signal_15297 ), .Q ( new_AGEMA_signal_15298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3802 ( .C ( clk ), .D ( new_AGEMA_signal_15301 ), .Q ( new_AGEMA_signal_15302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3806 ( .C ( clk ), .D ( new_AGEMA_signal_15305 ), .Q ( new_AGEMA_signal_15306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3808 ( .C ( clk ), .D ( new_AGEMA_signal_15307 ), .Q ( new_AGEMA_signal_15308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3810 ( .C ( clk ), .D ( new_AGEMA_signal_15309 ), .Q ( new_AGEMA_signal_15310 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3812 ( .C ( clk ), .D ( new_AGEMA_signal_15311 ), .Q ( new_AGEMA_signal_15312 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3814 ( .C ( clk ), .D ( new_AGEMA_signal_15313 ), .Q ( new_AGEMA_signal_15314 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3822 ( .C ( clk ), .D ( new_AGEMA_signal_15321 ), .Q ( new_AGEMA_signal_15322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3830 ( .C ( clk ), .D ( new_AGEMA_signal_15329 ), .Q ( new_AGEMA_signal_15330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3838 ( .C ( clk ), .D ( new_AGEMA_signal_15337 ), .Q ( new_AGEMA_signal_15338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3846 ( .C ( clk ), .D ( new_AGEMA_signal_15345 ), .Q ( new_AGEMA_signal_15346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3848 ( .C ( clk ), .D ( new_AGEMA_signal_15347 ), .Q ( new_AGEMA_signal_15348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3850 ( .C ( clk ), .D ( new_AGEMA_signal_15349 ), .Q ( new_AGEMA_signal_15350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3852 ( .C ( clk ), .D ( new_AGEMA_signal_15351 ), .Q ( new_AGEMA_signal_15352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3854 ( .C ( clk ), .D ( new_AGEMA_signal_15353 ), .Q ( new_AGEMA_signal_15354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3858 ( .C ( clk ), .D ( new_AGEMA_signal_15357 ), .Q ( new_AGEMA_signal_15358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3862 ( .C ( clk ), .D ( new_AGEMA_signal_15361 ), .Q ( new_AGEMA_signal_15362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3866 ( .C ( clk ), .D ( new_AGEMA_signal_15365 ), .Q ( new_AGEMA_signal_15366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3870 ( .C ( clk ), .D ( new_AGEMA_signal_15369 ), .Q ( new_AGEMA_signal_15370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3874 ( .C ( clk ), .D ( new_AGEMA_signal_15373 ), .Q ( new_AGEMA_signal_15374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3878 ( .C ( clk ), .D ( new_AGEMA_signal_15377 ), .Q ( new_AGEMA_signal_15378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3882 ( .C ( clk ), .D ( new_AGEMA_signal_15381 ), .Q ( new_AGEMA_signal_15382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3886 ( .C ( clk ), .D ( new_AGEMA_signal_15385 ), .Q ( new_AGEMA_signal_15386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3890 ( .C ( clk ), .D ( new_AGEMA_signal_15389 ), .Q ( new_AGEMA_signal_15390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3894 ( .C ( clk ), .D ( new_AGEMA_signal_15393 ), .Q ( new_AGEMA_signal_15394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3898 ( .C ( clk ), .D ( new_AGEMA_signal_15397 ), .Q ( new_AGEMA_signal_15398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3902 ( .C ( clk ), .D ( new_AGEMA_signal_15401 ), .Q ( new_AGEMA_signal_15402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3906 ( .C ( clk ), .D ( new_AGEMA_signal_15405 ), .Q ( new_AGEMA_signal_15406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3910 ( .C ( clk ), .D ( new_AGEMA_signal_15409 ), .Q ( new_AGEMA_signal_15410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3914 ( .C ( clk ), .D ( new_AGEMA_signal_15413 ), .Q ( new_AGEMA_signal_15414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3918 ( .C ( clk ), .D ( new_AGEMA_signal_15417 ), .Q ( new_AGEMA_signal_15418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3922 ( .C ( clk ), .D ( new_AGEMA_signal_15421 ), .Q ( new_AGEMA_signal_15422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3926 ( .C ( clk ), .D ( new_AGEMA_signal_15425 ), .Q ( new_AGEMA_signal_15426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3930 ( .C ( clk ), .D ( new_AGEMA_signal_15429 ), .Q ( new_AGEMA_signal_15430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3934 ( .C ( clk ), .D ( new_AGEMA_signal_15433 ), .Q ( new_AGEMA_signal_15434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3942 ( .C ( clk ), .D ( new_AGEMA_signal_15441 ), .Q ( new_AGEMA_signal_15442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3950 ( .C ( clk ), .D ( new_AGEMA_signal_15449 ), .Q ( new_AGEMA_signal_15450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3958 ( .C ( clk ), .D ( new_AGEMA_signal_15457 ), .Q ( new_AGEMA_signal_15458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3966 ( .C ( clk ), .D ( new_AGEMA_signal_15465 ), .Q ( new_AGEMA_signal_15466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3968 ( .C ( clk ), .D ( new_AGEMA_signal_15467 ), .Q ( new_AGEMA_signal_15468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3970 ( .C ( clk ), .D ( new_AGEMA_signal_15469 ), .Q ( new_AGEMA_signal_15470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3972 ( .C ( clk ), .D ( new_AGEMA_signal_15471 ), .Q ( new_AGEMA_signal_15472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3974 ( .C ( clk ), .D ( new_AGEMA_signal_15473 ), .Q ( new_AGEMA_signal_15474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3978 ( .C ( clk ), .D ( new_AGEMA_signal_15477 ), .Q ( new_AGEMA_signal_15478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3982 ( .C ( clk ), .D ( new_AGEMA_signal_15481 ), .Q ( new_AGEMA_signal_15482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3986 ( .C ( clk ), .D ( new_AGEMA_signal_15485 ), .Q ( new_AGEMA_signal_15486 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3990 ( .C ( clk ), .D ( new_AGEMA_signal_15489 ), .Q ( new_AGEMA_signal_15490 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3992 ( .C ( clk ), .D ( new_AGEMA_signal_15491 ), .Q ( new_AGEMA_signal_15492 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3994 ( .C ( clk ), .D ( new_AGEMA_signal_15493 ), .Q ( new_AGEMA_signal_15494 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3996 ( .C ( clk ), .D ( new_AGEMA_signal_15495 ), .Q ( new_AGEMA_signal_15496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3998 ( .C ( clk ), .D ( new_AGEMA_signal_15497 ), .Q ( new_AGEMA_signal_15498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4004 ( .C ( clk ), .D ( new_AGEMA_signal_15503 ), .Q ( new_AGEMA_signal_15504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4010 ( .C ( clk ), .D ( new_AGEMA_signal_15509 ), .Q ( new_AGEMA_signal_15510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4016 ( .C ( clk ), .D ( new_AGEMA_signal_15515 ), .Q ( new_AGEMA_signal_15516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4022 ( .C ( clk ), .D ( new_AGEMA_signal_15521 ), .Q ( new_AGEMA_signal_15522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4036 ( .C ( clk ), .D ( new_AGEMA_signal_15535 ), .Q ( new_AGEMA_signal_15536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4044 ( .C ( clk ), .D ( new_AGEMA_signal_15543 ), .Q ( new_AGEMA_signal_15544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4052 ( .C ( clk ), .D ( new_AGEMA_signal_15551 ), .Q ( new_AGEMA_signal_15552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4060 ( .C ( clk ), .D ( new_AGEMA_signal_15559 ), .Q ( new_AGEMA_signal_15560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4072 ( .C ( clk ), .D ( new_AGEMA_signal_15571 ), .Q ( new_AGEMA_signal_15572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4076 ( .C ( clk ), .D ( new_AGEMA_signal_15575 ), .Q ( new_AGEMA_signal_15576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4080 ( .C ( clk ), .D ( new_AGEMA_signal_15579 ), .Q ( new_AGEMA_signal_15580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4084 ( .C ( clk ), .D ( new_AGEMA_signal_15583 ), .Q ( new_AGEMA_signal_15584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4092 ( .C ( clk ), .D ( new_AGEMA_signal_15591 ), .Q ( new_AGEMA_signal_15592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4100 ( .C ( clk ), .D ( new_AGEMA_signal_15599 ), .Q ( new_AGEMA_signal_15600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4108 ( .C ( clk ), .D ( new_AGEMA_signal_15607 ), .Q ( new_AGEMA_signal_15608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4116 ( .C ( clk ), .D ( new_AGEMA_signal_15615 ), .Q ( new_AGEMA_signal_15616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4130 ( .C ( clk ), .D ( new_AGEMA_signal_15629 ), .Q ( new_AGEMA_signal_15630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4136 ( .C ( clk ), .D ( new_AGEMA_signal_15635 ), .Q ( new_AGEMA_signal_15636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4142 ( .C ( clk ), .D ( new_AGEMA_signal_15641 ), .Q ( new_AGEMA_signal_15642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4148 ( .C ( clk ), .D ( new_AGEMA_signal_15647 ), .Q ( new_AGEMA_signal_15648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4152 ( .C ( clk ), .D ( new_AGEMA_signal_15651 ), .Q ( new_AGEMA_signal_15652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4156 ( .C ( clk ), .D ( new_AGEMA_signal_15655 ), .Q ( new_AGEMA_signal_15656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4160 ( .C ( clk ), .D ( new_AGEMA_signal_15659 ), .Q ( new_AGEMA_signal_15660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4164 ( .C ( clk ), .D ( new_AGEMA_signal_15663 ), .Q ( new_AGEMA_signal_15664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4172 ( .C ( clk ), .D ( new_AGEMA_signal_15671 ), .Q ( new_AGEMA_signal_15672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4180 ( .C ( clk ), .D ( new_AGEMA_signal_15679 ), .Q ( new_AGEMA_signal_15680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4188 ( .C ( clk ), .D ( new_AGEMA_signal_15687 ), .Q ( new_AGEMA_signal_15688 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4196 ( .C ( clk ), .D ( new_AGEMA_signal_15695 ), .Q ( new_AGEMA_signal_15696 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4200 ( .C ( clk ), .D ( new_AGEMA_signal_15699 ), .Q ( new_AGEMA_signal_15700 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4204 ( .C ( clk ), .D ( new_AGEMA_signal_15703 ), .Q ( new_AGEMA_signal_15704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4208 ( .C ( clk ), .D ( new_AGEMA_signal_15707 ), .Q ( new_AGEMA_signal_15708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4212 ( .C ( clk ), .D ( new_AGEMA_signal_15711 ), .Q ( new_AGEMA_signal_15712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4218 ( .C ( clk ), .D ( new_AGEMA_signal_15717 ), .Q ( new_AGEMA_signal_15718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4224 ( .C ( clk ), .D ( new_AGEMA_signal_15723 ), .Q ( new_AGEMA_signal_15724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4230 ( .C ( clk ), .D ( new_AGEMA_signal_15729 ), .Q ( new_AGEMA_signal_15730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4236 ( .C ( clk ), .D ( new_AGEMA_signal_15735 ), .Q ( new_AGEMA_signal_15736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4242 ( .C ( clk ), .D ( new_AGEMA_signal_15741 ), .Q ( new_AGEMA_signal_15742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4248 ( .C ( clk ), .D ( new_AGEMA_signal_15747 ), .Q ( new_AGEMA_signal_15748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4254 ( .C ( clk ), .D ( new_AGEMA_signal_15753 ), .Q ( new_AGEMA_signal_15754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4260 ( .C ( clk ), .D ( new_AGEMA_signal_15759 ), .Q ( new_AGEMA_signal_15760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4266 ( .C ( clk ), .D ( new_AGEMA_signal_15765 ), .Q ( new_AGEMA_signal_15766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4272 ( .C ( clk ), .D ( new_AGEMA_signal_15771 ), .Q ( new_AGEMA_signal_15772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4278 ( .C ( clk ), .D ( new_AGEMA_signal_15777 ), .Q ( new_AGEMA_signal_15778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4284 ( .C ( clk ), .D ( new_AGEMA_signal_15783 ), .Q ( new_AGEMA_signal_15784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4290 ( .C ( clk ), .D ( new_AGEMA_signal_15789 ), .Q ( new_AGEMA_signal_15790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4296 ( .C ( clk ), .D ( new_AGEMA_signal_15795 ), .Q ( new_AGEMA_signal_15796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4302 ( .C ( clk ), .D ( new_AGEMA_signal_15801 ), .Q ( new_AGEMA_signal_15802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4308 ( .C ( clk ), .D ( new_AGEMA_signal_15807 ), .Q ( new_AGEMA_signal_15808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4314 ( .C ( clk ), .D ( new_AGEMA_signal_15813 ), .Q ( new_AGEMA_signal_15814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4320 ( .C ( clk ), .D ( new_AGEMA_signal_15819 ), .Q ( new_AGEMA_signal_15820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4326 ( .C ( clk ), .D ( new_AGEMA_signal_15825 ), .Q ( new_AGEMA_signal_15826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4332 ( .C ( clk ), .D ( new_AGEMA_signal_15831 ), .Q ( new_AGEMA_signal_15832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4336 ( .C ( clk ), .D ( new_AGEMA_signal_15835 ), .Q ( new_AGEMA_signal_15836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4340 ( .C ( clk ), .D ( new_AGEMA_signal_15839 ), .Q ( new_AGEMA_signal_15840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4344 ( .C ( clk ), .D ( new_AGEMA_signal_15843 ), .Q ( new_AGEMA_signal_15844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4348 ( .C ( clk ), .D ( new_AGEMA_signal_15847 ), .Q ( new_AGEMA_signal_15848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4356 ( .C ( clk ), .D ( new_AGEMA_signal_15855 ), .Q ( new_AGEMA_signal_15856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4364 ( .C ( clk ), .D ( new_AGEMA_signal_15863 ), .Q ( new_AGEMA_signal_15864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4372 ( .C ( clk ), .D ( new_AGEMA_signal_15871 ), .Q ( new_AGEMA_signal_15872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4380 ( .C ( clk ), .D ( new_AGEMA_signal_15879 ), .Q ( new_AGEMA_signal_15880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4384 ( .C ( clk ), .D ( new_AGEMA_signal_15883 ), .Q ( new_AGEMA_signal_15884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4388 ( .C ( clk ), .D ( new_AGEMA_signal_15887 ), .Q ( new_AGEMA_signal_15888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4392 ( .C ( clk ), .D ( new_AGEMA_signal_15891 ), .Q ( new_AGEMA_signal_15892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4396 ( .C ( clk ), .D ( new_AGEMA_signal_15895 ), .Q ( new_AGEMA_signal_15896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4402 ( .C ( clk ), .D ( new_AGEMA_signal_15901 ), .Q ( new_AGEMA_signal_15902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4408 ( .C ( clk ), .D ( new_AGEMA_signal_15907 ), .Q ( new_AGEMA_signal_15908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4414 ( .C ( clk ), .D ( new_AGEMA_signal_15913 ), .Q ( new_AGEMA_signal_15914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4420 ( .C ( clk ), .D ( new_AGEMA_signal_15919 ), .Q ( new_AGEMA_signal_15920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4428 ( .C ( clk ), .D ( new_AGEMA_signal_15927 ), .Q ( new_AGEMA_signal_15928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4436 ( .C ( clk ), .D ( new_AGEMA_signal_15935 ), .Q ( new_AGEMA_signal_15936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4444 ( .C ( clk ), .D ( new_AGEMA_signal_15943 ), .Q ( new_AGEMA_signal_15944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4452 ( .C ( clk ), .D ( new_AGEMA_signal_15951 ), .Q ( new_AGEMA_signal_15952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4466 ( .C ( clk ), .D ( new_AGEMA_signal_15965 ), .Q ( new_AGEMA_signal_15966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4472 ( .C ( clk ), .D ( new_AGEMA_signal_15971 ), .Q ( new_AGEMA_signal_15972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4478 ( .C ( clk ), .D ( new_AGEMA_signal_15977 ), .Q ( new_AGEMA_signal_15978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4484 ( .C ( clk ), .D ( new_AGEMA_signal_15983 ), .Q ( new_AGEMA_signal_15984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4506 ( .C ( clk ), .D ( new_AGEMA_signal_16005 ), .Q ( new_AGEMA_signal_16006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4512 ( .C ( clk ), .D ( new_AGEMA_signal_16011 ), .Q ( new_AGEMA_signal_16012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4518 ( .C ( clk ), .D ( new_AGEMA_signal_16017 ), .Q ( new_AGEMA_signal_16018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4524 ( .C ( clk ), .D ( new_AGEMA_signal_16023 ), .Q ( new_AGEMA_signal_16024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4530 ( .C ( clk ), .D ( new_AGEMA_signal_16029 ), .Q ( new_AGEMA_signal_16030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4536 ( .C ( clk ), .D ( new_AGEMA_signal_16035 ), .Q ( new_AGEMA_signal_16036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4542 ( .C ( clk ), .D ( new_AGEMA_signal_16041 ), .Q ( new_AGEMA_signal_16042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4548 ( .C ( clk ), .D ( new_AGEMA_signal_16047 ), .Q ( new_AGEMA_signal_16048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4556 ( .C ( clk ), .D ( new_AGEMA_signal_16055 ), .Q ( new_AGEMA_signal_16056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4564 ( .C ( clk ), .D ( new_AGEMA_signal_16063 ), .Q ( new_AGEMA_signal_16064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4572 ( .C ( clk ), .D ( new_AGEMA_signal_16071 ), .Q ( new_AGEMA_signal_16072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4580 ( .C ( clk ), .D ( new_AGEMA_signal_16079 ), .Q ( new_AGEMA_signal_16080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4588 ( .C ( clk ), .D ( new_AGEMA_signal_16087 ), .Q ( new_AGEMA_signal_16088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4596 ( .C ( clk ), .D ( new_AGEMA_signal_16095 ), .Q ( new_AGEMA_signal_16096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4604 ( .C ( clk ), .D ( new_AGEMA_signal_16103 ), .Q ( new_AGEMA_signal_16104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4612 ( .C ( clk ), .D ( new_AGEMA_signal_16111 ), .Q ( new_AGEMA_signal_16112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4618 ( .C ( clk ), .D ( new_AGEMA_signal_16117 ), .Q ( new_AGEMA_signal_16118 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4624 ( .C ( clk ), .D ( new_AGEMA_signal_16123 ), .Q ( new_AGEMA_signal_16124 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4630 ( .C ( clk ), .D ( new_AGEMA_signal_16129 ), .Q ( new_AGEMA_signal_16130 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4636 ( .C ( clk ), .D ( new_AGEMA_signal_16135 ), .Q ( new_AGEMA_signal_16136 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4642 ( .C ( clk ), .D ( new_AGEMA_signal_16141 ), .Q ( new_AGEMA_signal_16142 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4648 ( .C ( clk ), .D ( new_AGEMA_signal_16147 ), .Q ( new_AGEMA_signal_16148 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4654 ( .C ( clk ), .D ( new_AGEMA_signal_16153 ), .Q ( new_AGEMA_signal_16154 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4660 ( .C ( clk ), .D ( new_AGEMA_signal_16159 ), .Q ( new_AGEMA_signal_16160 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4672 ( .C ( clk ), .D ( new_AGEMA_signal_16171 ), .Q ( new_AGEMA_signal_16172 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4676 ( .C ( clk ), .D ( new_AGEMA_signal_16175 ), .Q ( new_AGEMA_signal_16176 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4680 ( .C ( clk ), .D ( new_AGEMA_signal_16179 ), .Q ( new_AGEMA_signal_16180 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4684 ( .C ( clk ), .D ( new_AGEMA_signal_16183 ), .Q ( new_AGEMA_signal_16184 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4688 ( .C ( clk ), .D ( new_AGEMA_signal_16187 ), .Q ( new_AGEMA_signal_16188 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4692 ( .C ( clk ), .D ( new_AGEMA_signal_16191 ), .Q ( new_AGEMA_signal_16192 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4696 ( .C ( clk ), .D ( new_AGEMA_signal_16195 ), .Q ( new_AGEMA_signal_16196 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4700 ( .C ( clk ), .D ( new_AGEMA_signal_16199 ), .Q ( new_AGEMA_signal_16200 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4704 ( .C ( clk ), .D ( new_AGEMA_signal_16203 ), .Q ( new_AGEMA_signal_16204 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4708 ( .C ( clk ), .D ( new_AGEMA_signal_16207 ), .Q ( new_AGEMA_signal_16208 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4712 ( .C ( clk ), .D ( new_AGEMA_signal_16211 ), .Q ( new_AGEMA_signal_16212 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4716 ( .C ( clk ), .D ( new_AGEMA_signal_16215 ), .Q ( new_AGEMA_signal_16216 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4728 ( .C ( clk ), .D ( new_AGEMA_signal_16227 ), .Q ( new_AGEMA_signal_16228 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4734 ( .C ( clk ), .D ( new_AGEMA_signal_16233 ), .Q ( new_AGEMA_signal_16234 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4740 ( .C ( clk ), .D ( new_AGEMA_signal_16239 ), .Q ( new_AGEMA_signal_16240 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4746 ( .C ( clk ), .D ( new_AGEMA_signal_16245 ), .Q ( new_AGEMA_signal_16246 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4778 ( .C ( clk ), .D ( new_AGEMA_signal_16277 ), .Q ( new_AGEMA_signal_16278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4786 ( .C ( clk ), .D ( new_AGEMA_signal_16285 ), .Q ( new_AGEMA_signal_16286 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4794 ( .C ( clk ), .D ( new_AGEMA_signal_16293 ), .Q ( new_AGEMA_signal_16294 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4802 ( .C ( clk ), .D ( new_AGEMA_signal_16301 ), .Q ( new_AGEMA_signal_16302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4810 ( .C ( clk ), .D ( new_AGEMA_signal_16309 ), .Q ( new_AGEMA_signal_16310 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4818 ( .C ( clk ), .D ( new_AGEMA_signal_16317 ), .Q ( new_AGEMA_signal_16318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4826 ( .C ( clk ), .D ( new_AGEMA_signal_16325 ), .Q ( new_AGEMA_signal_16326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4834 ( .C ( clk ), .D ( new_AGEMA_signal_16333 ), .Q ( new_AGEMA_signal_16334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4842 ( .C ( clk ), .D ( new_AGEMA_signal_16341 ), .Q ( new_AGEMA_signal_16342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4850 ( .C ( clk ), .D ( new_AGEMA_signal_16349 ), .Q ( new_AGEMA_signal_16350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4858 ( .C ( clk ), .D ( new_AGEMA_signal_16357 ), .Q ( new_AGEMA_signal_16358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4866 ( .C ( clk ), .D ( new_AGEMA_signal_16365 ), .Q ( new_AGEMA_signal_16366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4874 ( .C ( clk ), .D ( new_AGEMA_signal_16373 ), .Q ( new_AGEMA_signal_16374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4882 ( .C ( clk ), .D ( new_AGEMA_signal_16381 ), .Q ( new_AGEMA_signal_16382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4890 ( .C ( clk ), .D ( new_AGEMA_signal_16389 ), .Q ( new_AGEMA_signal_16390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4898 ( .C ( clk ), .D ( new_AGEMA_signal_16397 ), .Q ( new_AGEMA_signal_16398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4904 ( .C ( clk ), .D ( new_AGEMA_signal_16403 ), .Q ( new_AGEMA_signal_16404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4910 ( .C ( clk ), .D ( new_AGEMA_signal_16409 ), .Q ( new_AGEMA_signal_16410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4916 ( .C ( clk ), .D ( new_AGEMA_signal_16415 ), .Q ( new_AGEMA_signal_16416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4922 ( .C ( clk ), .D ( new_AGEMA_signal_16421 ), .Q ( new_AGEMA_signal_16422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4932 ( .C ( clk ), .D ( new_AGEMA_signal_16431 ), .Q ( new_AGEMA_signal_16432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4942 ( .C ( clk ), .D ( new_AGEMA_signal_16441 ), .Q ( new_AGEMA_signal_16442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4952 ( .C ( clk ), .D ( new_AGEMA_signal_16451 ), .Q ( new_AGEMA_signal_16452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4962 ( .C ( clk ), .D ( new_AGEMA_signal_16461 ), .Q ( new_AGEMA_signal_16462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4970 ( .C ( clk ), .D ( new_AGEMA_signal_16469 ), .Q ( new_AGEMA_signal_16470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4978 ( .C ( clk ), .D ( new_AGEMA_signal_16477 ), .Q ( new_AGEMA_signal_16478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4986 ( .C ( clk ), .D ( new_AGEMA_signal_16485 ), .Q ( new_AGEMA_signal_16486 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4994 ( .C ( clk ), .D ( new_AGEMA_signal_16493 ), .Q ( new_AGEMA_signal_16494 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5002 ( .C ( clk ), .D ( new_AGEMA_signal_16501 ), .Q ( new_AGEMA_signal_16502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5010 ( .C ( clk ), .D ( new_AGEMA_signal_16509 ), .Q ( new_AGEMA_signal_16510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5018 ( .C ( clk ), .D ( new_AGEMA_signal_16517 ), .Q ( new_AGEMA_signal_16518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5026 ( .C ( clk ), .D ( new_AGEMA_signal_16525 ), .Q ( new_AGEMA_signal_16526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5034 ( .C ( clk ), .D ( new_AGEMA_signal_16533 ), .Q ( new_AGEMA_signal_16534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5042 ( .C ( clk ), .D ( new_AGEMA_signal_16541 ), .Q ( new_AGEMA_signal_16542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5050 ( .C ( clk ), .D ( new_AGEMA_signal_16549 ), .Q ( new_AGEMA_signal_16550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5058 ( .C ( clk ), .D ( new_AGEMA_signal_16557 ), .Q ( new_AGEMA_signal_16558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5088 ( .C ( clk ), .D ( new_AGEMA_signal_16587 ), .Q ( new_AGEMA_signal_16588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5094 ( .C ( clk ), .D ( new_AGEMA_signal_16593 ), .Q ( new_AGEMA_signal_16594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5100 ( .C ( clk ), .D ( new_AGEMA_signal_16599 ), .Q ( new_AGEMA_signal_16600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5106 ( .C ( clk ), .D ( new_AGEMA_signal_16605 ), .Q ( new_AGEMA_signal_16606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5132 ( .C ( clk ), .D ( new_AGEMA_signal_16631 ), .Q ( new_AGEMA_signal_16632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5142 ( .C ( clk ), .D ( new_AGEMA_signal_16641 ), .Q ( new_AGEMA_signal_16642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5152 ( .C ( clk ), .D ( new_AGEMA_signal_16651 ), .Q ( new_AGEMA_signal_16652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5162 ( .C ( clk ), .D ( new_AGEMA_signal_16661 ), .Q ( new_AGEMA_signal_16662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5170 ( .C ( clk ), .D ( new_AGEMA_signal_16669 ), .Q ( new_AGEMA_signal_16670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5178 ( .C ( clk ), .D ( new_AGEMA_signal_16677 ), .Q ( new_AGEMA_signal_16678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5186 ( .C ( clk ), .D ( new_AGEMA_signal_16685 ), .Q ( new_AGEMA_signal_16686 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5194 ( .C ( clk ), .D ( new_AGEMA_signal_16693 ), .Q ( new_AGEMA_signal_16694 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5226 ( .C ( clk ), .D ( new_AGEMA_signal_16725 ), .Q ( new_AGEMA_signal_16726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5234 ( .C ( clk ), .D ( new_AGEMA_signal_16733 ), .Q ( new_AGEMA_signal_16734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5242 ( .C ( clk ), .D ( new_AGEMA_signal_16741 ), .Q ( new_AGEMA_signal_16742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5250 ( .C ( clk ), .D ( new_AGEMA_signal_16749 ), .Q ( new_AGEMA_signal_16750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5258 ( .C ( clk ), .D ( new_AGEMA_signal_16757 ), .Q ( new_AGEMA_signal_16758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5266 ( .C ( clk ), .D ( new_AGEMA_signal_16765 ), .Q ( new_AGEMA_signal_16766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5274 ( .C ( clk ), .D ( new_AGEMA_signal_16773 ), .Q ( new_AGEMA_signal_16774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5282 ( .C ( clk ), .D ( new_AGEMA_signal_16781 ), .Q ( new_AGEMA_signal_16782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5288 ( .C ( clk ), .D ( new_AGEMA_signal_16787 ), .Q ( new_AGEMA_signal_16788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5294 ( .C ( clk ), .D ( new_AGEMA_signal_16793 ), .Q ( new_AGEMA_signal_16794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5300 ( .C ( clk ), .D ( new_AGEMA_signal_16799 ), .Q ( new_AGEMA_signal_16800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5306 ( .C ( clk ), .D ( new_AGEMA_signal_16805 ), .Q ( new_AGEMA_signal_16806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5330 ( .C ( clk ), .D ( new_AGEMA_signal_16829 ), .Q ( new_AGEMA_signal_16830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5338 ( .C ( clk ), .D ( new_AGEMA_signal_16837 ), .Q ( new_AGEMA_signal_16838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5346 ( .C ( clk ), .D ( new_AGEMA_signal_16845 ), .Q ( new_AGEMA_signal_16846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5354 ( .C ( clk ), .D ( new_AGEMA_signal_16853 ), .Q ( new_AGEMA_signal_16854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5456 ( .C ( clk ), .D ( new_AGEMA_signal_16955 ), .Q ( new_AGEMA_signal_16956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5464 ( .C ( clk ), .D ( new_AGEMA_signal_16963 ), .Q ( new_AGEMA_signal_16964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5472 ( .C ( clk ), .D ( new_AGEMA_signal_16971 ), .Q ( new_AGEMA_signal_16972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5480 ( .C ( clk ), .D ( new_AGEMA_signal_16979 ), .Q ( new_AGEMA_signal_16980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5528 ( .C ( clk ), .D ( new_AGEMA_signal_17027 ), .Q ( new_AGEMA_signal_17028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5536 ( .C ( clk ), .D ( new_AGEMA_signal_17035 ), .Q ( new_AGEMA_signal_17036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5544 ( .C ( clk ), .D ( new_AGEMA_signal_17043 ), .Q ( new_AGEMA_signal_17044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5552 ( .C ( clk ), .D ( new_AGEMA_signal_17051 ), .Q ( new_AGEMA_signal_17052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5560 ( .C ( clk ), .D ( new_AGEMA_signal_17059 ), .Q ( new_AGEMA_signal_17060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5568 ( .C ( clk ), .D ( new_AGEMA_signal_17067 ), .Q ( new_AGEMA_signal_17068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5576 ( .C ( clk ), .D ( new_AGEMA_signal_17075 ), .Q ( new_AGEMA_signal_17076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5584 ( .C ( clk ), .D ( new_AGEMA_signal_17083 ), .Q ( new_AGEMA_signal_17084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5594 ( .C ( clk ), .D ( new_AGEMA_signal_17093 ), .Q ( new_AGEMA_signal_17094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5604 ( .C ( clk ), .D ( new_AGEMA_signal_17103 ), .Q ( new_AGEMA_signal_17104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5614 ( .C ( clk ), .D ( new_AGEMA_signal_17113 ), .Q ( new_AGEMA_signal_17114 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5624 ( .C ( clk ), .D ( new_AGEMA_signal_17123 ), .Q ( new_AGEMA_signal_17124 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5632 ( .C ( clk ), .D ( new_AGEMA_signal_17131 ), .Q ( new_AGEMA_signal_17132 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5640 ( .C ( clk ), .D ( new_AGEMA_signal_17139 ), .Q ( new_AGEMA_signal_17140 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5648 ( .C ( clk ), .D ( new_AGEMA_signal_17147 ), .Q ( new_AGEMA_signal_17148 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5656 ( .C ( clk ), .D ( new_AGEMA_signal_17155 ), .Q ( new_AGEMA_signal_17156 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5728 ( .C ( clk ), .D ( new_AGEMA_signal_17227 ), .Q ( new_AGEMA_signal_17228 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5736 ( .C ( clk ), .D ( new_AGEMA_signal_17235 ), .Q ( new_AGEMA_signal_17236 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5744 ( .C ( clk ), .D ( new_AGEMA_signal_17243 ), .Q ( new_AGEMA_signal_17244 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5752 ( .C ( clk ), .D ( new_AGEMA_signal_17251 ), .Q ( new_AGEMA_signal_17252 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5792 ( .C ( clk ), .D ( new_AGEMA_signal_17291 ), .Q ( new_AGEMA_signal_17292 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5800 ( .C ( clk ), .D ( new_AGEMA_signal_17299 ), .Q ( new_AGEMA_signal_17300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5808 ( .C ( clk ), .D ( new_AGEMA_signal_17307 ), .Q ( new_AGEMA_signal_17308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5816 ( .C ( clk ), .D ( new_AGEMA_signal_17315 ), .Q ( new_AGEMA_signal_17316 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5968 ( .C ( clk ), .D ( new_AGEMA_signal_17467 ), .Q ( new_AGEMA_signal_17468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5978 ( .C ( clk ), .D ( new_AGEMA_signal_17477 ), .Q ( new_AGEMA_signal_17478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5988 ( .C ( clk ), .D ( new_AGEMA_signal_17487 ), .Q ( new_AGEMA_signal_17488 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5998 ( .C ( clk ), .D ( new_AGEMA_signal_17497 ), .Q ( new_AGEMA_signal_17498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6328 ( .C ( clk ), .D ( new_AGEMA_signal_17827 ), .Q ( new_AGEMA_signal_17828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6340 ( .C ( clk ), .D ( new_AGEMA_signal_17839 ), .Q ( new_AGEMA_signal_17840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6352 ( .C ( clk ), .D ( new_AGEMA_signal_17851 ), .Q ( new_AGEMA_signal_17852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6364 ( .C ( clk ), .D ( new_AGEMA_signal_17863 ), .Q ( new_AGEMA_signal_17864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6378 ( .C ( clk ), .D ( new_AGEMA_signal_17877 ), .Q ( new_AGEMA_signal_17878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6392 ( .C ( clk ), .D ( new_AGEMA_signal_17891 ), .Q ( new_AGEMA_signal_17892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6406 ( .C ( clk ), .D ( new_AGEMA_signal_17905 ), .Q ( new_AGEMA_signal_17906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6420 ( .C ( clk ), .D ( new_AGEMA_signal_17919 ), .Q ( new_AGEMA_signal_17920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6466 ( .C ( clk ), .D ( new_AGEMA_signal_17965 ), .Q ( new_AGEMA_signal_17966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6480 ( .C ( clk ), .D ( new_AGEMA_signal_17979 ), .Q ( new_AGEMA_signal_17980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6494 ( .C ( clk ), .D ( new_AGEMA_signal_17993 ), .Q ( new_AGEMA_signal_17994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6508 ( .C ( clk ), .D ( new_AGEMA_signal_18007 ), .Q ( new_AGEMA_signal_18008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6610 ( .C ( clk ), .D ( new_AGEMA_signal_18109 ), .Q ( new_AGEMA_signal_18110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6626 ( .C ( clk ), .D ( new_AGEMA_signal_18125 ), .Q ( new_AGEMA_signal_18126 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6642 ( .C ( clk ), .D ( new_AGEMA_signal_18141 ), .Q ( new_AGEMA_signal_18142 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6658 ( .C ( clk ), .D ( new_AGEMA_signal_18157 ), .Q ( new_AGEMA_signal_18158 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6698 ( .C ( clk ), .D ( new_AGEMA_signal_18197 ), .Q ( new_AGEMA_signal_18198 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6714 ( .C ( clk ), .D ( new_AGEMA_signal_18213 ), .Q ( new_AGEMA_signal_18214 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6730 ( .C ( clk ), .D ( new_AGEMA_signal_18229 ), .Q ( new_AGEMA_signal_18230 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6746 ( .C ( clk ), .D ( new_AGEMA_signal_18245 ), .Q ( new_AGEMA_signal_18246 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6896 ( .C ( clk ), .D ( new_AGEMA_signal_18395 ), .Q ( new_AGEMA_signal_18396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6912 ( .C ( clk ), .D ( new_AGEMA_signal_18411 ), .Q ( new_AGEMA_signal_18412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6928 ( .C ( clk ), .D ( new_AGEMA_signal_18427 ), .Q ( new_AGEMA_signal_18428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6944 ( .C ( clk ), .D ( new_AGEMA_signal_18443 ), .Q ( new_AGEMA_signal_18444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7002 ( .C ( clk ), .D ( new_AGEMA_signal_18501 ), .Q ( new_AGEMA_signal_18502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7020 ( .C ( clk ), .D ( new_AGEMA_signal_18519 ), .Q ( new_AGEMA_signal_18520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7038 ( .C ( clk ), .D ( new_AGEMA_signal_18537 ), .Q ( new_AGEMA_signal_18538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7056 ( .C ( clk ), .D ( new_AGEMA_signal_18555 ), .Q ( new_AGEMA_signal_18556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7202 ( .C ( clk ), .D ( new_AGEMA_signal_18701 ), .Q ( new_AGEMA_signal_18702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7222 ( .C ( clk ), .D ( new_AGEMA_signal_18721 ), .Q ( new_AGEMA_signal_18722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7242 ( .C ( clk ), .D ( new_AGEMA_signal_18741 ), .Q ( new_AGEMA_signal_18742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7262 ( .C ( clk ), .D ( new_AGEMA_signal_18761 ), .Q ( new_AGEMA_signal_18762 ) ) ;

    /* cells in depth 11 */
    buf_clk new_AGEMA_reg_buffer_4023 ( .C ( clk ), .D ( n1934 ), .Q ( new_AGEMA_signal_15523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4025 ( .C ( clk ), .D ( new_AGEMA_signal_2871 ), .Q ( new_AGEMA_signal_15525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4027 ( .C ( clk ), .D ( new_AGEMA_signal_2872 ), .Q ( new_AGEMA_signal_15527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4029 ( .C ( clk ), .D ( new_AGEMA_signal_2873 ), .Q ( new_AGEMA_signal_15529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4037 ( .C ( clk ), .D ( new_AGEMA_signal_15536 ), .Q ( new_AGEMA_signal_15537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4045 ( .C ( clk ), .D ( new_AGEMA_signal_15544 ), .Q ( new_AGEMA_signal_15545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4053 ( .C ( clk ), .D ( new_AGEMA_signal_15552 ), .Q ( new_AGEMA_signal_15553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4061 ( .C ( clk ), .D ( new_AGEMA_signal_15560 ), .Q ( new_AGEMA_signal_15561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4063 ( .C ( clk ), .D ( n1981 ), .Q ( new_AGEMA_signal_15563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4065 ( .C ( clk ), .D ( new_AGEMA_signal_2895 ), .Q ( new_AGEMA_signal_15565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4067 ( .C ( clk ), .D ( new_AGEMA_signal_2896 ), .Q ( new_AGEMA_signal_15567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4069 ( .C ( clk ), .D ( new_AGEMA_signal_2897 ), .Q ( new_AGEMA_signal_15569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4073 ( .C ( clk ), .D ( new_AGEMA_signal_15572 ), .Q ( new_AGEMA_signal_15573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4077 ( .C ( clk ), .D ( new_AGEMA_signal_15576 ), .Q ( new_AGEMA_signal_15577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4081 ( .C ( clk ), .D ( new_AGEMA_signal_15580 ), .Q ( new_AGEMA_signal_15581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4085 ( .C ( clk ), .D ( new_AGEMA_signal_15584 ), .Q ( new_AGEMA_signal_15585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4093 ( .C ( clk ), .D ( new_AGEMA_signal_15592 ), .Q ( new_AGEMA_signal_15593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4101 ( .C ( clk ), .D ( new_AGEMA_signal_15600 ), .Q ( new_AGEMA_signal_15601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4109 ( .C ( clk ), .D ( new_AGEMA_signal_15608 ), .Q ( new_AGEMA_signal_15609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4117 ( .C ( clk ), .D ( new_AGEMA_signal_15616 ), .Q ( new_AGEMA_signal_15617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4119 ( .C ( clk ), .D ( new_AGEMA_signal_14674 ), .Q ( new_AGEMA_signal_15619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4121 ( .C ( clk ), .D ( new_AGEMA_signal_14682 ), .Q ( new_AGEMA_signal_15621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4123 ( .C ( clk ), .D ( new_AGEMA_signal_14690 ), .Q ( new_AGEMA_signal_15623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4125 ( .C ( clk ), .D ( new_AGEMA_signal_14698 ), .Q ( new_AGEMA_signal_15625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4131 ( .C ( clk ), .D ( new_AGEMA_signal_15630 ), .Q ( new_AGEMA_signal_15631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4137 ( .C ( clk ), .D ( new_AGEMA_signal_15636 ), .Q ( new_AGEMA_signal_15637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4143 ( .C ( clk ), .D ( new_AGEMA_signal_15642 ), .Q ( new_AGEMA_signal_15643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4149 ( .C ( clk ), .D ( new_AGEMA_signal_15648 ), .Q ( new_AGEMA_signal_15649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4153 ( .C ( clk ), .D ( new_AGEMA_signal_15652 ), .Q ( new_AGEMA_signal_15653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4157 ( .C ( clk ), .D ( new_AGEMA_signal_15656 ), .Q ( new_AGEMA_signal_15657 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4161 ( .C ( clk ), .D ( new_AGEMA_signal_15660 ), .Q ( new_AGEMA_signal_15661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4165 ( .C ( clk ), .D ( new_AGEMA_signal_15664 ), .Q ( new_AGEMA_signal_15665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4173 ( .C ( clk ), .D ( new_AGEMA_signal_15672 ), .Q ( new_AGEMA_signal_15673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4181 ( .C ( clk ), .D ( new_AGEMA_signal_15680 ), .Q ( new_AGEMA_signal_15681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4189 ( .C ( clk ), .D ( new_AGEMA_signal_15688 ), .Q ( new_AGEMA_signal_15689 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4197 ( .C ( clk ), .D ( new_AGEMA_signal_15696 ), .Q ( new_AGEMA_signal_15697 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4201 ( .C ( clk ), .D ( new_AGEMA_signal_15700 ), .Q ( new_AGEMA_signal_15701 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4205 ( .C ( clk ), .D ( new_AGEMA_signal_15704 ), .Q ( new_AGEMA_signal_15705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4209 ( .C ( clk ), .D ( new_AGEMA_signal_15708 ), .Q ( new_AGEMA_signal_15709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4213 ( .C ( clk ), .D ( new_AGEMA_signal_15712 ), .Q ( new_AGEMA_signal_15713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4219 ( .C ( clk ), .D ( new_AGEMA_signal_15718 ), .Q ( new_AGEMA_signal_15719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4225 ( .C ( clk ), .D ( new_AGEMA_signal_15724 ), .Q ( new_AGEMA_signal_15725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4231 ( .C ( clk ), .D ( new_AGEMA_signal_15730 ), .Q ( new_AGEMA_signal_15731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4237 ( .C ( clk ), .D ( new_AGEMA_signal_15736 ), .Q ( new_AGEMA_signal_15737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4243 ( .C ( clk ), .D ( new_AGEMA_signal_15742 ), .Q ( new_AGEMA_signal_15743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4249 ( .C ( clk ), .D ( new_AGEMA_signal_15748 ), .Q ( new_AGEMA_signal_15749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4255 ( .C ( clk ), .D ( new_AGEMA_signal_15754 ), .Q ( new_AGEMA_signal_15755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4261 ( .C ( clk ), .D ( new_AGEMA_signal_15760 ), .Q ( new_AGEMA_signal_15761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4267 ( .C ( clk ), .D ( new_AGEMA_signal_15766 ), .Q ( new_AGEMA_signal_15767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4273 ( .C ( clk ), .D ( new_AGEMA_signal_15772 ), .Q ( new_AGEMA_signal_15773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4279 ( .C ( clk ), .D ( new_AGEMA_signal_15778 ), .Q ( new_AGEMA_signal_15779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4285 ( .C ( clk ), .D ( new_AGEMA_signal_15784 ), .Q ( new_AGEMA_signal_15785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4291 ( .C ( clk ), .D ( new_AGEMA_signal_15790 ), .Q ( new_AGEMA_signal_15791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4297 ( .C ( clk ), .D ( new_AGEMA_signal_15796 ), .Q ( new_AGEMA_signal_15797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4303 ( .C ( clk ), .D ( new_AGEMA_signal_15802 ), .Q ( new_AGEMA_signal_15803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4309 ( .C ( clk ), .D ( new_AGEMA_signal_15808 ), .Q ( new_AGEMA_signal_15809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4315 ( .C ( clk ), .D ( new_AGEMA_signal_15814 ), .Q ( new_AGEMA_signal_15815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4321 ( .C ( clk ), .D ( new_AGEMA_signal_15820 ), .Q ( new_AGEMA_signal_15821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4327 ( .C ( clk ), .D ( new_AGEMA_signal_15826 ), .Q ( new_AGEMA_signal_15827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4333 ( .C ( clk ), .D ( new_AGEMA_signal_15832 ), .Q ( new_AGEMA_signal_15833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4337 ( .C ( clk ), .D ( new_AGEMA_signal_15836 ), .Q ( new_AGEMA_signal_15837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4341 ( .C ( clk ), .D ( new_AGEMA_signal_15840 ), .Q ( new_AGEMA_signal_15841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4345 ( .C ( clk ), .D ( new_AGEMA_signal_15844 ), .Q ( new_AGEMA_signal_15845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4349 ( .C ( clk ), .D ( new_AGEMA_signal_15848 ), .Q ( new_AGEMA_signal_15849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4357 ( .C ( clk ), .D ( new_AGEMA_signal_15856 ), .Q ( new_AGEMA_signal_15857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4365 ( .C ( clk ), .D ( new_AGEMA_signal_15864 ), .Q ( new_AGEMA_signal_15865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4373 ( .C ( clk ), .D ( new_AGEMA_signal_15872 ), .Q ( new_AGEMA_signal_15873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4381 ( .C ( clk ), .D ( new_AGEMA_signal_15880 ), .Q ( new_AGEMA_signal_15881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4385 ( .C ( clk ), .D ( new_AGEMA_signal_15884 ), .Q ( new_AGEMA_signal_15885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4389 ( .C ( clk ), .D ( new_AGEMA_signal_15888 ), .Q ( new_AGEMA_signal_15889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4393 ( .C ( clk ), .D ( new_AGEMA_signal_15892 ), .Q ( new_AGEMA_signal_15893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4397 ( .C ( clk ), .D ( new_AGEMA_signal_15896 ), .Q ( new_AGEMA_signal_15897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4403 ( .C ( clk ), .D ( new_AGEMA_signal_15902 ), .Q ( new_AGEMA_signal_15903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4409 ( .C ( clk ), .D ( new_AGEMA_signal_15908 ), .Q ( new_AGEMA_signal_15909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4415 ( .C ( clk ), .D ( new_AGEMA_signal_15914 ), .Q ( new_AGEMA_signal_15915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4421 ( .C ( clk ), .D ( new_AGEMA_signal_15920 ), .Q ( new_AGEMA_signal_15921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4429 ( .C ( clk ), .D ( new_AGEMA_signal_15928 ), .Q ( new_AGEMA_signal_15929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4437 ( .C ( clk ), .D ( new_AGEMA_signal_15936 ), .Q ( new_AGEMA_signal_15937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4445 ( .C ( clk ), .D ( new_AGEMA_signal_15944 ), .Q ( new_AGEMA_signal_15945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4453 ( .C ( clk ), .D ( new_AGEMA_signal_15952 ), .Q ( new_AGEMA_signal_15953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4455 ( .C ( clk ), .D ( new_AGEMA_signal_15236 ), .Q ( new_AGEMA_signal_15955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4457 ( .C ( clk ), .D ( new_AGEMA_signal_15238 ), .Q ( new_AGEMA_signal_15957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4459 ( .C ( clk ), .D ( new_AGEMA_signal_15240 ), .Q ( new_AGEMA_signal_15959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4461 ( .C ( clk ), .D ( new_AGEMA_signal_15242 ), .Q ( new_AGEMA_signal_15961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4467 ( .C ( clk ), .D ( new_AGEMA_signal_15966 ), .Q ( new_AGEMA_signal_15967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4473 ( .C ( clk ), .D ( new_AGEMA_signal_15972 ), .Q ( new_AGEMA_signal_15973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4479 ( .C ( clk ), .D ( new_AGEMA_signal_15978 ), .Q ( new_AGEMA_signal_15979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4485 ( .C ( clk ), .D ( new_AGEMA_signal_15984 ), .Q ( new_AGEMA_signal_15985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4487 ( .C ( clk ), .D ( n2410 ), .Q ( new_AGEMA_signal_15987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4489 ( .C ( clk ), .D ( new_AGEMA_signal_3012 ), .Q ( new_AGEMA_signal_15989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4491 ( .C ( clk ), .D ( new_AGEMA_signal_3013 ), .Q ( new_AGEMA_signal_15991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4493 ( .C ( clk ), .D ( new_AGEMA_signal_3014 ), .Q ( new_AGEMA_signal_15993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4495 ( .C ( clk ), .D ( n2421 ), .Q ( new_AGEMA_signal_15995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4497 ( .C ( clk ), .D ( new_AGEMA_signal_3015 ), .Q ( new_AGEMA_signal_15997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4499 ( .C ( clk ), .D ( new_AGEMA_signal_3016 ), .Q ( new_AGEMA_signal_15999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4501 ( .C ( clk ), .D ( new_AGEMA_signal_3017 ), .Q ( new_AGEMA_signal_16001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4507 ( .C ( clk ), .D ( new_AGEMA_signal_16006 ), .Q ( new_AGEMA_signal_16007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4513 ( .C ( clk ), .D ( new_AGEMA_signal_16012 ), .Q ( new_AGEMA_signal_16013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4519 ( .C ( clk ), .D ( new_AGEMA_signal_16018 ), .Q ( new_AGEMA_signal_16019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4525 ( .C ( clk ), .D ( new_AGEMA_signal_16024 ), .Q ( new_AGEMA_signal_16025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4531 ( .C ( clk ), .D ( new_AGEMA_signal_16030 ), .Q ( new_AGEMA_signal_16031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4537 ( .C ( clk ), .D ( new_AGEMA_signal_16036 ), .Q ( new_AGEMA_signal_16037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4543 ( .C ( clk ), .D ( new_AGEMA_signal_16042 ), .Q ( new_AGEMA_signal_16043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4549 ( .C ( clk ), .D ( new_AGEMA_signal_16048 ), .Q ( new_AGEMA_signal_16049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4557 ( .C ( clk ), .D ( new_AGEMA_signal_16056 ), .Q ( new_AGEMA_signal_16057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4565 ( .C ( clk ), .D ( new_AGEMA_signal_16064 ), .Q ( new_AGEMA_signal_16065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4573 ( .C ( clk ), .D ( new_AGEMA_signal_16072 ), .Q ( new_AGEMA_signal_16073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4581 ( .C ( clk ), .D ( new_AGEMA_signal_16080 ), .Q ( new_AGEMA_signal_16081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4589 ( .C ( clk ), .D ( new_AGEMA_signal_16088 ), .Q ( new_AGEMA_signal_16089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4597 ( .C ( clk ), .D ( new_AGEMA_signal_16096 ), .Q ( new_AGEMA_signal_16097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4605 ( .C ( clk ), .D ( new_AGEMA_signal_16104 ), .Q ( new_AGEMA_signal_16105 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4613 ( .C ( clk ), .D ( new_AGEMA_signal_16112 ), .Q ( new_AGEMA_signal_16113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4619 ( .C ( clk ), .D ( new_AGEMA_signal_16118 ), .Q ( new_AGEMA_signal_16119 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4625 ( .C ( clk ), .D ( new_AGEMA_signal_16124 ), .Q ( new_AGEMA_signal_16125 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4631 ( .C ( clk ), .D ( new_AGEMA_signal_16130 ), .Q ( new_AGEMA_signal_16131 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4637 ( .C ( clk ), .D ( new_AGEMA_signal_16136 ), .Q ( new_AGEMA_signal_16137 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4643 ( .C ( clk ), .D ( new_AGEMA_signal_16142 ), .Q ( new_AGEMA_signal_16143 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4649 ( .C ( clk ), .D ( new_AGEMA_signal_16148 ), .Q ( new_AGEMA_signal_16149 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4655 ( .C ( clk ), .D ( new_AGEMA_signal_16154 ), .Q ( new_AGEMA_signal_16155 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4661 ( .C ( clk ), .D ( new_AGEMA_signal_16160 ), .Q ( new_AGEMA_signal_16161 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4663 ( .C ( clk ), .D ( new_AGEMA_signal_15198 ), .Q ( new_AGEMA_signal_16163 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4665 ( .C ( clk ), .D ( new_AGEMA_signal_15202 ), .Q ( new_AGEMA_signal_16165 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4667 ( .C ( clk ), .D ( new_AGEMA_signal_15206 ), .Q ( new_AGEMA_signal_16167 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4669 ( .C ( clk ), .D ( new_AGEMA_signal_15210 ), .Q ( new_AGEMA_signal_16169 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4673 ( .C ( clk ), .D ( new_AGEMA_signal_16172 ), .Q ( new_AGEMA_signal_16173 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4677 ( .C ( clk ), .D ( new_AGEMA_signal_16176 ), .Q ( new_AGEMA_signal_16177 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4681 ( .C ( clk ), .D ( new_AGEMA_signal_16180 ), .Q ( new_AGEMA_signal_16181 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4685 ( .C ( clk ), .D ( new_AGEMA_signal_16184 ), .Q ( new_AGEMA_signal_16185 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4689 ( .C ( clk ), .D ( new_AGEMA_signal_16188 ), .Q ( new_AGEMA_signal_16189 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4693 ( .C ( clk ), .D ( new_AGEMA_signal_16192 ), .Q ( new_AGEMA_signal_16193 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4697 ( .C ( clk ), .D ( new_AGEMA_signal_16196 ), .Q ( new_AGEMA_signal_16197 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4701 ( .C ( clk ), .D ( new_AGEMA_signal_16200 ), .Q ( new_AGEMA_signal_16201 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4705 ( .C ( clk ), .D ( new_AGEMA_signal_16204 ), .Q ( new_AGEMA_signal_16205 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4709 ( .C ( clk ), .D ( new_AGEMA_signal_16208 ), .Q ( new_AGEMA_signal_16209 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4713 ( .C ( clk ), .D ( new_AGEMA_signal_16212 ), .Q ( new_AGEMA_signal_16213 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4717 ( .C ( clk ), .D ( new_AGEMA_signal_16216 ), .Q ( new_AGEMA_signal_16217 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4719 ( .C ( clk ), .D ( new_AGEMA_signal_14978 ), .Q ( new_AGEMA_signal_16219 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4721 ( .C ( clk ), .D ( new_AGEMA_signal_14986 ), .Q ( new_AGEMA_signal_16221 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4723 ( .C ( clk ), .D ( new_AGEMA_signal_14994 ), .Q ( new_AGEMA_signal_16223 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4725 ( .C ( clk ), .D ( new_AGEMA_signal_15002 ), .Q ( new_AGEMA_signal_16225 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4729 ( .C ( clk ), .D ( new_AGEMA_signal_16228 ), .Q ( new_AGEMA_signal_16229 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4735 ( .C ( clk ), .D ( new_AGEMA_signal_16234 ), .Q ( new_AGEMA_signal_16235 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4741 ( .C ( clk ), .D ( new_AGEMA_signal_16240 ), .Q ( new_AGEMA_signal_16241 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4747 ( .C ( clk ), .D ( new_AGEMA_signal_16246 ), .Q ( new_AGEMA_signal_16247 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4759 ( .C ( clk ), .D ( n1984 ), .Q ( new_AGEMA_signal_16259 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4763 ( .C ( clk ), .D ( new_AGEMA_signal_3123 ), .Q ( new_AGEMA_signal_16263 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4767 ( .C ( clk ), .D ( new_AGEMA_signal_3124 ), .Q ( new_AGEMA_signal_16267 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4771 ( .C ( clk ), .D ( new_AGEMA_signal_3125 ), .Q ( new_AGEMA_signal_16271 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4779 ( .C ( clk ), .D ( new_AGEMA_signal_16278 ), .Q ( new_AGEMA_signal_16279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4787 ( .C ( clk ), .D ( new_AGEMA_signal_16286 ), .Q ( new_AGEMA_signal_16287 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4795 ( .C ( clk ), .D ( new_AGEMA_signal_16294 ), .Q ( new_AGEMA_signal_16295 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4803 ( .C ( clk ), .D ( new_AGEMA_signal_16302 ), .Q ( new_AGEMA_signal_16303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4811 ( .C ( clk ), .D ( new_AGEMA_signal_16310 ), .Q ( new_AGEMA_signal_16311 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4819 ( .C ( clk ), .D ( new_AGEMA_signal_16318 ), .Q ( new_AGEMA_signal_16319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4827 ( .C ( clk ), .D ( new_AGEMA_signal_16326 ), .Q ( new_AGEMA_signal_16327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4835 ( .C ( clk ), .D ( new_AGEMA_signal_16334 ), .Q ( new_AGEMA_signal_16335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4843 ( .C ( clk ), .D ( new_AGEMA_signal_16342 ), .Q ( new_AGEMA_signal_16343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4851 ( .C ( clk ), .D ( new_AGEMA_signal_16350 ), .Q ( new_AGEMA_signal_16351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4859 ( .C ( clk ), .D ( new_AGEMA_signal_16358 ), .Q ( new_AGEMA_signal_16359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4867 ( .C ( clk ), .D ( new_AGEMA_signal_16366 ), .Q ( new_AGEMA_signal_16367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4875 ( .C ( clk ), .D ( new_AGEMA_signal_16374 ), .Q ( new_AGEMA_signal_16375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4883 ( .C ( clk ), .D ( new_AGEMA_signal_16382 ), .Q ( new_AGEMA_signal_16383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4891 ( .C ( clk ), .D ( new_AGEMA_signal_16390 ), .Q ( new_AGEMA_signal_16391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4899 ( .C ( clk ), .D ( new_AGEMA_signal_16398 ), .Q ( new_AGEMA_signal_16399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4905 ( .C ( clk ), .D ( new_AGEMA_signal_16404 ), .Q ( new_AGEMA_signal_16405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4911 ( .C ( clk ), .D ( new_AGEMA_signal_16410 ), .Q ( new_AGEMA_signal_16411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4917 ( .C ( clk ), .D ( new_AGEMA_signal_16416 ), .Q ( new_AGEMA_signal_16417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4923 ( .C ( clk ), .D ( new_AGEMA_signal_16422 ), .Q ( new_AGEMA_signal_16423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4933 ( .C ( clk ), .D ( new_AGEMA_signal_16432 ), .Q ( new_AGEMA_signal_16433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4943 ( .C ( clk ), .D ( new_AGEMA_signal_16442 ), .Q ( new_AGEMA_signal_16443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4953 ( .C ( clk ), .D ( new_AGEMA_signal_16452 ), .Q ( new_AGEMA_signal_16453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4963 ( .C ( clk ), .D ( new_AGEMA_signal_16462 ), .Q ( new_AGEMA_signal_16463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4971 ( .C ( clk ), .D ( new_AGEMA_signal_16470 ), .Q ( new_AGEMA_signal_16471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4979 ( .C ( clk ), .D ( new_AGEMA_signal_16478 ), .Q ( new_AGEMA_signal_16479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4987 ( .C ( clk ), .D ( new_AGEMA_signal_16486 ), .Q ( new_AGEMA_signal_16487 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4995 ( .C ( clk ), .D ( new_AGEMA_signal_16494 ), .Q ( new_AGEMA_signal_16495 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5003 ( .C ( clk ), .D ( new_AGEMA_signal_16502 ), .Q ( new_AGEMA_signal_16503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5011 ( .C ( clk ), .D ( new_AGEMA_signal_16510 ), .Q ( new_AGEMA_signal_16511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5019 ( .C ( clk ), .D ( new_AGEMA_signal_16518 ), .Q ( new_AGEMA_signal_16519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5027 ( .C ( clk ), .D ( new_AGEMA_signal_16526 ), .Q ( new_AGEMA_signal_16527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5035 ( .C ( clk ), .D ( new_AGEMA_signal_16534 ), .Q ( new_AGEMA_signal_16535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5043 ( .C ( clk ), .D ( new_AGEMA_signal_16542 ), .Q ( new_AGEMA_signal_16543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5051 ( .C ( clk ), .D ( new_AGEMA_signal_16550 ), .Q ( new_AGEMA_signal_16551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5059 ( .C ( clk ), .D ( new_AGEMA_signal_16558 ), .Q ( new_AGEMA_signal_16559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5071 ( .C ( clk ), .D ( new_AGEMA_signal_15222 ), .Q ( new_AGEMA_signal_16571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5075 ( .C ( clk ), .D ( new_AGEMA_signal_15226 ), .Q ( new_AGEMA_signal_16575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5079 ( .C ( clk ), .D ( new_AGEMA_signal_15230 ), .Q ( new_AGEMA_signal_16579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5083 ( .C ( clk ), .D ( new_AGEMA_signal_15234 ), .Q ( new_AGEMA_signal_16583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5089 ( .C ( clk ), .D ( new_AGEMA_signal_16588 ), .Q ( new_AGEMA_signal_16589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5095 ( .C ( clk ), .D ( new_AGEMA_signal_16594 ), .Q ( new_AGEMA_signal_16595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5101 ( .C ( clk ), .D ( new_AGEMA_signal_16600 ), .Q ( new_AGEMA_signal_16601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5107 ( .C ( clk ), .D ( new_AGEMA_signal_16606 ), .Q ( new_AGEMA_signal_16607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5111 ( .C ( clk ), .D ( new_AGEMA_signal_14776 ), .Q ( new_AGEMA_signal_16611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5115 ( .C ( clk ), .D ( new_AGEMA_signal_14782 ), .Q ( new_AGEMA_signal_16615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5119 ( .C ( clk ), .D ( new_AGEMA_signal_14788 ), .Q ( new_AGEMA_signal_16619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5123 ( .C ( clk ), .D ( new_AGEMA_signal_14794 ), .Q ( new_AGEMA_signal_16623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5133 ( .C ( clk ), .D ( new_AGEMA_signal_16632 ), .Q ( new_AGEMA_signal_16633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5143 ( .C ( clk ), .D ( new_AGEMA_signal_16642 ), .Q ( new_AGEMA_signal_16643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5153 ( .C ( clk ), .D ( new_AGEMA_signal_16652 ), .Q ( new_AGEMA_signal_16653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5163 ( .C ( clk ), .D ( new_AGEMA_signal_16662 ), .Q ( new_AGEMA_signal_16663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5171 ( .C ( clk ), .D ( new_AGEMA_signal_16670 ), .Q ( new_AGEMA_signal_16671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5179 ( .C ( clk ), .D ( new_AGEMA_signal_16678 ), .Q ( new_AGEMA_signal_16679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5187 ( .C ( clk ), .D ( new_AGEMA_signal_16686 ), .Q ( new_AGEMA_signal_16687 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5195 ( .C ( clk ), .D ( new_AGEMA_signal_16694 ), .Q ( new_AGEMA_signal_16695 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5199 ( .C ( clk ), .D ( n2478 ), .Q ( new_AGEMA_signal_16699 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5203 ( .C ( clk ), .D ( new_AGEMA_signal_2775 ), .Q ( new_AGEMA_signal_16703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5207 ( .C ( clk ), .D ( new_AGEMA_signal_2776 ), .Q ( new_AGEMA_signal_16707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5211 ( .C ( clk ), .D ( new_AGEMA_signal_2777 ), .Q ( new_AGEMA_signal_16711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5227 ( .C ( clk ), .D ( new_AGEMA_signal_16726 ), .Q ( new_AGEMA_signal_16727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5235 ( .C ( clk ), .D ( new_AGEMA_signal_16734 ), .Q ( new_AGEMA_signal_16735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5243 ( .C ( clk ), .D ( new_AGEMA_signal_16742 ), .Q ( new_AGEMA_signal_16743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5251 ( .C ( clk ), .D ( new_AGEMA_signal_16750 ), .Q ( new_AGEMA_signal_16751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5259 ( .C ( clk ), .D ( new_AGEMA_signal_16758 ), .Q ( new_AGEMA_signal_16759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5267 ( .C ( clk ), .D ( new_AGEMA_signal_16766 ), .Q ( new_AGEMA_signal_16767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5275 ( .C ( clk ), .D ( new_AGEMA_signal_16774 ), .Q ( new_AGEMA_signal_16775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5283 ( .C ( clk ), .D ( new_AGEMA_signal_16782 ), .Q ( new_AGEMA_signal_16783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5289 ( .C ( clk ), .D ( new_AGEMA_signal_16788 ), .Q ( new_AGEMA_signal_16789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5295 ( .C ( clk ), .D ( new_AGEMA_signal_16794 ), .Q ( new_AGEMA_signal_16795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5301 ( .C ( clk ), .D ( new_AGEMA_signal_16800 ), .Q ( new_AGEMA_signal_16801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5307 ( .C ( clk ), .D ( new_AGEMA_signal_16806 ), .Q ( new_AGEMA_signal_16807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5311 ( .C ( clk ), .D ( n2660 ), .Q ( new_AGEMA_signal_16811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5315 ( .C ( clk ), .D ( new_AGEMA_signal_3075 ), .Q ( new_AGEMA_signal_16815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5319 ( .C ( clk ), .D ( new_AGEMA_signal_3076 ), .Q ( new_AGEMA_signal_16819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5323 ( .C ( clk ), .D ( new_AGEMA_signal_3077 ), .Q ( new_AGEMA_signal_16823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5331 ( .C ( clk ), .D ( new_AGEMA_signal_16830 ), .Q ( new_AGEMA_signal_16831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5339 ( .C ( clk ), .D ( new_AGEMA_signal_16838 ), .Q ( new_AGEMA_signal_16839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5347 ( .C ( clk ), .D ( new_AGEMA_signal_16846 ), .Q ( new_AGEMA_signal_16847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5355 ( .C ( clk ), .D ( new_AGEMA_signal_16854 ), .Q ( new_AGEMA_signal_16855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5367 ( .C ( clk ), .D ( n1940 ), .Q ( new_AGEMA_signal_16867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5373 ( .C ( clk ), .D ( new_AGEMA_signal_2877 ), .Q ( new_AGEMA_signal_16873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5379 ( .C ( clk ), .D ( new_AGEMA_signal_2878 ), .Q ( new_AGEMA_signal_16879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5385 ( .C ( clk ), .D ( new_AGEMA_signal_2879 ), .Q ( new_AGEMA_signal_16885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5391 ( .C ( clk ), .D ( n1961 ), .Q ( new_AGEMA_signal_16891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5397 ( .C ( clk ), .D ( new_AGEMA_signal_2880 ), .Q ( new_AGEMA_signal_16897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5403 ( .C ( clk ), .D ( new_AGEMA_signal_2881 ), .Q ( new_AGEMA_signal_16903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5409 ( .C ( clk ), .D ( new_AGEMA_signal_2882 ), .Q ( new_AGEMA_signal_16909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5415 ( .C ( clk ), .D ( n1987 ), .Q ( new_AGEMA_signal_16915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5421 ( .C ( clk ), .D ( new_AGEMA_signal_2571 ), .Q ( new_AGEMA_signal_16921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5427 ( .C ( clk ), .D ( new_AGEMA_signal_2572 ), .Q ( new_AGEMA_signal_16927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5433 ( .C ( clk ), .D ( new_AGEMA_signal_2573 ), .Q ( new_AGEMA_signal_16933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5457 ( .C ( clk ), .D ( new_AGEMA_signal_16956 ), .Q ( new_AGEMA_signal_16957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5465 ( .C ( clk ), .D ( new_AGEMA_signal_16964 ), .Q ( new_AGEMA_signal_16965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5473 ( .C ( clk ), .D ( new_AGEMA_signal_16972 ), .Q ( new_AGEMA_signal_16973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5481 ( .C ( clk ), .D ( new_AGEMA_signal_16980 ), .Q ( new_AGEMA_signal_16981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5487 ( .C ( clk ), .D ( n2054 ), .Q ( new_AGEMA_signal_16987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5493 ( .C ( clk ), .D ( new_AGEMA_signal_2910 ), .Q ( new_AGEMA_signal_16993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5499 ( .C ( clk ), .D ( new_AGEMA_signal_2911 ), .Q ( new_AGEMA_signal_16999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5505 ( .C ( clk ), .D ( new_AGEMA_signal_2912 ), .Q ( new_AGEMA_signal_17005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5529 ( .C ( clk ), .D ( new_AGEMA_signal_17028 ), .Q ( new_AGEMA_signal_17029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5537 ( .C ( clk ), .D ( new_AGEMA_signal_17036 ), .Q ( new_AGEMA_signal_17037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5545 ( .C ( clk ), .D ( new_AGEMA_signal_17044 ), .Q ( new_AGEMA_signal_17045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5553 ( .C ( clk ), .D ( new_AGEMA_signal_17052 ), .Q ( new_AGEMA_signal_17053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5561 ( .C ( clk ), .D ( new_AGEMA_signal_17060 ), .Q ( new_AGEMA_signal_17061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5569 ( .C ( clk ), .D ( new_AGEMA_signal_17068 ), .Q ( new_AGEMA_signal_17069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5577 ( .C ( clk ), .D ( new_AGEMA_signal_17076 ), .Q ( new_AGEMA_signal_17077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5585 ( .C ( clk ), .D ( new_AGEMA_signal_17084 ), .Q ( new_AGEMA_signal_17085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5595 ( .C ( clk ), .D ( new_AGEMA_signal_17094 ), .Q ( new_AGEMA_signal_17095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5605 ( .C ( clk ), .D ( new_AGEMA_signal_17104 ), .Q ( new_AGEMA_signal_17105 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5615 ( .C ( clk ), .D ( new_AGEMA_signal_17114 ), .Q ( new_AGEMA_signal_17115 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5625 ( .C ( clk ), .D ( new_AGEMA_signal_17124 ), .Q ( new_AGEMA_signal_17125 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5633 ( .C ( clk ), .D ( new_AGEMA_signal_17132 ), .Q ( new_AGEMA_signal_17133 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5641 ( .C ( clk ), .D ( new_AGEMA_signal_17140 ), .Q ( new_AGEMA_signal_17141 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5649 ( .C ( clk ), .D ( new_AGEMA_signal_17148 ), .Q ( new_AGEMA_signal_17149 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5657 ( .C ( clk ), .D ( new_AGEMA_signal_17156 ), .Q ( new_AGEMA_signal_17157 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5663 ( .C ( clk ), .D ( n2255 ), .Q ( new_AGEMA_signal_17163 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5669 ( .C ( clk ), .D ( new_AGEMA_signal_2970 ), .Q ( new_AGEMA_signal_17169 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5675 ( .C ( clk ), .D ( new_AGEMA_signal_2971 ), .Q ( new_AGEMA_signal_17175 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5681 ( .C ( clk ), .D ( new_AGEMA_signal_2972 ), .Q ( new_AGEMA_signal_17181 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5703 ( .C ( clk ), .D ( n2304 ), .Q ( new_AGEMA_signal_17203 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5709 ( .C ( clk ), .D ( new_AGEMA_signal_2982 ), .Q ( new_AGEMA_signal_17209 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5715 ( .C ( clk ), .D ( new_AGEMA_signal_2983 ), .Q ( new_AGEMA_signal_17215 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5721 ( .C ( clk ), .D ( new_AGEMA_signal_2984 ), .Q ( new_AGEMA_signal_17221 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5729 ( .C ( clk ), .D ( new_AGEMA_signal_17228 ), .Q ( new_AGEMA_signal_17229 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5737 ( .C ( clk ), .D ( new_AGEMA_signal_17236 ), .Q ( new_AGEMA_signal_17237 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5745 ( .C ( clk ), .D ( new_AGEMA_signal_17244 ), .Q ( new_AGEMA_signal_17245 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5753 ( .C ( clk ), .D ( new_AGEMA_signal_17252 ), .Q ( new_AGEMA_signal_17253 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5759 ( .C ( clk ), .D ( n2450 ), .Q ( new_AGEMA_signal_17259 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5765 ( .C ( clk ), .D ( new_AGEMA_signal_3024 ), .Q ( new_AGEMA_signal_17265 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5771 ( .C ( clk ), .D ( new_AGEMA_signal_3025 ), .Q ( new_AGEMA_signal_17271 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5777 ( .C ( clk ), .D ( new_AGEMA_signal_3026 ), .Q ( new_AGEMA_signal_17277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5793 ( .C ( clk ), .D ( new_AGEMA_signal_17292 ), .Q ( new_AGEMA_signal_17293 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5801 ( .C ( clk ), .D ( new_AGEMA_signal_17300 ), .Q ( new_AGEMA_signal_17301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5809 ( .C ( clk ), .D ( new_AGEMA_signal_17308 ), .Q ( new_AGEMA_signal_17309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5817 ( .C ( clk ), .D ( new_AGEMA_signal_17316 ), .Q ( new_AGEMA_signal_17317 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5839 ( .C ( clk ), .D ( n2666 ), .Q ( new_AGEMA_signal_17339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5845 ( .C ( clk ), .D ( new_AGEMA_signal_3081 ), .Q ( new_AGEMA_signal_17345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5851 ( .C ( clk ), .D ( new_AGEMA_signal_3082 ), .Q ( new_AGEMA_signal_17351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5857 ( .C ( clk ), .D ( new_AGEMA_signal_3083 ), .Q ( new_AGEMA_signal_17357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5863 ( .C ( clk ), .D ( n2704 ), .Q ( new_AGEMA_signal_17363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5869 ( .C ( clk ), .D ( new_AGEMA_signal_3087 ), .Q ( new_AGEMA_signal_17369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5875 ( .C ( clk ), .D ( new_AGEMA_signal_3088 ), .Q ( new_AGEMA_signal_17375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5881 ( .C ( clk ), .D ( new_AGEMA_signal_3089 ), .Q ( new_AGEMA_signal_17381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5969 ( .C ( clk ), .D ( new_AGEMA_signal_17468 ), .Q ( new_AGEMA_signal_17469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5979 ( .C ( clk ), .D ( new_AGEMA_signal_17478 ), .Q ( new_AGEMA_signal_17479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5989 ( .C ( clk ), .D ( new_AGEMA_signal_17488 ), .Q ( new_AGEMA_signal_17489 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5999 ( .C ( clk ), .D ( new_AGEMA_signal_17498 ), .Q ( new_AGEMA_signal_17499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6087 ( .C ( clk ), .D ( n2280 ), .Q ( new_AGEMA_signal_17587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6095 ( .C ( clk ), .D ( new_AGEMA_signal_2694 ), .Q ( new_AGEMA_signal_17595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6103 ( .C ( clk ), .D ( new_AGEMA_signal_2695 ), .Q ( new_AGEMA_signal_17603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6111 ( .C ( clk ), .D ( new_AGEMA_signal_2696 ), .Q ( new_AGEMA_signal_17611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6143 ( .C ( clk ), .D ( new_AGEMA_signal_14764 ), .Q ( new_AGEMA_signal_17643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6151 ( .C ( clk ), .D ( new_AGEMA_signal_14766 ), .Q ( new_AGEMA_signal_17651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6159 ( .C ( clk ), .D ( new_AGEMA_signal_14768 ), .Q ( new_AGEMA_signal_17659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6167 ( .C ( clk ), .D ( new_AGEMA_signal_14770 ), .Q ( new_AGEMA_signal_17667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6175 ( .C ( clk ), .D ( n2456 ), .Q ( new_AGEMA_signal_17675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6183 ( .C ( clk ), .D ( new_AGEMA_signal_3027 ), .Q ( new_AGEMA_signal_17683 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6191 ( .C ( clk ), .D ( new_AGEMA_signal_3028 ), .Q ( new_AGEMA_signal_17691 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6199 ( .C ( clk ), .D ( new_AGEMA_signal_3029 ), .Q ( new_AGEMA_signal_17699 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6247 ( .C ( clk ), .D ( n2706 ), .Q ( new_AGEMA_signal_17747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6255 ( .C ( clk ), .D ( new_AGEMA_signal_3084 ), .Q ( new_AGEMA_signal_17755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6263 ( .C ( clk ), .D ( new_AGEMA_signal_3085 ), .Q ( new_AGEMA_signal_17763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6271 ( .C ( clk ), .D ( new_AGEMA_signal_3086 ), .Q ( new_AGEMA_signal_17771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6329 ( .C ( clk ), .D ( new_AGEMA_signal_17828 ), .Q ( new_AGEMA_signal_17829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6341 ( .C ( clk ), .D ( new_AGEMA_signal_17840 ), .Q ( new_AGEMA_signal_17841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6353 ( .C ( clk ), .D ( new_AGEMA_signal_17852 ), .Q ( new_AGEMA_signal_17853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6365 ( .C ( clk ), .D ( new_AGEMA_signal_17864 ), .Q ( new_AGEMA_signal_17865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6379 ( .C ( clk ), .D ( new_AGEMA_signal_17878 ), .Q ( new_AGEMA_signal_17879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6393 ( .C ( clk ), .D ( new_AGEMA_signal_17892 ), .Q ( new_AGEMA_signal_17893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6407 ( .C ( clk ), .D ( new_AGEMA_signal_17906 ), .Q ( new_AGEMA_signal_17907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6421 ( .C ( clk ), .D ( new_AGEMA_signal_17920 ), .Q ( new_AGEMA_signal_17921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6467 ( .C ( clk ), .D ( new_AGEMA_signal_17966 ), .Q ( new_AGEMA_signal_17967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6481 ( .C ( clk ), .D ( new_AGEMA_signal_17980 ), .Q ( new_AGEMA_signal_17981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6495 ( .C ( clk ), .D ( new_AGEMA_signal_17994 ), .Q ( new_AGEMA_signal_17995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6509 ( .C ( clk ), .D ( new_AGEMA_signal_18008 ), .Q ( new_AGEMA_signal_18009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6611 ( .C ( clk ), .D ( new_AGEMA_signal_18110 ), .Q ( new_AGEMA_signal_18111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6627 ( .C ( clk ), .D ( new_AGEMA_signal_18126 ), .Q ( new_AGEMA_signal_18127 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6643 ( .C ( clk ), .D ( new_AGEMA_signal_18142 ), .Q ( new_AGEMA_signal_18143 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6659 ( .C ( clk ), .D ( new_AGEMA_signal_18158 ), .Q ( new_AGEMA_signal_18159 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6699 ( .C ( clk ), .D ( new_AGEMA_signal_18198 ), .Q ( new_AGEMA_signal_18199 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6715 ( .C ( clk ), .D ( new_AGEMA_signal_18214 ), .Q ( new_AGEMA_signal_18215 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6731 ( .C ( clk ), .D ( new_AGEMA_signal_18230 ), .Q ( new_AGEMA_signal_18231 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6747 ( .C ( clk ), .D ( new_AGEMA_signal_18246 ), .Q ( new_AGEMA_signal_18247 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6897 ( .C ( clk ), .D ( new_AGEMA_signal_18396 ), .Q ( new_AGEMA_signal_18397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6913 ( .C ( clk ), .D ( new_AGEMA_signal_18412 ), .Q ( new_AGEMA_signal_18413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6929 ( .C ( clk ), .D ( new_AGEMA_signal_18428 ), .Q ( new_AGEMA_signal_18429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6945 ( .C ( clk ), .D ( new_AGEMA_signal_18444 ), .Q ( new_AGEMA_signal_18445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7003 ( .C ( clk ), .D ( new_AGEMA_signal_18502 ), .Q ( new_AGEMA_signal_18503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7021 ( .C ( clk ), .D ( new_AGEMA_signal_18520 ), .Q ( new_AGEMA_signal_18521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7039 ( .C ( clk ), .D ( new_AGEMA_signal_18538 ), .Q ( new_AGEMA_signal_18539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7057 ( .C ( clk ), .D ( new_AGEMA_signal_18556 ), .Q ( new_AGEMA_signal_18557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7203 ( .C ( clk ), .D ( new_AGEMA_signal_18702 ), .Q ( new_AGEMA_signal_18703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7223 ( .C ( clk ), .D ( new_AGEMA_signal_18722 ), .Q ( new_AGEMA_signal_18723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7243 ( .C ( clk ), .D ( new_AGEMA_signal_18742 ), .Q ( new_AGEMA_signal_18743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7263 ( .C ( clk ), .D ( new_AGEMA_signal_18762 ), .Q ( new_AGEMA_signal_18763 ) ) ;

    /* cells in depth 12 */
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2001 ( .ina ({new_AGEMA_signal_2876, new_AGEMA_signal_2875, new_AGEMA_signal_2874, n1932}), .inb ({new_AGEMA_signal_14610, new_AGEMA_signal_14606, new_AGEMA_signal_14602, new_AGEMA_signal_14598}), .clk ( clk ), .rnd ({Fresh[6609], Fresh[6608], Fresh[6607], Fresh[6606], Fresh[6605], Fresh[6604], Fresh[6603], Fresh[6602], Fresh[6601], Fresh[6600]}), .outt ({new_AGEMA_signal_3119, new_AGEMA_signal_3118, new_AGEMA_signal_3117, n1933}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2051 ( .ina ({new_AGEMA_signal_14626, new_AGEMA_signal_14622, new_AGEMA_signal_14618, new_AGEMA_signal_14614}), .inb ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, new_AGEMA_signal_2883, n1955}), .clk ( clk ), .rnd ({Fresh[6619], Fresh[6618], Fresh[6617], Fresh[6616], Fresh[6615], Fresh[6614], Fresh[6613], Fresh[6612], Fresh[6611], Fresh[6610]}), .outt ({new_AGEMA_signal_3122, new_AGEMA_signal_3121, new_AGEMA_signal_3120, n1958}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2067 ( .ina ({new_AGEMA_signal_2555, new_AGEMA_signal_2554, new_AGEMA_signal_2553, n1967}), .inb ({new_AGEMA_signal_14658, new_AGEMA_signal_14650, new_AGEMA_signal_14642, new_AGEMA_signal_14634}), .clk ( clk ), .rnd ({Fresh[6629], Fresh[6628], Fresh[6627], Fresh[6626], Fresh[6625], Fresh[6624], Fresh[6623], Fresh[6622], Fresh[6621], Fresh[6620]}), .outt ({new_AGEMA_signal_2888, new_AGEMA_signal_2887, new_AGEMA_signal_2886, n1990}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2104 ( .ina ({new_AGEMA_signal_14666, new_AGEMA_signal_14664, new_AGEMA_signal_14662, new_AGEMA_signal_14660}), .inb ({new_AGEMA_signal_2894, new_AGEMA_signal_2893, new_AGEMA_signal_2892, n1977}), .clk ( clk ), .rnd ({Fresh[6639], Fresh[6638], Fresh[6637], Fresh[6636], Fresh[6635], Fresh[6634], Fresh[6633], Fresh[6632], Fresh[6631], Fresh[6630]}), .outt ({new_AGEMA_signal_3128, new_AGEMA_signal_3127, new_AGEMA_signal_3126, n1982}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2128 ( .ina ({new_AGEMA_signal_14698, new_AGEMA_signal_14690, new_AGEMA_signal_14682, new_AGEMA_signal_14674}), .inb ({new_AGEMA_signal_2900, new_AGEMA_signal_2899, new_AGEMA_signal_2898, n1998}), .clk ( clk ), .rnd ({Fresh[6649], Fresh[6648], Fresh[6647], Fresh[6646], Fresh[6645], Fresh[6644], Fresh[6643], Fresh[6642], Fresh[6641], Fresh[6640]}), .outt ({new_AGEMA_signal_3131, new_AGEMA_signal_3130, new_AGEMA_signal_3129, n1999}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2148 ( .ina ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, new_AGEMA_signal_2901, n2010}), .inb ({new_AGEMA_signal_14722, new_AGEMA_signal_14716, new_AGEMA_signal_14710, new_AGEMA_signal_14704}), .clk ( clk ), .rnd ({Fresh[6659], Fresh[6658], Fresh[6657], Fresh[6656], Fresh[6655], Fresh[6654], Fresh[6653], Fresh[6652], Fresh[6651], Fresh[6650]}), .outt ({new_AGEMA_signal_3134, new_AGEMA_signal_3133, new_AGEMA_signal_3132, n2011}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2165 ( .ina ({new_AGEMA_signal_2585, new_AGEMA_signal_2584, new_AGEMA_signal_2583, n2024}), .inb ({new_AGEMA_signal_14738, new_AGEMA_signal_14734, new_AGEMA_signal_14730, new_AGEMA_signal_14726}), .clk ( clk ), .rnd ({Fresh[6669], Fresh[6668], Fresh[6667], Fresh[6666], Fresh[6665], Fresh[6664], Fresh[6663], Fresh[6662], Fresh[6661], Fresh[6660]}), .outt ({new_AGEMA_signal_2906, new_AGEMA_signal_2905, new_AGEMA_signal_2904, n2025}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2179 ( .ina ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, new_AGEMA_signal_2907, n2035}), .inb ({new_AGEMA_signal_14762, new_AGEMA_signal_14756, new_AGEMA_signal_14750, new_AGEMA_signal_14744}), .clk ( clk ), .rnd ({Fresh[6679], Fresh[6678], Fresh[6677], Fresh[6676], Fresh[6675], Fresh[6674], Fresh[6673], Fresh[6672], Fresh[6671], Fresh[6670]}), .outt ({new_AGEMA_signal_3140, new_AGEMA_signal_3139, new_AGEMA_signal_3138, n2036}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2196 ( .ina ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, new_AGEMA_signal_2913, n2048}), .inb ({new_AGEMA_signal_2918, new_AGEMA_signal_2917, new_AGEMA_signal_2916, n2047}), .clk ( clk ), .rnd ({Fresh[6689], Fresh[6688], Fresh[6687], Fresh[6686], Fresh[6685], Fresh[6684], Fresh[6683], Fresh[6682], Fresh[6681], Fresh[6680]}), .outt ({new_AGEMA_signal_3143, new_AGEMA_signal_3142, new_AGEMA_signal_3141, n2049}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2207 ( .ina ({new_AGEMA_signal_14770, new_AGEMA_signal_14768, new_AGEMA_signal_14766, new_AGEMA_signal_14764}), .inb ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, new_AGEMA_signal_2919, n2059}), .clk ( clk ), .rnd ({Fresh[6699], Fresh[6698], Fresh[6697], Fresh[6696], Fresh[6695], Fresh[6694], Fresh[6693], Fresh[6692], Fresh[6691], Fresh[6690]}), .outt ({new_AGEMA_signal_3146, new_AGEMA_signal_3145, new_AGEMA_signal_3144, n2072}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2214 ( .ina ({new_AGEMA_signal_14794, new_AGEMA_signal_14788, new_AGEMA_signal_14782, new_AGEMA_signal_14776}), .inb ({new_AGEMA_signal_2924, new_AGEMA_signal_2923, new_AGEMA_signal_2922, n2064}), .clk ( clk ), .rnd ({Fresh[6709], Fresh[6708], Fresh[6707], Fresh[6706], Fresh[6705], Fresh[6704], Fresh[6703], Fresh[6702], Fresh[6701], Fresh[6700]}), .outt ({new_AGEMA_signal_3149, new_AGEMA_signal_3148, new_AGEMA_signal_3147, n2067}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2230 ( .ina ({new_AGEMA_signal_14818, new_AGEMA_signal_14812, new_AGEMA_signal_14806, new_AGEMA_signal_14800}), .inb ({new_AGEMA_signal_2927, new_AGEMA_signal_2926, new_AGEMA_signal_2925, n2077}), .clk ( clk ), .rnd ({Fresh[6719], Fresh[6718], Fresh[6717], Fresh[6716], Fresh[6715], Fresh[6714], Fresh[6713], Fresh[6712], Fresh[6711], Fresh[6710]}), .outt ({new_AGEMA_signal_3152, new_AGEMA_signal_3151, new_AGEMA_signal_3150, n2078}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2250 ( .ina ({new_AGEMA_signal_14826, new_AGEMA_signal_14824, new_AGEMA_signal_14822, new_AGEMA_signal_14820}), .inb ({new_AGEMA_signal_2930, new_AGEMA_signal_2929, new_AGEMA_signal_2928, n2158}), .clk ( clk ), .rnd ({Fresh[6729], Fresh[6728], Fresh[6727], Fresh[6726], Fresh[6725], Fresh[6724], Fresh[6723], Fresh[6722], Fresh[6721], Fresh[6720]}), .outt ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, new_AGEMA_signal_3153, n2097}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2257 ( .ina ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, new_AGEMA_signal_2931, n2095}), .inb ({new_AGEMA_signal_14842, new_AGEMA_signal_14838, new_AGEMA_signal_14834, new_AGEMA_signal_14830}), .clk ( clk ), .rnd ({Fresh[6739], Fresh[6738], Fresh[6737], Fresh[6736], Fresh[6735], Fresh[6734], Fresh[6733], Fresh[6732], Fresh[6731], Fresh[6730]}), .outt ({new_AGEMA_signal_3158, new_AGEMA_signal_3157, new_AGEMA_signal_3156, n2096}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2275 ( .ina ({new_AGEMA_signal_14866, new_AGEMA_signal_14860, new_AGEMA_signal_14854, new_AGEMA_signal_14848}), .inb ({new_AGEMA_signal_3161, new_AGEMA_signal_3160, new_AGEMA_signal_3159, n2117}), .clk ( clk ), .rnd ({Fresh[6749], Fresh[6748], Fresh[6747], Fresh[6746], Fresh[6745], Fresh[6744], Fresh[6743], Fresh[6742], Fresh[6741], Fresh[6740]}), .outt ({new_AGEMA_signal_3323, new_AGEMA_signal_3322, new_AGEMA_signal_3321, n2128}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2285 ( .ina ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, new_AGEMA_signal_2937, n2123}), .inb ({new_AGEMA_signal_14890, new_AGEMA_signal_14884, new_AGEMA_signal_14878, new_AGEMA_signal_14872}), .clk ( clk ), .rnd ({Fresh[6759], Fresh[6758], Fresh[6757], Fresh[6756], Fresh[6755], Fresh[6754], Fresh[6753], Fresh[6752], Fresh[6751], Fresh[6750]}), .outt ({new_AGEMA_signal_3164, new_AGEMA_signal_3163, new_AGEMA_signal_3162, n2124}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2301 ( .ina ({new_AGEMA_signal_14898, new_AGEMA_signal_14896, new_AGEMA_signal_14894, new_AGEMA_signal_14892}), .inb ({new_AGEMA_signal_2639, new_AGEMA_signal_2638, new_AGEMA_signal_2637, n2135}), .clk ( clk ), .rnd ({Fresh[6769], Fresh[6768], Fresh[6767], Fresh[6766], Fresh[6765], Fresh[6764], Fresh[6763], Fresh[6762], Fresh[6761], Fresh[6760]}), .outt ({new_AGEMA_signal_2942, new_AGEMA_signal_2941, new_AGEMA_signal_2940, n2148}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2310 ( .ina ({new_AGEMA_signal_14922, new_AGEMA_signal_14916, new_AGEMA_signal_14910, new_AGEMA_signal_14904}), .inb ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, new_AGEMA_signal_2943, n2141}), .clk ( clk ), .rnd ({Fresh[6779], Fresh[6778], Fresh[6777], Fresh[6776], Fresh[6775], Fresh[6774], Fresh[6773], Fresh[6772], Fresh[6771], Fresh[6770]}), .outt ({new_AGEMA_signal_3167, new_AGEMA_signal_3166, new_AGEMA_signal_3165, n2142}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2325 ( .ina ({new_AGEMA_signal_14930, new_AGEMA_signal_14928, new_AGEMA_signal_14926, new_AGEMA_signal_14924}), .inb ({new_AGEMA_signal_2930, new_AGEMA_signal_2929, new_AGEMA_signal_2928, n2158}), .clk ( clk ), .rnd ({Fresh[6789], Fresh[6788], Fresh[6787], Fresh[6786], Fresh[6785], Fresh[6784], Fresh[6783], Fresh[6782], Fresh[6781], Fresh[6780]}), .outt ({new_AGEMA_signal_3170, new_AGEMA_signal_3169, new_AGEMA_signal_3168, n2168}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2332 ( .ina ({new_AGEMA_signal_2948, new_AGEMA_signal_2947, new_AGEMA_signal_2946, n2166}), .inb ({new_AGEMA_signal_2654, new_AGEMA_signal_2653, new_AGEMA_signal_2652, n2165}), .clk ( clk ), .rnd ({Fresh[6799], Fresh[6798], Fresh[6797], Fresh[6796], Fresh[6795], Fresh[6794], Fresh[6793], Fresh[6792], Fresh[6791], Fresh[6790]}), .outt ({new_AGEMA_signal_3173, new_AGEMA_signal_3172, new_AGEMA_signal_3171, n2167}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2347 ( .ina ({new_AGEMA_signal_14946, new_AGEMA_signal_14942, new_AGEMA_signal_14938, new_AGEMA_signal_14934}), .inb ({new_AGEMA_signal_2951, new_AGEMA_signal_2950, new_AGEMA_signal_2949, n2180}), .clk ( clk ), .rnd ({Fresh[6809], Fresh[6808], Fresh[6807], Fresh[6806], Fresh[6805], Fresh[6804], Fresh[6803], Fresh[6802], Fresh[6801], Fresh[6800]}), .outt ({new_AGEMA_signal_3176, new_AGEMA_signal_3175, new_AGEMA_signal_3174, n2184}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2361 ( .ina ({new_AGEMA_signal_14962, new_AGEMA_signal_14958, new_AGEMA_signal_14954, new_AGEMA_signal_14950}), .inb ({new_AGEMA_signal_2954, new_AGEMA_signal_2953, new_AGEMA_signal_2952, n2194}), .clk ( clk ), .rnd ({Fresh[6819], Fresh[6818], Fresh[6817], Fresh[6816], Fresh[6815], Fresh[6814], Fresh[6813], Fresh[6812], Fresh[6811], Fresh[6810]}), .outt ({new_AGEMA_signal_3179, new_AGEMA_signal_3178, new_AGEMA_signal_3177, n2197}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2373 ( .ina ({new_AGEMA_signal_14970, new_AGEMA_signal_14968, new_AGEMA_signal_14966, new_AGEMA_signal_14964}), .inb ({new_AGEMA_signal_3182, new_AGEMA_signal_3181, new_AGEMA_signal_3180, n2204}), .clk ( clk ), .rnd ({Fresh[6829], Fresh[6828], Fresh[6827], Fresh[6826], Fresh[6825], Fresh[6824], Fresh[6823], Fresh[6822], Fresh[6821], Fresh[6820]}), .outt ({new_AGEMA_signal_3341, new_AGEMA_signal_3340, new_AGEMA_signal_3339, n2205}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2390 ( .ina ({new_AGEMA_signal_15002, new_AGEMA_signal_14994, new_AGEMA_signal_14986, new_AGEMA_signal_14978}), .inb ({new_AGEMA_signal_2960, new_AGEMA_signal_2959, new_AGEMA_signal_2958, n2225}), .clk ( clk ), .rnd ({Fresh[6839], Fresh[6838], Fresh[6837], Fresh[6836], Fresh[6835], Fresh[6834], Fresh[6833], Fresh[6832], Fresh[6831], Fresh[6830]}), .outt ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, new_AGEMA_signal_3183, n2232}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2395 ( .ina ({new_AGEMA_signal_2675, new_AGEMA_signal_2674, new_AGEMA_signal_2673, n2230}), .inb ({new_AGEMA_signal_15026, new_AGEMA_signal_15020, new_AGEMA_signal_15014, new_AGEMA_signal_15008}), .clk ( clk ), .rnd ({Fresh[6849], Fresh[6848], Fresh[6847], Fresh[6846], Fresh[6845], Fresh[6844], Fresh[6843], Fresh[6842], Fresh[6841], Fresh[6840]}), .outt ({new_AGEMA_signal_2963, new_AGEMA_signal_2962, new_AGEMA_signal_2961, n2231}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2401 ( .ina ({new_AGEMA_signal_15042, new_AGEMA_signal_15038, new_AGEMA_signal_15034, new_AGEMA_signal_15030}), .inb ({new_AGEMA_signal_3188, new_AGEMA_signal_3187, new_AGEMA_signal_3186, n2236}), .clk ( clk ), .rnd ({Fresh[6859], Fresh[6858], Fresh[6857], Fresh[6856], Fresh[6855], Fresh[6854], Fresh[6853], Fresh[6852], Fresh[6851], Fresh[6850]}), .outt ({new_AGEMA_signal_3347, new_AGEMA_signal_3346, new_AGEMA_signal_3345, n2239}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2413 ( .ina ({new_AGEMA_signal_15058, new_AGEMA_signal_15054, new_AGEMA_signal_15050, new_AGEMA_signal_15046}), .inb ({new_AGEMA_signal_2969, new_AGEMA_signal_2968, new_AGEMA_signal_2967, n2247}), .clk ( clk ), .rnd ({Fresh[6869], Fresh[6868], Fresh[6867], Fresh[6866], Fresh[6865], Fresh[6864], Fresh[6863], Fresh[6862], Fresh[6861], Fresh[6860]}), .outt ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, new_AGEMA_signal_3189, n2250}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2428 ( .ina ({new_AGEMA_signal_14770, new_AGEMA_signal_14768, new_AGEMA_signal_14766, new_AGEMA_signal_14764}), .inb ({new_AGEMA_signal_2975, new_AGEMA_signal_2974, new_AGEMA_signal_2973, n2264}), .clk ( clk ), .rnd ({Fresh[6879], Fresh[6878], Fresh[6877], Fresh[6876], Fresh[6875], Fresh[6874], Fresh[6873], Fresh[6872], Fresh[6871], Fresh[6870]}), .outt ({new_AGEMA_signal_3194, new_AGEMA_signal_3193, new_AGEMA_signal_3192, n2276}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2439 ( .ina ({new_AGEMA_signal_2978, new_AGEMA_signal_2977, new_AGEMA_signal_2976, n2271}), .inb ({new_AGEMA_signal_15066, new_AGEMA_signal_15064, new_AGEMA_signal_15062, new_AGEMA_signal_15060}), .clk ( clk ), .rnd ({Fresh[6889], Fresh[6888], Fresh[6887], Fresh[6886], Fresh[6885], Fresh[6884], Fresh[6883], Fresh[6882], Fresh[6881], Fresh[6880]}), .outt ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, new_AGEMA_signal_3195, n2272}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2454 ( .ina ({new_AGEMA_signal_2699, new_AGEMA_signal_2698, new_AGEMA_signal_2697, n2286}), .inb ({new_AGEMA_signal_15074, new_AGEMA_signal_15072, new_AGEMA_signal_15070, new_AGEMA_signal_15068}), .clk ( clk ), .rnd ({Fresh[6899], Fresh[6898], Fresh[6897], Fresh[6896], Fresh[6895], Fresh[6894], Fresh[6893], Fresh[6892], Fresh[6891], Fresh[6890]}), .outt ({new_AGEMA_signal_2981, new_AGEMA_signal_2980, new_AGEMA_signal_2979, n2306}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2468 ( .ina ({new_AGEMA_signal_2987, new_AGEMA_signal_2986, new_AGEMA_signal_2985, n2295}), .inb ({new_AGEMA_signal_15090, new_AGEMA_signal_15086, new_AGEMA_signal_15082, new_AGEMA_signal_15078}), .clk ( clk ), .rnd ({Fresh[6909], Fresh[6908], Fresh[6907], Fresh[6906], Fresh[6905], Fresh[6904], Fresh[6903], Fresh[6902], Fresh[6901], Fresh[6900]}), .outt ({new_AGEMA_signal_3200, new_AGEMA_signal_3199, new_AGEMA_signal_3198, n2296}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2489 ( .ina ({new_AGEMA_signal_15106, new_AGEMA_signal_15102, new_AGEMA_signal_15098, new_AGEMA_signal_15094}), .inb ({new_AGEMA_signal_2990, new_AGEMA_signal_2989, new_AGEMA_signal_2988, n2322}), .clk ( clk ), .rnd ({Fresh[6919], Fresh[6918], Fresh[6917], Fresh[6916], Fresh[6915], Fresh[6914], Fresh[6913], Fresh[6912], Fresh[6911], Fresh[6910]}), .outt ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, new_AGEMA_signal_3201, n2324}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2500 ( .ina ({new_AGEMA_signal_15114, new_AGEMA_signal_15112, new_AGEMA_signal_15110, new_AGEMA_signal_15108}), .inb ({new_AGEMA_signal_2993, new_AGEMA_signal_2992, new_AGEMA_signal_2991, n2333}), .clk ( clk ), .rnd ({Fresh[6929], Fresh[6928], Fresh[6927], Fresh[6926], Fresh[6925], Fresh[6924], Fresh[6923], Fresh[6922], Fresh[6921], Fresh[6920]}), .outt ({new_AGEMA_signal_3206, new_AGEMA_signal_3205, new_AGEMA_signal_3204, n2337}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2511 ( .ina ({new_AGEMA_signal_2999, new_AGEMA_signal_2998, new_AGEMA_signal_2997, n2345}), .inb ({new_AGEMA_signal_15138, new_AGEMA_signal_15132, new_AGEMA_signal_15126, new_AGEMA_signal_15120}), .clk ( clk ), .rnd ({Fresh[6939], Fresh[6938], Fresh[6937], Fresh[6936], Fresh[6935], Fresh[6934], Fresh[6933], Fresh[6932], Fresh[6931], Fresh[6930]}), .outt ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, new_AGEMA_signal_3207, n2350}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2528 ( .ina ({new_AGEMA_signal_3002, new_AGEMA_signal_3001, new_AGEMA_signal_3000, n2361}), .inb ({new_AGEMA_signal_15154, new_AGEMA_signal_15150, new_AGEMA_signal_15146, new_AGEMA_signal_15142}), .clk ( clk ), .rnd ({Fresh[6949], Fresh[6948], Fresh[6947], Fresh[6946], Fresh[6945], Fresh[6944], Fresh[6943], Fresh[6942], Fresh[6941], Fresh[6940]}), .outt ({new_AGEMA_signal_3212, new_AGEMA_signal_3211, new_AGEMA_signal_3210, n2362}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2550 ( .ina ({new_AGEMA_signal_15162, new_AGEMA_signal_15160, new_AGEMA_signal_15158, new_AGEMA_signal_15156}), .inb ({new_AGEMA_signal_2741, new_AGEMA_signal_2740, new_AGEMA_signal_2739, n2388}), .clk ( clk ), .rnd ({Fresh[6959], Fresh[6958], Fresh[6957], Fresh[6956], Fresh[6955], Fresh[6954], Fresh[6953], Fresh[6952], Fresh[6951], Fresh[6950]}), .outt ({new_AGEMA_signal_3005, new_AGEMA_signal_3004, new_AGEMA_signal_3003, n2389}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2557 ( .ina ({new_AGEMA_signal_15178, new_AGEMA_signal_15174, new_AGEMA_signal_15170, new_AGEMA_signal_15166}), .inb ({new_AGEMA_signal_3008, new_AGEMA_signal_3007, new_AGEMA_signal_3006, n2393}), .clk ( clk ), .rnd ({Fresh[6969], Fresh[6968], Fresh[6967], Fresh[6966], Fresh[6965], Fresh[6964], Fresh[6963], Fresh[6962], Fresh[6961], Fresh[6960]}), .outt ({new_AGEMA_signal_3218, new_AGEMA_signal_3217, new_AGEMA_signal_3216, n2397}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2568 ( .ina ({new_AGEMA_signal_15194, new_AGEMA_signal_15190, new_AGEMA_signal_15186, new_AGEMA_signal_15182}), .inb ({new_AGEMA_signal_2747, new_AGEMA_signal_2746, new_AGEMA_signal_2745, n2405}), .clk ( clk ), .rnd ({Fresh[6979], Fresh[6978], Fresh[6977], Fresh[6976], Fresh[6975], Fresh[6974], Fresh[6973], Fresh[6972], Fresh[6971], Fresh[6970]}), .outt ({new_AGEMA_signal_3011, new_AGEMA_signal_3010, new_AGEMA_signal_3009, n2411}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2580 ( .ina ({new_AGEMA_signal_15210, new_AGEMA_signal_15206, new_AGEMA_signal_15202, new_AGEMA_signal_15198}), .inb ({new_AGEMA_signal_2756, new_AGEMA_signal_2755, new_AGEMA_signal_2754, n2419}), .clk ( clk ), .rnd ({Fresh[6989], Fresh[6988], Fresh[6987], Fresh[6986], Fresh[6985], Fresh[6984], Fresh[6983], Fresh[6982], Fresh[6981], Fresh[6980]}), .outt ({new_AGEMA_signal_3020, new_AGEMA_signal_3019, new_AGEMA_signal_3018, n2420}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2593 ( .ina ({new_AGEMA_signal_3023, new_AGEMA_signal_3022, new_AGEMA_signal_3021, n2436}), .inb ({new_AGEMA_signal_15218, new_AGEMA_signal_15216, new_AGEMA_signal_15214, new_AGEMA_signal_15212}), .clk ( clk ), .rnd ({Fresh[6999], Fresh[6998], Fresh[6997], Fresh[6996], Fresh[6995], Fresh[6994], Fresh[6993], Fresh[6992], Fresh[6991], Fresh[6990]}), .outt ({new_AGEMA_signal_3227, new_AGEMA_signal_3226, new_AGEMA_signal_3225, n2440}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2614 ( .ina ({new_AGEMA_signal_15234, new_AGEMA_signal_15230, new_AGEMA_signal_15226, new_AGEMA_signal_15222}), .inb ({new_AGEMA_signal_3032, new_AGEMA_signal_3031, new_AGEMA_signal_3030, n2461}), .clk ( clk ), .rnd ({Fresh[7009], Fresh[7008], Fresh[7007], Fresh[7006], Fresh[7005], Fresh[7004], Fresh[7003], Fresh[7002], Fresh[7001], Fresh[7000]}), .outt ({new_AGEMA_signal_3230, new_AGEMA_signal_3229, new_AGEMA_signal_3228, n2516}) ) ;
    mux2_HPC1 #(.security_order(3), .pipeline(1)) U2621 ( .ins ({new_AGEMA_signal_15242, new_AGEMA_signal_15240, new_AGEMA_signal_15238, new_AGEMA_signal_15236}), .inb ({new_AGEMA_signal_2774, new_AGEMA_signal_2773, new_AGEMA_signal_2772, n2469}), .ina ({new_AGEMA_signal_15266, new_AGEMA_signal_15260, new_AGEMA_signal_15254, new_AGEMA_signal_15248}), .clk ( clk ), .rnd ({Fresh[7019], Fresh[7018], Fresh[7017], Fresh[7016], Fresh[7015], Fresh[7014], Fresh[7013], Fresh[7012], Fresh[7011], Fresh[7010]}), .outt ({new_AGEMA_signal_3035, new_AGEMA_signal_3034, new_AGEMA_signal_3033, n2471}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2636 ( .ina ({new_AGEMA_signal_15290, new_AGEMA_signal_15284, new_AGEMA_signal_15278, new_AGEMA_signal_15272}), .inb ({new_AGEMA_signal_3038, new_AGEMA_signal_3037, new_AGEMA_signal_3036, n2484}), .clk ( clk ), .rnd ({Fresh[7029], Fresh[7028], Fresh[7027], Fresh[7026], Fresh[7025], Fresh[7024], Fresh[7023], Fresh[7022], Fresh[7021], Fresh[7020]}), .outt ({new_AGEMA_signal_3236, new_AGEMA_signal_3235, new_AGEMA_signal_3234, n2485}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2644 ( .ina ({new_AGEMA_signal_14794, new_AGEMA_signal_14788, new_AGEMA_signal_14782, new_AGEMA_signal_14776}), .inb ({new_AGEMA_signal_2783, new_AGEMA_signal_2782, new_AGEMA_signal_2781, n2491}), .clk ( clk ), .rnd ({Fresh[7039], Fresh[7038], Fresh[7037], Fresh[7036], Fresh[7035], Fresh[7034], Fresh[7033], Fresh[7032], Fresh[7031], Fresh[7030]}), .outt ({new_AGEMA_signal_3041, new_AGEMA_signal_3040, new_AGEMA_signal_3039, n2502}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2651 ( .ina ({new_AGEMA_signal_3044, new_AGEMA_signal_3043, new_AGEMA_signal_3042, n2500}), .inb ({new_AGEMA_signal_15306, new_AGEMA_signal_15302, new_AGEMA_signal_15298, new_AGEMA_signal_15294}), .clk ( clk ), .rnd ({Fresh[7049], Fresh[7048], Fresh[7047], Fresh[7046], Fresh[7045], Fresh[7044], Fresh[7043], Fresh[7042], Fresh[7041], Fresh[7040]}), .outt ({new_AGEMA_signal_3239, new_AGEMA_signal_3238, new_AGEMA_signal_3237, n2501}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2657 ( .ina ({new_AGEMA_signal_15210, new_AGEMA_signal_15206, new_AGEMA_signal_15202, new_AGEMA_signal_15198}), .inb ({new_AGEMA_signal_3242, new_AGEMA_signal_3241, new_AGEMA_signal_3240, n2508}), .clk ( clk ), .rnd ({Fresh[7059], Fresh[7058], Fresh[7057], Fresh[7056], Fresh[7055], Fresh[7054], Fresh[7053], Fresh[7052], Fresh[7051], Fresh[7050]}), .outt ({new_AGEMA_signal_3389, new_AGEMA_signal_3388, new_AGEMA_signal_3387, n2509}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2671 ( .ina ({new_AGEMA_signal_15314, new_AGEMA_signal_15312, new_AGEMA_signal_15310, new_AGEMA_signal_15308}), .inb ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, new_AGEMA_signal_3243, n2526}), .clk ( clk ), .rnd ({Fresh[7069], Fresh[7068], Fresh[7067], Fresh[7066], Fresh[7065], Fresh[7064], Fresh[7063], Fresh[7062], Fresh[7061], Fresh[7060]}), .outt ({new_AGEMA_signal_3392, new_AGEMA_signal_3391, new_AGEMA_signal_3390, n2527}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2680 ( .ina ({new_AGEMA_signal_3053, new_AGEMA_signal_3052, new_AGEMA_signal_3051, n2539}), .inb ({new_AGEMA_signal_15346, new_AGEMA_signal_15338, new_AGEMA_signal_15330, new_AGEMA_signal_15322}), .clk ( clk ), .rnd ({Fresh[7079], Fresh[7078], Fresh[7077], Fresh[7076], Fresh[7075], Fresh[7074], Fresh[7073], Fresh[7072], Fresh[7071], Fresh[7070]}), .outt ({new_AGEMA_signal_3248, new_AGEMA_signal_3247, new_AGEMA_signal_3246, n2550}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2685 ( .ina ({new_AGEMA_signal_3056, new_AGEMA_signal_3055, new_AGEMA_signal_3054, n2548}), .inb ({new_AGEMA_signal_15354, new_AGEMA_signal_15352, new_AGEMA_signal_15350, new_AGEMA_signal_15348}), .clk ( clk ), .rnd ({Fresh[7089], Fresh[7088], Fresh[7087], Fresh[7086], Fresh[7085], Fresh[7084], Fresh[7083], Fresh[7082], Fresh[7081], Fresh[7080]}), .outt ({new_AGEMA_signal_3251, new_AGEMA_signal_3250, new_AGEMA_signal_3249, n2549}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2701 ( .ina ({new_AGEMA_signal_3059, new_AGEMA_signal_3058, new_AGEMA_signal_3057, n2568}), .inb ({new_AGEMA_signal_3062, new_AGEMA_signal_3061, new_AGEMA_signal_3060, n2567}), .clk ( clk ), .rnd ({Fresh[7099], Fresh[7098], Fresh[7097], Fresh[7096], Fresh[7095], Fresh[7094], Fresh[7093], Fresh[7092], Fresh[7091], Fresh[7090]}), .outt ({new_AGEMA_signal_3254, new_AGEMA_signal_3253, new_AGEMA_signal_3252, n2569}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2712 ( .ina ({new_AGEMA_signal_3065, new_AGEMA_signal_3064, new_AGEMA_signal_3063, n2583}), .inb ({new_AGEMA_signal_15370, new_AGEMA_signal_15366, new_AGEMA_signal_15362, new_AGEMA_signal_15358}), .clk ( clk ), .rnd ({Fresh[7109], Fresh[7108], Fresh[7107], Fresh[7106], Fresh[7105], Fresh[7104], Fresh[7103], Fresh[7102], Fresh[7101], Fresh[7100]}), .outt ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, new_AGEMA_signal_3255, n2584}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2729 ( .ina ({new_AGEMA_signal_15386, new_AGEMA_signal_15382, new_AGEMA_signal_15378, new_AGEMA_signal_15374}), .inb ({new_AGEMA_signal_2816, new_AGEMA_signal_2815, new_AGEMA_signal_2814, n2604}), .clk ( clk ), .rnd ({Fresh[7119], Fresh[7118], Fresh[7117], Fresh[7116], Fresh[7115], Fresh[7114], Fresh[7113], Fresh[7112], Fresh[7111], Fresh[7110]}), .outt ({new_AGEMA_signal_3068, new_AGEMA_signal_3067, new_AGEMA_signal_3066, n2606}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2740 ( .ina ({new_AGEMA_signal_14794, new_AGEMA_signal_14788, new_AGEMA_signal_14782, new_AGEMA_signal_14776}), .inb ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, new_AGEMA_signal_3069, n2621}), .clk ( clk ), .rnd ({Fresh[7129], Fresh[7128], Fresh[7127], Fresh[7126], Fresh[7125], Fresh[7124], Fresh[7123], Fresh[7122], Fresh[7121], Fresh[7120]}), .outt ({new_AGEMA_signal_3263, new_AGEMA_signal_3262, new_AGEMA_signal_3261, n2622}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2747 ( .ina ({new_AGEMA_signal_3074, new_AGEMA_signal_3073, new_AGEMA_signal_3072, n2633}), .inb ({new_AGEMA_signal_15402, new_AGEMA_signal_15398, new_AGEMA_signal_15394, new_AGEMA_signal_15390}), .clk ( clk ), .rnd ({Fresh[7139], Fresh[7138], Fresh[7137], Fresh[7136], Fresh[7135], Fresh[7134], Fresh[7133], Fresh[7132], Fresh[7131], Fresh[7130]}), .outt ({new_AGEMA_signal_3266, new_AGEMA_signal_3265, new_AGEMA_signal_3264, n2634}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2761 ( .ina ({new_AGEMA_signal_3080, new_AGEMA_signal_3079, new_AGEMA_signal_3078, n2656}), .inb ({new_AGEMA_signal_15418, new_AGEMA_signal_15414, new_AGEMA_signal_15410, new_AGEMA_signal_15406}), .clk ( clk ), .rnd ({Fresh[7149], Fresh[7148], Fresh[7147], Fresh[7146], Fresh[7145], Fresh[7144], Fresh[7143], Fresh[7142], Fresh[7141], Fresh[7140]}), .outt ({new_AGEMA_signal_3269, new_AGEMA_signal_3268, new_AGEMA_signal_3267, n2657}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2783 ( .ina ({new_AGEMA_signal_3092, new_AGEMA_signal_3091, new_AGEMA_signal_3090, n2696}), .inb ({new_AGEMA_signal_15434, new_AGEMA_signal_15430, new_AGEMA_signal_15426, new_AGEMA_signal_15422}), .clk ( clk ), .rnd ({Fresh[7159], Fresh[7158], Fresh[7157], Fresh[7156], Fresh[7155], Fresh[7154], Fresh[7153], Fresh[7152], Fresh[7151], Fresh[7150]}), .outt ({new_AGEMA_signal_3272, new_AGEMA_signal_3271, new_AGEMA_signal_3270, n2697}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2795 ( .ina ({new_AGEMA_signal_14770, new_AGEMA_signal_14768, new_AGEMA_signal_14766, new_AGEMA_signal_14764}), .inb ({new_AGEMA_signal_3095, new_AGEMA_signal_3094, new_AGEMA_signal_3093, n2718}), .clk ( clk ), .rnd ({Fresh[7169], Fresh[7168], Fresh[7167], Fresh[7166], Fresh[7165], Fresh[7164], Fresh[7163], Fresh[7162], Fresh[7161], Fresh[7160]}), .outt ({new_AGEMA_signal_3275, new_AGEMA_signal_3274, new_AGEMA_signal_3273, n2808}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2802 ( .ina ({new_AGEMA_signal_3098, new_AGEMA_signal_3097, new_AGEMA_signal_3096, n2730}), .inb ({new_AGEMA_signal_15466, new_AGEMA_signal_15458, new_AGEMA_signal_15450, new_AGEMA_signal_15442}), .clk ( clk ), .rnd ({Fresh[7179], Fresh[7178], Fresh[7177], Fresh[7176], Fresh[7175], Fresh[7174], Fresh[7173], Fresh[7172], Fresh[7171], Fresh[7170]}), .outt ({new_AGEMA_signal_3278, new_AGEMA_signal_3277, new_AGEMA_signal_3276, n2747}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2810 ( .ina ({new_AGEMA_signal_3101, new_AGEMA_signal_3100, new_AGEMA_signal_3099, n2745}), .inb ({new_AGEMA_signal_3104, new_AGEMA_signal_3103, new_AGEMA_signal_3102, n2744}), .clk ( clk ), .rnd ({Fresh[7189], Fresh[7188], Fresh[7187], Fresh[7186], Fresh[7185], Fresh[7184], Fresh[7183], Fresh[7182], Fresh[7181], Fresh[7180]}), .outt ({new_AGEMA_signal_3281, new_AGEMA_signal_3280, new_AGEMA_signal_3279, n2746}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2818 ( .ina ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, new_AGEMA_signal_3105, n2759}), .inb ({new_AGEMA_signal_15474, new_AGEMA_signal_15472, new_AGEMA_signal_15470, new_AGEMA_signal_15468}), .clk ( clk ), .rnd ({Fresh[7199], Fresh[7198], Fresh[7197], Fresh[7196], Fresh[7195], Fresh[7194], Fresh[7193], Fresh[7192], Fresh[7191], Fresh[7190]}), .outt ({new_AGEMA_signal_3284, new_AGEMA_signal_3283, new_AGEMA_signal_3282, n2804}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2824 ( .ina ({new_AGEMA_signal_3110, new_AGEMA_signal_3109, new_AGEMA_signal_3108, n2771}), .inb ({new_AGEMA_signal_15490, new_AGEMA_signal_15486, new_AGEMA_signal_15482, new_AGEMA_signal_15478}), .clk ( clk ), .rnd ({Fresh[7209], Fresh[7208], Fresh[7207], Fresh[7206], Fresh[7205], Fresh[7204], Fresh[7203], Fresh[7202], Fresh[7201], Fresh[7200]}), .outt ({new_AGEMA_signal_3287, new_AGEMA_signal_3286, new_AGEMA_signal_3285, n2802}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2838 ( .ina ({new_AGEMA_signal_2864, new_AGEMA_signal_2863, new_AGEMA_signal_2862, n2798}), .inb ({new_AGEMA_signal_15498, new_AGEMA_signal_15496, new_AGEMA_signal_15494, new_AGEMA_signal_15492}), .clk ( clk ), .rnd ({Fresh[7219], Fresh[7218], Fresh[7217], Fresh[7216], Fresh[7215], Fresh[7214], Fresh[7213], Fresh[7212], Fresh[7211], Fresh[7210]}), .outt ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, new_AGEMA_signal_3111, n2799}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2852 ( .ina ({new_AGEMA_signal_3116, new_AGEMA_signal_3115, new_AGEMA_signal_3114, n2826}), .inb ({new_AGEMA_signal_15522, new_AGEMA_signal_15516, new_AGEMA_signal_15510, new_AGEMA_signal_15504}), .clk ( clk ), .rnd ({Fresh[7229], Fresh[7228], Fresh[7227], Fresh[7226], Fresh[7225], Fresh[7224], Fresh[7223], Fresh[7222], Fresh[7221], Fresh[7220]}), .outt ({new_AGEMA_signal_3293, new_AGEMA_signal_3292, new_AGEMA_signal_3291, n2827}) ) ;
    buf_clk new_AGEMA_reg_buffer_4024 ( .C ( clk ), .D ( new_AGEMA_signal_15523 ), .Q ( new_AGEMA_signal_15524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4026 ( .C ( clk ), .D ( new_AGEMA_signal_15525 ), .Q ( new_AGEMA_signal_15526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4028 ( .C ( clk ), .D ( new_AGEMA_signal_15527 ), .Q ( new_AGEMA_signal_15528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4030 ( .C ( clk ), .D ( new_AGEMA_signal_15529 ), .Q ( new_AGEMA_signal_15530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4038 ( .C ( clk ), .D ( new_AGEMA_signal_15537 ), .Q ( new_AGEMA_signal_15538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4046 ( .C ( clk ), .D ( new_AGEMA_signal_15545 ), .Q ( new_AGEMA_signal_15546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4054 ( .C ( clk ), .D ( new_AGEMA_signal_15553 ), .Q ( new_AGEMA_signal_15554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4062 ( .C ( clk ), .D ( new_AGEMA_signal_15561 ), .Q ( new_AGEMA_signal_15562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4064 ( .C ( clk ), .D ( new_AGEMA_signal_15563 ), .Q ( new_AGEMA_signal_15564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4066 ( .C ( clk ), .D ( new_AGEMA_signal_15565 ), .Q ( new_AGEMA_signal_15566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4068 ( .C ( clk ), .D ( new_AGEMA_signal_15567 ), .Q ( new_AGEMA_signal_15568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4070 ( .C ( clk ), .D ( new_AGEMA_signal_15569 ), .Q ( new_AGEMA_signal_15570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4074 ( .C ( clk ), .D ( new_AGEMA_signal_15573 ), .Q ( new_AGEMA_signal_15574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4078 ( .C ( clk ), .D ( new_AGEMA_signal_15577 ), .Q ( new_AGEMA_signal_15578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4082 ( .C ( clk ), .D ( new_AGEMA_signal_15581 ), .Q ( new_AGEMA_signal_15582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4086 ( .C ( clk ), .D ( new_AGEMA_signal_15585 ), .Q ( new_AGEMA_signal_15586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4094 ( .C ( clk ), .D ( new_AGEMA_signal_15593 ), .Q ( new_AGEMA_signal_15594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4102 ( .C ( clk ), .D ( new_AGEMA_signal_15601 ), .Q ( new_AGEMA_signal_15602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4110 ( .C ( clk ), .D ( new_AGEMA_signal_15609 ), .Q ( new_AGEMA_signal_15610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4118 ( .C ( clk ), .D ( new_AGEMA_signal_15617 ), .Q ( new_AGEMA_signal_15618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4120 ( .C ( clk ), .D ( new_AGEMA_signal_15619 ), .Q ( new_AGEMA_signal_15620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4122 ( .C ( clk ), .D ( new_AGEMA_signal_15621 ), .Q ( new_AGEMA_signal_15622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4124 ( .C ( clk ), .D ( new_AGEMA_signal_15623 ), .Q ( new_AGEMA_signal_15624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4126 ( .C ( clk ), .D ( new_AGEMA_signal_15625 ), .Q ( new_AGEMA_signal_15626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4132 ( .C ( clk ), .D ( new_AGEMA_signal_15631 ), .Q ( new_AGEMA_signal_15632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4138 ( .C ( clk ), .D ( new_AGEMA_signal_15637 ), .Q ( new_AGEMA_signal_15638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4144 ( .C ( clk ), .D ( new_AGEMA_signal_15643 ), .Q ( new_AGEMA_signal_15644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4150 ( .C ( clk ), .D ( new_AGEMA_signal_15649 ), .Q ( new_AGEMA_signal_15650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4154 ( .C ( clk ), .D ( new_AGEMA_signal_15653 ), .Q ( new_AGEMA_signal_15654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4158 ( .C ( clk ), .D ( new_AGEMA_signal_15657 ), .Q ( new_AGEMA_signal_15658 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4162 ( .C ( clk ), .D ( new_AGEMA_signal_15661 ), .Q ( new_AGEMA_signal_15662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4166 ( .C ( clk ), .D ( new_AGEMA_signal_15665 ), .Q ( new_AGEMA_signal_15666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4174 ( .C ( clk ), .D ( new_AGEMA_signal_15673 ), .Q ( new_AGEMA_signal_15674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4182 ( .C ( clk ), .D ( new_AGEMA_signal_15681 ), .Q ( new_AGEMA_signal_15682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4190 ( .C ( clk ), .D ( new_AGEMA_signal_15689 ), .Q ( new_AGEMA_signal_15690 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4198 ( .C ( clk ), .D ( new_AGEMA_signal_15697 ), .Q ( new_AGEMA_signal_15698 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4202 ( .C ( clk ), .D ( new_AGEMA_signal_15701 ), .Q ( new_AGEMA_signal_15702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4206 ( .C ( clk ), .D ( new_AGEMA_signal_15705 ), .Q ( new_AGEMA_signal_15706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4210 ( .C ( clk ), .D ( new_AGEMA_signal_15709 ), .Q ( new_AGEMA_signal_15710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4214 ( .C ( clk ), .D ( new_AGEMA_signal_15713 ), .Q ( new_AGEMA_signal_15714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4220 ( .C ( clk ), .D ( new_AGEMA_signal_15719 ), .Q ( new_AGEMA_signal_15720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4226 ( .C ( clk ), .D ( new_AGEMA_signal_15725 ), .Q ( new_AGEMA_signal_15726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4232 ( .C ( clk ), .D ( new_AGEMA_signal_15731 ), .Q ( new_AGEMA_signal_15732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4238 ( .C ( clk ), .D ( new_AGEMA_signal_15737 ), .Q ( new_AGEMA_signal_15738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4244 ( .C ( clk ), .D ( new_AGEMA_signal_15743 ), .Q ( new_AGEMA_signal_15744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4250 ( .C ( clk ), .D ( new_AGEMA_signal_15749 ), .Q ( new_AGEMA_signal_15750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4256 ( .C ( clk ), .D ( new_AGEMA_signal_15755 ), .Q ( new_AGEMA_signal_15756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4262 ( .C ( clk ), .D ( new_AGEMA_signal_15761 ), .Q ( new_AGEMA_signal_15762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4268 ( .C ( clk ), .D ( new_AGEMA_signal_15767 ), .Q ( new_AGEMA_signal_15768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4274 ( .C ( clk ), .D ( new_AGEMA_signal_15773 ), .Q ( new_AGEMA_signal_15774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4280 ( .C ( clk ), .D ( new_AGEMA_signal_15779 ), .Q ( new_AGEMA_signal_15780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4286 ( .C ( clk ), .D ( new_AGEMA_signal_15785 ), .Q ( new_AGEMA_signal_15786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4292 ( .C ( clk ), .D ( new_AGEMA_signal_15791 ), .Q ( new_AGEMA_signal_15792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4298 ( .C ( clk ), .D ( new_AGEMA_signal_15797 ), .Q ( new_AGEMA_signal_15798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4304 ( .C ( clk ), .D ( new_AGEMA_signal_15803 ), .Q ( new_AGEMA_signal_15804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4310 ( .C ( clk ), .D ( new_AGEMA_signal_15809 ), .Q ( new_AGEMA_signal_15810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4316 ( .C ( clk ), .D ( new_AGEMA_signal_15815 ), .Q ( new_AGEMA_signal_15816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4322 ( .C ( clk ), .D ( new_AGEMA_signal_15821 ), .Q ( new_AGEMA_signal_15822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4328 ( .C ( clk ), .D ( new_AGEMA_signal_15827 ), .Q ( new_AGEMA_signal_15828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4334 ( .C ( clk ), .D ( new_AGEMA_signal_15833 ), .Q ( new_AGEMA_signal_15834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4338 ( .C ( clk ), .D ( new_AGEMA_signal_15837 ), .Q ( new_AGEMA_signal_15838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4342 ( .C ( clk ), .D ( new_AGEMA_signal_15841 ), .Q ( new_AGEMA_signal_15842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4346 ( .C ( clk ), .D ( new_AGEMA_signal_15845 ), .Q ( new_AGEMA_signal_15846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4350 ( .C ( clk ), .D ( new_AGEMA_signal_15849 ), .Q ( new_AGEMA_signal_15850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4358 ( .C ( clk ), .D ( new_AGEMA_signal_15857 ), .Q ( new_AGEMA_signal_15858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4366 ( .C ( clk ), .D ( new_AGEMA_signal_15865 ), .Q ( new_AGEMA_signal_15866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4374 ( .C ( clk ), .D ( new_AGEMA_signal_15873 ), .Q ( new_AGEMA_signal_15874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4382 ( .C ( clk ), .D ( new_AGEMA_signal_15881 ), .Q ( new_AGEMA_signal_15882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4386 ( .C ( clk ), .D ( new_AGEMA_signal_15885 ), .Q ( new_AGEMA_signal_15886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4390 ( .C ( clk ), .D ( new_AGEMA_signal_15889 ), .Q ( new_AGEMA_signal_15890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4394 ( .C ( clk ), .D ( new_AGEMA_signal_15893 ), .Q ( new_AGEMA_signal_15894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4398 ( .C ( clk ), .D ( new_AGEMA_signal_15897 ), .Q ( new_AGEMA_signal_15898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4404 ( .C ( clk ), .D ( new_AGEMA_signal_15903 ), .Q ( new_AGEMA_signal_15904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4410 ( .C ( clk ), .D ( new_AGEMA_signal_15909 ), .Q ( new_AGEMA_signal_15910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4416 ( .C ( clk ), .D ( new_AGEMA_signal_15915 ), .Q ( new_AGEMA_signal_15916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4422 ( .C ( clk ), .D ( new_AGEMA_signal_15921 ), .Q ( new_AGEMA_signal_15922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4430 ( .C ( clk ), .D ( new_AGEMA_signal_15929 ), .Q ( new_AGEMA_signal_15930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4438 ( .C ( clk ), .D ( new_AGEMA_signal_15937 ), .Q ( new_AGEMA_signal_15938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4446 ( .C ( clk ), .D ( new_AGEMA_signal_15945 ), .Q ( new_AGEMA_signal_15946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4454 ( .C ( clk ), .D ( new_AGEMA_signal_15953 ), .Q ( new_AGEMA_signal_15954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4456 ( .C ( clk ), .D ( new_AGEMA_signal_15955 ), .Q ( new_AGEMA_signal_15956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4458 ( .C ( clk ), .D ( new_AGEMA_signal_15957 ), .Q ( new_AGEMA_signal_15958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4460 ( .C ( clk ), .D ( new_AGEMA_signal_15959 ), .Q ( new_AGEMA_signal_15960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4462 ( .C ( clk ), .D ( new_AGEMA_signal_15961 ), .Q ( new_AGEMA_signal_15962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4468 ( .C ( clk ), .D ( new_AGEMA_signal_15967 ), .Q ( new_AGEMA_signal_15968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4474 ( .C ( clk ), .D ( new_AGEMA_signal_15973 ), .Q ( new_AGEMA_signal_15974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4480 ( .C ( clk ), .D ( new_AGEMA_signal_15979 ), .Q ( new_AGEMA_signal_15980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4486 ( .C ( clk ), .D ( new_AGEMA_signal_15985 ), .Q ( new_AGEMA_signal_15986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4488 ( .C ( clk ), .D ( new_AGEMA_signal_15987 ), .Q ( new_AGEMA_signal_15988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4490 ( .C ( clk ), .D ( new_AGEMA_signal_15989 ), .Q ( new_AGEMA_signal_15990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4492 ( .C ( clk ), .D ( new_AGEMA_signal_15991 ), .Q ( new_AGEMA_signal_15992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4494 ( .C ( clk ), .D ( new_AGEMA_signal_15993 ), .Q ( new_AGEMA_signal_15994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4496 ( .C ( clk ), .D ( new_AGEMA_signal_15995 ), .Q ( new_AGEMA_signal_15996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4498 ( .C ( clk ), .D ( new_AGEMA_signal_15997 ), .Q ( new_AGEMA_signal_15998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4500 ( .C ( clk ), .D ( new_AGEMA_signal_15999 ), .Q ( new_AGEMA_signal_16000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4502 ( .C ( clk ), .D ( new_AGEMA_signal_16001 ), .Q ( new_AGEMA_signal_16002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4508 ( .C ( clk ), .D ( new_AGEMA_signal_16007 ), .Q ( new_AGEMA_signal_16008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4514 ( .C ( clk ), .D ( new_AGEMA_signal_16013 ), .Q ( new_AGEMA_signal_16014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4520 ( .C ( clk ), .D ( new_AGEMA_signal_16019 ), .Q ( new_AGEMA_signal_16020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4526 ( .C ( clk ), .D ( new_AGEMA_signal_16025 ), .Q ( new_AGEMA_signal_16026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4532 ( .C ( clk ), .D ( new_AGEMA_signal_16031 ), .Q ( new_AGEMA_signal_16032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4538 ( .C ( clk ), .D ( new_AGEMA_signal_16037 ), .Q ( new_AGEMA_signal_16038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4544 ( .C ( clk ), .D ( new_AGEMA_signal_16043 ), .Q ( new_AGEMA_signal_16044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4550 ( .C ( clk ), .D ( new_AGEMA_signal_16049 ), .Q ( new_AGEMA_signal_16050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4558 ( .C ( clk ), .D ( new_AGEMA_signal_16057 ), .Q ( new_AGEMA_signal_16058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4566 ( .C ( clk ), .D ( new_AGEMA_signal_16065 ), .Q ( new_AGEMA_signal_16066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4574 ( .C ( clk ), .D ( new_AGEMA_signal_16073 ), .Q ( new_AGEMA_signal_16074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4582 ( .C ( clk ), .D ( new_AGEMA_signal_16081 ), .Q ( new_AGEMA_signal_16082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4590 ( .C ( clk ), .D ( new_AGEMA_signal_16089 ), .Q ( new_AGEMA_signal_16090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4598 ( .C ( clk ), .D ( new_AGEMA_signal_16097 ), .Q ( new_AGEMA_signal_16098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4606 ( .C ( clk ), .D ( new_AGEMA_signal_16105 ), .Q ( new_AGEMA_signal_16106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4614 ( .C ( clk ), .D ( new_AGEMA_signal_16113 ), .Q ( new_AGEMA_signal_16114 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4620 ( .C ( clk ), .D ( new_AGEMA_signal_16119 ), .Q ( new_AGEMA_signal_16120 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4626 ( .C ( clk ), .D ( new_AGEMA_signal_16125 ), .Q ( new_AGEMA_signal_16126 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4632 ( .C ( clk ), .D ( new_AGEMA_signal_16131 ), .Q ( new_AGEMA_signal_16132 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4638 ( .C ( clk ), .D ( new_AGEMA_signal_16137 ), .Q ( new_AGEMA_signal_16138 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4644 ( .C ( clk ), .D ( new_AGEMA_signal_16143 ), .Q ( new_AGEMA_signal_16144 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4650 ( .C ( clk ), .D ( new_AGEMA_signal_16149 ), .Q ( new_AGEMA_signal_16150 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4656 ( .C ( clk ), .D ( new_AGEMA_signal_16155 ), .Q ( new_AGEMA_signal_16156 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4662 ( .C ( clk ), .D ( new_AGEMA_signal_16161 ), .Q ( new_AGEMA_signal_16162 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4664 ( .C ( clk ), .D ( new_AGEMA_signal_16163 ), .Q ( new_AGEMA_signal_16164 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4666 ( .C ( clk ), .D ( new_AGEMA_signal_16165 ), .Q ( new_AGEMA_signal_16166 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4668 ( .C ( clk ), .D ( new_AGEMA_signal_16167 ), .Q ( new_AGEMA_signal_16168 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4670 ( .C ( clk ), .D ( new_AGEMA_signal_16169 ), .Q ( new_AGEMA_signal_16170 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4674 ( .C ( clk ), .D ( new_AGEMA_signal_16173 ), .Q ( new_AGEMA_signal_16174 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4678 ( .C ( clk ), .D ( new_AGEMA_signal_16177 ), .Q ( new_AGEMA_signal_16178 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4682 ( .C ( clk ), .D ( new_AGEMA_signal_16181 ), .Q ( new_AGEMA_signal_16182 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4686 ( .C ( clk ), .D ( new_AGEMA_signal_16185 ), .Q ( new_AGEMA_signal_16186 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4690 ( .C ( clk ), .D ( new_AGEMA_signal_16189 ), .Q ( new_AGEMA_signal_16190 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4694 ( .C ( clk ), .D ( new_AGEMA_signal_16193 ), .Q ( new_AGEMA_signal_16194 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4698 ( .C ( clk ), .D ( new_AGEMA_signal_16197 ), .Q ( new_AGEMA_signal_16198 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4702 ( .C ( clk ), .D ( new_AGEMA_signal_16201 ), .Q ( new_AGEMA_signal_16202 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4706 ( .C ( clk ), .D ( new_AGEMA_signal_16205 ), .Q ( new_AGEMA_signal_16206 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4710 ( .C ( clk ), .D ( new_AGEMA_signal_16209 ), .Q ( new_AGEMA_signal_16210 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4714 ( .C ( clk ), .D ( new_AGEMA_signal_16213 ), .Q ( new_AGEMA_signal_16214 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4718 ( .C ( clk ), .D ( new_AGEMA_signal_16217 ), .Q ( new_AGEMA_signal_16218 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4720 ( .C ( clk ), .D ( new_AGEMA_signal_16219 ), .Q ( new_AGEMA_signal_16220 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4722 ( .C ( clk ), .D ( new_AGEMA_signal_16221 ), .Q ( new_AGEMA_signal_16222 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4724 ( .C ( clk ), .D ( new_AGEMA_signal_16223 ), .Q ( new_AGEMA_signal_16224 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4726 ( .C ( clk ), .D ( new_AGEMA_signal_16225 ), .Q ( new_AGEMA_signal_16226 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4730 ( .C ( clk ), .D ( new_AGEMA_signal_16229 ), .Q ( new_AGEMA_signal_16230 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4736 ( .C ( clk ), .D ( new_AGEMA_signal_16235 ), .Q ( new_AGEMA_signal_16236 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4742 ( .C ( clk ), .D ( new_AGEMA_signal_16241 ), .Q ( new_AGEMA_signal_16242 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4748 ( .C ( clk ), .D ( new_AGEMA_signal_16247 ), .Q ( new_AGEMA_signal_16248 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4760 ( .C ( clk ), .D ( new_AGEMA_signal_16259 ), .Q ( new_AGEMA_signal_16260 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4764 ( .C ( clk ), .D ( new_AGEMA_signal_16263 ), .Q ( new_AGEMA_signal_16264 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4768 ( .C ( clk ), .D ( new_AGEMA_signal_16267 ), .Q ( new_AGEMA_signal_16268 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4772 ( .C ( clk ), .D ( new_AGEMA_signal_16271 ), .Q ( new_AGEMA_signal_16272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4780 ( .C ( clk ), .D ( new_AGEMA_signal_16279 ), .Q ( new_AGEMA_signal_16280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4788 ( .C ( clk ), .D ( new_AGEMA_signal_16287 ), .Q ( new_AGEMA_signal_16288 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4796 ( .C ( clk ), .D ( new_AGEMA_signal_16295 ), .Q ( new_AGEMA_signal_16296 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4804 ( .C ( clk ), .D ( new_AGEMA_signal_16303 ), .Q ( new_AGEMA_signal_16304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4812 ( .C ( clk ), .D ( new_AGEMA_signal_16311 ), .Q ( new_AGEMA_signal_16312 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4820 ( .C ( clk ), .D ( new_AGEMA_signal_16319 ), .Q ( new_AGEMA_signal_16320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4828 ( .C ( clk ), .D ( new_AGEMA_signal_16327 ), .Q ( new_AGEMA_signal_16328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4836 ( .C ( clk ), .D ( new_AGEMA_signal_16335 ), .Q ( new_AGEMA_signal_16336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4844 ( .C ( clk ), .D ( new_AGEMA_signal_16343 ), .Q ( new_AGEMA_signal_16344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4852 ( .C ( clk ), .D ( new_AGEMA_signal_16351 ), .Q ( new_AGEMA_signal_16352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4860 ( .C ( clk ), .D ( new_AGEMA_signal_16359 ), .Q ( new_AGEMA_signal_16360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4868 ( .C ( clk ), .D ( new_AGEMA_signal_16367 ), .Q ( new_AGEMA_signal_16368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4876 ( .C ( clk ), .D ( new_AGEMA_signal_16375 ), .Q ( new_AGEMA_signal_16376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4884 ( .C ( clk ), .D ( new_AGEMA_signal_16383 ), .Q ( new_AGEMA_signal_16384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4892 ( .C ( clk ), .D ( new_AGEMA_signal_16391 ), .Q ( new_AGEMA_signal_16392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4900 ( .C ( clk ), .D ( new_AGEMA_signal_16399 ), .Q ( new_AGEMA_signal_16400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4906 ( .C ( clk ), .D ( new_AGEMA_signal_16405 ), .Q ( new_AGEMA_signal_16406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4912 ( .C ( clk ), .D ( new_AGEMA_signal_16411 ), .Q ( new_AGEMA_signal_16412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4918 ( .C ( clk ), .D ( new_AGEMA_signal_16417 ), .Q ( new_AGEMA_signal_16418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4924 ( .C ( clk ), .D ( new_AGEMA_signal_16423 ), .Q ( new_AGEMA_signal_16424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4934 ( .C ( clk ), .D ( new_AGEMA_signal_16433 ), .Q ( new_AGEMA_signal_16434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4944 ( .C ( clk ), .D ( new_AGEMA_signal_16443 ), .Q ( new_AGEMA_signal_16444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4954 ( .C ( clk ), .D ( new_AGEMA_signal_16453 ), .Q ( new_AGEMA_signal_16454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4964 ( .C ( clk ), .D ( new_AGEMA_signal_16463 ), .Q ( new_AGEMA_signal_16464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4972 ( .C ( clk ), .D ( new_AGEMA_signal_16471 ), .Q ( new_AGEMA_signal_16472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4980 ( .C ( clk ), .D ( new_AGEMA_signal_16479 ), .Q ( new_AGEMA_signal_16480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4988 ( .C ( clk ), .D ( new_AGEMA_signal_16487 ), .Q ( new_AGEMA_signal_16488 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4996 ( .C ( clk ), .D ( new_AGEMA_signal_16495 ), .Q ( new_AGEMA_signal_16496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5004 ( .C ( clk ), .D ( new_AGEMA_signal_16503 ), .Q ( new_AGEMA_signal_16504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5012 ( .C ( clk ), .D ( new_AGEMA_signal_16511 ), .Q ( new_AGEMA_signal_16512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5020 ( .C ( clk ), .D ( new_AGEMA_signal_16519 ), .Q ( new_AGEMA_signal_16520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5028 ( .C ( clk ), .D ( new_AGEMA_signal_16527 ), .Q ( new_AGEMA_signal_16528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5036 ( .C ( clk ), .D ( new_AGEMA_signal_16535 ), .Q ( new_AGEMA_signal_16536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5044 ( .C ( clk ), .D ( new_AGEMA_signal_16543 ), .Q ( new_AGEMA_signal_16544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5052 ( .C ( clk ), .D ( new_AGEMA_signal_16551 ), .Q ( new_AGEMA_signal_16552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5060 ( .C ( clk ), .D ( new_AGEMA_signal_16559 ), .Q ( new_AGEMA_signal_16560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5072 ( .C ( clk ), .D ( new_AGEMA_signal_16571 ), .Q ( new_AGEMA_signal_16572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5076 ( .C ( clk ), .D ( new_AGEMA_signal_16575 ), .Q ( new_AGEMA_signal_16576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5080 ( .C ( clk ), .D ( new_AGEMA_signal_16579 ), .Q ( new_AGEMA_signal_16580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5084 ( .C ( clk ), .D ( new_AGEMA_signal_16583 ), .Q ( new_AGEMA_signal_16584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5090 ( .C ( clk ), .D ( new_AGEMA_signal_16589 ), .Q ( new_AGEMA_signal_16590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5096 ( .C ( clk ), .D ( new_AGEMA_signal_16595 ), .Q ( new_AGEMA_signal_16596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5102 ( .C ( clk ), .D ( new_AGEMA_signal_16601 ), .Q ( new_AGEMA_signal_16602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5108 ( .C ( clk ), .D ( new_AGEMA_signal_16607 ), .Q ( new_AGEMA_signal_16608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5112 ( .C ( clk ), .D ( new_AGEMA_signal_16611 ), .Q ( new_AGEMA_signal_16612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5116 ( .C ( clk ), .D ( new_AGEMA_signal_16615 ), .Q ( new_AGEMA_signal_16616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5120 ( .C ( clk ), .D ( new_AGEMA_signal_16619 ), .Q ( new_AGEMA_signal_16620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5124 ( .C ( clk ), .D ( new_AGEMA_signal_16623 ), .Q ( new_AGEMA_signal_16624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5134 ( .C ( clk ), .D ( new_AGEMA_signal_16633 ), .Q ( new_AGEMA_signal_16634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5144 ( .C ( clk ), .D ( new_AGEMA_signal_16643 ), .Q ( new_AGEMA_signal_16644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5154 ( .C ( clk ), .D ( new_AGEMA_signal_16653 ), .Q ( new_AGEMA_signal_16654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5164 ( .C ( clk ), .D ( new_AGEMA_signal_16663 ), .Q ( new_AGEMA_signal_16664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5172 ( .C ( clk ), .D ( new_AGEMA_signal_16671 ), .Q ( new_AGEMA_signal_16672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5180 ( .C ( clk ), .D ( new_AGEMA_signal_16679 ), .Q ( new_AGEMA_signal_16680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5188 ( .C ( clk ), .D ( new_AGEMA_signal_16687 ), .Q ( new_AGEMA_signal_16688 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5196 ( .C ( clk ), .D ( new_AGEMA_signal_16695 ), .Q ( new_AGEMA_signal_16696 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5200 ( .C ( clk ), .D ( new_AGEMA_signal_16699 ), .Q ( new_AGEMA_signal_16700 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5204 ( .C ( clk ), .D ( new_AGEMA_signal_16703 ), .Q ( new_AGEMA_signal_16704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5208 ( .C ( clk ), .D ( new_AGEMA_signal_16707 ), .Q ( new_AGEMA_signal_16708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5212 ( .C ( clk ), .D ( new_AGEMA_signal_16711 ), .Q ( new_AGEMA_signal_16712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5228 ( .C ( clk ), .D ( new_AGEMA_signal_16727 ), .Q ( new_AGEMA_signal_16728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5236 ( .C ( clk ), .D ( new_AGEMA_signal_16735 ), .Q ( new_AGEMA_signal_16736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5244 ( .C ( clk ), .D ( new_AGEMA_signal_16743 ), .Q ( new_AGEMA_signal_16744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5252 ( .C ( clk ), .D ( new_AGEMA_signal_16751 ), .Q ( new_AGEMA_signal_16752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5260 ( .C ( clk ), .D ( new_AGEMA_signal_16759 ), .Q ( new_AGEMA_signal_16760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5268 ( .C ( clk ), .D ( new_AGEMA_signal_16767 ), .Q ( new_AGEMA_signal_16768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5276 ( .C ( clk ), .D ( new_AGEMA_signal_16775 ), .Q ( new_AGEMA_signal_16776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5284 ( .C ( clk ), .D ( new_AGEMA_signal_16783 ), .Q ( new_AGEMA_signal_16784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5290 ( .C ( clk ), .D ( new_AGEMA_signal_16789 ), .Q ( new_AGEMA_signal_16790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5296 ( .C ( clk ), .D ( new_AGEMA_signal_16795 ), .Q ( new_AGEMA_signal_16796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5302 ( .C ( clk ), .D ( new_AGEMA_signal_16801 ), .Q ( new_AGEMA_signal_16802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5308 ( .C ( clk ), .D ( new_AGEMA_signal_16807 ), .Q ( new_AGEMA_signal_16808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5312 ( .C ( clk ), .D ( new_AGEMA_signal_16811 ), .Q ( new_AGEMA_signal_16812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5316 ( .C ( clk ), .D ( new_AGEMA_signal_16815 ), .Q ( new_AGEMA_signal_16816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5320 ( .C ( clk ), .D ( new_AGEMA_signal_16819 ), .Q ( new_AGEMA_signal_16820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5324 ( .C ( clk ), .D ( new_AGEMA_signal_16823 ), .Q ( new_AGEMA_signal_16824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5332 ( .C ( clk ), .D ( new_AGEMA_signal_16831 ), .Q ( new_AGEMA_signal_16832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5340 ( .C ( clk ), .D ( new_AGEMA_signal_16839 ), .Q ( new_AGEMA_signal_16840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5348 ( .C ( clk ), .D ( new_AGEMA_signal_16847 ), .Q ( new_AGEMA_signal_16848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5356 ( .C ( clk ), .D ( new_AGEMA_signal_16855 ), .Q ( new_AGEMA_signal_16856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5368 ( .C ( clk ), .D ( new_AGEMA_signal_16867 ), .Q ( new_AGEMA_signal_16868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5374 ( .C ( clk ), .D ( new_AGEMA_signal_16873 ), .Q ( new_AGEMA_signal_16874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5380 ( .C ( clk ), .D ( new_AGEMA_signal_16879 ), .Q ( new_AGEMA_signal_16880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5386 ( .C ( clk ), .D ( new_AGEMA_signal_16885 ), .Q ( new_AGEMA_signal_16886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5392 ( .C ( clk ), .D ( new_AGEMA_signal_16891 ), .Q ( new_AGEMA_signal_16892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5398 ( .C ( clk ), .D ( new_AGEMA_signal_16897 ), .Q ( new_AGEMA_signal_16898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5404 ( .C ( clk ), .D ( new_AGEMA_signal_16903 ), .Q ( new_AGEMA_signal_16904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5410 ( .C ( clk ), .D ( new_AGEMA_signal_16909 ), .Q ( new_AGEMA_signal_16910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5416 ( .C ( clk ), .D ( new_AGEMA_signal_16915 ), .Q ( new_AGEMA_signal_16916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5422 ( .C ( clk ), .D ( new_AGEMA_signal_16921 ), .Q ( new_AGEMA_signal_16922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5428 ( .C ( clk ), .D ( new_AGEMA_signal_16927 ), .Q ( new_AGEMA_signal_16928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5434 ( .C ( clk ), .D ( new_AGEMA_signal_16933 ), .Q ( new_AGEMA_signal_16934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5458 ( .C ( clk ), .D ( new_AGEMA_signal_16957 ), .Q ( new_AGEMA_signal_16958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5466 ( .C ( clk ), .D ( new_AGEMA_signal_16965 ), .Q ( new_AGEMA_signal_16966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5474 ( .C ( clk ), .D ( new_AGEMA_signal_16973 ), .Q ( new_AGEMA_signal_16974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5482 ( .C ( clk ), .D ( new_AGEMA_signal_16981 ), .Q ( new_AGEMA_signal_16982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5488 ( .C ( clk ), .D ( new_AGEMA_signal_16987 ), .Q ( new_AGEMA_signal_16988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5494 ( .C ( clk ), .D ( new_AGEMA_signal_16993 ), .Q ( new_AGEMA_signal_16994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5500 ( .C ( clk ), .D ( new_AGEMA_signal_16999 ), .Q ( new_AGEMA_signal_17000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5506 ( .C ( clk ), .D ( new_AGEMA_signal_17005 ), .Q ( new_AGEMA_signal_17006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5530 ( .C ( clk ), .D ( new_AGEMA_signal_17029 ), .Q ( new_AGEMA_signal_17030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5538 ( .C ( clk ), .D ( new_AGEMA_signal_17037 ), .Q ( new_AGEMA_signal_17038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5546 ( .C ( clk ), .D ( new_AGEMA_signal_17045 ), .Q ( new_AGEMA_signal_17046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5554 ( .C ( clk ), .D ( new_AGEMA_signal_17053 ), .Q ( new_AGEMA_signal_17054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5562 ( .C ( clk ), .D ( new_AGEMA_signal_17061 ), .Q ( new_AGEMA_signal_17062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5570 ( .C ( clk ), .D ( new_AGEMA_signal_17069 ), .Q ( new_AGEMA_signal_17070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5578 ( .C ( clk ), .D ( new_AGEMA_signal_17077 ), .Q ( new_AGEMA_signal_17078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5586 ( .C ( clk ), .D ( new_AGEMA_signal_17085 ), .Q ( new_AGEMA_signal_17086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5596 ( .C ( clk ), .D ( new_AGEMA_signal_17095 ), .Q ( new_AGEMA_signal_17096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5606 ( .C ( clk ), .D ( new_AGEMA_signal_17105 ), .Q ( new_AGEMA_signal_17106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5616 ( .C ( clk ), .D ( new_AGEMA_signal_17115 ), .Q ( new_AGEMA_signal_17116 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5626 ( .C ( clk ), .D ( new_AGEMA_signal_17125 ), .Q ( new_AGEMA_signal_17126 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5634 ( .C ( clk ), .D ( new_AGEMA_signal_17133 ), .Q ( new_AGEMA_signal_17134 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5642 ( .C ( clk ), .D ( new_AGEMA_signal_17141 ), .Q ( new_AGEMA_signal_17142 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5650 ( .C ( clk ), .D ( new_AGEMA_signal_17149 ), .Q ( new_AGEMA_signal_17150 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5658 ( .C ( clk ), .D ( new_AGEMA_signal_17157 ), .Q ( new_AGEMA_signal_17158 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5664 ( .C ( clk ), .D ( new_AGEMA_signal_17163 ), .Q ( new_AGEMA_signal_17164 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5670 ( .C ( clk ), .D ( new_AGEMA_signal_17169 ), .Q ( new_AGEMA_signal_17170 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5676 ( .C ( clk ), .D ( new_AGEMA_signal_17175 ), .Q ( new_AGEMA_signal_17176 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5682 ( .C ( clk ), .D ( new_AGEMA_signal_17181 ), .Q ( new_AGEMA_signal_17182 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5704 ( .C ( clk ), .D ( new_AGEMA_signal_17203 ), .Q ( new_AGEMA_signal_17204 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5710 ( .C ( clk ), .D ( new_AGEMA_signal_17209 ), .Q ( new_AGEMA_signal_17210 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5716 ( .C ( clk ), .D ( new_AGEMA_signal_17215 ), .Q ( new_AGEMA_signal_17216 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5722 ( .C ( clk ), .D ( new_AGEMA_signal_17221 ), .Q ( new_AGEMA_signal_17222 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5730 ( .C ( clk ), .D ( new_AGEMA_signal_17229 ), .Q ( new_AGEMA_signal_17230 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5738 ( .C ( clk ), .D ( new_AGEMA_signal_17237 ), .Q ( new_AGEMA_signal_17238 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5746 ( .C ( clk ), .D ( new_AGEMA_signal_17245 ), .Q ( new_AGEMA_signal_17246 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5754 ( .C ( clk ), .D ( new_AGEMA_signal_17253 ), .Q ( new_AGEMA_signal_17254 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5760 ( .C ( clk ), .D ( new_AGEMA_signal_17259 ), .Q ( new_AGEMA_signal_17260 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5766 ( .C ( clk ), .D ( new_AGEMA_signal_17265 ), .Q ( new_AGEMA_signal_17266 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5772 ( .C ( clk ), .D ( new_AGEMA_signal_17271 ), .Q ( new_AGEMA_signal_17272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5778 ( .C ( clk ), .D ( new_AGEMA_signal_17277 ), .Q ( new_AGEMA_signal_17278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5794 ( .C ( clk ), .D ( new_AGEMA_signal_17293 ), .Q ( new_AGEMA_signal_17294 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5802 ( .C ( clk ), .D ( new_AGEMA_signal_17301 ), .Q ( new_AGEMA_signal_17302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5810 ( .C ( clk ), .D ( new_AGEMA_signal_17309 ), .Q ( new_AGEMA_signal_17310 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5818 ( .C ( clk ), .D ( new_AGEMA_signal_17317 ), .Q ( new_AGEMA_signal_17318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5840 ( .C ( clk ), .D ( new_AGEMA_signal_17339 ), .Q ( new_AGEMA_signal_17340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5846 ( .C ( clk ), .D ( new_AGEMA_signal_17345 ), .Q ( new_AGEMA_signal_17346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5852 ( .C ( clk ), .D ( new_AGEMA_signal_17351 ), .Q ( new_AGEMA_signal_17352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5858 ( .C ( clk ), .D ( new_AGEMA_signal_17357 ), .Q ( new_AGEMA_signal_17358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5864 ( .C ( clk ), .D ( new_AGEMA_signal_17363 ), .Q ( new_AGEMA_signal_17364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5870 ( .C ( clk ), .D ( new_AGEMA_signal_17369 ), .Q ( new_AGEMA_signal_17370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5876 ( .C ( clk ), .D ( new_AGEMA_signal_17375 ), .Q ( new_AGEMA_signal_17376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5882 ( .C ( clk ), .D ( new_AGEMA_signal_17381 ), .Q ( new_AGEMA_signal_17382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5970 ( .C ( clk ), .D ( new_AGEMA_signal_17469 ), .Q ( new_AGEMA_signal_17470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5980 ( .C ( clk ), .D ( new_AGEMA_signal_17479 ), .Q ( new_AGEMA_signal_17480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5990 ( .C ( clk ), .D ( new_AGEMA_signal_17489 ), .Q ( new_AGEMA_signal_17490 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6000 ( .C ( clk ), .D ( new_AGEMA_signal_17499 ), .Q ( new_AGEMA_signal_17500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6088 ( .C ( clk ), .D ( new_AGEMA_signal_17587 ), .Q ( new_AGEMA_signal_17588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6096 ( .C ( clk ), .D ( new_AGEMA_signal_17595 ), .Q ( new_AGEMA_signal_17596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6104 ( .C ( clk ), .D ( new_AGEMA_signal_17603 ), .Q ( new_AGEMA_signal_17604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6112 ( .C ( clk ), .D ( new_AGEMA_signal_17611 ), .Q ( new_AGEMA_signal_17612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6144 ( .C ( clk ), .D ( new_AGEMA_signal_17643 ), .Q ( new_AGEMA_signal_17644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6152 ( .C ( clk ), .D ( new_AGEMA_signal_17651 ), .Q ( new_AGEMA_signal_17652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6160 ( .C ( clk ), .D ( new_AGEMA_signal_17659 ), .Q ( new_AGEMA_signal_17660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6168 ( .C ( clk ), .D ( new_AGEMA_signal_17667 ), .Q ( new_AGEMA_signal_17668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6176 ( .C ( clk ), .D ( new_AGEMA_signal_17675 ), .Q ( new_AGEMA_signal_17676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6184 ( .C ( clk ), .D ( new_AGEMA_signal_17683 ), .Q ( new_AGEMA_signal_17684 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6192 ( .C ( clk ), .D ( new_AGEMA_signal_17691 ), .Q ( new_AGEMA_signal_17692 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6200 ( .C ( clk ), .D ( new_AGEMA_signal_17699 ), .Q ( new_AGEMA_signal_17700 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6248 ( .C ( clk ), .D ( new_AGEMA_signal_17747 ), .Q ( new_AGEMA_signal_17748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6256 ( .C ( clk ), .D ( new_AGEMA_signal_17755 ), .Q ( new_AGEMA_signal_17756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6264 ( .C ( clk ), .D ( new_AGEMA_signal_17763 ), .Q ( new_AGEMA_signal_17764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6272 ( .C ( clk ), .D ( new_AGEMA_signal_17771 ), .Q ( new_AGEMA_signal_17772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6330 ( .C ( clk ), .D ( new_AGEMA_signal_17829 ), .Q ( new_AGEMA_signal_17830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6342 ( .C ( clk ), .D ( new_AGEMA_signal_17841 ), .Q ( new_AGEMA_signal_17842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6354 ( .C ( clk ), .D ( new_AGEMA_signal_17853 ), .Q ( new_AGEMA_signal_17854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6366 ( .C ( clk ), .D ( new_AGEMA_signal_17865 ), .Q ( new_AGEMA_signal_17866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6380 ( .C ( clk ), .D ( new_AGEMA_signal_17879 ), .Q ( new_AGEMA_signal_17880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6394 ( .C ( clk ), .D ( new_AGEMA_signal_17893 ), .Q ( new_AGEMA_signal_17894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6408 ( .C ( clk ), .D ( new_AGEMA_signal_17907 ), .Q ( new_AGEMA_signal_17908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6422 ( .C ( clk ), .D ( new_AGEMA_signal_17921 ), .Q ( new_AGEMA_signal_17922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6468 ( .C ( clk ), .D ( new_AGEMA_signal_17967 ), .Q ( new_AGEMA_signal_17968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6482 ( .C ( clk ), .D ( new_AGEMA_signal_17981 ), .Q ( new_AGEMA_signal_17982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6496 ( .C ( clk ), .D ( new_AGEMA_signal_17995 ), .Q ( new_AGEMA_signal_17996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6510 ( .C ( clk ), .D ( new_AGEMA_signal_18009 ), .Q ( new_AGEMA_signal_18010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6612 ( .C ( clk ), .D ( new_AGEMA_signal_18111 ), .Q ( new_AGEMA_signal_18112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6628 ( .C ( clk ), .D ( new_AGEMA_signal_18127 ), .Q ( new_AGEMA_signal_18128 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6644 ( .C ( clk ), .D ( new_AGEMA_signal_18143 ), .Q ( new_AGEMA_signal_18144 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6660 ( .C ( clk ), .D ( new_AGEMA_signal_18159 ), .Q ( new_AGEMA_signal_18160 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6700 ( .C ( clk ), .D ( new_AGEMA_signal_18199 ), .Q ( new_AGEMA_signal_18200 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6716 ( .C ( clk ), .D ( new_AGEMA_signal_18215 ), .Q ( new_AGEMA_signal_18216 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6732 ( .C ( clk ), .D ( new_AGEMA_signal_18231 ), .Q ( new_AGEMA_signal_18232 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6748 ( .C ( clk ), .D ( new_AGEMA_signal_18247 ), .Q ( new_AGEMA_signal_18248 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6898 ( .C ( clk ), .D ( new_AGEMA_signal_18397 ), .Q ( new_AGEMA_signal_18398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6914 ( .C ( clk ), .D ( new_AGEMA_signal_18413 ), .Q ( new_AGEMA_signal_18414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6930 ( .C ( clk ), .D ( new_AGEMA_signal_18429 ), .Q ( new_AGEMA_signal_18430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6946 ( .C ( clk ), .D ( new_AGEMA_signal_18445 ), .Q ( new_AGEMA_signal_18446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7004 ( .C ( clk ), .D ( new_AGEMA_signal_18503 ), .Q ( new_AGEMA_signal_18504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7022 ( .C ( clk ), .D ( new_AGEMA_signal_18521 ), .Q ( new_AGEMA_signal_18522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7040 ( .C ( clk ), .D ( new_AGEMA_signal_18539 ), .Q ( new_AGEMA_signal_18540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7058 ( .C ( clk ), .D ( new_AGEMA_signal_18557 ), .Q ( new_AGEMA_signal_18558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7204 ( .C ( clk ), .D ( new_AGEMA_signal_18703 ), .Q ( new_AGEMA_signal_18704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7224 ( .C ( clk ), .D ( new_AGEMA_signal_18723 ), .Q ( new_AGEMA_signal_18724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7244 ( .C ( clk ), .D ( new_AGEMA_signal_18743 ), .Q ( new_AGEMA_signal_18744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7264 ( .C ( clk ), .D ( new_AGEMA_signal_18763 ), .Q ( new_AGEMA_signal_18764 ) ) ;

    /* cells in depth 13 */
    buf_clk new_AGEMA_reg_buffer_4731 ( .C ( clk ), .D ( new_AGEMA_signal_16230 ), .Q ( new_AGEMA_signal_16231 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4737 ( .C ( clk ), .D ( new_AGEMA_signal_16236 ), .Q ( new_AGEMA_signal_16237 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4743 ( .C ( clk ), .D ( new_AGEMA_signal_16242 ), .Q ( new_AGEMA_signal_16243 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4749 ( .C ( clk ), .D ( new_AGEMA_signal_16248 ), .Q ( new_AGEMA_signal_16249 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4751 ( .C ( clk ), .D ( new_AGEMA_signal_16174 ), .Q ( new_AGEMA_signal_16251 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4753 ( .C ( clk ), .D ( new_AGEMA_signal_16178 ), .Q ( new_AGEMA_signal_16253 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4755 ( .C ( clk ), .D ( new_AGEMA_signal_16182 ), .Q ( new_AGEMA_signal_16255 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4757 ( .C ( clk ), .D ( new_AGEMA_signal_16186 ), .Q ( new_AGEMA_signal_16257 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4761 ( .C ( clk ), .D ( new_AGEMA_signal_16260 ), .Q ( new_AGEMA_signal_16261 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4765 ( .C ( clk ), .D ( new_AGEMA_signal_16264 ), .Q ( new_AGEMA_signal_16265 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4769 ( .C ( clk ), .D ( new_AGEMA_signal_16268 ), .Q ( new_AGEMA_signal_16269 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4773 ( .C ( clk ), .D ( new_AGEMA_signal_16272 ), .Q ( new_AGEMA_signal_16273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4781 ( .C ( clk ), .D ( new_AGEMA_signal_16280 ), .Q ( new_AGEMA_signal_16281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4789 ( .C ( clk ), .D ( new_AGEMA_signal_16288 ), .Q ( new_AGEMA_signal_16289 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4797 ( .C ( clk ), .D ( new_AGEMA_signal_16296 ), .Q ( new_AGEMA_signal_16297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4805 ( .C ( clk ), .D ( new_AGEMA_signal_16304 ), .Q ( new_AGEMA_signal_16305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4813 ( .C ( clk ), .D ( new_AGEMA_signal_16312 ), .Q ( new_AGEMA_signal_16313 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4821 ( .C ( clk ), .D ( new_AGEMA_signal_16320 ), .Q ( new_AGEMA_signal_16321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4829 ( .C ( clk ), .D ( new_AGEMA_signal_16328 ), .Q ( new_AGEMA_signal_16329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4837 ( .C ( clk ), .D ( new_AGEMA_signal_16336 ), .Q ( new_AGEMA_signal_16337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4845 ( .C ( clk ), .D ( new_AGEMA_signal_16344 ), .Q ( new_AGEMA_signal_16345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4853 ( .C ( clk ), .D ( new_AGEMA_signal_16352 ), .Q ( new_AGEMA_signal_16353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4861 ( .C ( clk ), .D ( new_AGEMA_signal_16360 ), .Q ( new_AGEMA_signal_16361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4869 ( .C ( clk ), .D ( new_AGEMA_signal_16368 ), .Q ( new_AGEMA_signal_16369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4877 ( .C ( clk ), .D ( new_AGEMA_signal_16376 ), .Q ( new_AGEMA_signal_16377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4885 ( .C ( clk ), .D ( new_AGEMA_signal_16384 ), .Q ( new_AGEMA_signal_16385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4893 ( .C ( clk ), .D ( new_AGEMA_signal_16392 ), .Q ( new_AGEMA_signal_16393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4901 ( .C ( clk ), .D ( new_AGEMA_signal_16400 ), .Q ( new_AGEMA_signal_16401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4907 ( .C ( clk ), .D ( new_AGEMA_signal_16406 ), .Q ( new_AGEMA_signal_16407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4913 ( .C ( clk ), .D ( new_AGEMA_signal_16412 ), .Q ( new_AGEMA_signal_16413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4919 ( .C ( clk ), .D ( new_AGEMA_signal_16418 ), .Q ( new_AGEMA_signal_16419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4925 ( .C ( clk ), .D ( new_AGEMA_signal_16424 ), .Q ( new_AGEMA_signal_16425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4935 ( .C ( clk ), .D ( new_AGEMA_signal_16434 ), .Q ( new_AGEMA_signal_16435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4945 ( .C ( clk ), .D ( new_AGEMA_signal_16444 ), .Q ( new_AGEMA_signal_16445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4955 ( .C ( clk ), .D ( new_AGEMA_signal_16454 ), .Q ( new_AGEMA_signal_16455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4965 ( .C ( clk ), .D ( new_AGEMA_signal_16464 ), .Q ( new_AGEMA_signal_16465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4973 ( .C ( clk ), .D ( new_AGEMA_signal_16472 ), .Q ( new_AGEMA_signal_16473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4981 ( .C ( clk ), .D ( new_AGEMA_signal_16480 ), .Q ( new_AGEMA_signal_16481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4989 ( .C ( clk ), .D ( new_AGEMA_signal_16488 ), .Q ( new_AGEMA_signal_16489 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4997 ( .C ( clk ), .D ( new_AGEMA_signal_16496 ), .Q ( new_AGEMA_signal_16497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5005 ( .C ( clk ), .D ( new_AGEMA_signal_16504 ), .Q ( new_AGEMA_signal_16505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5013 ( .C ( clk ), .D ( new_AGEMA_signal_16512 ), .Q ( new_AGEMA_signal_16513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5021 ( .C ( clk ), .D ( new_AGEMA_signal_16520 ), .Q ( new_AGEMA_signal_16521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5029 ( .C ( clk ), .D ( new_AGEMA_signal_16528 ), .Q ( new_AGEMA_signal_16529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5037 ( .C ( clk ), .D ( new_AGEMA_signal_16536 ), .Q ( new_AGEMA_signal_16537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5045 ( .C ( clk ), .D ( new_AGEMA_signal_16544 ), .Q ( new_AGEMA_signal_16545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5053 ( .C ( clk ), .D ( new_AGEMA_signal_16552 ), .Q ( new_AGEMA_signal_16553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5061 ( .C ( clk ), .D ( new_AGEMA_signal_16560 ), .Q ( new_AGEMA_signal_16561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5063 ( .C ( clk ), .D ( new_AGEMA_signal_15620 ), .Q ( new_AGEMA_signal_16563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5065 ( .C ( clk ), .D ( new_AGEMA_signal_15622 ), .Q ( new_AGEMA_signal_16565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5067 ( .C ( clk ), .D ( new_AGEMA_signal_15624 ), .Q ( new_AGEMA_signal_16567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5069 ( .C ( clk ), .D ( new_AGEMA_signal_15626 ), .Q ( new_AGEMA_signal_16569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5073 ( .C ( clk ), .D ( new_AGEMA_signal_16572 ), .Q ( new_AGEMA_signal_16573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5077 ( .C ( clk ), .D ( new_AGEMA_signal_16576 ), .Q ( new_AGEMA_signal_16577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5081 ( .C ( clk ), .D ( new_AGEMA_signal_16580 ), .Q ( new_AGEMA_signal_16581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5085 ( .C ( clk ), .D ( new_AGEMA_signal_16584 ), .Q ( new_AGEMA_signal_16585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5091 ( .C ( clk ), .D ( new_AGEMA_signal_16590 ), .Q ( new_AGEMA_signal_16591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5097 ( .C ( clk ), .D ( new_AGEMA_signal_16596 ), .Q ( new_AGEMA_signal_16597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5103 ( .C ( clk ), .D ( new_AGEMA_signal_16602 ), .Q ( new_AGEMA_signal_16603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5109 ( .C ( clk ), .D ( new_AGEMA_signal_16608 ), .Q ( new_AGEMA_signal_16609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5113 ( .C ( clk ), .D ( new_AGEMA_signal_16612 ), .Q ( new_AGEMA_signal_16613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5117 ( .C ( clk ), .D ( new_AGEMA_signal_16616 ), .Q ( new_AGEMA_signal_16617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5121 ( .C ( clk ), .D ( new_AGEMA_signal_16620 ), .Q ( new_AGEMA_signal_16621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5125 ( .C ( clk ), .D ( new_AGEMA_signal_16624 ), .Q ( new_AGEMA_signal_16625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5135 ( .C ( clk ), .D ( new_AGEMA_signal_16634 ), .Q ( new_AGEMA_signal_16635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5145 ( .C ( clk ), .D ( new_AGEMA_signal_16644 ), .Q ( new_AGEMA_signal_16645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5155 ( .C ( clk ), .D ( new_AGEMA_signal_16654 ), .Q ( new_AGEMA_signal_16655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5165 ( .C ( clk ), .D ( new_AGEMA_signal_16664 ), .Q ( new_AGEMA_signal_16665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5173 ( .C ( clk ), .D ( new_AGEMA_signal_16672 ), .Q ( new_AGEMA_signal_16673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5181 ( .C ( clk ), .D ( new_AGEMA_signal_16680 ), .Q ( new_AGEMA_signal_16681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5189 ( .C ( clk ), .D ( new_AGEMA_signal_16688 ), .Q ( new_AGEMA_signal_16689 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5197 ( .C ( clk ), .D ( new_AGEMA_signal_16696 ), .Q ( new_AGEMA_signal_16697 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5201 ( .C ( clk ), .D ( new_AGEMA_signal_16700 ), .Q ( new_AGEMA_signal_16701 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5205 ( .C ( clk ), .D ( new_AGEMA_signal_16704 ), .Q ( new_AGEMA_signal_16705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5209 ( .C ( clk ), .D ( new_AGEMA_signal_16708 ), .Q ( new_AGEMA_signal_16709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5213 ( .C ( clk ), .D ( new_AGEMA_signal_16712 ), .Q ( new_AGEMA_signal_16713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5215 ( .C ( clk ), .D ( n2509 ), .Q ( new_AGEMA_signal_16715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5217 ( .C ( clk ), .D ( new_AGEMA_signal_3387 ), .Q ( new_AGEMA_signal_16717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5219 ( .C ( clk ), .D ( new_AGEMA_signal_3388 ), .Q ( new_AGEMA_signal_16719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5221 ( .C ( clk ), .D ( new_AGEMA_signal_3389 ), .Q ( new_AGEMA_signal_16721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5229 ( .C ( clk ), .D ( new_AGEMA_signal_16728 ), .Q ( new_AGEMA_signal_16729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5237 ( .C ( clk ), .D ( new_AGEMA_signal_16736 ), .Q ( new_AGEMA_signal_16737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5245 ( .C ( clk ), .D ( new_AGEMA_signal_16744 ), .Q ( new_AGEMA_signal_16745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5253 ( .C ( clk ), .D ( new_AGEMA_signal_16752 ), .Q ( new_AGEMA_signal_16753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5261 ( .C ( clk ), .D ( new_AGEMA_signal_16760 ), .Q ( new_AGEMA_signal_16761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5269 ( .C ( clk ), .D ( new_AGEMA_signal_16768 ), .Q ( new_AGEMA_signal_16769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5277 ( .C ( clk ), .D ( new_AGEMA_signal_16776 ), .Q ( new_AGEMA_signal_16777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5285 ( .C ( clk ), .D ( new_AGEMA_signal_16784 ), .Q ( new_AGEMA_signal_16785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5291 ( .C ( clk ), .D ( new_AGEMA_signal_16790 ), .Q ( new_AGEMA_signal_16791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5297 ( .C ( clk ), .D ( new_AGEMA_signal_16796 ), .Q ( new_AGEMA_signal_16797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5303 ( .C ( clk ), .D ( new_AGEMA_signal_16802 ), .Q ( new_AGEMA_signal_16803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5309 ( .C ( clk ), .D ( new_AGEMA_signal_16808 ), .Q ( new_AGEMA_signal_16809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5313 ( .C ( clk ), .D ( new_AGEMA_signal_16812 ), .Q ( new_AGEMA_signal_16813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5317 ( .C ( clk ), .D ( new_AGEMA_signal_16816 ), .Q ( new_AGEMA_signal_16817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5321 ( .C ( clk ), .D ( new_AGEMA_signal_16820 ), .Q ( new_AGEMA_signal_16821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5325 ( .C ( clk ), .D ( new_AGEMA_signal_16824 ), .Q ( new_AGEMA_signal_16825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5333 ( .C ( clk ), .D ( new_AGEMA_signal_16832 ), .Q ( new_AGEMA_signal_16833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5341 ( .C ( clk ), .D ( new_AGEMA_signal_16840 ), .Q ( new_AGEMA_signal_16841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5349 ( .C ( clk ), .D ( new_AGEMA_signal_16848 ), .Q ( new_AGEMA_signal_16849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5357 ( .C ( clk ), .D ( new_AGEMA_signal_16856 ), .Q ( new_AGEMA_signal_16857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5359 ( .C ( clk ), .D ( n2802 ), .Q ( new_AGEMA_signal_16859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5361 ( .C ( clk ), .D ( new_AGEMA_signal_3285 ), .Q ( new_AGEMA_signal_16861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5363 ( .C ( clk ), .D ( new_AGEMA_signal_3286 ), .Q ( new_AGEMA_signal_16863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5365 ( .C ( clk ), .D ( new_AGEMA_signal_3287 ), .Q ( new_AGEMA_signal_16865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5369 ( .C ( clk ), .D ( new_AGEMA_signal_16868 ), .Q ( new_AGEMA_signal_16869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5375 ( .C ( clk ), .D ( new_AGEMA_signal_16874 ), .Q ( new_AGEMA_signal_16875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5381 ( .C ( clk ), .D ( new_AGEMA_signal_16880 ), .Q ( new_AGEMA_signal_16881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5387 ( .C ( clk ), .D ( new_AGEMA_signal_16886 ), .Q ( new_AGEMA_signal_16887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5393 ( .C ( clk ), .D ( new_AGEMA_signal_16892 ), .Q ( new_AGEMA_signal_16893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5399 ( .C ( clk ), .D ( new_AGEMA_signal_16898 ), .Q ( new_AGEMA_signal_16899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5405 ( .C ( clk ), .D ( new_AGEMA_signal_16904 ), .Q ( new_AGEMA_signal_16905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5411 ( .C ( clk ), .D ( new_AGEMA_signal_16910 ), .Q ( new_AGEMA_signal_16911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5417 ( .C ( clk ), .D ( new_AGEMA_signal_16916 ), .Q ( new_AGEMA_signal_16917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5423 ( .C ( clk ), .D ( new_AGEMA_signal_16922 ), .Q ( new_AGEMA_signal_16923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5429 ( .C ( clk ), .D ( new_AGEMA_signal_16928 ), .Q ( new_AGEMA_signal_16929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5435 ( .C ( clk ), .D ( new_AGEMA_signal_16934 ), .Q ( new_AGEMA_signal_16935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5439 ( .C ( clk ), .D ( new_AGEMA_signal_16220 ), .Q ( new_AGEMA_signal_16939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5443 ( .C ( clk ), .D ( new_AGEMA_signal_16222 ), .Q ( new_AGEMA_signal_16943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5447 ( .C ( clk ), .D ( new_AGEMA_signal_16224 ), .Q ( new_AGEMA_signal_16947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5451 ( .C ( clk ), .D ( new_AGEMA_signal_16226 ), .Q ( new_AGEMA_signal_16951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5459 ( .C ( clk ), .D ( new_AGEMA_signal_16958 ), .Q ( new_AGEMA_signal_16959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5467 ( .C ( clk ), .D ( new_AGEMA_signal_16966 ), .Q ( new_AGEMA_signal_16967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5475 ( .C ( clk ), .D ( new_AGEMA_signal_16974 ), .Q ( new_AGEMA_signal_16975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5483 ( .C ( clk ), .D ( new_AGEMA_signal_16982 ), .Q ( new_AGEMA_signal_16983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5489 ( .C ( clk ), .D ( new_AGEMA_signal_16988 ), .Q ( new_AGEMA_signal_16989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5495 ( .C ( clk ), .D ( new_AGEMA_signal_16994 ), .Q ( new_AGEMA_signal_16995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5501 ( .C ( clk ), .D ( new_AGEMA_signal_17000 ), .Q ( new_AGEMA_signal_17001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5507 ( .C ( clk ), .D ( new_AGEMA_signal_17006 ), .Q ( new_AGEMA_signal_17007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5511 ( .C ( clk ), .D ( n2072 ), .Q ( new_AGEMA_signal_17011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5515 ( .C ( clk ), .D ( new_AGEMA_signal_3144 ), .Q ( new_AGEMA_signal_17015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5519 ( .C ( clk ), .D ( new_AGEMA_signal_3145 ), .Q ( new_AGEMA_signal_17019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5523 ( .C ( clk ), .D ( new_AGEMA_signal_3146 ), .Q ( new_AGEMA_signal_17023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5531 ( .C ( clk ), .D ( new_AGEMA_signal_17030 ), .Q ( new_AGEMA_signal_17031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5539 ( .C ( clk ), .D ( new_AGEMA_signal_17038 ), .Q ( new_AGEMA_signal_17039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5547 ( .C ( clk ), .D ( new_AGEMA_signal_17046 ), .Q ( new_AGEMA_signal_17047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5555 ( .C ( clk ), .D ( new_AGEMA_signal_17054 ), .Q ( new_AGEMA_signal_17055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5563 ( .C ( clk ), .D ( new_AGEMA_signal_17062 ), .Q ( new_AGEMA_signal_17063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5571 ( .C ( clk ), .D ( new_AGEMA_signal_17070 ), .Q ( new_AGEMA_signal_17071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5579 ( .C ( clk ), .D ( new_AGEMA_signal_17078 ), .Q ( new_AGEMA_signal_17079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5587 ( .C ( clk ), .D ( new_AGEMA_signal_17086 ), .Q ( new_AGEMA_signal_17087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5597 ( .C ( clk ), .D ( new_AGEMA_signal_17096 ), .Q ( new_AGEMA_signal_17097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5607 ( .C ( clk ), .D ( new_AGEMA_signal_17106 ), .Q ( new_AGEMA_signal_17107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5617 ( .C ( clk ), .D ( new_AGEMA_signal_17116 ), .Q ( new_AGEMA_signal_17117 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5627 ( .C ( clk ), .D ( new_AGEMA_signal_17126 ), .Q ( new_AGEMA_signal_17127 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5635 ( .C ( clk ), .D ( new_AGEMA_signal_17134 ), .Q ( new_AGEMA_signal_17135 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5643 ( .C ( clk ), .D ( new_AGEMA_signal_17142 ), .Q ( new_AGEMA_signal_17143 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5651 ( .C ( clk ), .D ( new_AGEMA_signal_17150 ), .Q ( new_AGEMA_signal_17151 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5659 ( .C ( clk ), .D ( new_AGEMA_signal_17158 ), .Q ( new_AGEMA_signal_17159 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5665 ( .C ( clk ), .D ( new_AGEMA_signal_17164 ), .Q ( new_AGEMA_signal_17165 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5671 ( .C ( clk ), .D ( new_AGEMA_signal_17170 ), .Q ( new_AGEMA_signal_17171 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5677 ( .C ( clk ), .D ( new_AGEMA_signal_17176 ), .Q ( new_AGEMA_signal_17177 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5683 ( .C ( clk ), .D ( new_AGEMA_signal_17182 ), .Q ( new_AGEMA_signal_17183 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5687 ( .C ( clk ), .D ( n2276 ), .Q ( new_AGEMA_signal_17187 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5691 ( .C ( clk ), .D ( new_AGEMA_signal_3192 ), .Q ( new_AGEMA_signal_17191 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5695 ( .C ( clk ), .D ( new_AGEMA_signal_3193 ), .Q ( new_AGEMA_signal_17195 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5699 ( .C ( clk ), .D ( new_AGEMA_signal_3194 ), .Q ( new_AGEMA_signal_17199 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5705 ( .C ( clk ), .D ( new_AGEMA_signal_17204 ), .Q ( new_AGEMA_signal_17205 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5711 ( .C ( clk ), .D ( new_AGEMA_signal_17210 ), .Q ( new_AGEMA_signal_17211 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5717 ( .C ( clk ), .D ( new_AGEMA_signal_17216 ), .Q ( new_AGEMA_signal_17217 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5723 ( .C ( clk ), .D ( new_AGEMA_signal_17222 ), .Q ( new_AGEMA_signal_17223 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5731 ( .C ( clk ), .D ( new_AGEMA_signal_17230 ), .Q ( new_AGEMA_signal_17231 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5739 ( .C ( clk ), .D ( new_AGEMA_signal_17238 ), .Q ( new_AGEMA_signal_17239 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5747 ( .C ( clk ), .D ( new_AGEMA_signal_17246 ), .Q ( new_AGEMA_signal_17247 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5755 ( .C ( clk ), .D ( new_AGEMA_signal_17254 ), .Q ( new_AGEMA_signal_17255 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5761 ( .C ( clk ), .D ( new_AGEMA_signal_17260 ), .Q ( new_AGEMA_signal_17261 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5767 ( .C ( clk ), .D ( new_AGEMA_signal_17266 ), .Q ( new_AGEMA_signal_17267 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5773 ( .C ( clk ), .D ( new_AGEMA_signal_17272 ), .Q ( new_AGEMA_signal_17273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5779 ( .C ( clk ), .D ( new_AGEMA_signal_17278 ), .Q ( new_AGEMA_signal_17279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5795 ( .C ( clk ), .D ( new_AGEMA_signal_17294 ), .Q ( new_AGEMA_signal_17295 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5803 ( .C ( clk ), .D ( new_AGEMA_signal_17302 ), .Q ( new_AGEMA_signal_17303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5811 ( .C ( clk ), .D ( new_AGEMA_signal_17310 ), .Q ( new_AGEMA_signal_17311 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5819 ( .C ( clk ), .D ( new_AGEMA_signal_17318 ), .Q ( new_AGEMA_signal_17319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5823 ( .C ( clk ), .D ( n2622 ), .Q ( new_AGEMA_signal_17323 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5827 ( .C ( clk ), .D ( new_AGEMA_signal_3261 ), .Q ( new_AGEMA_signal_17327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5831 ( .C ( clk ), .D ( new_AGEMA_signal_3262 ), .Q ( new_AGEMA_signal_17331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5835 ( .C ( clk ), .D ( new_AGEMA_signal_3263 ), .Q ( new_AGEMA_signal_17335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5841 ( .C ( clk ), .D ( new_AGEMA_signal_17340 ), .Q ( new_AGEMA_signal_17341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5847 ( .C ( clk ), .D ( new_AGEMA_signal_17346 ), .Q ( new_AGEMA_signal_17347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5853 ( .C ( clk ), .D ( new_AGEMA_signal_17352 ), .Q ( new_AGEMA_signal_17353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5859 ( .C ( clk ), .D ( new_AGEMA_signal_17358 ), .Q ( new_AGEMA_signal_17359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5865 ( .C ( clk ), .D ( new_AGEMA_signal_17364 ), .Q ( new_AGEMA_signal_17365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5871 ( .C ( clk ), .D ( new_AGEMA_signal_17370 ), .Q ( new_AGEMA_signal_17371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5877 ( .C ( clk ), .D ( new_AGEMA_signal_17376 ), .Q ( new_AGEMA_signal_17377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5883 ( .C ( clk ), .D ( new_AGEMA_signal_17382 ), .Q ( new_AGEMA_signal_17383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5887 ( .C ( clk ), .D ( n2804 ), .Q ( new_AGEMA_signal_17387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5891 ( .C ( clk ), .D ( new_AGEMA_signal_3282 ), .Q ( new_AGEMA_signal_17391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5895 ( .C ( clk ), .D ( new_AGEMA_signal_3283 ), .Q ( new_AGEMA_signal_17395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5899 ( .C ( clk ), .D ( new_AGEMA_signal_3284 ), .Q ( new_AGEMA_signal_17399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5903 ( .C ( clk ), .D ( n1990 ), .Q ( new_AGEMA_signal_17403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5909 ( .C ( clk ), .D ( new_AGEMA_signal_2886 ), .Q ( new_AGEMA_signal_17409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5915 ( .C ( clk ), .D ( new_AGEMA_signal_2887 ), .Q ( new_AGEMA_signal_17415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5921 ( .C ( clk ), .D ( new_AGEMA_signal_2888 ), .Q ( new_AGEMA_signal_17421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5943 ( .C ( clk ), .D ( n2078 ), .Q ( new_AGEMA_signal_17443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5949 ( .C ( clk ), .D ( new_AGEMA_signal_3150 ), .Q ( new_AGEMA_signal_17449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5955 ( .C ( clk ), .D ( new_AGEMA_signal_3151 ), .Q ( new_AGEMA_signal_17455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5961 ( .C ( clk ), .D ( new_AGEMA_signal_3152 ), .Q ( new_AGEMA_signal_17461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5971 ( .C ( clk ), .D ( new_AGEMA_signal_17470 ), .Q ( new_AGEMA_signal_17471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5981 ( .C ( clk ), .D ( new_AGEMA_signal_17480 ), .Q ( new_AGEMA_signal_17481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5991 ( .C ( clk ), .D ( new_AGEMA_signal_17490 ), .Q ( new_AGEMA_signal_17491 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6001 ( .C ( clk ), .D ( new_AGEMA_signal_17500 ), .Q ( new_AGEMA_signal_17501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6007 ( .C ( clk ), .D ( n2128 ), .Q ( new_AGEMA_signal_17507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6013 ( .C ( clk ), .D ( new_AGEMA_signal_3321 ), .Q ( new_AGEMA_signal_17513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6019 ( .C ( clk ), .D ( new_AGEMA_signal_3322 ), .Q ( new_AGEMA_signal_17519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6025 ( .C ( clk ), .D ( new_AGEMA_signal_3323 ), .Q ( new_AGEMA_signal_17525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6031 ( .C ( clk ), .D ( n2148 ), .Q ( new_AGEMA_signal_17531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6037 ( .C ( clk ), .D ( new_AGEMA_signal_2940 ), .Q ( new_AGEMA_signal_17537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6043 ( .C ( clk ), .D ( new_AGEMA_signal_2941 ), .Q ( new_AGEMA_signal_17543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6049 ( .C ( clk ), .D ( new_AGEMA_signal_2942 ), .Q ( new_AGEMA_signal_17549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6089 ( .C ( clk ), .D ( new_AGEMA_signal_17588 ), .Q ( new_AGEMA_signal_17589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6097 ( .C ( clk ), .D ( new_AGEMA_signal_17596 ), .Q ( new_AGEMA_signal_17597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6105 ( .C ( clk ), .D ( new_AGEMA_signal_17604 ), .Q ( new_AGEMA_signal_17605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6113 ( .C ( clk ), .D ( new_AGEMA_signal_17612 ), .Q ( new_AGEMA_signal_17613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6119 ( .C ( clk ), .D ( n2306 ), .Q ( new_AGEMA_signal_17619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6125 ( .C ( clk ), .D ( new_AGEMA_signal_2979 ), .Q ( new_AGEMA_signal_17625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6131 ( .C ( clk ), .D ( new_AGEMA_signal_2980 ), .Q ( new_AGEMA_signal_17631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6137 ( .C ( clk ), .D ( new_AGEMA_signal_2981 ), .Q ( new_AGEMA_signal_17637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6145 ( .C ( clk ), .D ( new_AGEMA_signal_17644 ), .Q ( new_AGEMA_signal_17645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6153 ( .C ( clk ), .D ( new_AGEMA_signal_17652 ), .Q ( new_AGEMA_signal_17653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6161 ( .C ( clk ), .D ( new_AGEMA_signal_17660 ), .Q ( new_AGEMA_signal_17661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6169 ( .C ( clk ), .D ( new_AGEMA_signal_17668 ), .Q ( new_AGEMA_signal_17669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6177 ( .C ( clk ), .D ( new_AGEMA_signal_17676 ), .Q ( new_AGEMA_signal_17677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6185 ( .C ( clk ), .D ( new_AGEMA_signal_17684 ), .Q ( new_AGEMA_signal_17685 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6193 ( .C ( clk ), .D ( new_AGEMA_signal_17692 ), .Q ( new_AGEMA_signal_17693 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6201 ( .C ( clk ), .D ( new_AGEMA_signal_17700 ), .Q ( new_AGEMA_signal_17701 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6249 ( .C ( clk ), .D ( new_AGEMA_signal_17748 ), .Q ( new_AGEMA_signal_17749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6257 ( .C ( clk ), .D ( new_AGEMA_signal_17756 ), .Q ( new_AGEMA_signal_17757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6265 ( .C ( clk ), .D ( new_AGEMA_signal_17764 ), .Q ( new_AGEMA_signal_17765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6273 ( .C ( clk ), .D ( new_AGEMA_signal_17772 ), .Q ( new_AGEMA_signal_17773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6295 ( .C ( clk ), .D ( n1999 ), .Q ( new_AGEMA_signal_17795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6303 ( .C ( clk ), .D ( new_AGEMA_signal_3129 ), .Q ( new_AGEMA_signal_17803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6311 ( .C ( clk ), .D ( new_AGEMA_signal_3130 ), .Q ( new_AGEMA_signal_17811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6319 ( .C ( clk ), .D ( new_AGEMA_signal_3131 ), .Q ( new_AGEMA_signal_17819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6331 ( .C ( clk ), .D ( new_AGEMA_signal_17830 ), .Q ( new_AGEMA_signal_17831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6343 ( .C ( clk ), .D ( new_AGEMA_signal_17842 ), .Q ( new_AGEMA_signal_17843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6355 ( .C ( clk ), .D ( new_AGEMA_signal_17854 ), .Q ( new_AGEMA_signal_17855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6367 ( .C ( clk ), .D ( new_AGEMA_signal_17866 ), .Q ( new_AGEMA_signal_17867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6381 ( .C ( clk ), .D ( new_AGEMA_signal_17880 ), .Q ( new_AGEMA_signal_17881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6395 ( .C ( clk ), .D ( new_AGEMA_signal_17894 ), .Q ( new_AGEMA_signal_17895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6409 ( .C ( clk ), .D ( new_AGEMA_signal_17908 ), .Q ( new_AGEMA_signal_17909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6423 ( .C ( clk ), .D ( new_AGEMA_signal_17922 ), .Q ( new_AGEMA_signal_17923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6431 ( .C ( clk ), .D ( n2205 ), .Q ( new_AGEMA_signal_17931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6439 ( .C ( clk ), .D ( new_AGEMA_signal_3339 ), .Q ( new_AGEMA_signal_17939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6447 ( .C ( clk ), .D ( new_AGEMA_signal_3340 ), .Q ( new_AGEMA_signal_17947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6455 ( .C ( clk ), .D ( new_AGEMA_signal_3341 ), .Q ( new_AGEMA_signal_17955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6469 ( .C ( clk ), .D ( new_AGEMA_signal_17968 ), .Q ( new_AGEMA_signal_17969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6483 ( .C ( clk ), .D ( new_AGEMA_signal_17982 ), .Q ( new_AGEMA_signal_17983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6497 ( .C ( clk ), .D ( new_AGEMA_signal_17996 ), .Q ( new_AGEMA_signal_17997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6511 ( .C ( clk ), .D ( new_AGEMA_signal_18010 ), .Q ( new_AGEMA_signal_18011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6519 ( .C ( clk ), .D ( n2516 ), .Q ( new_AGEMA_signal_18019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6527 ( .C ( clk ), .D ( new_AGEMA_signal_3228 ), .Q ( new_AGEMA_signal_18027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6535 ( .C ( clk ), .D ( new_AGEMA_signal_3229 ), .Q ( new_AGEMA_signal_18035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6543 ( .C ( clk ), .D ( new_AGEMA_signal_3230 ), .Q ( new_AGEMA_signal_18043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6551 ( .C ( clk ), .D ( n2808 ), .Q ( new_AGEMA_signal_18051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6559 ( .C ( clk ), .D ( new_AGEMA_signal_3273 ), .Q ( new_AGEMA_signal_18059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6567 ( .C ( clk ), .D ( new_AGEMA_signal_3274 ), .Q ( new_AGEMA_signal_18067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6575 ( .C ( clk ), .D ( new_AGEMA_signal_3275 ), .Q ( new_AGEMA_signal_18075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6613 ( .C ( clk ), .D ( new_AGEMA_signal_18112 ), .Q ( new_AGEMA_signal_18113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6629 ( .C ( clk ), .D ( new_AGEMA_signal_18128 ), .Q ( new_AGEMA_signal_18129 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6645 ( .C ( clk ), .D ( new_AGEMA_signal_18144 ), .Q ( new_AGEMA_signal_18145 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6661 ( .C ( clk ), .D ( new_AGEMA_signal_18160 ), .Q ( new_AGEMA_signal_18161 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6701 ( .C ( clk ), .D ( new_AGEMA_signal_18200 ), .Q ( new_AGEMA_signal_18201 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6717 ( .C ( clk ), .D ( new_AGEMA_signal_18216 ), .Q ( new_AGEMA_signal_18217 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6733 ( .C ( clk ), .D ( new_AGEMA_signal_18232 ), .Q ( new_AGEMA_signal_18233 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6749 ( .C ( clk ), .D ( new_AGEMA_signal_18248 ), .Q ( new_AGEMA_signal_18249 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6759 ( .C ( clk ), .D ( n2527 ), .Q ( new_AGEMA_signal_18259 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6769 ( .C ( clk ), .D ( new_AGEMA_signal_3390 ), .Q ( new_AGEMA_signal_18269 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6779 ( .C ( clk ), .D ( new_AGEMA_signal_3391 ), .Q ( new_AGEMA_signal_18279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6789 ( .C ( clk ), .D ( new_AGEMA_signal_3392 ), .Q ( new_AGEMA_signal_18289 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6899 ( .C ( clk ), .D ( new_AGEMA_signal_18398 ), .Q ( new_AGEMA_signal_18399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6915 ( .C ( clk ), .D ( new_AGEMA_signal_18414 ), .Q ( new_AGEMA_signal_18415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6931 ( .C ( clk ), .D ( new_AGEMA_signal_18430 ), .Q ( new_AGEMA_signal_18431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6947 ( .C ( clk ), .D ( new_AGEMA_signal_18446 ), .Q ( new_AGEMA_signal_18447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7005 ( .C ( clk ), .D ( new_AGEMA_signal_18504 ), .Q ( new_AGEMA_signal_18505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7023 ( .C ( clk ), .D ( new_AGEMA_signal_18522 ), .Q ( new_AGEMA_signal_18523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7041 ( .C ( clk ), .D ( new_AGEMA_signal_18540 ), .Q ( new_AGEMA_signal_18541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7059 ( .C ( clk ), .D ( new_AGEMA_signal_18558 ), .Q ( new_AGEMA_signal_18559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7205 ( .C ( clk ), .D ( new_AGEMA_signal_18704 ), .Q ( new_AGEMA_signal_18705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7225 ( .C ( clk ), .D ( new_AGEMA_signal_18724 ), .Q ( new_AGEMA_signal_18725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7245 ( .C ( clk ), .D ( new_AGEMA_signal_18744 ), .Q ( new_AGEMA_signal_18745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7265 ( .C ( clk ), .D ( new_AGEMA_signal_18764 ), .Q ( new_AGEMA_signal_18765 ) ) ;

    /* cells in depth 14 */
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2002 ( .ina ({new_AGEMA_signal_15530, new_AGEMA_signal_15528, new_AGEMA_signal_15526, new_AGEMA_signal_15524}), .inb ({new_AGEMA_signal_3119, new_AGEMA_signal_3118, new_AGEMA_signal_3117, n1933}), .clk ( clk ), .rnd ({Fresh[7239], Fresh[7238], Fresh[7237], Fresh[7236], Fresh[7235], Fresh[7234], Fresh[7233], Fresh[7232], Fresh[7231], Fresh[7230]}), .outt ({new_AGEMA_signal_3296, new_AGEMA_signal_3295, new_AGEMA_signal_3294, n1935}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2054 ( .ina ({new_AGEMA_signal_3122, new_AGEMA_signal_3121, new_AGEMA_signal_3120, n1958}), .inb ({new_AGEMA_signal_15562, new_AGEMA_signal_15554, new_AGEMA_signal_15546, new_AGEMA_signal_15538}), .clk ( clk ), .rnd ({Fresh[7249], Fresh[7248], Fresh[7247], Fresh[7246], Fresh[7245], Fresh[7244], Fresh[7243], Fresh[7242], Fresh[7241], Fresh[7240]}), .outt ({new_AGEMA_signal_3299, new_AGEMA_signal_3298, new_AGEMA_signal_3297, n1959}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2109 ( .ina ({new_AGEMA_signal_3128, new_AGEMA_signal_3127, new_AGEMA_signal_3126, n1982}), .inb ({new_AGEMA_signal_15570, new_AGEMA_signal_15568, new_AGEMA_signal_15566, new_AGEMA_signal_15564}), .clk ( clk ), .rnd ({Fresh[7259], Fresh[7258], Fresh[7257], Fresh[7256], Fresh[7255], Fresh[7254], Fresh[7253], Fresh[7252], Fresh[7251], Fresh[7250]}), .outt ({new_AGEMA_signal_3302, new_AGEMA_signal_3301, new_AGEMA_signal_3300, n1983}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2149 ( .ina ({new_AGEMA_signal_15586, new_AGEMA_signal_15582, new_AGEMA_signal_15578, new_AGEMA_signal_15574}), .inb ({new_AGEMA_signal_3134, new_AGEMA_signal_3133, new_AGEMA_signal_3132, n2011}), .clk ( clk ), .rnd ({Fresh[7269], Fresh[7268], Fresh[7267], Fresh[7266], Fresh[7265], Fresh[7264], Fresh[7263], Fresh[7262], Fresh[7261], Fresh[7260]}), .outt ({new_AGEMA_signal_3305, new_AGEMA_signal_3304, new_AGEMA_signal_3303, n2014}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2166 ( .ina ({new_AGEMA_signal_15618, new_AGEMA_signal_15610, new_AGEMA_signal_15602, new_AGEMA_signal_15594}), .inb ({new_AGEMA_signal_2906, new_AGEMA_signal_2905, new_AGEMA_signal_2904, n2025}), .clk ( clk ), .rnd ({Fresh[7279], Fresh[7278], Fresh[7277], Fresh[7276], Fresh[7275], Fresh[7274], Fresh[7273], Fresh[7272], Fresh[7271], Fresh[7270]}), .outt ({new_AGEMA_signal_3137, new_AGEMA_signal_3136, new_AGEMA_signal_3135, n2029}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2180 ( .ina ({new_AGEMA_signal_15626, new_AGEMA_signal_15624, new_AGEMA_signal_15622, new_AGEMA_signal_15620}), .inb ({new_AGEMA_signal_3140, new_AGEMA_signal_3139, new_AGEMA_signal_3138, n2036}), .clk ( clk ), .rnd ({Fresh[7289], Fresh[7288], Fresh[7287], Fresh[7286], Fresh[7285], Fresh[7284], Fresh[7283], Fresh[7282], Fresh[7281], Fresh[7280]}), .outt ({new_AGEMA_signal_3311, new_AGEMA_signal_3310, new_AGEMA_signal_3309, n2037}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2197 ( .ina ({new_AGEMA_signal_15650, new_AGEMA_signal_15644, new_AGEMA_signal_15638, new_AGEMA_signal_15632}), .inb ({new_AGEMA_signal_3143, new_AGEMA_signal_3142, new_AGEMA_signal_3141, n2049}), .clk ( clk ), .rnd ({Fresh[7299], Fresh[7298], Fresh[7297], Fresh[7296], Fresh[7295], Fresh[7294], Fresh[7293], Fresh[7292], Fresh[7291], Fresh[7290]}), .outt ({new_AGEMA_signal_3314, new_AGEMA_signal_3313, new_AGEMA_signal_3312, n2052}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2219 ( .ina ({new_AGEMA_signal_3149, new_AGEMA_signal_3148, new_AGEMA_signal_3147, n2067}), .inb ({new_AGEMA_signal_15666, new_AGEMA_signal_15662, new_AGEMA_signal_15658, new_AGEMA_signal_15654}), .clk ( clk ), .rnd ({Fresh[7309], Fresh[7308], Fresh[7307], Fresh[7306], Fresh[7305], Fresh[7304], Fresh[7303], Fresh[7302], Fresh[7301], Fresh[7300]}), .outt ({new_AGEMA_signal_3317, new_AGEMA_signal_3316, new_AGEMA_signal_3315, n2070}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2258 ( .ina ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, new_AGEMA_signal_3153, n2097}), .inb ({new_AGEMA_signal_3158, new_AGEMA_signal_3157, new_AGEMA_signal_3156, n2096}), .clk ( clk ), .rnd ({Fresh[7319], Fresh[7318], Fresh[7317], Fresh[7316], Fresh[7315], Fresh[7314], Fresh[7313], Fresh[7312], Fresh[7311], Fresh[7310]}), .outt ({new_AGEMA_signal_3320, new_AGEMA_signal_3319, new_AGEMA_signal_3318, n2098}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2287 ( .ina ({new_AGEMA_signal_3164, new_AGEMA_signal_3163, new_AGEMA_signal_3162, n2124}), .inb ({new_AGEMA_signal_15698, new_AGEMA_signal_15690, new_AGEMA_signal_15682, new_AGEMA_signal_15674}), .clk ( clk ), .rnd ({Fresh[7329], Fresh[7328], Fresh[7327], Fresh[7326], Fresh[7325], Fresh[7324], Fresh[7323], Fresh[7322], Fresh[7321], Fresh[7320]}), .outt ({new_AGEMA_signal_3326, new_AGEMA_signal_3325, new_AGEMA_signal_3324, n2125}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2311 ( .ina ({new_AGEMA_signal_15714, new_AGEMA_signal_15710, new_AGEMA_signal_15706, new_AGEMA_signal_15702}), .inb ({new_AGEMA_signal_3167, new_AGEMA_signal_3166, new_AGEMA_signal_3165, n2142}), .clk ( clk ), .rnd ({Fresh[7339], Fresh[7338], Fresh[7337], Fresh[7336], Fresh[7335], Fresh[7334], Fresh[7333], Fresh[7332], Fresh[7331], Fresh[7330]}), .outt ({new_AGEMA_signal_3329, new_AGEMA_signal_3328, new_AGEMA_signal_3327, n2145}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2333 ( .ina ({new_AGEMA_signal_3170, new_AGEMA_signal_3169, new_AGEMA_signal_3168, n2168}), .inb ({new_AGEMA_signal_3173, new_AGEMA_signal_3172, new_AGEMA_signal_3171, n2167}), .clk ( clk ), .rnd ({Fresh[7349], Fresh[7348], Fresh[7347], Fresh[7346], Fresh[7345], Fresh[7344], Fresh[7343], Fresh[7342], Fresh[7341], Fresh[7340]}), .outt ({new_AGEMA_signal_3332, new_AGEMA_signal_3331, new_AGEMA_signal_3330, n2169}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2350 ( .ina ({new_AGEMA_signal_3176, new_AGEMA_signal_3175, new_AGEMA_signal_3174, n2184}), .inb ({new_AGEMA_signal_15738, new_AGEMA_signal_15732, new_AGEMA_signal_15726, new_AGEMA_signal_15720}), .clk ( clk ), .rnd ({Fresh[7359], Fresh[7358], Fresh[7357], Fresh[7356], Fresh[7355], Fresh[7354], Fresh[7353], Fresh[7352], Fresh[7351], Fresh[7350]}), .outt ({new_AGEMA_signal_3335, new_AGEMA_signal_3334, new_AGEMA_signal_3333, n2185}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2365 ( .ina ({new_AGEMA_signal_3179, new_AGEMA_signal_3178, new_AGEMA_signal_3177, n2197}), .inb ({new_AGEMA_signal_15762, new_AGEMA_signal_15756, new_AGEMA_signal_15750, new_AGEMA_signal_15744}), .clk ( clk ), .rnd ({Fresh[7369], Fresh[7368], Fresh[7367], Fresh[7366], Fresh[7365], Fresh[7364], Fresh[7363], Fresh[7362], Fresh[7361], Fresh[7360]}), .outt ({new_AGEMA_signal_3338, new_AGEMA_signal_3337, new_AGEMA_signal_3336, n2198}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2396 ( .ina ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, new_AGEMA_signal_3183, n2232}), .inb ({new_AGEMA_signal_2963, new_AGEMA_signal_2962, new_AGEMA_signal_2961, n2231}), .clk ( clk ), .rnd ({Fresh[7379], Fresh[7378], Fresh[7377], Fresh[7376], Fresh[7375], Fresh[7374], Fresh[7373], Fresh[7372], Fresh[7371], Fresh[7370]}), .outt ({new_AGEMA_signal_3344, new_AGEMA_signal_3343, new_AGEMA_signal_3342, n2312}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2404 ( .ina ({new_AGEMA_signal_3347, new_AGEMA_signal_3346, new_AGEMA_signal_3345, n2239}), .inb ({new_AGEMA_signal_15786, new_AGEMA_signal_15780, new_AGEMA_signal_15774, new_AGEMA_signal_15768}), .clk ( clk ), .rnd ({Fresh[7389], Fresh[7388], Fresh[7387], Fresh[7386], Fresh[7385], Fresh[7384], Fresh[7383], Fresh[7382], Fresh[7381], Fresh[7380]}), .outt ({new_AGEMA_signal_3461, new_AGEMA_signal_3460, new_AGEMA_signal_3459, n2258}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2415 ( .ina ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, new_AGEMA_signal_3189, n2250}), .inb ({new_AGEMA_signal_15810, new_AGEMA_signal_15804, new_AGEMA_signal_15798, new_AGEMA_signal_15792}), .clk ( clk ), .rnd ({Fresh[7399], Fresh[7398], Fresh[7397], Fresh[7396], Fresh[7395], Fresh[7394], Fresh[7393], Fresh[7392], Fresh[7391], Fresh[7390]}), .outt ({new_AGEMA_signal_3350, new_AGEMA_signal_3349, new_AGEMA_signal_3348, n2251}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2440 ( .ina ({new_AGEMA_signal_15834, new_AGEMA_signal_15828, new_AGEMA_signal_15822, new_AGEMA_signal_15816}), .inb ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, new_AGEMA_signal_3195, n2272}), .clk ( clk ), .rnd ({Fresh[7409], Fresh[7408], Fresh[7407], Fresh[7406], Fresh[7405], Fresh[7404], Fresh[7403], Fresh[7402], Fresh[7401], Fresh[7400]}), .outt ({new_AGEMA_signal_3353, new_AGEMA_signal_3352, new_AGEMA_signal_3351, n2274}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2469 ( .ina ({new_AGEMA_signal_15850, new_AGEMA_signal_15846, new_AGEMA_signal_15842, new_AGEMA_signal_15838}), .inb ({new_AGEMA_signal_3200, new_AGEMA_signal_3199, new_AGEMA_signal_3198, n2296}), .clk ( clk ), .rnd ({Fresh[7419], Fresh[7418], Fresh[7417], Fresh[7416], Fresh[7415], Fresh[7414], Fresh[7413], Fresh[7412], Fresh[7411], Fresh[7410]}), .outt ({new_AGEMA_signal_3356, new_AGEMA_signal_3355, new_AGEMA_signal_3354, n2302}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2490 ( .ina ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, new_AGEMA_signal_3201, n2324}), .inb ({new_AGEMA_signal_15882, new_AGEMA_signal_15874, new_AGEMA_signal_15866, new_AGEMA_signal_15858}), .clk ( clk ), .rnd ({Fresh[7429], Fresh[7428], Fresh[7427], Fresh[7426], Fresh[7425], Fresh[7424], Fresh[7423], Fresh[7422], Fresh[7421], Fresh[7420]}), .outt ({new_AGEMA_signal_3359, new_AGEMA_signal_3358, new_AGEMA_signal_3357, n2339}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2503 ( .ina ({new_AGEMA_signal_3206, new_AGEMA_signal_3205, new_AGEMA_signal_3204, n2337}), .inb ({new_AGEMA_signal_15898, new_AGEMA_signal_15894, new_AGEMA_signal_15890, new_AGEMA_signal_15886}), .clk ( clk ), .rnd ({Fresh[7439], Fresh[7438], Fresh[7437], Fresh[7436], Fresh[7435], Fresh[7434], Fresh[7433], Fresh[7432], Fresh[7431], Fresh[7430]}), .outt ({new_AGEMA_signal_3362, new_AGEMA_signal_3361, new_AGEMA_signal_3360, n2338}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2515 ( .ina ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, new_AGEMA_signal_3207, n2350}), .inb ({new_AGEMA_signal_15922, new_AGEMA_signal_15916, new_AGEMA_signal_15910, new_AGEMA_signal_15904}), .clk ( clk ), .rnd ({Fresh[7449], Fresh[7448], Fresh[7447], Fresh[7446], Fresh[7445], Fresh[7444], Fresh[7443], Fresh[7442], Fresh[7441], Fresh[7440]}), .outt ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, new_AGEMA_signal_3363, n2351}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2529 ( .ina ({new_AGEMA_signal_15954, new_AGEMA_signal_15946, new_AGEMA_signal_15938, new_AGEMA_signal_15930}), .inb ({new_AGEMA_signal_3212, new_AGEMA_signal_3211, new_AGEMA_signal_3210, n2362}), .clk ( clk ), .rnd ({Fresh[7459], Fresh[7458], Fresh[7457], Fresh[7456], Fresh[7455], Fresh[7454], Fresh[7453], Fresh[7452], Fresh[7451], Fresh[7450]}), .outt ({new_AGEMA_signal_3368, new_AGEMA_signal_3367, new_AGEMA_signal_3366, n2365}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2551 ( .ina ({new_AGEMA_signal_3005, new_AGEMA_signal_3004, new_AGEMA_signal_3003, n2389}), .inb ({new_AGEMA_signal_15962, new_AGEMA_signal_15960, new_AGEMA_signal_15958, new_AGEMA_signal_15956}), .clk ( clk ), .rnd ({Fresh[7469], Fresh[7468], Fresh[7467], Fresh[7466], Fresh[7465], Fresh[7464], Fresh[7463], Fresh[7462], Fresh[7461], Fresh[7460]}), .outt ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, new_AGEMA_signal_3213, n2399}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2560 ( .ina ({new_AGEMA_signal_3218, new_AGEMA_signal_3217, new_AGEMA_signal_3216, n2397}), .inb ({new_AGEMA_signal_15986, new_AGEMA_signal_15980, new_AGEMA_signal_15974, new_AGEMA_signal_15968}), .clk ( clk ), .rnd ({Fresh[7479], Fresh[7478], Fresh[7477], Fresh[7476], Fresh[7475], Fresh[7474], Fresh[7473], Fresh[7472], Fresh[7471], Fresh[7470]}), .outt ({new_AGEMA_signal_3371, new_AGEMA_signal_3370, new_AGEMA_signal_3369, n2398}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2572 ( .ina ({new_AGEMA_signal_3011, new_AGEMA_signal_3010, new_AGEMA_signal_3009, n2411}), .inb ({new_AGEMA_signal_15994, new_AGEMA_signal_15992, new_AGEMA_signal_15990, new_AGEMA_signal_15988}), .clk ( clk ), .rnd ({Fresh[7489], Fresh[7488], Fresh[7487], Fresh[7486], Fresh[7485], Fresh[7484], Fresh[7483], Fresh[7482], Fresh[7481], Fresh[7480]}), .outt ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, new_AGEMA_signal_3219, n2423}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2581 ( .ina ({new_AGEMA_signal_16002, new_AGEMA_signal_16000, new_AGEMA_signal_15998, new_AGEMA_signal_15996}), .inb ({new_AGEMA_signal_3020, new_AGEMA_signal_3019, new_AGEMA_signal_3018, n2420}), .clk ( clk ), .rnd ({Fresh[7499], Fresh[7498], Fresh[7497], Fresh[7496], Fresh[7495], Fresh[7494], Fresh[7493], Fresh[7492], Fresh[7491], Fresh[7490]}), .outt ({new_AGEMA_signal_3224, new_AGEMA_signal_3223, new_AGEMA_signal_3222, n2422}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2596 ( .ina ({new_AGEMA_signal_3227, new_AGEMA_signal_3226, new_AGEMA_signal_3225, n2440}), .inb ({new_AGEMA_signal_16026, new_AGEMA_signal_16020, new_AGEMA_signal_16014, new_AGEMA_signal_16008}), .clk ( clk ), .rnd ({Fresh[7509], Fresh[7508], Fresh[7507], Fresh[7506], Fresh[7505], Fresh[7504], Fresh[7503], Fresh[7502], Fresh[7501], Fresh[7500]}), .outt ({new_AGEMA_signal_3377, new_AGEMA_signal_3376, new_AGEMA_signal_3375, n2441}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2623 ( .ina ({new_AGEMA_signal_3035, new_AGEMA_signal_3034, new_AGEMA_signal_3033, n2471}), .inb ({new_AGEMA_signal_16050, new_AGEMA_signal_16044, new_AGEMA_signal_16038, new_AGEMA_signal_16032}), .clk ( clk ), .rnd ({Fresh[7519], Fresh[7518], Fresh[7517], Fresh[7516], Fresh[7515], Fresh[7514], Fresh[7513], Fresh[7512], Fresh[7511], Fresh[7510]}), .outt ({new_AGEMA_signal_3233, new_AGEMA_signal_3232, new_AGEMA_signal_3231, n2479}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2637 ( .ina ({new_AGEMA_signal_3236, new_AGEMA_signal_3235, new_AGEMA_signal_3234, n2485}), .inb ({new_AGEMA_signal_16082, new_AGEMA_signal_16074, new_AGEMA_signal_16066, new_AGEMA_signal_16058}), .clk ( clk ), .rnd ({Fresh[7529], Fresh[7528], Fresh[7527], Fresh[7526], Fresh[7525], Fresh[7524], Fresh[7523], Fresh[7522], Fresh[7521], Fresh[7520]}), .outt ({new_AGEMA_signal_3383, new_AGEMA_signal_3382, new_AGEMA_signal_3381, n2512}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2652 ( .ina ({new_AGEMA_signal_3041, new_AGEMA_signal_3040, new_AGEMA_signal_3039, n2502}), .inb ({new_AGEMA_signal_3239, new_AGEMA_signal_3238, new_AGEMA_signal_3237, n2501}), .clk ( clk ), .rnd ({Fresh[7539], Fresh[7538], Fresh[7537], Fresh[7536], Fresh[7535], Fresh[7534], Fresh[7533], Fresh[7532], Fresh[7531], Fresh[7530]}), .outt ({new_AGEMA_signal_3386, new_AGEMA_signal_3385, new_AGEMA_signal_3384, n2510}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2686 ( .ina ({new_AGEMA_signal_3248, new_AGEMA_signal_3247, new_AGEMA_signal_3246, n2550}), .inb ({new_AGEMA_signal_3251, new_AGEMA_signal_3250, new_AGEMA_signal_3249, n2549}), .clk ( clk ), .rnd ({Fresh[7549], Fresh[7548], Fresh[7547], Fresh[7546], Fresh[7545], Fresh[7544], Fresh[7543], Fresh[7542], Fresh[7541], Fresh[7540]}), .outt ({new_AGEMA_signal_3395, new_AGEMA_signal_3394, new_AGEMA_signal_3393, n2552}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2702 ( .ina ({new_AGEMA_signal_16114, new_AGEMA_signal_16106, new_AGEMA_signal_16098, new_AGEMA_signal_16090}), .inb ({new_AGEMA_signal_3254, new_AGEMA_signal_3253, new_AGEMA_signal_3252, n2569}), .clk ( clk ), .rnd ({Fresh[7559], Fresh[7558], Fresh[7557], Fresh[7556], Fresh[7555], Fresh[7554], Fresh[7553], Fresh[7552], Fresh[7551], Fresh[7550]}), .outt ({new_AGEMA_signal_3398, new_AGEMA_signal_3397, new_AGEMA_signal_3396, n2593}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2713 ( .ina ({new_AGEMA_signal_16138, new_AGEMA_signal_16132, new_AGEMA_signal_16126, new_AGEMA_signal_16120}), .inb ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, new_AGEMA_signal_3255, n2584}), .clk ( clk ), .rnd ({Fresh[7569], Fresh[7568], Fresh[7567], Fresh[7566], Fresh[7565], Fresh[7564], Fresh[7563], Fresh[7562], Fresh[7561], Fresh[7560]}), .outt ({new_AGEMA_signal_3401, new_AGEMA_signal_3400, new_AGEMA_signal_3399, n2589}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2730 ( .ina ({new_AGEMA_signal_16162, new_AGEMA_signal_16156, new_AGEMA_signal_16150, new_AGEMA_signal_16144}), .inb ({new_AGEMA_signal_3068, new_AGEMA_signal_3067, new_AGEMA_signal_3066, n2606}), .clk ( clk ), .rnd ({Fresh[7579], Fresh[7578], Fresh[7577], Fresh[7576], Fresh[7575], Fresh[7574], Fresh[7573], Fresh[7572], Fresh[7571], Fresh[7570]}), .outt ({new_AGEMA_signal_3260, new_AGEMA_signal_3259, new_AGEMA_signal_3258, n2608}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2748 ( .ina ({new_AGEMA_signal_16170, new_AGEMA_signal_16168, new_AGEMA_signal_16166, new_AGEMA_signal_16164}), .inb ({new_AGEMA_signal_3266, new_AGEMA_signal_3265, new_AGEMA_signal_3264, n2634}), .clk ( clk ), .rnd ({Fresh[7589], Fresh[7588], Fresh[7587], Fresh[7586], Fresh[7585], Fresh[7584], Fresh[7583], Fresh[7582], Fresh[7581], Fresh[7580]}), .outt ({new_AGEMA_signal_3407, new_AGEMA_signal_3406, new_AGEMA_signal_3405, n2636}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2762 ( .ina ({new_AGEMA_signal_16186, new_AGEMA_signal_16182, new_AGEMA_signal_16178, new_AGEMA_signal_16174}), .inb ({new_AGEMA_signal_3269, new_AGEMA_signal_3268, new_AGEMA_signal_3267, n2657}), .clk ( clk ), .rnd ({Fresh[7599], Fresh[7598], Fresh[7597], Fresh[7596], Fresh[7595], Fresh[7594], Fresh[7593], Fresh[7592], Fresh[7591], Fresh[7590]}), .outt ({new_AGEMA_signal_3410, new_AGEMA_signal_3409, new_AGEMA_signal_3408, n2659}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2784 ( .ina ({new_AGEMA_signal_16202, new_AGEMA_signal_16198, new_AGEMA_signal_16194, new_AGEMA_signal_16190}), .inb ({new_AGEMA_signal_3272, new_AGEMA_signal_3271, new_AGEMA_signal_3270, n2697}), .clk ( clk ), .rnd ({Fresh[7609], Fresh[7608], Fresh[7607], Fresh[7606], Fresh[7605], Fresh[7604], Fresh[7603], Fresh[7602], Fresh[7601], Fresh[7600]}), .outt ({new_AGEMA_signal_3413, new_AGEMA_signal_3412, new_AGEMA_signal_3411, n2702}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2811 ( .ina ({new_AGEMA_signal_3278, new_AGEMA_signal_3277, new_AGEMA_signal_3276, n2747}), .inb ({new_AGEMA_signal_3281, new_AGEMA_signal_3280, new_AGEMA_signal_3279, n2746}), .clk ( clk ), .rnd ({Fresh[7619], Fresh[7618], Fresh[7617], Fresh[7616], Fresh[7615], Fresh[7614], Fresh[7613], Fresh[7612], Fresh[7611], Fresh[7610]}), .outt ({new_AGEMA_signal_3416, new_AGEMA_signal_3415, new_AGEMA_signal_3414, n2806}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2839 ( .ina ({new_AGEMA_signal_16218, new_AGEMA_signal_16214, new_AGEMA_signal_16210, new_AGEMA_signal_16206}), .inb ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, new_AGEMA_signal_3111, n2799}), .clk ( clk ), .rnd ({Fresh[7629], Fresh[7628], Fresh[7627], Fresh[7626], Fresh[7625], Fresh[7624], Fresh[7623], Fresh[7622], Fresh[7621], Fresh[7620]}), .outt ({new_AGEMA_signal_3290, new_AGEMA_signal_3289, new_AGEMA_signal_3288, n2801}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2853 ( .ina ({new_AGEMA_signal_16226, new_AGEMA_signal_16224, new_AGEMA_signal_16222, new_AGEMA_signal_16220}), .inb ({new_AGEMA_signal_3293, new_AGEMA_signal_3292, new_AGEMA_signal_3291, n2827}), .clk ( clk ), .rnd ({Fresh[7639], Fresh[7638], Fresh[7637], Fresh[7636], Fresh[7635], Fresh[7634], Fresh[7633], Fresh[7632], Fresh[7631], Fresh[7630]}), .outt ({new_AGEMA_signal_3422, new_AGEMA_signal_3421, new_AGEMA_signal_3420, n2829}) ) ;
    buf_clk new_AGEMA_reg_buffer_4732 ( .C ( clk ), .D ( new_AGEMA_signal_16231 ), .Q ( new_AGEMA_signal_16232 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4738 ( .C ( clk ), .D ( new_AGEMA_signal_16237 ), .Q ( new_AGEMA_signal_16238 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4744 ( .C ( clk ), .D ( new_AGEMA_signal_16243 ), .Q ( new_AGEMA_signal_16244 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4750 ( .C ( clk ), .D ( new_AGEMA_signal_16249 ), .Q ( new_AGEMA_signal_16250 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4752 ( .C ( clk ), .D ( new_AGEMA_signal_16251 ), .Q ( new_AGEMA_signal_16252 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4754 ( .C ( clk ), .D ( new_AGEMA_signal_16253 ), .Q ( new_AGEMA_signal_16254 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4756 ( .C ( clk ), .D ( new_AGEMA_signal_16255 ), .Q ( new_AGEMA_signal_16256 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4758 ( .C ( clk ), .D ( new_AGEMA_signal_16257 ), .Q ( new_AGEMA_signal_16258 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4762 ( .C ( clk ), .D ( new_AGEMA_signal_16261 ), .Q ( new_AGEMA_signal_16262 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4766 ( .C ( clk ), .D ( new_AGEMA_signal_16265 ), .Q ( new_AGEMA_signal_16266 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4770 ( .C ( clk ), .D ( new_AGEMA_signal_16269 ), .Q ( new_AGEMA_signal_16270 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4774 ( .C ( clk ), .D ( new_AGEMA_signal_16273 ), .Q ( new_AGEMA_signal_16274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4782 ( .C ( clk ), .D ( new_AGEMA_signal_16281 ), .Q ( new_AGEMA_signal_16282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4790 ( .C ( clk ), .D ( new_AGEMA_signal_16289 ), .Q ( new_AGEMA_signal_16290 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4798 ( .C ( clk ), .D ( new_AGEMA_signal_16297 ), .Q ( new_AGEMA_signal_16298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4806 ( .C ( clk ), .D ( new_AGEMA_signal_16305 ), .Q ( new_AGEMA_signal_16306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4814 ( .C ( clk ), .D ( new_AGEMA_signal_16313 ), .Q ( new_AGEMA_signal_16314 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4822 ( .C ( clk ), .D ( new_AGEMA_signal_16321 ), .Q ( new_AGEMA_signal_16322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4830 ( .C ( clk ), .D ( new_AGEMA_signal_16329 ), .Q ( new_AGEMA_signal_16330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4838 ( .C ( clk ), .D ( new_AGEMA_signal_16337 ), .Q ( new_AGEMA_signal_16338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4846 ( .C ( clk ), .D ( new_AGEMA_signal_16345 ), .Q ( new_AGEMA_signal_16346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4854 ( .C ( clk ), .D ( new_AGEMA_signal_16353 ), .Q ( new_AGEMA_signal_16354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4862 ( .C ( clk ), .D ( new_AGEMA_signal_16361 ), .Q ( new_AGEMA_signal_16362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4870 ( .C ( clk ), .D ( new_AGEMA_signal_16369 ), .Q ( new_AGEMA_signal_16370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4878 ( .C ( clk ), .D ( new_AGEMA_signal_16377 ), .Q ( new_AGEMA_signal_16378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4886 ( .C ( clk ), .D ( new_AGEMA_signal_16385 ), .Q ( new_AGEMA_signal_16386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4894 ( .C ( clk ), .D ( new_AGEMA_signal_16393 ), .Q ( new_AGEMA_signal_16394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4902 ( .C ( clk ), .D ( new_AGEMA_signal_16401 ), .Q ( new_AGEMA_signal_16402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4908 ( .C ( clk ), .D ( new_AGEMA_signal_16407 ), .Q ( new_AGEMA_signal_16408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4914 ( .C ( clk ), .D ( new_AGEMA_signal_16413 ), .Q ( new_AGEMA_signal_16414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4920 ( .C ( clk ), .D ( new_AGEMA_signal_16419 ), .Q ( new_AGEMA_signal_16420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4926 ( .C ( clk ), .D ( new_AGEMA_signal_16425 ), .Q ( new_AGEMA_signal_16426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4936 ( .C ( clk ), .D ( new_AGEMA_signal_16435 ), .Q ( new_AGEMA_signal_16436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4946 ( .C ( clk ), .D ( new_AGEMA_signal_16445 ), .Q ( new_AGEMA_signal_16446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4956 ( .C ( clk ), .D ( new_AGEMA_signal_16455 ), .Q ( new_AGEMA_signal_16456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4966 ( .C ( clk ), .D ( new_AGEMA_signal_16465 ), .Q ( new_AGEMA_signal_16466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4974 ( .C ( clk ), .D ( new_AGEMA_signal_16473 ), .Q ( new_AGEMA_signal_16474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4982 ( .C ( clk ), .D ( new_AGEMA_signal_16481 ), .Q ( new_AGEMA_signal_16482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4990 ( .C ( clk ), .D ( new_AGEMA_signal_16489 ), .Q ( new_AGEMA_signal_16490 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4998 ( .C ( clk ), .D ( new_AGEMA_signal_16497 ), .Q ( new_AGEMA_signal_16498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5006 ( .C ( clk ), .D ( new_AGEMA_signal_16505 ), .Q ( new_AGEMA_signal_16506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5014 ( .C ( clk ), .D ( new_AGEMA_signal_16513 ), .Q ( new_AGEMA_signal_16514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5022 ( .C ( clk ), .D ( new_AGEMA_signal_16521 ), .Q ( new_AGEMA_signal_16522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5030 ( .C ( clk ), .D ( new_AGEMA_signal_16529 ), .Q ( new_AGEMA_signal_16530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5038 ( .C ( clk ), .D ( new_AGEMA_signal_16537 ), .Q ( new_AGEMA_signal_16538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5046 ( .C ( clk ), .D ( new_AGEMA_signal_16545 ), .Q ( new_AGEMA_signal_16546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5054 ( .C ( clk ), .D ( new_AGEMA_signal_16553 ), .Q ( new_AGEMA_signal_16554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5062 ( .C ( clk ), .D ( new_AGEMA_signal_16561 ), .Q ( new_AGEMA_signal_16562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5064 ( .C ( clk ), .D ( new_AGEMA_signal_16563 ), .Q ( new_AGEMA_signal_16564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5066 ( .C ( clk ), .D ( new_AGEMA_signal_16565 ), .Q ( new_AGEMA_signal_16566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5068 ( .C ( clk ), .D ( new_AGEMA_signal_16567 ), .Q ( new_AGEMA_signal_16568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5070 ( .C ( clk ), .D ( new_AGEMA_signal_16569 ), .Q ( new_AGEMA_signal_16570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5074 ( .C ( clk ), .D ( new_AGEMA_signal_16573 ), .Q ( new_AGEMA_signal_16574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5078 ( .C ( clk ), .D ( new_AGEMA_signal_16577 ), .Q ( new_AGEMA_signal_16578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5082 ( .C ( clk ), .D ( new_AGEMA_signal_16581 ), .Q ( new_AGEMA_signal_16582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5086 ( .C ( clk ), .D ( new_AGEMA_signal_16585 ), .Q ( new_AGEMA_signal_16586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5092 ( .C ( clk ), .D ( new_AGEMA_signal_16591 ), .Q ( new_AGEMA_signal_16592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5098 ( .C ( clk ), .D ( new_AGEMA_signal_16597 ), .Q ( new_AGEMA_signal_16598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5104 ( .C ( clk ), .D ( new_AGEMA_signal_16603 ), .Q ( new_AGEMA_signal_16604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5110 ( .C ( clk ), .D ( new_AGEMA_signal_16609 ), .Q ( new_AGEMA_signal_16610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5114 ( .C ( clk ), .D ( new_AGEMA_signal_16613 ), .Q ( new_AGEMA_signal_16614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5118 ( .C ( clk ), .D ( new_AGEMA_signal_16617 ), .Q ( new_AGEMA_signal_16618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5122 ( .C ( clk ), .D ( new_AGEMA_signal_16621 ), .Q ( new_AGEMA_signal_16622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5126 ( .C ( clk ), .D ( new_AGEMA_signal_16625 ), .Q ( new_AGEMA_signal_16626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5136 ( .C ( clk ), .D ( new_AGEMA_signal_16635 ), .Q ( new_AGEMA_signal_16636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5146 ( .C ( clk ), .D ( new_AGEMA_signal_16645 ), .Q ( new_AGEMA_signal_16646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5156 ( .C ( clk ), .D ( new_AGEMA_signal_16655 ), .Q ( new_AGEMA_signal_16656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5166 ( .C ( clk ), .D ( new_AGEMA_signal_16665 ), .Q ( new_AGEMA_signal_16666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5174 ( .C ( clk ), .D ( new_AGEMA_signal_16673 ), .Q ( new_AGEMA_signal_16674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5182 ( .C ( clk ), .D ( new_AGEMA_signal_16681 ), .Q ( new_AGEMA_signal_16682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5190 ( .C ( clk ), .D ( new_AGEMA_signal_16689 ), .Q ( new_AGEMA_signal_16690 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5198 ( .C ( clk ), .D ( new_AGEMA_signal_16697 ), .Q ( new_AGEMA_signal_16698 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5202 ( .C ( clk ), .D ( new_AGEMA_signal_16701 ), .Q ( new_AGEMA_signal_16702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5206 ( .C ( clk ), .D ( new_AGEMA_signal_16705 ), .Q ( new_AGEMA_signal_16706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5210 ( .C ( clk ), .D ( new_AGEMA_signal_16709 ), .Q ( new_AGEMA_signal_16710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5214 ( .C ( clk ), .D ( new_AGEMA_signal_16713 ), .Q ( new_AGEMA_signal_16714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5216 ( .C ( clk ), .D ( new_AGEMA_signal_16715 ), .Q ( new_AGEMA_signal_16716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5218 ( .C ( clk ), .D ( new_AGEMA_signal_16717 ), .Q ( new_AGEMA_signal_16718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5220 ( .C ( clk ), .D ( new_AGEMA_signal_16719 ), .Q ( new_AGEMA_signal_16720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5222 ( .C ( clk ), .D ( new_AGEMA_signal_16721 ), .Q ( new_AGEMA_signal_16722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5230 ( .C ( clk ), .D ( new_AGEMA_signal_16729 ), .Q ( new_AGEMA_signal_16730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5238 ( .C ( clk ), .D ( new_AGEMA_signal_16737 ), .Q ( new_AGEMA_signal_16738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5246 ( .C ( clk ), .D ( new_AGEMA_signal_16745 ), .Q ( new_AGEMA_signal_16746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5254 ( .C ( clk ), .D ( new_AGEMA_signal_16753 ), .Q ( new_AGEMA_signal_16754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5262 ( .C ( clk ), .D ( new_AGEMA_signal_16761 ), .Q ( new_AGEMA_signal_16762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5270 ( .C ( clk ), .D ( new_AGEMA_signal_16769 ), .Q ( new_AGEMA_signal_16770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5278 ( .C ( clk ), .D ( new_AGEMA_signal_16777 ), .Q ( new_AGEMA_signal_16778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5286 ( .C ( clk ), .D ( new_AGEMA_signal_16785 ), .Q ( new_AGEMA_signal_16786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5292 ( .C ( clk ), .D ( new_AGEMA_signal_16791 ), .Q ( new_AGEMA_signal_16792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5298 ( .C ( clk ), .D ( new_AGEMA_signal_16797 ), .Q ( new_AGEMA_signal_16798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5304 ( .C ( clk ), .D ( new_AGEMA_signal_16803 ), .Q ( new_AGEMA_signal_16804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5310 ( .C ( clk ), .D ( new_AGEMA_signal_16809 ), .Q ( new_AGEMA_signal_16810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5314 ( .C ( clk ), .D ( new_AGEMA_signal_16813 ), .Q ( new_AGEMA_signal_16814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5318 ( .C ( clk ), .D ( new_AGEMA_signal_16817 ), .Q ( new_AGEMA_signal_16818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5322 ( .C ( clk ), .D ( new_AGEMA_signal_16821 ), .Q ( new_AGEMA_signal_16822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5326 ( .C ( clk ), .D ( new_AGEMA_signal_16825 ), .Q ( new_AGEMA_signal_16826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5334 ( .C ( clk ), .D ( new_AGEMA_signal_16833 ), .Q ( new_AGEMA_signal_16834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5342 ( .C ( clk ), .D ( new_AGEMA_signal_16841 ), .Q ( new_AGEMA_signal_16842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5350 ( .C ( clk ), .D ( new_AGEMA_signal_16849 ), .Q ( new_AGEMA_signal_16850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5358 ( .C ( clk ), .D ( new_AGEMA_signal_16857 ), .Q ( new_AGEMA_signal_16858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5360 ( .C ( clk ), .D ( new_AGEMA_signal_16859 ), .Q ( new_AGEMA_signal_16860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5362 ( .C ( clk ), .D ( new_AGEMA_signal_16861 ), .Q ( new_AGEMA_signal_16862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5364 ( .C ( clk ), .D ( new_AGEMA_signal_16863 ), .Q ( new_AGEMA_signal_16864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5366 ( .C ( clk ), .D ( new_AGEMA_signal_16865 ), .Q ( new_AGEMA_signal_16866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5370 ( .C ( clk ), .D ( new_AGEMA_signal_16869 ), .Q ( new_AGEMA_signal_16870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5376 ( .C ( clk ), .D ( new_AGEMA_signal_16875 ), .Q ( new_AGEMA_signal_16876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5382 ( .C ( clk ), .D ( new_AGEMA_signal_16881 ), .Q ( new_AGEMA_signal_16882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5388 ( .C ( clk ), .D ( new_AGEMA_signal_16887 ), .Q ( new_AGEMA_signal_16888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5394 ( .C ( clk ), .D ( new_AGEMA_signal_16893 ), .Q ( new_AGEMA_signal_16894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5400 ( .C ( clk ), .D ( new_AGEMA_signal_16899 ), .Q ( new_AGEMA_signal_16900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5406 ( .C ( clk ), .D ( new_AGEMA_signal_16905 ), .Q ( new_AGEMA_signal_16906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5412 ( .C ( clk ), .D ( new_AGEMA_signal_16911 ), .Q ( new_AGEMA_signal_16912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5418 ( .C ( clk ), .D ( new_AGEMA_signal_16917 ), .Q ( new_AGEMA_signal_16918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5424 ( .C ( clk ), .D ( new_AGEMA_signal_16923 ), .Q ( new_AGEMA_signal_16924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5430 ( .C ( clk ), .D ( new_AGEMA_signal_16929 ), .Q ( new_AGEMA_signal_16930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5436 ( .C ( clk ), .D ( new_AGEMA_signal_16935 ), .Q ( new_AGEMA_signal_16936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5440 ( .C ( clk ), .D ( new_AGEMA_signal_16939 ), .Q ( new_AGEMA_signal_16940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5444 ( .C ( clk ), .D ( new_AGEMA_signal_16943 ), .Q ( new_AGEMA_signal_16944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5448 ( .C ( clk ), .D ( new_AGEMA_signal_16947 ), .Q ( new_AGEMA_signal_16948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5452 ( .C ( clk ), .D ( new_AGEMA_signal_16951 ), .Q ( new_AGEMA_signal_16952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5460 ( .C ( clk ), .D ( new_AGEMA_signal_16959 ), .Q ( new_AGEMA_signal_16960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5468 ( .C ( clk ), .D ( new_AGEMA_signal_16967 ), .Q ( new_AGEMA_signal_16968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5476 ( .C ( clk ), .D ( new_AGEMA_signal_16975 ), .Q ( new_AGEMA_signal_16976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5484 ( .C ( clk ), .D ( new_AGEMA_signal_16983 ), .Q ( new_AGEMA_signal_16984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5490 ( .C ( clk ), .D ( new_AGEMA_signal_16989 ), .Q ( new_AGEMA_signal_16990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5496 ( .C ( clk ), .D ( new_AGEMA_signal_16995 ), .Q ( new_AGEMA_signal_16996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5502 ( .C ( clk ), .D ( new_AGEMA_signal_17001 ), .Q ( new_AGEMA_signal_17002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5508 ( .C ( clk ), .D ( new_AGEMA_signal_17007 ), .Q ( new_AGEMA_signal_17008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5512 ( .C ( clk ), .D ( new_AGEMA_signal_17011 ), .Q ( new_AGEMA_signal_17012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5516 ( .C ( clk ), .D ( new_AGEMA_signal_17015 ), .Q ( new_AGEMA_signal_17016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5520 ( .C ( clk ), .D ( new_AGEMA_signal_17019 ), .Q ( new_AGEMA_signal_17020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5524 ( .C ( clk ), .D ( new_AGEMA_signal_17023 ), .Q ( new_AGEMA_signal_17024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5532 ( .C ( clk ), .D ( new_AGEMA_signal_17031 ), .Q ( new_AGEMA_signal_17032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5540 ( .C ( clk ), .D ( new_AGEMA_signal_17039 ), .Q ( new_AGEMA_signal_17040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5548 ( .C ( clk ), .D ( new_AGEMA_signal_17047 ), .Q ( new_AGEMA_signal_17048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5556 ( .C ( clk ), .D ( new_AGEMA_signal_17055 ), .Q ( new_AGEMA_signal_17056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5564 ( .C ( clk ), .D ( new_AGEMA_signal_17063 ), .Q ( new_AGEMA_signal_17064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5572 ( .C ( clk ), .D ( new_AGEMA_signal_17071 ), .Q ( new_AGEMA_signal_17072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5580 ( .C ( clk ), .D ( new_AGEMA_signal_17079 ), .Q ( new_AGEMA_signal_17080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5588 ( .C ( clk ), .D ( new_AGEMA_signal_17087 ), .Q ( new_AGEMA_signal_17088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5598 ( .C ( clk ), .D ( new_AGEMA_signal_17097 ), .Q ( new_AGEMA_signal_17098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5608 ( .C ( clk ), .D ( new_AGEMA_signal_17107 ), .Q ( new_AGEMA_signal_17108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5618 ( .C ( clk ), .D ( new_AGEMA_signal_17117 ), .Q ( new_AGEMA_signal_17118 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5628 ( .C ( clk ), .D ( new_AGEMA_signal_17127 ), .Q ( new_AGEMA_signal_17128 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5636 ( .C ( clk ), .D ( new_AGEMA_signal_17135 ), .Q ( new_AGEMA_signal_17136 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5644 ( .C ( clk ), .D ( new_AGEMA_signal_17143 ), .Q ( new_AGEMA_signal_17144 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5652 ( .C ( clk ), .D ( new_AGEMA_signal_17151 ), .Q ( new_AGEMA_signal_17152 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5660 ( .C ( clk ), .D ( new_AGEMA_signal_17159 ), .Q ( new_AGEMA_signal_17160 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5666 ( .C ( clk ), .D ( new_AGEMA_signal_17165 ), .Q ( new_AGEMA_signal_17166 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5672 ( .C ( clk ), .D ( new_AGEMA_signal_17171 ), .Q ( new_AGEMA_signal_17172 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5678 ( .C ( clk ), .D ( new_AGEMA_signal_17177 ), .Q ( new_AGEMA_signal_17178 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5684 ( .C ( clk ), .D ( new_AGEMA_signal_17183 ), .Q ( new_AGEMA_signal_17184 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5688 ( .C ( clk ), .D ( new_AGEMA_signal_17187 ), .Q ( new_AGEMA_signal_17188 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5692 ( .C ( clk ), .D ( new_AGEMA_signal_17191 ), .Q ( new_AGEMA_signal_17192 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5696 ( .C ( clk ), .D ( new_AGEMA_signal_17195 ), .Q ( new_AGEMA_signal_17196 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5700 ( .C ( clk ), .D ( new_AGEMA_signal_17199 ), .Q ( new_AGEMA_signal_17200 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5706 ( .C ( clk ), .D ( new_AGEMA_signal_17205 ), .Q ( new_AGEMA_signal_17206 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5712 ( .C ( clk ), .D ( new_AGEMA_signal_17211 ), .Q ( new_AGEMA_signal_17212 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5718 ( .C ( clk ), .D ( new_AGEMA_signal_17217 ), .Q ( new_AGEMA_signal_17218 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5724 ( .C ( clk ), .D ( new_AGEMA_signal_17223 ), .Q ( new_AGEMA_signal_17224 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5732 ( .C ( clk ), .D ( new_AGEMA_signal_17231 ), .Q ( new_AGEMA_signal_17232 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5740 ( .C ( clk ), .D ( new_AGEMA_signal_17239 ), .Q ( new_AGEMA_signal_17240 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5748 ( .C ( clk ), .D ( new_AGEMA_signal_17247 ), .Q ( new_AGEMA_signal_17248 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5756 ( .C ( clk ), .D ( new_AGEMA_signal_17255 ), .Q ( new_AGEMA_signal_17256 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5762 ( .C ( clk ), .D ( new_AGEMA_signal_17261 ), .Q ( new_AGEMA_signal_17262 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5768 ( .C ( clk ), .D ( new_AGEMA_signal_17267 ), .Q ( new_AGEMA_signal_17268 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5774 ( .C ( clk ), .D ( new_AGEMA_signal_17273 ), .Q ( new_AGEMA_signal_17274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5780 ( .C ( clk ), .D ( new_AGEMA_signal_17279 ), .Q ( new_AGEMA_signal_17280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5796 ( .C ( clk ), .D ( new_AGEMA_signal_17295 ), .Q ( new_AGEMA_signal_17296 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5804 ( .C ( clk ), .D ( new_AGEMA_signal_17303 ), .Q ( new_AGEMA_signal_17304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5812 ( .C ( clk ), .D ( new_AGEMA_signal_17311 ), .Q ( new_AGEMA_signal_17312 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5820 ( .C ( clk ), .D ( new_AGEMA_signal_17319 ), .Q ( new_AGEMA_signal_17320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5824 ( .C ( clk ), .D ( new_AGEMA_signal_17323 ), .Q ( new_AGEMA_signal_17324 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5828 ( .C ( clk ), .D ( new_AGEMA_signal_17327 ), .Q ( new_AGEMA_signal_17328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5832 ( .C ( clk ), .D ( new_AGEMA_signal_17331 ), .Q ( new_AGEMA_signal_17332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5836 ( .C ( clk ), .D ( new_AGEMA_signal_17335 ), .Q ( new_AGEMA_signal_17336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5842 ( .C ( clk ), .D ( new_AGEMA_signal_17341 ), .Q ( new_AGEMA_signal_17342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5848 ( .C ( clk ), .D ( new_AGEMA_signal_17347 ), .Q ( new_AGEMA_signal_17348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5854 ( .C ( clk ), .D ( new_AGEMA_signal_17353 ), .Q ( new_AGEMA_signal_17354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5860 ( .C ( clk ), .D ( new_AGEMA_signal_17359 ), .Q ( new_AGEMA_signal_17360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5866 ( .C ( clk ), .D ( new_AGEMA_signal_17365 ), .Q ( new_AGEMA_signal_17366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5872 ( .C ( clk ), .D ( new_AGEMA_signal_17371 ), .Q ( new_AGEMA_signal_17372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5878 ( .C ( clk ), .D ( new_AGEMA_signal_17377 ), .Q ( new_AGEMA_signal_17378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5884 ( .C ( clk ), .D ( new_AGEMA_signal_17383 ), .Q ( new_AGEMA_signal_17384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5888 ( .C ( clk ), .D ( new_AGEMA_signal_17387 ), .Q ( new_AGEMA_signal_17388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5892 ( .C ( clk ), .D ( new_AGEMA_signal_17391 ), .Q ( new_AGEMA_signal_17392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5896 ( .C ( clk ), .D ( new_AGEMA_signal_17395 ), .Q ( new_AGEMA_signal_17396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5900 ( .C ( clk ), .D ( new_AGEMA_signal_17399 ), .Q ( new_AGEMA_signal_17400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5904 ( .C ( clk ), .D ( new_AGEMA_signal_17403 ), .Q ( new_AGEMA_signal_17404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5910 ( .C ( clk ), .D ( new_AGEMA_signal_17409 ), .Q ( new_AGEMA_signal_17410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5916 ( .C ( clk ), .D ( new_AGEMA_signal_17415 ), .Q ( new_AGEMA_signal_17416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5922 ( .C ( clk ), .D ( new_AGEMA_signal_17421 ), .Q ( new_AGEMA_signal_17422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5944 ( .C ( clk ), .D ( new_AGEMA_signal_17443 ), .Q ( new_AGEMA_signal_17444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5950 ( .C ( clk ), .D ( new_AGEMA_signal_17449 ), .Q ( new_AGEMA_signal_17450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5956 ( .C ( clk ), .D ( new_AGEMA_signal_17455 ), .Q ( new_AGEMA_signal_17456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5962 ( .C ( clk ), .D ( new_AGEMA_signal_17461 ), .Q ( new_AGEMA_signal_17462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5972 ( .C ( clk ), .D ( new_AGEMA_signal_17471 ), .Q ( new_AGEMA_signal_17472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5982 ( .C ( clk ), .D ( new_AGEMA_signal_17481 ), .Q ( new_AGEMA_signal_17482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5992 ( .C ( clk ), .D ( new_AGEMA_signal_17491 ), .Q ( new_AGEMA_signal_17492 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6002 ( .C ( clk ), .D ( new_AGEMA_signal_17501 ), .Q ( new_AGEMA_signal_17502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6008 ( .C ( clk ), .D ( new_AGEMA_signal_17507 ), .Q ( new_AGEMA_signal_17508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6014 ( .C ( clk ), .D ( new_AGEMA_signal_17513 ), .Q ( new_AGEMA_signal_17514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6020 ( .C ( clk ), .D ( new_AGEMA_signal_17519 ), .Q ( new_AGEMA_signal_17520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6026 ( .C ( clk ), .D ( new_AGEMA_signal_17525 ), .Q ( new_AGEMA_signal_17526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6032 ( .C ( clk ), .D ( new_AGEMA_signal_17531 ), .Q ( new_AGEMA_signal_17532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6038 ( .C ( clk ), .D ( new_AGEMA_signal_17537 ), .Q ( new_AGEMA_signal_17538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6044 ( .C ( clk ), .D ( new_AGEMA_signal_17543 ), .Q ( new_AGEMA_signal_17544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6050 ( .C ( clk ), .D ( new_AGEMA_signal_17549 ), .Q ( new_AGEMA_signal_17550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6090 ( .C ( clk ), .D ( new_AGEMA_signal_17589 ), .Q ( new_AGEMA_signal_17590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6098 ( .C ( clk ), .D ( new_AGEMA_signal_17597 ), .Q ( new_AGEMA_signal_17598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6106 ( .C ( clk ), .D ( new_AGEMA_signal_17605 ), .Q ( new_AGEMA_signal_17606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6114 ( .C ( clk ), .D ( new_AGEMA_signal_17613 ), .Q ( new_AGEMA_signal_17614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6120 ( .C ( clk ), .D ( new_AGEMA_signal_17619 ), .Q ( new_AGEMA_signal_17620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6126 ( .C ( clk ), .D ( new_AGEMA_signal_17625 ), .Q ( new_AGEMA_signal_17626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6132 ( .C ( clk ), .D ( new_AGEMA_signal_17631 ), .Q ( new_AGEMA_signal_17632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6138 ( .C ( clk ), .D ( new_AGEMA_signal_17637 ), .Q ( new_AGEMA_signal_17638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6146 ( .C ( clk ), .D ( new_AGEMA_signal_17645 ), .Q ( new_AGEMA_signal_17646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6154 ( .C ( clk ), .D ( new_AGEMA_signal_17653 ), .Q ( new_AGEMA_signal_17654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6162 ( .C ( clk ), .D ( new_AGEMA_signal_17661 ), .Q ( new_AGEMA_signal_17662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6170 ( .C ( clk ), .D ( new_AGEMA_signal_17669 ), .Q ( new_AGEMA_signal_17670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6178 ( .C ( clk ), .D ( new_AGEMA_signal_17677 ), .Q ( new_AGEMA_signal_17678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6186 ( .C ( clk ), .D ( new_AGEMA_signal_17685 ), .Q ( new_AGEMA_signal_17686 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6194 ( .C ( clk ), .D ( new_AGEMA_signal_17693 ), .Q ( new_AGEMA_signal_17694 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6202 ( .C ( clk ), .D ( new_AGEMA_signal_17701 ), .Q ( new_AGEMA_signal_17702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6250 ( .C ( clk ), .D ( new_AGEMA_signal_17749 ), .Q ( new_AGEMA_signal_17750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6258 ( .C ( clk ), .D ( new_AGEMA_signal_17757 ), .Q ( new_AGEMA_signal_17758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6266 ( .C ( clk ), .D ( new_AGEMA_signal_17765 ), .Q ( new_AGEMA_signal_17766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6274 ( .C ( clk ), .D ( new_AGEMA_signal_17773 ), .Q ( new_AGEMA_signal_17774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6296 ( .C ( clk ), .D ( new_AGEMA_signal_17795 ), .Q ( new_AGEMA_signal_17796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6304 ( .C ( clk ), .D ( new_AGEMA_signal_17803 ), .Q ( new_AGEMA_signal_17804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6312 ( .C ( clk ), .D ( new_AGEMA_signal_17811 ), .Q ( new_AGEMA_signal_17812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6320 ( .C ( clk ), .D ( new_AGEMA_signal_17819 ), .Q ( new_AGEMA_signal_17820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6332 ( .C ( clk ), .D ( new_AGEMA_signal_17831 ), .Q ( new_AGEMA_signal_17832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6344 ( .C ( clk ), .D ( new_AGEMA_signal_17843 ), .Q ( new_AGEMA_signal_17844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6356 ( .C ( clk ), .D ( new_AGEMA_signal_17855 ), .Q ( new_AGEMA_signal_17856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6368 ( .C ( clk ), .D ( new_AGEMA_signal_17867 ), .Q ( new_AGEMA_signal_17868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6382 ( .C ( clk ), .D ( new_AGEMA_signal_17881 ), .Q ( new_AGEMA_signal_17882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6396 ( .C ( clk ), .D ( new_AGEMA_signal_17895 ), .Q ( new_AGEMA_signal_17896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6410 ( .C ( clk ), .D ( new_AGEMA_signal_17909 ), .Q ( new_AGEMA_signal_17910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6424 ( .C ( clk ), .D ( new_AGEMA_signal_17923 ), .Q ( new_AGEMA_signal_17924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6432 ( .C ( clk ), .D ( new_AGEMA_signal_17931 ), .Q ( new_AGEMA_signal_17932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6440 ( .C ( clk ), .D ( new_AGEMA_signal_17939 ), .Q ( new_AGEMA_signal_17940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6448 ( .C ( clk ), .D ( new_AGEMA_signal_17947 ), .Q ( new_AGEMA_signal_17948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6456 ( .C ( clk ), .D ( new_AGEMA_signal_17955 ), .Q ( new_AGEMA_signal_17956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6470 ( .C ( clk ), .D ( new_AGEMA_signal_17969 ), .Q ( new_AGEMA_signal_17970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6484 ( .C ( clk ), .D ( new_AGEMA_signal_17983 ), .Q ( new_AGEMA_signal_17984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6498 ( .C ( clk ), .D ( new_AGEMA_signal_17997 ), .Q ( new_AGEMA_signal_17998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6512 ( .C ( clk ), .D ( new_AGEMA_signal_18011 ), .Q ( new_AGEMA_signal_18012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6520 ( .C ( clk ), .D ( new_AGEMA_signal_18019 ), .Q ( new_AGEMA_signal_18020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6528 ( .C ( clk ), .D ( new_AGEMA_signal_18027 ), .Q ( new_AGEMA_signal_18028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6536 ( .C ( clk ), .D ( new_AGEMA_signal_18035 ), .Q ( new_AGEMA_signal_18036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6544 ( .C ( clk ), .D ( new_AGEMA_signal_18043 ), .Q ( new_AGEMA_signal_18044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6552 ( .C ( clk ), .D ( new_AGEMA_signal_18051 ), .Q ( new_AGEMA_signal_18052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6560 ( .C ( clk ), .D ( new_AGEMA_signal_18059 ), .Q ( new_AGEMA_signal_18060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6568 ( .C ( clk ), .D ( new_AGEMA_signal_18067 ), .Q ( new_AGEMA_signal_18068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6576 ( .C ( clk ), .D ( new_AGEMA_signal_18075 ), .Q ( new_AGEMA_signal_18076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6614 ( .C ( clk ), .D ( new_AGEMA_signal_18113 ), .Q ( new_AGEMA_signal_18114 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6630 ( .C ( clk ), .D ( new_AGEMA_signal_18129 ), .Q ( new_AGEMA_signal_18130 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6646 ( .C ( clk ), .D ( new_AGEMA_signal_18145 ), .Q ( new_AGEMA_signal_18146 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6662 ( .C ( clk ), .D ( new_AGEMA_signal_18161 ), .Q ( new_AGEMA_signal_18162 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6702 ( .C ( clk ), .D ( new_AGEMA_signal_18201 ), .Q ( new_AGEMA_signal_18202 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6718 ( .C ( clk ), .D ( new_AGEMA_signal_18217 ), .Q ( new_AGEMA_signal_18218 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6734 ( .C ( clk ), .D ( new_AGEMA_signal_18233 ), .Q ( new_AGEMA_signal_18234 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6750 ( .C ( clk ), .D ( new_AGEMA_signal_18249 ), .Q ( new_AGEMA_signal_18250 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6760 ( .C ( clk ), .D ( new_AGEMA_signal_18259 ), .Q ( new_AGEMA_signal_18260 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6770 ( .C ( clk ), .D ( new_AGEMA_signal_18269 ), .Q ( new_AGEMA_signal_18270 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6780 ( .C ( clk ), .D ( new_AGEMA_signal_18279 ), .Q ( new_AGEMA_signal_18280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6790 ( .C ( clk ), .D ( new_AGEMA_signal_18289 ), .Q ( new_AGEMA_signal_18290 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6900 ( .C ( clk ), .D ( new_AGEMA_signal_18399 ), .Q ( new_AGEMA_signal_18400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6916 ( .C ( clk ), .D ( new_AGEMA_signal_18415 ), .Q ( new_AGEMA_signal_18416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6932 ( .C ( clk ), .D ( new_AGEMA_signal_18431 ), .Q ( new_AGEMA_signal_18432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6948 ( .C ( clk ), .D ( new_AGEMA_signal_18447 ), .Q ( new_AGEMA_signal_18448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7006 ( .C ( clk ), .D ( new_AGEMA_signal_18505 ), .Q ( new_AGEMA_signal_18506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7024 ( .C ( clk ), .D ( new_AGEMA_signal_18523 ), .Q ( new_AGEMA_signal_18524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7042 ( .C ( clk ), .D ( new_AGEMA_signal_18541 ), .Q ( new_AGEMA_signal_18542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7060 ( .C ( clk ), .D ( new_AGEMA_signal_18559 ), .Q ( new_AGEMA_signal_18560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7206 ( .C ( clk ), .D ( new_AGEMA_signal_18705 ), .Q ( new_AGEMA_signal_18706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7226 ( .C ( clk ), .D ( new_AGEMA_signal_18725 ), .Q ( new_AGEMA_signal_18726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7246 ( .C ( clk ), .D ( new_AGEMA_signal_18745 ), .Q ( new_AGEMA_signal_18746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7266 ( .C ( clk ), .D ( new_AGEMA_signal_18765 ), .Q ( new_AGEMA_signal_18766 ) ) ;

    /* cells in depth 15 */
    buf_clk new_AGEMA_reg_buffer_5371 ( .C ( clk ), .D ( new_AGEMA_signal_16870 ), .Q ( new_AGEMA_signal_16871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5377 ( .C ( clk ), .D ( new_AGEMA_signal_16876 ), .Q ( new_AGEMA_signal_16877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5383 ( .C ( clk ), .D ( new_AGEMA_signal_16882 ), .Q ( new_AGEMA_signal_16883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5389 ( .C ( clk ), .D ( new_AGEMA_signal_16888 ), .Q ( new_AGEMA_signal_16889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5395 ( .C ( clk ), .D ( new_AGEMA_signal_16894 ), .Q ( new_AGEMA_signal_16895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5401 ( .C ( clk ), .D ( new_AGEMA_signal_16900 ), .Q ( new_AGEMA_signal_16901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5407 ( .C ( clk ), .D ( new_AGEMA_signal_16906 ), .Q ( new_AGEMA_signal_16907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5413 ( .C ( clk ), .D ( new_AGEMA_signal_16912 ), .Q ( new_AGEMA_signal_16913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5419 ( .C ( clk ), .D ( new_AGEMA_signal_16918 ), .Q ( new_AGEMA_signal_16919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5425 ( .C ( clk ), .D ( new_AGEMA_signal_16924 ), .Q ( new_AGEMA_signal_16925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5431 ( .C ( clk ), .D ( new_AGEMA_signal_16930 ), .Q ( new_AGEMA_signal_16931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5437 ( .C ( clk ), .D ( new_AGEMA_signal_16936 ), .Q ( new_AGEMA_signal_16937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5441 ( .C ( clk ), .D ( new_AGEMA_signal_16940 ), .Q ( new_AGEMA_signal_16941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5445 ( .C ( clk ), .D ( new_AGEMA_signal_16944 ), .Q ( new_AGEMA_signal_16945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5449 ( .C ( clk ), .D ( new_AGEMA_signal_16948 ), .Q ( new_AGEMA_signal_16949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5453 ( .C ( clk ), .D ( new_AGEMA_signal_16952 ), .Q ( new_AGEMA_signal_16953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5461 ( .C ( clk ), .D ( new_AGEMA_signal_16960 ), .Q ( new_AGEMA_signal_16961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5469 ( .C ( clk ), .D ( new_AGEMA_signal_16968 ), .Q ( new_AGEMA_signal_16969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5477 ( .C ( clk ), .D ( new_AGEMA_signal_16976 ), .Q ( new_AGEMA_signal_16977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5485 ( .C ( clk ), .D ( new_AGEMA_signal_16984 ), .Q ( new_AGEMA_signal_16985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5491 ( .C ( clk ), .D ( new_AGEMA_signal_16990 ), .Q ( new_AGEMA_signal_16991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5497 ( .C ( clk ), .D ( new_AGEMA_signal_16996 ), .Q ( new_AGEMA_signal_16997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5503 ( .C ( clk ), .D ( new_AGEMA_signal_17002 ), .Q ( new_AGEMA_signal_17003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5509 ( .C ( clk ), .D ( new_AGEMA_signal_17008 ), .Q ( new_AGEMA_signal_17009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5513 ( .C ( clk ), .D ( new_AGEMA_signal_17012 ), .Q ( new_AGEMA_signal_17013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5517 ( .C ( clk ), .D ( new_AGEMA_signal_17016 ), .Q ( new_AGEMA_signal_17017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5521 ( .C ( clk ), .D ( new_AGEMA_signal_17020 ), .Q ( new_AGEMA_signal_17021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5525 ( .C ( clk ), .D ( new_AGEMA_signal_17024 ), .Q ( new_AGEMA_signal_17025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5533 ( .C ( clk ), .D ( new_AGEMA_signal_17032 ), .Q ( new_AGEMA_signal_17033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5541 ( .C ( clk ), .D ( new_AGEMA_signal_17040 ), .Q ( new_AGEMA_signal_17041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5549 ( .C ( clk ), .D ( new_AGEMA_signal_17048 ), .Q ( new_AGEMA_signal_17049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5557 ( .C ( clk ), .D ( new_AGEMA_signal_17056 ), .Q ( new_AGEMA_signal_17057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5565 ( .C ( clk ), .D ( new_AGEMA_signal_17064 ), .Q ( new_AGEMA_signal_17065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5573 ( .C ( clk ), .D ( new_AGEMA_signal_17072 ), .Q ( new_AGEMA_signal_17073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5581 ( .C ( clk ), .D ( new_AGEMA_signal_17080 ), .Q ( new_AGEMA_signal_17081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5589 ( .C ( clk ), .D ( new_AGEMA_signal_17088 ), .Q ( new_AGEMA_signal_17089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5599 ( .C ( clk ), .D ( new_AGEMA_signal_17098 ), .Q ( new_AGEMA_signal_17099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5609 ( .C ( clk ), .D ( new_AGEMA_signal_17108 ), .Q ( new_AGEMA_signal_17109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5619 ( .C ( clk ), .D ( new_AGEMA_signal_17118 ), .Q ( new_AGEMA_signal_17119 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5629 ( .C ( clk ), .D ( new_AGEMA_signal_17128 ), .Q ( new_AGEMA_signal_17129 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5637 ( .C ( clk ), .D ( new_AGEMA_signal_17136 ), .Q ( new_AGEMA_signal_17137 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5645 ( .C ( clk ), .D ( new_AGEMA_signal_17144 ), .Q ( new_AGEMA_signal_17145 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5653 ( .C ( clk ), .D ( new_AGEMA_signal_17152 ), .Q ( new_AGEMA_signal_17153 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5661 ( .C ( clk ), .D ( new_AGEMA_signal_17160 ), .Q ( new_AGEMA_signal_17161 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5667 ( .C ( clk ), .D ( new_AGEMA_signal_17166 ), .Q ( new_AGEMA_signal_17167 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5673 ( .C ( clk ), .D ( new_AGEMA_signal_17172 ), .Q ( new_AGEMA_signal_17173 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5679 ( .C ( clk ), .D ( new_AGEMA_signal_17178 ), .Q ( new_AGEMA_signal_17179 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5685 ( .C ( clk ), .D ( new_AGEMA_signal_17184 ), .Q ( new_AGEMA_signal_17185 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5689 ( .C ( clk ), .D ( new_AGEMA_signal_17188 ), .Q ( new_AGEMA_signal_17189 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5693 ( .C ( clk ), .D ( new_AGEMA_signal_17192 ), .Q ( new_AGEMA_signal_17193 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5697 ( .C ( clk ), .D ( new_AGEMA_signal_17196 ), .Q ( new_AGEMA_signal_17197 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5701 ( .C ( clk ), .D ( new_AGEMA_signal_17200 ), .Q ( new_AGEMA_signal_17201 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5707 ( .C ( clk ), .D ( new_AGEMA_signal_17206 ), .Q ( new_AGEMA_signal_17207 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5713 ( .C ( clk ), .D ( new_AGEMA_signal_17212 ), .Q ( new_AGEMA_signal_17213 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5719 ( .C ( clk ), .D ( new_AGEMA_signal_17218 ), .Q ( new_AGEMA_signal_17219 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5725 ( .C ( clk ), .D ( new_AGEMA_signal_17224 ), .Q ( new_AGEMA_signal_17225 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5733 ( .C ( clk ), .D ( new_AGEMA_signal_17232 ), .Q ( new_AGEMA_signal_17233 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5741 ( .C ( clk ), .D ( new_AGEMA_signal_17240 ), .Q ( new_AGEMA_signal_17241 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5749 ( .C ( clk ), .D ( new_AGEMA_signal_17248 ), .Q ( new_AGEMA_signal_17249 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5757 ( .C ( clk ), .D ( new_AGEMA_signal_17256 ), .Q ( new_AGEMA_signal_17257 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5763 ( .C ( clk ), .D ( new_AGEMA_signal_17262 ), .Q ( new_AGEMA_signal_17263 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5769 ( .C ( clk ), .D ( new_AGEMA_signal_17268 ), .Q ( new_AGEMA_signal_17269 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5775 ( .C ( clk ), .D ( new_AGEMA_signal_17274 ), .Q ( new_AGEMA_signal_17275 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5781 ( .C ( clk ), .D ( new_AGEMA_signal_17280 ), .Q ( new_AGEMA_signal_17281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5783 ( .C ( clk ), .D ( n2512 ), .Q ( new_AGEMA_signal_17283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5785 ( .C ( clk ), .D ( new_AGEMA_signal_3381 ), .Q ( new_AGEMA_signal_17285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5787 ( .C ( clk ), .D ( new_AGEMA_signal_3382 ), .Q ( new_AGEMA_signal_17287 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5789 ( .C ( clk ), .D ( new_AGEMA_signal_3383 ), .Q ( new_AGEMA_signal_17289 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5797 ( .C ( clk ), .D ( new_AGEMA_signal_17296 ), .Q ( new_AGEMA_signal_17297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5805 ( .C ( clk ), .D ( new_AGEMA_signal_17304 ), .Q ( new_AGEMA_signal_17305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5813 ( .C ( clk ), .D ( new_AGEMA_signal_17312 ), .Q ( new_AGEMA_signal_17313 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5821 ( .C ( clk ), .D ( new_AGEMA_signal_17320 ), .Q ( new_AGEMA_signal_17321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5825 ( .C ( clk ), .D ( new_AGEMA_signal_17324 ), .Q ( new_AGEMA_signal_17325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5829 ( .C ( clk ), .D ( new_AGEMA_signal_17328 ), .Q ( new_AGEMA_signal_17329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5833 ( .C ( clk ), .D ( new_AGEMA_signal_17332 ), .Q ( new_AGEMA_signal_17333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5837 ( .C ( clk ), .D ( new_AGEMA_signal_17336 ), .Q ( new_AGEMA_signal_17337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5843 ( .C ( clk ), .D ( new_AGEMA_signal_17342 ), .Q ( new_AGEMA_signal_17343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5849 ( .C ( clk ), .D ( new_AGEMA_signal_17348 ), .Q ( new_AGEMA_signal_17349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5855 ( .C ( clk ), .D ( new_AGEMA_signal_17354 ), .Q ( new_AGEMA_signal_17355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5861 ( .C ( clk ), .D ( new_AGEMA_signal_17360 ), .Q ( new_AGEMA_signal_17361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5867 ( .C ( clk ), .D ( new_AGEMA_signal_17366 ), .Q ( new_AGEMA_signal_17367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5873 ( .C ( clk ), .D ( new_AGEMA_signal_17372 ), .Q ( new_AGEMA_signal_17373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5879 ( .C ( clk ), .D ( new_AGEMA_signal_17378 ), .Q ( new_AGEMA_signal_17379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5885 ( .C ( clk ), .D ( new_AGEMA_signal_17384 ), .Q ( new_AGEMA_signal_17385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5889 ( .C ( clk ), .D ( new_AGEMA_signal_17388 ), .Q ( new_AGEMA_signal_17389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5893 ( .C ( clk ), .D ( new_AGEMA_signal_17392 ), .Q ( new_AGEMA_signal_17393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5897 ( .C ( clk ), .D ( new_AGEMA_signal_17396 ), .Q ( new_AGEMA_signal_17397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5901 ( .C ( clk ), .D ( new_AGEMA_signal_17400 ), .Q ( new_AGEMA_signal_17401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5905 ( .C ( clk ), .D ( new_AGEMA_signal_17404 ), .Q ( new_AGEMA_signal_17405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5911 ( .C ( clk ), .D ( new_AGEMA_signal_17410 ), .Q ( new_AGEMA_signal_17411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5917 ( .C ( clk ), .D ( new_AGEMA_signal_17416 ), .Q ( new_AGEMA_signal_17417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5923 ( .C ( clk ), .D ( new_AGEMA_signal_17422 ), .Q ( new_AGEMA_signal_17423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5927 ( .C ( clk ), .D ( n2037 ), .Q ( new_AGEMA_signal_17427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5931 ( .C ( clk ), .D ( new_AGEMA_signal_3309 ), .Q ( new_AGEMA_signal_17431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5935 ( .C ( clk ), .D ( new_AGEMA_signal_3310 ), .Q ( new_AGEMA_signal_17435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5939 ( .C ( clk ), .D ( new_AGEMA_signal_3311 ), .Q ( new_AGEMA_signal_17439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5945 ( .C ( clk ), .D ( new_AGEMA_signal_17444 ), .Q ( new_AGEMA_signal_17445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5951 ( .C ( clk ), .D ( new_AGEMA_signal_17450 ), .Q ( new_AGEMA_signal_17451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5957 ( .C ( clk ), .D ( new_AGEMA_signal_17456 ), .Q ( new_AGEMA_signal_17457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5963 ( .C ( clk ), .D ( new_AGEMA_signal_17462 ), .Q ( new_AGEMA_signal_17463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5973 ( .C ( clk ), .D ( new_AGEMA_signal_17472 ), .Q ( new_AGEMA_signal_17473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5983 ( .C ( clk ), .D ( new_AGEMA_signal_17482 ), .Q ( new_AGEMA_signal_17483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5993 ( .C ( clk ), .D ( new_AGEMA_signal_17492 ), .Q ( new_AGEMA_signal_17493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6003 ( .C ( clk ), .D ( new_AGEMA_signal_17502 ), .Q ( new_AGEMA_signal_17503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6009 ( .C ( clk ), .D ( new_AGEMA_signal_17508 ), .Q ( new_AGEMA_signal_17509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6015 ( .C ( clk ), .D ( new_AGEMA_signal_17514 ), .Q ( new_AGEMA_signal_17515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6021 ( .C ( clk ), .D ( new_AGEMA_signal_17520 ), .Q ( new_AGEMA_signal_17521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6027 ( .C ( clk ), .D ( new_AGEMA_signal_17526 ), .Q ( new_AGEMA_signal_17527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6033 ( .C ( clk ), .D ( new_AGEMA_signal_17532 ), .Q ( new_AGEMA_signal_17533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6039 ( .C ( clk ), .D ( new_AGEMA_signal_17538 ), .Q ( new_AGEMA_signal_17539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6045 ( .C ( clk ), .D ( new_AGEMA_signal_17544 ), .Q ( new_AGEMA_signal_17545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6051 ( .C ( clk ), .D ( new_AGEMA_signal_17550 ), .Q ( new_AGEMA_signal_17551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6055 ( .C ( clk ), .D ( n2198 ), .Q ( new_AGEMA_signal_17555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6059 ( .C ( clk ), .D ( new_AGEMA_signal_3336 ), .Q ( new_AGEMA_signal_17559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6063 ( .C ( clk ), .D ( new_AGEMA_signal_3337 ), .Q ( new_AGEMA_signal_17563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6067 ( .C ( clk ), .D ( new_AGEMA_signal_3338 ), .Q ( new_AGEMA_signal_17567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6071 ( .C ( clk ), .D ( n2258 ), .Q ( new_AGEMA_signal_17571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6075 ( .C ( clk ), .D ( new_AGEMA_signal_3459 ), .Q ( new_AGEMA_signal_17575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6079 ( .C ( clk ), .D ( new_AGEMA_signal_3460 ), .Q ( new_AGEMA_signal_17579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6083 ( .C ( clk ), .D ( new_AGEMA_signal_3461 ), .Q ( new_AGEMA_signal_17583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6091 ( .C ( clk ), .D ( new_AGEMA_signal_17590 ), .Q ( new_AGEMA_signal_17591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6099 ( .C ( clk ), .D ( new_AGEMA_signal_17598 ), .Q ( new_AGEMA_signal_17599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6107 ( .C ( clk ), .D ( new_AGEMA_signal_17606 ), .Q ( new_AGEMA_signal_17607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6115 ( .C ( clk ), .D ( new_AGEMA_signal_17614 ), .Q ( new_AGEMA_signal_17615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6121 ( .C ( clk ), .D ( new_AGEMA_signal_17620 ), .Q ( new_AGEMA_signal_17621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6127 ( .C ( clk ), .D ( new_AGEMA_signal_17626 ), .Q ( new_AGEMA_signal_17627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6133 ( .C ( clk ), .D ( new_AGEMA_signal_17632 ), .Q ( new_AGEMA_signal_17633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6139 ( .C ( clk ), .D ( new_AGEMA_signal_17638 ), .Q ( new_AGEMA_signal_17639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6147 ( .C ( clk ), .D ( new_AGEMA_signal_17646 ), .Q ( new_AGEMA_signal_17647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6155 ( .C ( clk ), .D ( new_AGEMA_signal_17654 ), .Q ( new_AGEMA_signal_17655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6163 ( .C ( clk ), .D ( new_AGEMA_signal_17662 ), .Q ( new_AGEMA_signal_17663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6171 ( .C ( clk ), .D ( new_AGEMA_signal_17670 ), .Q ( new_AGEMA_signal_17671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6179 ( .C ( clk ), .D ( new_AGEMA_signal_17678 ), .Q ( new_AGEMA_signal_17679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6187 ( .C ( clk ), .D ( new_AGEMA_signal_17686 ), .Q ( new_AGEMA_signal_17687 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6195 ( .C ( clk ), .D ( new_AGEMA_signal_17694 ), .Q ( new_AGEMA_signal_17695 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6203 ( .C ( clk ), .D ( new_AGEMA_signal_17702 ), .Q ( new_AGEMA_signal_17703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6215 ( .C ( clk ), .D ( n2593 ), .Q ( new_AGEMA_signal_17715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6219 ( .C ( clk ), .D ( new_AGEMA_signal_3396 ), .Q ( new_AGEMA_signal_17719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6223 ( .C ( clk ), .D ( new_AGEMA_signal_3397 ), .Q ( new_AGEMA_signal_17723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6227 ( .C ( clk ), .D ( new_AGEMA_signal_3398 ), .Q ( new_AGEMA_signal_17727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6231 ( .C ( clk ), .D ( n2636 ), .Q ( new_AGEMA_signal_17731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6235 ( .C ( clk ), .D ( new_AGEMA_signal_3405 ), .Q ( new_AGEMA_signal_17735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6239 ( .C ( clk ), .D ( new_AGEMA_signal_3406 ), .Q ( new_AGEMA_signal_17739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6243 ( .C ( clk ), .D ( new_AGEMA_signal_3407 ), .Q ( new_AGEMA_signal_17743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6251 ( .C ( clk ), .D ( new_AGEMA_signal_17750 ), .Q ( new_AGEMA_signal_17751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6259 ( .C ( clk ), .D ( new_AGEMA_signal_17758 ), .Q ( new_AGEMA_signal_17759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6267 ( .C ( clk ), .D ( new_AGEMA_signal_17766 ), .Q ( new_AGEMA_signal_17767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6275 ( .C ( clk ), .D ( new_AGEMA_signal_17774 ), .Q ( new_AGEMA_signal_17775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6279 ( .C ( clk ), .D ( n2806 ), .Q ( new_AGEMA_signal_17779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6283 ( .C ( clk ), .D ( new_AGEMA_signal_3414 ), .Q ( new_AGEMA_signal_17783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6287 ( .C ( clk ), .D ( new_AGEMA_signal_3415 ), .Q ( new_AGEMA_signal_17787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6291 ( .C ( clk ), .D ( new_AGEMA_signal_3416 ), .Q ( new_AGEMA_signal_17791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6297 ( .C ( clk ), .D ( new_AGEMA_signal_17796 ), .Q ( new_AGEMA_signal_17797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6305 ( .C ( clk ), .D ( new_AGEMA_signal_17804 ), .Q ( new_AGEMA_signal_17805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6313 ( .C ( clk ), .D ( new_AGEMA_signal_17812 ), .Q ( new_AGEMA_signal_17813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6321 ( .C ( clk ), .D ( new_AGEMA_signal_17820 ), .Q ( new_AGEMA_signal_17821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6333 ( .C ( clk ), .D ( new_AGEMA_signal_17832 ), .Q ( new_AGEMA_signal_17833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6345 ( .C ( clk ), .D ( new_AGEMA_signal_17844 ), .Q ( new_AGEMA_signal_17845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6357 ( .C ( clk ), .D ( new_AGEMA_signal_17856 ), .Q ( new_AGEMA_signal_17857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6369 ( .C ( clk ), .D ( new_AGEMA_signal_17868 ), .Q ( new_AGEMA_signal_17869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6383 ( .C ( clk ), .D ( new_AGEMA_signal_17882 ), .Q ( new_AGEMA_signal_17883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6397 ( .C ( clk ), .D ( new_AGEMA_signal_17896 ), .Q ( new_AGEMA_signal_17897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6411 ( .C ( clk ), .D ( new_AGEMA_signal_17910 ), .Q ( new_AGEMA_signal_17911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6425 ( .C ( clk ), .D ( new_AGEMA_signal_17924 ), .Q ( new_AGEMA_signal_17925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6433 ( .C ( clk ), .D ( new_AGEMA_signal_17932 ), .Q ( new_AGEMA_signal_17933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6441 ( .C ( clk ), .D ( new_AGEMA_signal_17940 ), .Q ( new_AGEMA_signal_17941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6449 ( .C ( clk ), .D ( new_AGEMA_signal_17948 ), .Q ( new_AGEMA_signal_17949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6457 ( .C ( clk ), .D ( new_AGEMA_signal_17956 ), .Q ( new_AGEMA_signal_17957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6471 ( .C ( clk ), .D ( new_AGEMA_signal_17970 ), .Q ( new_AGEMA_signal_17971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6485 ( .C ( clk ), .D ( new_AGEMA_signal_17984 ), .Q ( new_AGEMA_signal_17985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6499 ( .C ( clk ), .D ( new_AGEMA_signal_17998 ), .Q ( new_AGEMA_signal_17999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6513 ( .C ( clk ), .D ( new_AGEMA_signal_18012 ), .Q ( new_AGEMA_signal_18013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6521 ( .C ( clk ), .D ( new_AGEMA_signal_18020 ), .Q ( new_AGEMA_signal_18021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6529 ( .C ( clk ), .D ( new_AGEMA_signal_18028 ), .Q ( new_AGEMA_signal_18029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6537 ( .C ( clk ), .D ( new_AGEMA_signal_18036 ), .Q ( new_AGEMA_signal_18037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6545 ( .C ( clk ), .D ( new_AGEMA_signal_18044 ), .Q ( new_AGEMA_signal_18045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6553 ( .C ( clk ), .D ( new_AGEMA_signal_18052 ), .Q ( new_AGEMA_signal_18053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6561 ( .C ( clk ), .D ( new_AGEMA_signal_18060 ), .Q ( new_AGEMA_signal_18061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6569 ( .C ( clk ), .D ( new_AGEMA_signal_18068 ), .Q ( new_AGEMA_signal_18069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6577 ( .C ( clk ), .D ( new_AGEMA_signal_18076 ), .Q ( new_AGEMA_signal_18077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6615 ( .C ( clk ), .D ( new_AGEMA_signal_18114 ), .Q ( new_AGEMA_signal_18115 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6631 ( .C ( clk ), .D ( new_AGEMA_signal_18130 ), .Q ( new_AGEMA_signal_18131 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6647 ( .C ( clk ), .D ( new_AGEMA_signal_18146 ), .Q ( new_AGEMA_signal_18147 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6663 ( .C ( clk ), .D ( new_AGEMA_signal_18162 ), .Q ( new_AGEMA_signal_18163 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6703 ( .C ( clk ), .D ( new_AGEMA_signal_18202 ), .Q ( new_AGEMA_signal_18203 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6719 ( .C ( clk ), .D ( new_AGEMA_signal_18218 ), .Q ( new_AGEMA_signal_18219 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6735 ( .C ( clk ), .D ( new_AGEMA_signal_18234 ), .Q ( new_AGEMA_signal_18235 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6751 ( .C ( clk ), .D ( new_AGEMA_signal_18250 ), .Q ( new_AGEMA_signal_18251 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6761 ( .C ( clk ), .D ( new_AGEMA_signal_18260 ), .Q ( new_AGEMA_signal_18261 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6771 ( .C ( clk ), .D ( new_AGEMA_signal_18270 ), .Q ( new_AGEMA_signal_18271 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6781 ( .C ( clk ), .D ( new_AGEMA_signal_18280 ), .Q ( new_AGEMA_signal_18281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6791 ( .C ( clk ), .D ( new_AGEMA_signal_18290 ), .Q ( new_AGEMA_signal_18291 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6815 ( .C ( clk ), .D ( n2829 ), .Q ( new_AGEMA_signal_18315 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6823 ( .C ( clk ), .D ( new_AGEMA_signal_3420 ), .Q ( new_AGEMA_signal_18323 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6831 ( .C ( clk ), .D ( new_AGEMA_signal_3421 ), .Q ( new_AGEMA_signal_18331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6839 ( .C ( clk ), .D ( new_AGEMA_signal_3422 ), .Q ( new_AGEMA_signal_18339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6901 ( .C ( clk ), .D ( new_AGEMA_signal_18400 ), .Q ( new_AGEMA_signal_18401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6917 ( .C ( clk ), .D ( new_AGEMA_signal_18416 ), .Q ( new_AGEMA_signal_18417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6933 ( .C ( clk ), .D ( new_AGEMA_signal_18432 ), .Q ( new_AGEMA_signal_18433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6949 ( .C ( clk ), .D ( new_AGEMA_signal_18448 ), .Q ( new_AGEMA_signal_18449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6959 ( .C ( clk ), .D ( n2312 ), .Q ( new_AGEMA_signal_18459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6969 ( .C ( clk ), .D ( new_AGEMA_signal_3342 ), .Q ( new_AGEMA_signal_18469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6979 ( .C ( clk ), .D ( new_AGEMA_signal_3343 ), .Q ( new_AGEMA_signal_18479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6989 ( .C ( clk ), .D ( new_AGEMA_signal_3344 ), .Q ( new_AGEMA_signal_18489 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7007 ( .C ( clk ), .D ( new_AGEMA_signal_18506 ), .Q ( new_AGEMA_signal_18507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7025 ( .C ( clk ), .D ( new_AGEMA_signal_18524 ), .Q ( new_AGEMA_signal_18525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7043 ( .C ( clk ), .D ( new_AGEMA_signal_18542 ), .Q ( new_AGEMA_signal_18543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7061 ( .C ( clk ), .D ( new_AGEMA_signal_18560 ), .Q ( new_AGEMA_signal_18561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7207 ( .C ( clk ), .D ( new_AGEMA_signal_18706 ), .Q ( new_AGEMA_signal_18707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7227 ( .C ( clk ), .D ( new_AGEMA_signal_18726 ), .Q ( new_AGEMA_signal_18727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7247 ( .C ( clk ), .D ( new_AGEMA_signal_18746 ), .Q ( new_AGEMA_signal_18747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7267 ( .C ( clk ), .D ( new_AGEMA_signal_18766 ), .Q ( new_AGEMA_signal_18767 ) ) ;

    /* cells in depth 16 */
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2003 ( .ina ({new_AGEMA_signal_16250, new_AGEMA_signal_16244, new_AGEMA_signal_16238, new_AGEMA_signal_16232}), .inb ({new_AGEMA_signal_3296, new_AGEMA_signal_3295, new_AGEMA_signal_3294, n1935}), .clk ( clk ), .rnd ({Fresh[7649], Fresh[7648], Fresh[7647], Fresh[7646], Fresh[7645], Fresh[7644], Fresh[7643], Fresh[7642], Fresh[7641], Fresh[7640]}), .outt ({new_AGEMA_signal_3425, new_AGEMA_signal_3424, new_AGEMA_signal_3423, n1941}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2059 ( .ina ({new_AGEMA_signal_3299, new_AGEMA_signal_3298, new_AGEMA_signal_3297, n1959}), .inb ({new_AGEMA_signal_16258, new_AGEMA_signal_16256, new_AGEMA_signal_16254, new_AGEMA_signal_16252}), .clk ( clk ), .rnd ({Fresh[7659], Fresh[7658], Fresh[7657], Fresh[7656], Fresh[7655], Fresh[7654], Fresh[7653], Fresh[7652], Fresh[7651], Fresh[7650]}), .outt ({new_AGEMA_signal_3428, new_AGEMA_signal_3427, new_AGEMA_signal_3426, n1960}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2110 ( .ina ({new_AGEMA_signal_16274, new_AGEMA_signal_16270, new_AGEMA_signal_16266, new_AGEMA_signal_16262}), .inb ({new_AGEMA_signal_3302, new_AGEMA_signal_3301, new_AGEMA_signal_3300, n1983}), .clk ( clk ), .rnd ({Fresh[7669], Fresh[7668], Fresh[7667], Fresh[7666], Fresh[7665], Fresh[7664], Fresh[7663], Fresh[7662], Fresh[7661], Fresh[7660]}), .outt ({new_AGEMA_signal_3431, new_AGEMA_signal_3430, new_AGEMA_signal_3429, n1988}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2153 ( .ina ({new_AGEMA_signal_3305, new_AGEMA_signal_3304, new_AGEMA_signal_3303, n2014}), .inb ({new_AGEMA_signal_16306, new_AGEMA_signal_16298, new_AGEMA_signal_16290, new_AGEMA_signal_16282}), .clk ( clk ), .rnd ({Fresh[7679], Fresh[7678], Fresh[7677], Fresh[7676], Fresh[7675], Fresh[7674], Fresh[7673], Fresh[7672], Fresh[7671], Fresh[7670]}), .outt ({new_AGEMA_signal_3434, new_AGEMA_signal_3433, new_AGEMA_signal_3432, n2015}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2169 ( .ina ({new_AGEMA_signal_3137, new_AGEMA_signal_3136, new_AGEMA_signal_3135, n2029}), .inb ({new_AGEMA_signal_16338, new_AGEMA_signal_16330, new_AGEMA_signal_16322, new_AGEMA_signal_16314}), .clk ( clk ), .rnd ({Fresh[7689], Fresh[7688], Fresh[7687], Fresh[7686], Fresh[7685], Fresh[7684], Fresh[7683], Fresh[7682], Fresh[7681], Fresh[7680]}), .outt ({new_AGEMA_signal_3308, new_AGEMA_signal_3307, new_AGEMA_signal_3306, n2030}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2200 ( .ina ({new_AGEMA_signal_3314, new_AGEMA_signal_3313, new_AGEMA_signal_3312, n2052}), .inb ({new_AGEMA_signal_16370, new_AGEMA_signal_16362, new_AGEMA_signal_16354, new_AGEMA_signal_16346}), .clk ( clk ), .rnd ({Fresh[7699], Fresh[7698], Fresh[7697], Fresh[7696], Fresh[7695], Fresh[7694], Fresh[7693], Fresh[7692], Fresh[7691], Fresh[7690]}), .outt ({new_AGEMA_signal_3440, new_AGEMA_signal_3439, new_AGEMA_signal_3438, n2053}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2222 ( .ina ({new_AGEMA_signal_3317, new_AGEMA_signal_3316, new_AGEMA_signal_3315, n2070}), .inb ({new_AGEMA_signal_16402, new_AGEMA_signal_16394, new_AGEMA_signal_16386, new_AGEMA_signal_16378}), .clk ( clk ), .rnd ({Fresh[7709], Fresh[7708], Fresh[7707], Fresh[7706], Fresh[7705], Fresh[7704], Fresh[7703], Fresh[7702], Fresh[7701], Fresh[7700]}), .outt ({new_AGEMA_signal_3443, new_AGEMA_signal_3442, new_AGEMA_signal_3441, n2071}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2259 ( .ina ({new_AGEMA_signal_16426, new_AGEMA_signal_16420, new_AGEMA_signal_16414, new_AGEMA_signal_16408}), .inb ({new_AGEMA_signal_3320, new_AGEMA_signal_3319, new_AGEMA_signal_3318, n2098}), .clk ( clk ), .rnd ({Fresh[7719], Fresh[7718], Fresh[7717], Fresh[7716], Fresh[7715], Fresh[7714], Fresh[7713], Fresh[7712], Fresh[7711], Fresh[7710]}), .outt ({new_AGEMA_signal_3446, new_AGEMA_signal_3445, new_AGEMA_signal_3444, n2103}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2288 ( .ina ({new_AGEMA_signal_16466, new_AGEMA_signal_16456, new_AGEMA_signal_16446, new_AGEMA_signal_16436}), .inb ({new_AGEMA_signal_3326, new_AGEMA_signal_3325, new_AGEMA_signal_3324, n2125}), .clk ( clk ), .rnd ({Fresh[7729], Fresh[7728], Fresh[7727], Fresh[7726], Fresh[7725], Fresh[7724], Fresh[7723], Fresh[7722], Fresh[7721], Fresh[7720]}), .outt ({new_AGEMA_signal_3449, new_AGEMA_signal_3448, new_AGEMA_signal_3447, n2126}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2314 ( .ina ({new_AGEMA_signal_3329, new_AGEMA_signal_3328, new_AGEMA_signal_3327, n2145}), .inb ({new_AGEMA_signal_16498, new_AGEMA_signal_16490, new_AGEMA_signal_16482, new_AGEMA_signal_16474}), .clk ( clk ), .rnd ({Fresh[7739], Fresh[7738], Fresh[7737], Fresh[7736], Fresh[7735], Fresh[7734], Fresh[7733], Fresh[7732], Fresh[7731], Fresh[7730]}), .outt ({new_AGEMA_signal_3452, new_AGEMA_signal_3451, new_AGEMA_signal_3450, n2146}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2334 ( .ina ({new_AGEMA_signal_16530, new_AGEMA_signal_16522, new_AGEMA_signal_16514, new_AGEMA_signal_16506}), .inb ({new_AGEMA_signal_3332, new_AGEMA_signal_3331, new_AGEMA_signal_3330, n2169}), .clk ( clk ), .rnd ({Fresh[7749], Fresh[7748], Fresh[7747], Fresh[7746], Fresh[7745], Fresh[7744], Fresh[7743], Fresh[7742], Fresh[7741], Fresh[7740]}), .outt ({new_AGEMA_signal_3455, new_AGEMA_signal_3454, new_AGEMA_signal_3453, n2173}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2351 ( .ina ({new_AGEMA_signal_16562, new_AGEMA_signal_16554, new_AGEMA_signal_16546, new_AGEMA_signal_16538}), .inb ({new_AGEMA_signal_3335, new_AGEMA_signal_3334, new_AGEMA_signal_3333, n2185}), .clk ( clk ), .rnd ({Fresh[7759], Fresh[7758], Fresh[7757], Fresh[7756], Fresh[7755], Fresh[7754], Fresh[7753], Fresh[7752], Fresh[7751], Fresh[7750]}), .outt ({new_AGEMA_signal_3458, new_AGEMA_signal_3457, new_AGEMA_signal_3456, n2187}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2416 ( .ina ({new_AGEMA_signal_16570, new_AGEMA_signal_16568, new_AGEMA_signal_16566, new_AGEMA_signal_16564}), .inb ({new_AGEMA_signal_3350, new_AGEMA_signal_3349, new_AGEMA_signal_3348, n2251}), .clk ( clk ), .rnd ({Fresh[7769], Fresh[7768], Fresh[7767], Fresh[7766], Fresh[7765], Fresh[7764], Fresh[7763], Fresh[7762], Fresh[7761], Fresh[7760]}), .outt ({new_AGEMA_signal_3464, new_AGEMA_signal_3463, new_AGEMA_signal_3462, n2256}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2441 ( .ina ({new_AGEMA_signal_3353, new_AGEMA_signal_3352, new_AGEMA_signal_3351, n2274}), .inb ({new_AGEMA_signal_16586, new_AGEMA_signal_16582, new_AGEMA_signal_16578, new_AGEMA_signal_16574}), .clk ( clk ), .rnd ({Fresh[7779], Fresh[7778], Fresh[7777], Fresh[7776], Fresh[7775], Fresh[7774], Fresh[7773], Fresh[7772], Fresh[7771], Fresh[7770]}), .outt ({new_AGEMA_signal_3467, new_AGEMA_signal_3466, new_AGEMA_signal_3465, n2275}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2474 ( .ina ({new_AGEMA_signal_3356, new_AGEMA_signal_3355, new_AGEMA_signal_3354, n2302}), .inb ({new_AGEMA_signal_16610, new_AGEMA_signal_16604, new_AGEMA_signal_16598, new_AGEMA_signal_16592}), .clk ( clk ), .rnd ({Fresh[7789], Fresh[7788], Fresh[7787], Fresh[7786], Fresh[7785], Fresh[7784], Fresh[7783], Fresh[7782], Fresh[7781], Fresh[7780]}), .outt ({new_AGEMA_signal_3470, new_AGEMA_signal_3469, new_AGEMA_signal_3468, n2303}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2504 ( .ina ({new_AGEMA_signal_3359, new_AGEMA_signal_3358, new_AGEMA_signal_3357, n2339}), .inb ({new_AGEMA_signal_3362, new_AGEMA_signal_3361, new_AGEMA_signal_3360, n2338}), .clk ( clk ), .rnd ({Fresh[7799], Fresh[7798], Fresh[7797], Fresh[7796], Fresh[7795], Fresh[7794], Fresh[7793], Fresh[7792], Fresh[7791], Fresh[7790]}), .outt ({new_AGEMA_signal_3473, new_AGEMA_signal_3472, new_AGEMA_signal_3471, n2382}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2516 ( .ina ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, new_AGEMA_signal_3363, n2351}), .inb ({new_AGEMA_signal_16626, new_AGEMA_signal_16622, new_AGEMA_signal_16618, new_AGEMA_signal_16614}), .clk ( clk ), .rnd ({Fresh[7809], Fresh[7808], Fresh[7807], Fresh[7806], Fresh[7805], Fresh[7804], Fresh[7803], Fresh[7802], Fresh[7801], Fresh[7800]}), .outt ({new_AGEMA_signal_3476, new_AGEMA_signal_3475, new_AGEMA_signal_3474, n2380}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2531 ( .ina ({new_AGEMA_signal_3368, new_AGEMA_signal_3367, new_AGEMA_signal_3366, n2365}), .inb ({new_AGEMA_signal_16666, new_AGEMA_signal_16656, new_AGEMA_signal_16646, new_AGEMA_signal_16636}), .clk ( clk ), .rnd ({Fresh[7819], Fresh[7818], Fresh[7817], Fresh[7816], Fresh[7815], Fresh[7814], Fresh[7813], Fresh[7812], Fresh[7811], Fresh[7810]}), .outt ({new_AGEMA_signal_3479, new_AGEMA_signal_3478, new_AGEMA_signal_3477, n2366}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2561 ( .ina ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, new_AGEMA_signal_3213, n2399}), .inb ({new_AGEMA_signal_3371, new_AGEMA_signal_3370, new_AGEMA_signal_3369, n2398}), .clk ( clk ), .rnd ({Fresh[7829], Fresh[7828], Fresh[7827], Fresh[7826], Fresh[7825], Fresh[7824], Fresh[7823], Fresh[7822], Fresh[7821], Fresh[7820]}), .outt ({new_AGEMA_signal_3482, new_AGEMA_signal_3481, new_AGEMA_signal_3480, n2425}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2582 ( .ina ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, new_AGEMA_signal_3219, n2423}), .inb ({new_AGEMA_signal_3224, new_AGEMA_signal_3223, new_AGEMA_signal_3222, n2422}), .clk ( clk ), .rnd ({Fresh[7839], Fresh[7838], Fresh[7837], Fresh[7836], Fresh[7835], Fresh[7834], Fresh[7833], Fresh[7832], Fresh[7831], Fresh[7830]}), .outt ({new_AGEMA_signal_3374, new_AGEMA_signal_3373, new_AGEMA_signal_3372, n2424}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2597 ( .ina ({new_AGEMA_signal_16698, new_AGEMA_signal_16690, new_AGEMA_signal_16682, new_AGEMA_signal_16674}), .inb ({new_AGEMA_signal_3377, new_AGEMA_signal_3376, new_AGEMA_signal_3375, n2441}), .clk ( clk ), .rnd ({Fresh[7849], Fresh[7848], Fresh[7847], Fresh[7846], Fresh[7845], Fresh[7844], Fresh[7843], Fresh[7842], Fresh[7841], Fresh[7840]}), .outt ({new_AGEMA_signal_3485, new_AGEMA_signal_3484, new_AGEMA_signal_3483, n2451}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2631 ( .ina ({new_AGEMA_signal_3233, new_AGEMA_signal_3232, new_AGEMA_signal_3231, n2479}), .inb ({new_AGEMA_signal_16714, new_AGEMA_signal_16710, new_AGEMA_signal_16706, new_AGEMA_signal_16702}), .clk ( clk ), .rnd ({Fresh[7859], Fresh[7858], Fresh[7857], Fresh[7856], Fresh[7855], Fresh[7854], Fresh[7853], Fresh[7852], Fresh[7851], Fresh[7850]}), .outt ({new_AGEMA_signal_3380, new_AGEMA_signal_3379, new_AGEMA_signal_3378, n2514}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2658 ( .ina ({new_AGEMA_signal_3386, new_AGEMA_signal_3385, new_AGEMA_signal_3384, n2510}), .inb ({new_AGEMA_signal_16722, new_AGEMA_signal_16720, new_AGEMA_signal_16718, new_AGEMA_signal_16716}), .clk ( clk ), .rnd ({Fresh[7869], Fresh[7868], Fresh[7867], Fresh[7866], Fresh[7865], Fresh[7864], Fresh[7863], Fresh[7862], Fresh[7861], Fresh[7860]}), .outt ({new_AGEMA_signal_3488, new_AGEMA_signal_3487, new_AGEMA_signal_3486, n2511}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2688 ( .ina ({new_AGEMA_signal_3395, new_AGEMA_signal_3394, new_AGEMA_signal_3393, n2552}), .inb ({new_AGEMA_signal_16754, new_AGEMA_signal_16746, new_AGEMA_signal_16738, new_AGEMA_signal_16730}), .clk ( clk ), .rnd ({Fresh[7879], Fresh[7878], Fresh[7877], Fresh[7876], Fresh[7875], Fresh[7874], Fresh[7873], Fresh[7872], Fresh[7871], Fresh[7870]}), .outt ({new_AGEMA_signal_3491, new_AGEMA_signal_3490, new_AGEMA_signal_3489, n2671}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2716 ( .ina ({new_AGEMA_signal_3401, new_AGEMA_signal_3400, new_AGEMA_signal_3399, n2589}), .inb ({new_AGEMA_signal_16786, new_AGEMA_signal_16778, new_AGEMA_signal_16770, new_AGEMA_signal_16762}), .clk ( clk ), .rnd ({Fresh[7889], Fresh[7888], Fresh[7887], Fresh[7886], Fresh[7885], Fresh[7884], Fresh[7883], Fresh[7882], Fresh[7881], Fresh[7880]}), .outt ({new_AGEMA_signal_3494, new_AGEMA_signal_3493, new_AGEMA_signal_3492, n2590}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2731 ( .ina ({new_AGEMA_signal_3260, new_AGEMA_signal_3259, new_AGEMA_signal_3258, n2608}), .inb ({new_AGEMA_signal_16810, new_AGEMA_signal_16804, new_AGEMA_signal_16798, new_AGEMA_signal_16792}), .clk ( clk ), .rnd ({Fresh[7899], Fresh[7898], Fresh[7897], Fresh[7896], Fresh[7895], Fresh[7894], Fresh[7893], Fresh[7892], Fresh[7891], Fresh[7890]}), .outt ({new_AGEMA_signal_3404, new_AGEMA_signal_3403, new_AGEMA_signal_3402, n2623}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2763 ( .ina ({new_AGEMA_signal_16826, new_AGEMA_signal_16822, new_AGEMA_signal_16818, new_AGEMA_signal_16814}), .inb ({new_AGEMA_signal_3410, new_AGEMA_signal_3409, new_AGEMA_signal_3408, n2659}), .clk ( clk ), .rnd ({Fresh[7909], Fresh[7908], Fresh[7907], Fresh[7906], Fresh[7905], Fresh[7904], Fresh[7903], Fresh[7902], Fresh[7901], Fresh[7900]}), .outt ({new_AGEMA_signal_3500, new_AGEMA_signal_3499, new_AGEMA_signal_3498, n2667}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2786 ( .ina ({new_AGEMA_signal_3413, new_AGEMA_signal_3412, new_AGEMA_signal_3411, n2702}), .inb ({new_AGEMA_signal_16858, new_AGEMA_signal_16850, new_AGEMA_signal_16842, new_AGEMA_signal_16834}), .clk ( clk ), .rnd ({Fresh[7919], Fresh[7918], Fresh[7917], Fresh[7916], Fresh[7915], Fresh[7914], Fresh[7913], Fresh[7912], Fresh[7911], Fresh[7910]}), .outt ({new_AGEMA_signal_3503, new_AGEMA_signal_3502, new_AGEMA_signal_3501, n2703}) ) ;
    mux2_HPC1 #(.security_order(3), .pipeline(1)) U2840 ( .ins ({new_AGEMA_signal_16586, new_AGEMA_signal_16582, new_AGEMA_signal_16578, new_AGEMA_signal_16574}), .inb ({new_AGEMA_signal_16866, new_AGEMA_signal_16864, new_AGEMA_signal_16862, new_AGEMA_signal_16860}), .ina ({new_AGEMA_signal_3290, new_AGEMA_signal_3289, new_AGEMA_signal_3288, n2801}), .clk ( clk ), .rnd ({Fresh[7929], Fresh[7928], Fresh[7927], Fresh[7926], Fresh[7925], Fresh[7924], Fresh[7923], Fresh[7922], Fresh[7921], Fresh[7920]}), .outt ({new_AGEMA_signal_3419, new_AGEMA_signal_3418, new_AGEMA_signal_3417, n2803}) ) ;
    buf_clk new_AGEMA_reg_buffer_5372 ( .C ( clk ), .D ( new_AGEMA_signal_16871 ), .Q ( new_AGEMA_signal_16872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5378 ( .C ( clk ), .D ( new_AGEMA_signal_16877 ), .Q ( new_AGEMA_signal_16878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5384 ( .C ( clk ), .D ( new_AGEMA_signal_16883 ), .Q ( new_AGEMA_signal_16884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5390 ( .C ( clk ), .D ( new_AGEMA_signal_16889 ), .Q ( new_AGEMA_signal_16890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5396 ( .C ( clk ), .D ( new_AGEMA_signal_16895 ), .Q ( new_AGEMA_signal_16896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5402 ( .C ( clk ), .D ( new_AGEMA_signal_16901 ), .Q ( new_AGEMA_signal_16902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5408 ( .C ( clk ), .D ( new_AGEMA_signal_16907 ), .Q ( new_AGEMA_signal_16908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5414 ( .C ( clk ), .D ( new_AGEMA_signal_16913 ), .Q ( new_AGEMA_signal_16914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5420 ( .C ( clk ), .D ( new_AGEMA_signal_16919 ), .Q ( new_AGEMA_signal_16920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5426 ( .C ( clk ), .D ( new_AGEMA_signal_16925 ), .Q ( new_AGEMA_signal_16926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5432 ( .C ( clk ), .D ( new_AGEMA_signal_16931 ), .Q ( new_AGEMA_signal_16932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5438 ( .C ( clk ), .D ( new_AGEMA_signal_16937 ), .Q ( new_AGEMA_signal_16938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5442 ( .C ( clk ), .D ( new_AGEMA_signal_16941 ), .Q ( new_AGEMA_signal_16942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5446 ( .C ( clk ), .D ( new_AGEMA_signal_16945 ), .Q ( new_AGEMA_signal_16946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5450 ( .C ( clk ), .D ( new_AGEMA_signal_16949 ), .Q ( new_AGEMA_signal_16950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5454 ( .C ( clk ), .D ( new_AGEMA_signal_16953 ), .Q ( new_AGEMA_signal_16954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5462 ( .C ( clk ), .D ( new_AGEMA_signal_16961 ), .Q ( new_AGEMA_signal_16962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5470 ( .C ( clk ), .D ( new_AGEMA_signal_16969 ), .Q ( new_AGEMA_signal_16970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5478 ( .C ( clk ), .D ( new_AGEMA_signal_16977 ), .Q ( new_AGEMA_signal_16978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5486 ( .C ( clk ), .D ( new_AGEMA_signal_16985 ), .Q ( new_AGEMA_signal_16986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5492 ( .C ( clk ), .D ( new_AGEMA_signal_16991 ), .Q ( new_AGEMA_signal_16992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5498 ( .C ( clk ), .D ( new_AGEMA_signal_16997 ), .Q ( new_AGEMA_signal_16998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5504 ( .C ( clk ), .D ( new_AGEMA_signal_17003 ), .Q ( new_AGEMA_signal_17004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5510 ( .C ( clk ), .D ( new_AGEMA_signal_17009 ), .Q ( new_AGEMA_signal_17010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5514 ( .C ( clk ), .D ( new_AGEMA_signal_17013 ), .Q ( new_AGEMA_signal_17014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5518 ( .C ( clk ), .D ( new_AGEMA_signal_17017 ), .Q ( new_AGEMA_signal_17018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5522 ( .C ( clk ), .D ( new_AGEMA_signal_17021 ), .Q ( new_AGEMA_signal_17022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5526 ( .C ( clk ), .D ( new_AGEMA_signal_17025 ), .Q ( new_AGEMA_signal_17026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5534 ( .C ( clk ), .D ( new_AGEMA_signal_17033 ), .Q ( new_AGEMA_signal_17034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5542 ( .C ( clk ), .D ( new_AGEMA_signal_17041 ), .Q ( new_AGEMA_signal_17042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5550 ( .C ( clk ), .D ( new_AGEMA_signal_17049 ), .Q ( new_AGEMA_signal_17050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5558 ( .C ( clk ), .D ( new_AGEMA_signal_17057 ), .Q ( new_AGEMA_signal_17058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5566 ( .C ( clk ), .D ( new_AGEMA_signal_17065 ), .Q ( new_AGEMA_signal_17066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5574 ( .C ( clk ), .D ( new_AGEMA_signal_17073 ), .Q ( new_AGEMA_signal_17074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5582 ( .C ( clk ), .D ( new_AGEMA_signal_17081 ), .Q ( new_AGEMA_signal_17082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5590 ( .C ( clk ), .D ( new_AGEMA_signal_17089 ), .Q ( new_AGEMA_signal_17090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5600 ( .C ( clk ), .D ( new_AGEMA_signal_17099 ), .Q ( new_AGEMA_signal_17100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5610 ( .C ( clk ), .D ( new_AGEMA_signal_17109 ), .Q ( new_AGEMA_signal_17110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5620 ( .C ( clk ), .D ( new_AGEMA_signal_17119 ), .Q ( new_AGEMA_signal_17120 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5630 ( .C ( clk ), .D ( new_AGEMA_signal_17129 ), .Q ( new_AGEMA_signal_17130 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5638 ( .C ( clk ), .D ( new_AGEMA_signal_17137 ), .Q ( new_AGEMA_signal_17138 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5646 ( .C ( clk ), .D ( new_AGEMA_signal_17145 ), .Q ( new_AGEMA_signal_17146 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5654 ( .C ( clk ), .D ( new_AGEMA_signal_17153 ), .Q ( new_AGEMA_signal_17154 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5662 ( .C ( clk ), .D ( new_AGEMA_signal_17161 ), .Q ( new_AGEMA_signal_17162 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5668 ( .C ( clk ), .D ( new_AGEMA_signal_17167 ), .Q ( new_AGEMA_signal_17168 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5674 ( .C ( clk ), .D ( new_AGEMA_signal_17173 ), .Q ( new_AGEMA_signal_17174 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5680 ( .C ( clk ), .D ( new_AGEMA_signal_17179 ), .Q ( new_AGEMA_signal_17180 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5686 ( .C ( clk ), .D ( new_AGEMA_signal_17185 ), .Q ( new_AGEMA_signal_17186 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5690 ( .C ( clk ), .D ( new_AGEMA_signal_17189 ), .Q ( new_AGEMA_signal_17190 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5694 ( .C ( clk ), .D ( new_AGEMA_signal_17193 ), .Q ( new_AGEMA_signal_17194 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5698 ( .C ( clk ), .D ( new_AGEMA_signal_17197 ), .Q ( new_AGEMA_signal_17198 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5702 ( .C ( clk ), .D ( new_AGEMA_signal_17201 ), .Q ( new_AGEMA_signal_17202 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5708 ( .C ( clk ), .D ( new_AGEMA_signal_17207 ), .Q ( new_AGEMA_signal_17208 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5714 ( .C ( clk ), .D ( new_AGEMA_signal_17213 ), .Q ( new_AGEMA_signal_17214 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5720 ( .C ( clk ), .D ( new_AGEMA_signal_17219 ), .Q ( new_AGEMA_signal_17220 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5726 ( .C ( clk ), .D ( new_AGEMA_signal_17225 ), .Q ( new_AGEMA_signal_17226 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5734 ( .C ( clk ), .D ( new_AGEMA_signal_17233 ), .Q ( new_AGEMA_signal_17234 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5742 ( .C ( clk ), .D ( new_AGEMA_signal_17241 ), .Q ( new_AGEMA_signal_17242 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5750 ( .C ( clk ), .D ( new_AGEMA_signal_17249 ), .Q ( new_AGEMA_signal_17250 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5758 ( .C ( clk ), .D ( new_AGEMA_signal_17257 ), .Q ( new_AGEMA_signal_17258 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5764 ( .C ( clk ), .D ( new_AGEMA_signal_17263 ), .Q ( new_AGEMA_signal_17264 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5770 ( .C ( clk ), .D ( new_AGEMA_signal_17269 ), .Q ( new_AGEMA_signal_17270 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5776 ( .C ( clk ), .D ( new_AGEMA_signal_17275 ), .Q ( new_AGEMA_signal_17276 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5782 ( .C ( clk ), .D ( new_AGEMA_signal_17281 ), .Q ( new_AGEMA_signal_17282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5784 ( .C ( clk ), .D ( new_AGEMA_signal_17283 ), .Q ( new_AGEMA_signal_17284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5786 ( .C ( clk ), .D ( new_AGEMA_signal_17285 ), .Q ( new_AGEMA_signal_17286 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5788 ( .C ( clk ), .D ( new_AGEMA_signal_17287 ), .Q ( new_AGEMA_signal_17288 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5790 ( .C ( clk ), .D ( new_AGEMA_signal_17289 ), .Q ( new_AGEMA_signal_17290 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5798 ( .C ( clk ), .D ( new_AGEMA_signal_17297 ), .Q ( new_AGEMA_signal_17298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5806 ( .C ( clk ), .D ( new_AGEMA_signal_17305 ), .Q ( new_AGEMA_signal_17306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5814 ( .C ( clk ), .D ( new_AGEMA_signal_17313 ), .Q ( new_AGEMA_signal_17314 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5822 ( .C ( clk ), .D ( new_AGEMA_signal_17321 ), .Q ( new_AGEMA_signal_17322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5826 ( .C ( clk ), .D ( new_AGEMA_signal_17325 ), .Q ( new_AGEMA_signal_17326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5830 ( .C ( clk ), .D ( new_AGEMA_signal_17329 ), .Q ( new_AGEMA_signal_17330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5834 ( .C ( clk ), .D ( new_AGEMA_signal_17333 ), .Q ( new_AGEMA_signal_17334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5838 ( .C ( clk ), .D ( new_AGEMA_signal_17337 ), .Q ( new_AGEMA_signal_17338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5844 ( .C ( clk ), .D ( new_AGEMA_signal_17343 ), .Q ( new_AGEMA_signal_17344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5850 ( .C ( clk ), .D ( new_AGEMA_signal_17349 ), .Q ( new_AGEMA_signal_17350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5856 ( .C ( clk ), .D ( new_AGEMA_signal_17355 ), .Q ( new_AGEMA_signal_17356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5862 ( .C ( clk ), .D ( new_AGEMA_signal_17361 ), .Q ( new_AGEMA_signal_17362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5868 ( .C ( clk ), .D ( new_AGEMA_signal_17367 ), .Q ( new_AGEMA_signal_17368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5874 ( .C ( clk ), .D ( new_AGEMA_signal_17373 ), .Q ( new_AGEMA_signal_17374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5880 ( .C ( clk ), .D ( new_AGEMA_signal_17379 ), .Q ( new_AGEMA_signal_17380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5886 ( .C ( clk ), .D ( new_AGEMA_signal_17385 ), .Q ( new_AGEMA_signal_17386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5890 ( .C ( clk ), .D ( new_AGEMA_signal_17389 ), .Q ( new_AGEMA_signal_17390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5894 ( .C ( clk ), .D ( new_AGEMA_signal_17393 ), .Q ( new_AGEMA_signal_17394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5898 ( .C ( clk ), .D ( new_AGEMA_signal_17397 ), .Q ( new_AGEMA_signal_17398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5902 ( .C ( clk ), .D ( new_AGEMA_signal_17401 ), .Q ( new_AGEMA_signal_17402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5906 ( .C ( clk ), .D ( new_AGEMA_signal_17405 ), .Q ( new_AGEMA_signal_17406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5912 ( .C ( clk ), .D ( new_AGEMA_signal_17411 ), .Q ( new_AGEMA_signal_17412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5918 ( .C ( clk ), .D ( new_AGEMA_signal_17417 ), .Q ( new_AGEMA_signal_17418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5924 ( .C ( clk ), .D ( new_AGEMA_signal_17423 ), .Q ( new_AGEMA_signal_17424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5928 ( .C ( clk ), .D ( new_AGEMA_signal_17427 ), .Q ( new_AGEMA_signal_17428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5932 ( .C ( clk ), .D ( new_AGEMA_signal_17431 ), .Q ( new_AGEMA_signal_17432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5936 ( .C ( clk ), .D ( new_AGEMA_signal_17435 ), .Q ( new_AGEMA_signal_17436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5940 ( .C ( clk ), .D ( new_AGEMA_signal_17439 ), .Q ( new_AGEMA_signal_17440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5946 ( .C ( clk ), .D ( new_AGEMA_signal_17445 ), .Q ( new_AGEMA_signal_17446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5952 ( .C ( clk ), .D ( new_AGEMA_signal_17451 ), .Q ( new_AGEMA_signal_17452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5958 ( .C ( clk ), .D ( new_AGEMA_signal_17457 ), .Q ( new_AGEMA_signal_17458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5964 ( .C ( clk ), .D ( new_AGEMA_signal_17463 ), .Q ( new_AGEMA_signal_17464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5974 ( .C ( clk ), .D ( new_AGEMA_signal_17473 ), .Q ( new_AGEMA_signal_17474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5984 ( .C ( clk ), .D ( new_AGEMA_signal_17483 ), .Q ( new_AGEMA_signal_17484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5994 ( .C ( clk ), .D ( new_AGEMA_signal_17493 ), .Q ( new_AGEMA_signal_17494 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6004 ( .C ( clk ), .D ( new_AGEMA_signal_17503 ), .Q ( new_AGEMA_signal_17504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6010 ( .C ( clk ), .D ( new_AGEMA_signal_17509 ), .Q ( new_AGEMA_signal_17510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6016 ( .C ( clk ), .D ( new_AGEMA_signal_17515 ), .Q ( new_AGEMA_signal_17516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6022 ( .C ( clk ), .D ( new_AGEMA_signal_17521 ), .Q ( new_AGEMA_signal_17522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6028 ( .C ( clk ), .D ( new_AGEMA_signal_17527 ), .Q ( new_AGEMA_signal_17528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6034 ( .C ( clk ), .D ( new_AGEMA_signal_17533 ), .Q ( new_AGEMA_signal_17534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6040 ( .C ( clk ), .D ( new_AGEMA_signal_17539 ), .Q ( new_AGEMA_signal_17540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6046 ( .C ( clk ), .D ( new_AGEMA_signal_17545 ), .Q ( new_AGEMA_signal_17546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6052 ( .C ( clk ), .D ( new_AGEMA_signal_17551 ), .Q ( new_AGEMA_signal_17552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6056 ( .C ( clk ), .D ( new_AGEMA_signal_17555 ), .Q ( new_AGEMA_signal_17556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6060 ( .C ( clk ), .D ( new_AGEMA_signal_17559 ), .Q ( new_AGEMA_signal_17560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6064 ( .C ( clk ), .D ( new_AGEMA_signal_17563 ), .Q ( new_AGEMA_signal_17564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6068 ( .C ( clk ), .D ( new_AGEMA_signal_17567 ), .Q ( new_AGEMA_signal_17568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6072 ( .C ( clk ), .D ( new_AGEMA_signal_17571 ), .Q ( new_AGEMA_signal_17572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6076 ( .C ( clk ), .D ( new_AGEMA_signal_17575 ), .Q ( new_AGEMA_signal_17576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6080 ( .C ( clk ), .D ( new_AGEMA_signal_17579 ), .Q ( new_AGEMA_signal_17580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6084 ( .C ( clk ), .D ( new_AGEMA_signal_17583 ), .Q ( new_AGEMA_signal_17584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6092 ( .C ( clk ), .D ( new_AGEMA_signal_17591 ), .Q ( new_AGEMA_signal_17592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6100 ( .C ( clk ), .D ( new_AGEMA_signal_17599 ), .Q ( new_AGEMA_signal_17600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6108 ( .C ( clk ), .D ( new_AGEMA_signal_17607 ), .Q ( new_AGEMA_signal_17608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6116 ( .C ( clk ), .D ( new_AGEMA_signal_17615 ), .Q ( new_AGEMA_signal_17616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6122 ( .C ( clk ), .D ( new_AGEMA_signal_17621 ), .Q ( new_AGEMA_signal_17622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6128 ( .C ( clk ), .D ( new_AGEMA_signal_17627 ), .Q ( new_AGEMA_signal_17628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6134 ( .C ( clk ), .D ( new_AGEMA_signal_17633 ), .Q ( new_AGEMA_signal_17634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6140 ( .C ( clk ), .D ( new_AGEMA_signal_17639 ), .Q ( new_AGEMA_signal_17640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6148 ( .C ( clk ), .D ( new_AGEMA_signal_17647 ), .Q ( new_AGEMA_signal_17648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6156 ( .C ( clk ), .D ( new_AGEMA_signal_17655 ), .Q ( new_AGEMA_signal_17656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6164 ( .C ( clk ), .D ( new_AGEMA_signal_17663 ), .Q ( new_AGEMA_signal_17664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6172 ( .C ( clk ), .D ( new_AGEMA_signal_17671 ), .Q ( new_AGEMA_signal_17672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6180 ( .C ( clk ), .D ( new_AGEMA_signal_17679 ), .Q ( new_AGEMA_signal_17680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6188 ( .C ( clk ), .D ( new_AGEMA_signal_17687 ), .Q ( new_AGEMA_signal_17688 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6196 ( .C ( clk ), .D ( new_AGEMA_signal_17695 ), .Q ( new_AGEMA_signal_17696 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6204 ( .C ( clk ), .D ( new_AGEMA_signal_17703 ), .Q ( new_AGEMA_signal_17704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6216 ( .C ( clk ), .D ( new_AGEMA_signal_17715 ), .Q ( new_AGEMA_signal_17716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6220 ( .C ( clk ), .D ( new_AGEMA_signal_17719 ), .Q ( new_AGEMA_signal_17720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6224 ( .C ( clk ), .D ( new_AGEMA_signal_17723 ), .Q ( new_AGEMA_signal_17724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6228 ( .C ( clk ), .D ( new_AGEMA_signal_17727 ), .Q ( new_AGEMA_signal_17728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6232 ( .C ( clk ), .D ( new_AGEMA_signal_17731 ), .Q ( new_AGEMA_signal_17732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6236 ( .C ( clk ), .D ( new_AGEMA_signal_17735 ), .Q ( new_AGEMA_signal_17736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6240 ( .C ( clk ), .D ( new_AGEMA_signal_17739 ), .Q ( new_AGEMA_signal_17740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6244 ( .C ( clk ), .D ( new_AGEMA_signal_17743 ), .Q ( new_AGEMA_signal_17744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6252 ( .C ( clk ), .D ( new_AGEMA_signal_17751 ), .Q ( new_AGEMA_signal_17752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6260 ( .C ( clk ), .D ( new_AGEMA_signal_17759 ), .Q ( new_AGEMA_signal_17760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6268 ( .C ( clk ), .D ( new_AGEMA_signal_17767 ), .Q ( new_AGEMA_signal_17768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6276 ( .C ( clk ), .D ( new_AGEMA_signal_17775 ), .Q ( new_AGEMA_signal_17776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6280 ( .C ( clk ), .D ( new_AGEMA_signal_17779 ), .Q ( new_AGEMA_signal_17780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6284 ( .C ( clk ), .D ( new_AGEMA_signal_17783 ), .Q ( new_AGEMA_signal_17784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6288 ( .C ( clk ), .D ( new_AGEMA_signal_17787 ), .Q ( new_AGEMA_signal_17788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6292 ( .C ( clk ), .D ( new_AGEMA_signal_17791 ), .Q ( new_AGEMA_signal_17792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6298 ( .C ( clk ), .D ( new_AGEMA_signal_17797 ), .Q ( new_AGEMA_signal_17798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6306 ( .C ( clk ), .D ( new_AGEMA_signal_17805 ), .Q ( new_AGEMA_signal_17806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6314 ( .C ( clk ), .D ( new_AGEMA_signal_17813 ), .Q ( new_AGEMA_signal_17814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6322 ( .C ( clk ), .D ( new_AGEMA_signal_17821 ), .Q ( new_AGEMA_signal_17822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6334 ( .C ( clk ), .D ( new_AGEMA_signal_17833 ), .Q ( new_AGEMA_signal_17834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6346 ( .C ( clk ), .D ( new_AGEMA_signal_17845 ), .Q ( new_AGEMA_signal_17846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6358 ( .C ( clk ), .D ( new_AGEMA_signal_17857 ), .Q ( new_AGEMA_signal_17858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6370 ( .C ( clk ), .D ( new_AGEMA_signal_17869 ), .Q ( new_AGEMA_signal_17870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6384 ( .C ( clk ), .D ( new_AGEMA_signal_17883 ), .Q ( new_AGEMA_signal_17884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6398 ( .C ( clk ), .D ( new_AGEMA_signal_17897 ), .Q ( new_AGEMA_signal_17898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6412 ( .C ( clk ), .D ( new_AGEMA_signal_17911 ), .Q ( new_AGEMA_signal_17912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6426 ( .C ( clk ), .D ( new_AGEMA_signal_17925 ), .Q ( new_AGEMA_signal_17926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6434 ( .C ( clk ), .D ( new_AGEMA_signal_17933 ), .Q ( new_AGEMA_signal_17934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6442 ( .C ( clk ), .D ( new_AGEMA_signal_17941 ), .Q ( new_AGEMA_signal_17942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6450 ( .C ( clk ), .D ( new_AGEMA_signal_17949 ), .Q ( new_AGEMA_signal_17950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6458 ( .C ( clk ), .D ( new_AGEMA_signal_17957 ), .Q ( new_AGEMA_signal_17958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6472 ( .C ( clk ), .D ( new_AGEMA_signal_17971 ), .Q ( new_AGEMA_signal_17972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6486 ( .C ( clk ), .D ( new_AGEMA_signal_17985 ), .Q ( new_AGEMA_signal_17986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6500 ( .C ( clk ), .D ( new_AGEMA_signal_17999 ), .Q ( new_AGEMA_signal_18000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6514 ( .C ( clk ), .D ( new_AGEMA_signal_18013 ), .Q ( new_AGEMA_signal_18014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6522 ( .C ( clk ), .D ( new_AGEMA_signal_18021 ), .Q ( new_AGEMA_signal_18022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6530 ( .C ( clk ), .D ( new_AGEMA_signal_18029 ), .Q ( new_AGEMA_signal_18030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6538 ( .C ( clk ), .D ( new_AGEMA_signal_18037 ), .Q ( new_AGEMA_signal_18038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6546 ( .C ( clk ), .D ( new_AGEMA_signal_18045 ), .Q ( new_AGEMA_signal_18046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6554 ( .C ( clk ), .D ( new_AGEMA_signal_18053 ), .Q ( new_AGEMA_signal_18054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6562 ( .C ( clk ), .D ( new_AGEMA_signal_18061 ), .Q ( new_AGEMA_signal_18062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6570 ( .C ( clk ), .D ( new_AGEMA_signal_18069 ), .Q ( new_AGEMA_signal_18070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6578 ( .C ( clk ), .D ( new_AGEMA_signal_18077 ), .Q ( new_AGEMA_signal_18078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6616 ( .C ( clk ), .D ( new_AGEMA_signal_18115 ), .Q ( new_AGEMA_signal_18116 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6632 ( .C ( clk ), .D ( new_AGEMA_signal_18131 ), .Q ( new_AGEMA_signal_18132 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6648 ( .C ( clk ), .D ( new_AGEMA_signal_18147 ), .Q ( new_AGEMA_signal_18148 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6664 ( .C ( clk ), .D ( new_AGEMA_signal_18163 ), .Q ( new_AGEMA_signal_18164 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6704 ( .C ( clk ), .D ( new_AGEMA_signal_18203 ), .Q ( new_AGEMA_signal_18204 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6720 ( .C ( clk ), .D ( new_AGEMA_signal_18219 ), .Q ( new_AGEMA_signal_18220 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6736 ( .C ( clk ), .D ( new_AGEMA_signal_18235 ), .Q ( new_AGEMA_signal_18236 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6752 ( .C ( clk ), .D ( new_AGEMA_signal_18251 ), .Q ( new_AGEMA_signal_18252 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6762 ( .C ( clk ), .D ( new_AGEMA_signal_18261 ), .Q ( new_AGEMA_signal_18262 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6772 ( .C ( clk ), .D ( new_AGEMA_signal_18271 ), .Q ( new_AGEMA_signal_18272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6782 ( .C ( clk ), .D ( new_AGEMA_signal_18281 ), .Q ( new_AGEMA_signal_18282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6792 ( .C ( clk ), .D ( new_AGEMA_signal_18291 ), .Q ( new_AGEMA_signal_18292 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6816 ( .C ( clk ), .D ( new_AGEMA_signal_18315 ), .Q ( new_AGEMA_signal_18316 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6824 ( .C ( clk ), .D ( new_AGEMA_signal_18323 ), .Q ( new_AGEMA_signal_18324 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6832 ( .C ( clk ), .D ( new_AGEMA_signal_18331 ), .Q ( new_AGEMA_signal_18332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6840 ( .C ( clk ), .D ( new_AGEMA_signal_18339 ), .Q ( new_AGEMA_signal_18340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6902 ( .C ( clk ), .D ( new_AGEMA_signal_18401 ), .Q ( new_AGEMA_signal_18402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6918 ( .C ( clk ), .D ( new_AGEMA_signal_18417 ), .Q ( new_AGEMA_signal_18418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6934 ( .C ( clk ), .D ( new_AGEMA_signal_18433 ), .Q ( new_AGEMA_signal_18434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6950 ( .C ( clk ), .D ( new_AGEMA_signal_18449 ), .Q ( new_AGEMA_signal_18450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6960 ( .C ( clk ), .D ( new_AGEMA_signal_18459 ), .Q ( new_AGEMA_signal_18460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6970 ( .C ( clk ), .D ( new_AGEMA_signal_18469 ), .Q ( new_AGEMA_signal_18470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6980 ( .C ( clk ), .D ( new_AGEMA_signal_18479 ), .Q ( new_AGEMA_signal_18480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6990 ( .C ( clk ), .D ( new_AGEMA_signal_18489 ), .Q ( new_AGEMA_signal_18490 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7008 ( .C ( clk ), .D ( new_AGEMA_signal_18507 ), .Q ( new_AGEMA_signal_18508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7026 ( .C ( clk ), .D ( new_AGEMA_signal_18525 ), .Q ( new_AGEMA_signal_18526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7044 ( .C ( clk ), .D ( new_AGEMA_signal_18543 ), .Q ( new_AGEMA_signal_18544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7062 ( .C ( clk ), .D ( new_AGEMA_signal_18561 ), .Q ( new_AGEMA_signal_18562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7208 ( .C ( clk ), .D ( new_AGEMA_signal_18707 ), .Q ( new_AGEMA_signal_18708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7228 ( .C ( clk ), .D ( new_AGEMA_signal_18727 ), .Q ( new_AGEMA_signal_18728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7248 ( .C ( clk ), .D ( new_AGEMA_signal_18747 ), .Q ( new_AGEMA_signal_18748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7268 ( .C ( clk ), .D ( new_AGEMA_signal_18767 ), .Q ( new_AGEMA_signal_18768 ) ) ;

    /* cells in depth 17 */
    buf_clk new_AGEMA_reg_buffer_5907 ( .C ( clk ), .D ( new_AGEMA_signal_17406 ), .Q ( new_AGEMA_signal_17407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5913 ( .C ( clk ), .D ( new_AGEMA_signal_17412 ), .Q ( new_AGEMA_signal_17413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5919 ( .C ( clk ), .D ( new_AGEMA_signal_17418 ), .Q ( new_AGEMA_signal_17419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5925 ( .C ( clk ), .D ( new_AGEMA_signal_17424 ), .Q ( new_AGEMA_signal_17425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5929 ( .C ( clk ), .D ( new_AGEMA_signal_17428 ), .Q ( new_AGEMA_signal_17429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5933 ( .C ( clk ), .D ( new_AGEMA_signal_17432 ), .Q ( new_AGEMA_signal_17433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5937 ( .C ( clk ), .D ( new_AGEMA_signal_17436 ), .Q ( new_AGEMA_signal_17437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5941 ( .C ( clk ), .D ( new_AGEMA_signal_17440 ), .Q ( new_AGEMA_signal_17441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5947 ( .C ( clk ), .D ( new_AGEMA_signal_17446 ), .Q ( new_AGEMA_signal_17447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5953 ( .C ( clk ), .D ( new_AGEMA_signal_17452 ), .Q ( new_AGEMA_signal_17453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5959 ( .C ( clk ), .D ( new_AGEMA_signal_17458 ), .Q ( new_AGEMA_signal_17459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5965 ( .C ( clk ), .D ( new_AGEMA_signal_17464 ), .Q ( new_AGEMA_signal_17465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5975 ( .C ( clk ), .D ( new_AGEMA_signal_17474 ), .Q ( new_AGEMA_signal_17475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5985 ( .C ( clk ), .D ( new_AGEMA_signal_17484 ), .Q ( new_AGEMA_signal_17485 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5995 ( .C ( clk ), .D ( new_AGEMA_signal_17494 ), .Q ( new_AGEMA_signal_17495 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6005 ( .C ( clk ), .D ( new_AGEMA_signal_17504 ), .Q ( new_AGEMA_signal_17505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6011 ( .C ( clk ), .D ( new_AGEMA_signal_17510 ), .Q ( new_AGEMA_signal_17511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6017 ( .C ( clk ), .D ( new_AGEMA_signal_17516 ), .Q ( new_AGEMA_signal_17517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6023 ( .C ( clk ), .D ( new_AGEMA_signal_17522 ), .Q ( new_AGEMA_signal_17523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6029 ( .C ( clk ), .D ( new_AGEMA_signal_17528 ), .Q ( new_AGEMA_signal_17529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6035 ( .C ( clk ), .D ( new_AGEMA_signal_17534 ), .Q ( new_AGEMA_signal_17535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6041 ( .C ( clk ), .D ( new_AGEMA_signal_17540 ), .Q ( new_AGEMA_signal_17541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6047 ( .C ( clk ), .D ( new_AGEMA_signal_17546 ), .Q ( new_AGEMA_signal_17547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6053 ( .C ( clk ), .D ( new_AGEMA_signal_17552 ), .Q ( new_AGEMA_signal_17553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6057 ( .C ( clk ), .D ( new_AGEMA_signal_17556 ), .Q ( new_AGEMA_signal_17557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6061 ( .C ( clk ), .D ( new_AGEMA_signal_17560 ), .Q ( new_AGEMA_signal_17561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6065 ( .C ( clk ), .D ( new_AGEMA_signal_17564 ), .Q ( new_AGEMA_signal_17565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6069 ( .C ( clk ), .D ( new_AGEMA_signal_17568 ), .Q ( new_AGEMA_signal_17569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6073 ( .C ( clk ), .D ( new_AGEMA_signal_17572 ), .Q ( new_AGEMA_signal_17573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6077 ( .C ( clk ), .D ( new_AGEMA_signal_17576 ), .Q ( new_AGEMA_signal_17577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6081 ( .C ( clk ), .D ( new_AGEMA_signal_17580 ), .Q ( new_AGEMA_signal_17581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6085 ( .C ( clk ), .D ( new_AGEMA_signal_17584 ), .Q ( new_AGEMA_signal_17585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6093 ( .C ( clk ), .D ( new_AGEMA_signal_17592 ), .Q ( new_AGEMA_signal_17593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6101 ( .C ( clk ), .D ( new_AGEMA_signal_17600 ), .Q ( new_AGEMA_signal_17601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6109 ( .C ( clk ), .D ( new_AGEMA_signal_17608 ), .Q ( new_AGEMA_signal_17609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6117 ( .C ( clk ), .D ( new_AGEMA_signal_17616 ), .Q ( new_AGEMA_signal_17617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6123 ( .C ( clk ), .D ( new_AGEMA_signal_17622 ), .Q ( new_AGEMA_signal_17623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6129 ( .C ( clk ), .D ( new_AGEMA_signal_17628 ), .Q ( new_AGEMA_signal_17629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6135 ( .C ( clk ), .D ( new_AGEMA_signal_17634 ), .Q ( new_AGEMA_signal_17635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6141 ( .C ( clk ), .D ( new_AGEMA_signal_17640 ), .Q ( new_AGEMA_signal_17641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6149 ( .C ( clk ), .D ( new_AGEMA_signal_17648 ), .Q ( new_AGEMA_signal_17649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6157 ( .C ( clk ), .D ( new_AGEMA_signal_17656 ), .Q ( new_AGEMA_signal_17657 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6165 ( .C ( clk ), .D ( new_AGEMA_signal_17664 ), .Q ( new_AGEMA_signal_17665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6173 ( .C ( clk ), .D ( new_AGEMA_signal_17672 ), .Q ( new_AGEMA_signal_17673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6181 ( .C ( clk ), .D ( new_AGEMA_signal_17680 ), .Q ( new_AGEMA_signal_17681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6189 ( .C ( clk ), .D ( new_AGEMA_signal_17688 ), .Q ( new_AGEMA_signal_17689 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6197 ( .C ( clk ), .D ( new_AGEMA_signal_17696 ), .Q ( new_AGEMA_signal_17697 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6205 ( .C ( clk ), .D ( new_AGEMA_signal_17704 ), .Q ( new_AGEMA_signal_17705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6207 ( .C ( clk ), .D ( n2514 ), .Q ( new_AGEMA_signal_17707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6209 ( .C ( clk ), .D ( new_AGEMA_signal_3378 ), .Q ( new_AGEMA_signal_17709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6211 ( .C ( clk ), .D ( new_AGEMA_signal_3379 ), .Q ( new_AGEMA_signal_17711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6213 ( .C ( clk ), .D ( new_AGEMA_signal_3380 ), .Q ( new_AGEMA_signal_17713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6217 ( .C ( clk ), .D ( new_AGEMA_signal_17716 ), .Q ( new_AGEMA_signal_17717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6221 ( .C ( clk ), .D ( new_AGEMA_signal_17720 ), .Q ( new_AGEMA_signal_17721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6225 ( .C ( clk ), .D ( new_AGEMA_signal_17724 ), .Q ( new_AGEMA_signal_17725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6229 ( .C ( clk ), .D ( new_AGEMA_signal_17728 ), .Q ( new_AGEMA_signal_17729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6233 ( .C ( clk ), .D ( new_AGEMA_signal_17732 ), .Q ( new_AGEMA_signal_17733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6237 ( .C ( clk ), .D ( new_AGEMA_signal_17736 ), .Q ( new_AGEMA_signal_17737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6241 ( .C ( clk ), .D ( new_AGEMA_signal_17740 ), .Q ( new_AGEMA_signal_17741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6245 ( .C ( clk ), .D ( new_AGEMA_signal_17744 ), .Q ( new_AGEMA_signal_17745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6253 ( .C ( clk ), .D ( new_AGEMA_signal_17752 ), .Q ( new_AGEMA_signal_17753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6261 ( .C ( clk ), .D ( new_AGEMA_signal_17760 ), .Q ( new_AGEMA_signal_17761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6269 ( .C ( clk ), .D ( new_AGEMA_signal_17768 ), .Q ( new_AGEMA_signal_17769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6277 ( .C ( clk ), .D ( new_AGEMA_signal_17776 ), .Q ( new_AGEMA_signal_17777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6281 ( .C ( clk ), .D ( new_AGEMA_signal_17780 ), .Q ( new_AGEMA_signal_17781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6285 ( .C ( clk ), .D ( new_AGEMA_signal_17784 ), .Q ( new_AGEMA_signal_17785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6289 ( .C ( clk ), .D ( new_AGEMA_signal_17788 ), .Q ( new_AGEMA_signal_17789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6293 ( .C ( clk ), .D ( new_AGEMA_signal_17792 ), .Q ( new_AGEMA_signal_17793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6299 ( .C ( clk ), .D ( new_AGEMA_signal_17798 ), .Q ( new_AGEMA_signal_17799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6307 ( .C ( clk ), .D ( new_AGEMA_signal_17806 ), .Q ( new_AGEMA_signal_17807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6315 ( .C ( clk ), .D ( new_AGEMA_signal_17814 ), .Q ( new_AGEMA_signal_17815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6323 ( .C ( clk ), .D ( new_AGEMA_signal_17822 ), .Q ( new_AGEMA_signal_17823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6335 ( .C ( clk ), .D ( new_AGEMA_signal_17834 ), .Q ( new_AGEMA_signal_17835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6347 ( .C ( clk ), .D ( new_AGEMA_signal_17846 ), .Q ( new_AGEMA_signal_17847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6359 ( .C ( clk ), .D ( new_AGEMA_signal_17858 ), .Q ( new_AGEMA_signal_17859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6371 ( .C ( clk ), .D ( new_AGEMA_signal_17870 ), .Q ( new_AGEMA_signal_17871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6385 ( .C ( clk ), .D ( new_AGEMA_signal_17884 ), .Q ( new_AGEMA_signal_17885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6399 ( .C ( clk ), .D ( new_AGEMA_signal_17898 ), .Q ( new_AGEMA_signal_17899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6413 ( .C ( clk ), .D ( new_AGEMA_signal_17912 ), .Q ( new_AGEMA_signal_17913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6427 ( .C ( clk ), .D ( new_AGEMA_signal_17926 ), .Q ( new_AGEMA_signal_17927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6435 ( .C ( clk ), .D ( new_AGEMA_signal_17934 ), .Q ( new_AGEMA_signal_17935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6443 ( .C ( clk ), .D ( new_AGEMA_signal_17942 ), .Q ( new_AGEMA_signal_17943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6451 ( .C ( clk ), .D ( new_AGEMA_signal_17950 ), .Q ( new_AGEMA_signal_17951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6459 ( .C ( clk ), .D ( new_AGEMA_signal_17958 ), .Q ( new_AGEMA_signal_17959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6473 ( .C ( clk ), .D ( new_AGEMA_signal_17972 ), .Q ( new_AGEMA_signal_17973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6487 ( .C ( clk ), .D ( new_AGEMA_signal_17986 ), .Q ( new_AGEMA_signal_17987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6501 ( .C ( clk ), .D ( new_AGEMA_signal_18000 ), .Q ( new_AGEMA_signal_18001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6515 ( .C ( clk ), .D ( new_AGEMA_signal_18014 ), .Q ( new_AGEMA_signal_18015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6523 ( .C ( clk ), .D ( new_AGEMA_signal_18022 ), .Q ( new_AGEMA_signal_18023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6531 ( .C ( clk ), .D ( new_AGEMA_signal_18030 ), .Q ( new_AGEMA_signal_18031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6539 ( .C ( clk ), .D ( new_AGEMA_signal_18038 ), .Q ( new_AGEMA_signal_18039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6547 ( .C ( clk ), .D ( new_AGEMA_signal_18046 ), .Q ( new_AGEMA_signal_18047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6555 ( .C ( clk ), .D ( new_AGEMA_signal_18054 ), .Q ( new_AGEMA_signal_18055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6563 ( .C ( clk ), .D ( new_AGEMA_signal_18062 ), .Q ( new_AGEMA_signal_18063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6571 ( .C ( clk ), .D ( new_AGEMA_signal_18070 ), .Q ( new_AGEMA_signal_18071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6579 ( .C ( clk ), .D ( new_AGEMA_signal_18078 ), .Q ( new_AGEMA_signal_18079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6617 ( .C ( clk ), .D ( new_AGEMA_signal_18116 ), .Q ( new_AGEMA_signal_18117 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6633 ( .C ( clk ), .D ( new_AGEMA_signal_18132 ), .Q ( new_AGEMA_signal_18133 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6649 ( .C ( clk ), .D ( new_AGEMA_signal_18148 ), .Q ( new_AGEMA_signal_18149 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6665 ( .C ( clk ), .D ( new_AGEMA_signal_18164 ), .Q ( new_AGEMA_signal_18165 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6705 ( .C ( clk ), .D ( new_AGEMA_signal_18204 ), .Q ( new_AGEMA_signal_18205 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6721 ( .C ( clk ), .D ( new_AGEMA_signal_18220 ), .Q ( new_AGEMA_signal_18221 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6737 ( .C ( clk ), .D ( new_AGEMA_signal_18236 ), .Q ( new_AGEMA_signal_18237 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6753 ( .C ( clk ), .D ( new_AGEMA_signal_18252 ), .Q ( new_AGEMA_signal_18253 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6763 ( .C ( clk ), .D ( new_AGEMA_signal_18262 ), .Q ( new_AGEMA_signal_18263 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6773 ( .C ( clk ), .D ( new_AGEMA_signal_18272 ), .Q ( new_AGEMA_signal_18273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6783 ( .C ( clk ), .D ( new_AGEMA_signal_18282 ), .Q ( new_AGEMA_signal_18283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6793 ( .C ( clk ), .D ( new_AGEMA_signal_18292 ), .Q ( new_AGEMA_signal_18293 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6817 ( .C ( clk ), .D ( new_AGEMA_signal_18316 ), .Q ( new_AGEMA_signal_18317 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6825 ( .C ( clk ), .D ( new_AGEMA_signal_18324 ), .Q ( new_AGEMA_signal_18325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6833 ( .C ( clk ), .D ( new_AGEMA_signal_18332 ), .Q ( new_AGEMA_signal_18333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6841 ( .C ( clk ), .D ( new_AGEMA_signal_18340 ), .Q ( new_AGEMA_signal_18341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6903 ( .C ( clk ), .D ( new_AGEMA_signal_18402 ), .Q ( new_AGEMA_signal_18403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6919 ( .C ( clk ), .D ( new_AGEMA_signal_18418 ), .Q ( new_AGEMA_signal_18419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6935 ( .C ( clk ), .D ( new_AGEMA_signal_18434 ), .Q ( new_AGEMA_signal_18435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6951 ( .C ( clk ), .D ( new_AGEMA_signal_18450 ), .Q ( new_AGEMA_signal_18451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6961 ( .C ( clk ), .D ( new_AGEMA_signal_18460 ), .Q ( new_AGEMA_signal_18461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6971 ( .C ( clk ), .D ( new_AGEMA_signal_18470 ), .Q ( new_AGEMA_signal_18471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6981 ( .C ( clk ), .D ( new_AGEMA_signal_18480 ), .Q ( new_AGEMA_signal_18481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6991 ( .C ( clk ), .D ( new_AGEMA_signal_18490 ), .Q ( new_AGEMA_signal_18491 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7009 ( .C ( clk ), .D ( new_AGEMA_signal_18508 ), .Q ( new_AGEMA_signal_18509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7027 ( .C ( clk ), .D ( new_AGEMA_signal_18526 ), .Q ( new_AGEMA_signal_18527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7045 ( .C ( clk ), .D ( new_AGEMA_signal_18544 ), .Q ( new_AGEMA_signal_18545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7063 ( .C ( clk ), .D ( new_AGEMA_signal_18562 ), .Q ( new_AGEMA_signal_18563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7087 ( .C ( clk ), .D ( n2671 ), .Q ( new_AGEMA_signal_18587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7095 ( .C ( clk ), .D ( new_AGEMA_signal_3489 ), .Q ( new_AGEMA_signal_18595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7103 ( .C ( clk ), .D ( new_AGEMA_signal_3490 ), .Q ( new_AGEMA_signal_18603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7111 ( .C ( clk ), .D ( new_AGEMA_signal_3491 ), .Q ( new_AGEMA_signal_18611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7209 ( .C ( clk ), .D ( new_AGEMA_signal_18708 ), .Q ( new_AGEMA_signal_18709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7229 ( .C ( clk ), .D ( new_AGEMA_signal_18728 ), .Q ( new_AGEMA_signal_18729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7249 ( .C ( clk ), .D ( new_AGEMA_signal_18748 ), .Q ( new_AGEMA_signal_18749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7269 ( .C ( clk ), .D ( new_AGEMA_signal_18768 ), .Q ( new_AGEMA_signal_18769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7311 ( .C ( clk ), .D ( n2380 ), .Q ( new_AGEMA_signal_18811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7323 ( .C ( clk ), .D ( new_AGEMA_signal_3474 ), .Q ( new_AGEMA_signal_18823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7335 ( .C ( clk ), .D ( new_AGEMA_signal_3475 ), .Q ( new_AGEMA_signal_18835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7347 ( .C ( clk ), .D ( new_AGEMA_signal_3476 ), .Q ( new_AGEMA_signal_18847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7359 ( .C ( clk ), .D ( n2382 ), .Q ( new_AGEMA_signal_18859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7373 ( .C ( clk ), .D ( new_AGEMA_signal_3471 ), .Q ( new_AGEMA_signal_18873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7387 ( .C ( clk ), .D ( new_AGEMA_signal_3472 ), .Q ( new_AGEMA_signal_18887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7401 ( .C ( clk ), .D ( new_AGEMA_signal_3473 ), .Q ( new_AGEMA_signal_18901 ) ) ;

    /* cells in depth 18 */
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2016 ( .ina ({new_AGEMA_signal_3425, new_AGEMA_signal_3424, new_AGEMA_signal_3423, n1941}), .inb ({new_AGEMA_signal_16890, new_AGEMA_signal_16884, new_AGEMA_signal_16878, new_AGEMA_signal_16872}), .clk ( clk ), .rnd ({Fresh[7939], Fresh[7938], Fresh[7937], Fresh[7936], Fresh[7935], Fresh[7934], Fresh[7933], Fresh[7932], Fresh[7931], Fresh[7930]}), .outt ({new_AGEMA_signal_3509, new_AGEMA_signal_3508, new_AGEMA_signal_3507, n2019}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2060 ( .ina ({new_AGEMA_signal_16914, new_AGEMA_signal_16908, new_AGEMA_signal_16902, new_AGEMA_signal_16896}), .inb ({new_AGEMA_signal_3428, new_AGEMA_signal_3427, new_AGEMA_signal_3426, n1960}), .clk ( clk ), .rnd ({Fresh[7949], Fresh[7948], Fresh[7947], Fresh[7946], Fresh[7945], Fresh[7944], Fresh[7943], Fresh[7942], Fresh[7941], Fresh[7940]}), .outt ({new_AGEMA_signal_3512, new_AGEMA_signal_3511, new_AGEMA_signal_3510, n2002}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2116 ( .ina ({new_AGEMA_signal_3431, new_AGEMA_signal_3430, new_AGEMA_signal_3429, n1988}), .inb ({new_AGEMA_signal_16938, new_AGEMA_signal_16932, new_AGEMA_signal_16926, new_AGEMA_signal_16920}), .clk ( clk ), .rnd ({Fresh[7959], Fresh[7958], Fresh[7957], Fresh[7956], Fresh[7955], Fresh[7954], Fresh[7953], Fresh[7952], Fresh[7951], Fresh[7950]}), .outt ({new_AGEMA_signal_3515, new_AGEMA_signal_3514, new_AGEMA_signal_3513, n1989}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2154 ( .ina ({new_AGEMA_signal_16954, new_AGEMA_signal_16950, new_AGEMA_signal_16946, new_AGEMA_signal_16942}), .inb ({new_AGEMA_signal_3434, new_AGEMA_signal_3433, new_AGEMA_signal_3432, n2015}), .clk ( clk ), .rnd ({Fresh[7969], Fresh[7968], Fresh[7967], Fresh[7966], Fresh[7965], Fresh[7964], Fresh[7963], Fresh[7962], Fresh[7961], Fresh[7960]}), .outt ({new_AGEMA_signal_3518, new_AGEMA_signal_3517, new_AGEMA_signal_3516, n2016}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2170 ( .ina ({new_AGEMA_signal_16986, new_AGEMA_signal_16978, new_AGEMA_signal_16970, new_AGEMA_signal_16962}), .inb ({new_AGEMA_signal_3308, new_AGEMA_signal_3307, new_AGEMA_signal_3306, n2030}), .clk ( clk ), .rnd ({Fresh[7979], Fresh[7978], Fresh[7977], Fresh[7976], Fresh[7975], Fresh[7974], Fresh[7973], Fresh[7972], Fresh[7971], Fresh[7970]}), .outt ({new_AGEMA_signal_3437, new_AGEMA_signal_3436, new_AGEMA_signal_3435, n2038}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2201 ( .ina ({new_AGEMA_signal_17010, new_AGEMA_signal_17004, new_AGEMA_signal_16998, new_AGEMA_signal_16992}), .inb ({new_AGEMA_signal_3440, new_AGEMA_signal_3439, new_AGEMA_signal_3438, n2053}), .clk ( clk ), .rnd ({Fresh[7989], Fresh[7988], Fresh[7987], Fresh[7986], Fresh[7985], Fresh[7984], Fresh[7983], Fresh[7982], Fresh[7981], Fresh[7980]}), .outt ({new_AGEMA_signal_3524, new_AGEMA_signal_3523, new_AGEMA_signal_3522, n2111}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2223 ( .ina ({new_AGEMA_signal_17026, new_AGEMA_signal_17022, new_AGEMA_signal_17018, new_AGEMA_signal_17014}), .inb ({new_AGEMA_signal_3443, new_AGEMA_signal_3442, new_AGEMA_signal_3441, n2071}), .clk ( clk ), .rnd ({Fresh[7999], Fresh[7998], Fresh[7997], Fresh[7996], Fresh[7995], Fresh[7994], Fresh[7993], Fresh[7992], Fresh[7991], Fresh[7990]}), .outt ({new_AGEMA_signal_3527, new_AGEMA_signal_3526, new_AGEMA_signal_3525, n2079}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2263 ( .ina ({new_AGEMA_signal_3446, new_AGEMA_signal_3445, new_AGEMA_signal_3444, n2103}), .inb ({new_AGEMA_signal_17058, new_AGEMA_signal_17050, new_AGEMA_signal_17042, new_AGEMA_signal_17034}), .clk ( clk ), .rnd ({Fresh[8009], Fresh[8008], Fresh[8007], Fresh[8006], Fresh[8005], Fresh[8004], Fresh[8003], Fresh[8002], Fresh[8001], Fresh[8000]}), .outt ({new_AGEMA_signal_3530, new_AGEMA_signal_3529, new_AGEMA_signal_3528, n2104}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2289 ( .ina ({new_AGEMA_signal_17090, new_AGEMA_signal_17082, new_AGEMA_signal_17074, new_AGEMA_signal_17066}), .inb ({new_AGEMA_signal_3449, new_AGEMA_signal_3448, new_AGEMA_signal_3447, n2126}), .clk ( clk ), .rnd ({Fresh[8019], Fresh[8018], Fresh[8017], Fresh[8016], Fresh[8015], Fresh[8014], Fresh[8013], Fresh[8012], Fresh[8011], Fresh[8010]}), .outt ({new_AGEMA_signal_3533, new_AGEMA_signal_3532, new_AGEMA_signal_3531, n2127}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2315 ( .ina ({new_AGEMA_signal_16954, new_AGEMA_signal_16950, new_AGEMA_signal_16946, new_AGEMA_signal_16942}), .inb ({new_AGEMA_signal_3452, new_AGEMA_signal_3451, new_AGEMA_signal_3450, n2146}), .clk ( clk ), .rnd ({Fresh[8029], Fresh[8028], Fresh[8027], Fresh[8026], Fresh[8025], Fresh[8024], Fresh[8023], Fresh[8022], Fresh[8021], Fresh[8020]}), .outt ({new_AGEMA_signal_3536, new_AGEMA_signal_3535, new_AGEMA_signal_3534, n2147}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2336 ( .ina ({new_AGEMA_signal_3455, new_AGEMA_signal_3454, new_AGEMA_signal_3453, n2173}), .inb ({new_AGEMA_signal_17130, new_AGEMA_signal_17120, new_AGEMA_signal_17110, new_AGEMA_signal_17100}), .clk ( clk ), .rnd ({Fresh[8039], Fresh[8038], Fresh[8037], Fresh[8036], Fresh[8035], Fresh[8034], Fresh[8033], Fresh[8032], Fresh[8031], Fresh[8030]}), .outt ({new_AGEMA_signal_3539, new_AGEMA_signal_3538, new_AGEMA_signal_3537, n2208}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2352 ( .ina ({new_AGEMA_signal_3458, new_AGEMA_signal_3457, new_AGEMA_signal_3456, n2187}), .inb ({new_AGEMA_signal_17162, new_AGEMA_signal_17154, new_AGEMA_signal_17146, new_AGEMA_signal_17138}), .clk ( clk ), .rnd ({Fresh[8049], Fresh[8048], Fresh[8047], Fresh[8046], Fresh[8045], Fresh[8044], Fresh[8043], Fresh[8042], Fresh[8041], Fresh[8040]}), .outt ({new_AGEMA_signal_3542, new_AGEMA_signal_3541, new_AGEMA_signal_3540, n2199}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2420 ( .ina ({new_AGEMA_signal_3464, new_AGEMA_signal_3463, new_AGEMA_signal_3462, n2256}), .inb ({new_AGEMA_signal_17186, new_AGEMA_signal_17180, new_AGEMA_signal_17174, new_AGEMA_signal_17168}), .clk ( clk ), .rnd ({Fresh[8059], Fresh[8058], Fresh[8057], Fresh[8056], Fresh[8055], Fresh[8054], Fresh[8053], Fresh[8052], Fresh[8051], Fresh[8050]}), .outt ({new_AGEMA_signal_3545, new_AGEMA_signal_3544, new_AGEMA_signal_3543, n2257}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2442 ( .ina ({new_AGEMA_signal_17202, new_AGEMA_signal_17198, new_AGEMA_signal_17194, new_AGEMA_signal_17190}), .inb ({new_AGEMA_signal_3467, new_AGEMA_signal_3466, new_AGEMA_signal_3465, n2275}), .clk ( clk ), .rnd ({Fresh[8069], Fresh[8068], Fresh[8067], Fresh[8066], Fresh[8065], Fresh[8064], Fresh[8063], Fresh[8062], Fresh[8061], Fresh[8060]}), .outt ({new_AGEMA_signal_3548, new_AGEMA_signal_3547, new_AGEMA_signal_3546, n2281}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2475 ( .ina ({new_AGEMA_signal_17226, new_AGEMA_signal_17220, new_AGEMA_signal_17214, new_AGEMA_signal_17208}), .inb ({new_AGEMA_signal_3470, new_AGEMA_signal_3469, new_AGEMA_signal_3468, n2303}), .clk ( clk ), .rnd ({Fresh[8079], Fresh[8078], Fresh[8077], Fresh[8076], Fresh[8075], Fresh[8074], Fresh[8073], Fresh[8072], Fresh[8071], Fresh[8070]}), .outt ({new_AGEMA_signal_3551, new_AGEMA_signal_3550, new_AGEMA_signal_3549, n2305}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2532 ( .ina ({new_AGEMA_signal_17258, new_AGEMA_signal_17250, new_AGEMA_signal_17242, new_AGEMA_signal_17234}), .inb ({new_AGEMA_signal_3479, new_AGEMA_signal_3478, new_AGEMA_signal_3477, n2366}), .clk ( clk ), .rnd ({Fresh[8089], Fresh[8088], Fresh[8087], Fresh[8086], Fresh[8085], Fresh[8084], Fresh[8083], Fresh[8082], Fresh[8081], Fresh[8080]}), .outt ({new_AGEMA_signal_3554, new_AGEMA_signal_3553, new_AGEMA_signal_3552, n2368}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2583 ( .ina ({new_AGEMA_signal_3482, new_AGEMA_signal_3481, new_AGEMA_signal_3480, n2425}), .inb ({new_AGEMA_signal_3374, new_AGEMA_signal_3373, new_AGEMA_signal_3372, n2424}), .clk ( clk ), .rnd ({Fresh[8099], Fresh[8098], Fresh[8097], Fresh[8096], Fresh[8095], Fresh[8094], Fresh[8093], Fresh[8092], Fresh[8091], Fresh[8090]}), .outt ({new_AGEMA_signal_3557, new_AGEMA_signal_3556, new_AGEMA_signal_3555, n2426}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2605 ( .ina ({new_AGEMA_signal_3485, new_AGEMA_signal_3484, new_AGEMA_signal_3483, n2451}), .inb ({new_AGEMA_signal_17282, new_AGEMA_signal_17276, new_AGEMA_signal_17270, new_AGEMA_signal_17264}), .clk ( clk ), .rnd ({Fresh[8109], Fresh[8108], Fresh[8107], Fresh[8106], Fresh[8105], Fresh[8104], Fresh[8103], Fresh[8102], Fresh[8101], Fresh[8100]}), .outt ({new_AGEMA_signal_3560, new_AGEMA_signal_3559, new_AGEMA_signal_3558, n2457}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2659 ( .ina ({new_AGEMA_signal_17290, new_AGEMA_signal_17288, new_AGEMA_signal_17286, new_AGEMA_signal_17284}), .inb ({new_AGEMA_signal_3488, new_AGEMA_signal_3487, new_AGEMA_signal_3486, n2511}), .clk ( clk ), .rnd ({Fresh[8119], Fresh[8118], Fresh[8117], Fresh[8116], Fresh[8115], Fresh[8114], Fresh[8113], Fresh[8112], Fresh[8111], Fresh[8110]}), .outt ({new_AGEMA_signal_3563, new_AGEMA_signal_3562, new_AGEMA_signal_3561, n2513}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2717 ( .ina ({new_AGEMA_signal_17322, new_AGEMA_signal_17314, new_AGEMA_signal_17306, new_AGEMA_signal_17298}), .inb ({new_AGEMA_signal_3494, new_AGEMA_signal_3493, new_AGEMA_signal_3492, n2590}), .clk ( clk ), .rnd ({Fresh[8129], Fresh[8128], Fresh[8127], Fresh[8126], Fresh[8125], Fresh[8124], Fresh[8123], Fresh[8122], Fresh[8121], Fresh[8120]}), .outt ({new_AGEMA_signal_3566, new_AGEMA_signal_3565, new_AGEMA_signal_3564, n2592}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2741 ( .ina ({new_AGEMA_signal_3404, new_AGEMA_signal_3403, new_AGEMA_signal_3402, n2623}), .inb ({new_AGEMA_signal_17338, new_AGEMA_signal_17334, new_AGEMA_signal_17330, new_AGEMA_signal_17326}), .clk ( clk ), .rnd ({Fresh[8139], Fresh[8138], Fresh[8137], Fresh[8136], Fresh[8135], Fresh[8134], Fresh[8133], Fresh[8132], Fresh[8131], Fresh[8130]}), .outt ({new_AGEMA_signal_3497, new_AGEMA_signal_3496, new_AGEMA_signal_3495, n2637}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2767 ( .ina ({new_AGEMA_signal_3500, new_AGEMA_signal_3499, new_AGEMA_signal_3498, n2667}), .inb ({new_AGEMA_signal_17362, new_AGEMA_signal_17356, new_AGEMA_signal_17350, new_AGEMA_signal_17344}), .clk ( clk ), .rnd ({Fresh[8149], Fresh[8148], Fresh[8147], Fresh[8146], Fresh[8145], Fresh[8144], Fresh[8143], Fresh[8142], Fresh[8141], Fresh[8140]}), .outt ({new_AGEMA_signal_3572, new_AGEMA_signal_3571, new_AGEMA_signal_3570, n2668}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2787 ( .ina ({new_AGEMA_signal_17386, new_AGEMA_signal_17380, new_AGEMA_signal_17374, new_AGEMA_signal_17368}), .inb ({new_AGEMA_signal_3503, new_AGEMA_signal_3502, new_AGEMA_signal_3501, n2703}), .clk ( clk ), .rnd ({Fresh[8159], Fresh[8158], Fresh[8157], Fresh[8156], Fresh[8155], Fresh[8154], Fresh[8153], Fresh[8152], Fresh[8151], Fresh[8150]}), .outt ({new_AGEMA_signal_3575, new_AGEMA_signal_3574, new_AGEMA_signal_3573, n2705}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2841 ( .ina ({new_AGEMA_signal_17402, new_AGEMA_signal_17398, new_AGEMA_signal_17394, new_AGEMA_signal_17390}), .inb ({new_AGEMA_signal_3419, new_AGEMA_signal_3418, new_AGEMA_signal_3417, n2803}), .clk ( clk ), .rnd ({Fresh[8169], Fresh[8168], Fresh[8167], Fresh[8166], Fresh[8165], Fresh[8164], Fresh[8163], Fresh[8162], Fresh[8161], Fresh[8160]}), .outt ({new_AGEMA_signal_3506, new_AGEMA_signal_3505, new_AGEMA_signal_3504, n2805}) ) ;
    buf_clk new_AGEMA_reg_buffer_5908 ( .C ( clk ), .D ( new_AGEMA_signal_17407 ), .Q ( new_AGEMA_signal_17408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5914 ( .C ( clk ), .D ( new_AGEMA_signal_17413 ), .Q ( new_AGEMA_signal_17414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5920 ( .C ( clk ), .D ( new_AGEMA_signal_17419 ), .Q ( new_AGEMA_signal_17420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5926 ( .C ( clk ), .D ( new_AGEMA_signal_17425 ), .Q ( new_AGEMA_signal_17426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5930 ( .C ( clk ), .D ( new_AGEMA_signal_17429 ), .Q ( new_AGEMA_signal_17430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5934 ( .C ( clk ), .D ( new_AGEMA_signal_17433 ), .Q ( new_AGEMA_signal_17434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5938 ( .C ( clk ), .D ( new_AGEMA_signal_17437 ), .Q ( new_AGEMA_signal_17438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5942 ( .C ( clk ), .D ( new_AGEMA_signal_17441 ), .Q ( new_AGEMA_signal_17442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5948 ( .C ( clk ), .D ( new_AGEMA_signal_17447 ), .Q ( new_AGEMA_signal_17448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5954 ( .C ( clk ), .D ( new_AGEMA_signal_17453 ), .Q ( new_AGEMA_signal_17454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5960 ( .C ( clk ), .D ( new_AGEMA_signal_17459 ), .Q ( new_AGEMA_signal_17460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5966 ( .C ( clk ), .D ( new_AGEMA_signal_17465 ), .Q ( new_AGEMA_signal_17466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5976 ( .C ( clk ), .D ( new_AGEMA_signal_17475 ), .Q ( new_AGEMA_signal_17476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5986 ( .C ( clk ), .D ( new_AGEMA_signal_17485 ), .Q ( new_AGEMA_signal_17486 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5996 ( .C ( clk ), .D ( new_AGEMA_signal_17495 ), .Q ( new_AGEMA_signal_17496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6006 ( .C ( clk ), .D ( new_AGEMA_signal_17505 ), .Q ( new_AGEMA_signal_17506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6012 ( .C ( clk ), .D ( new_AGEMA_signal_17511 ), .Q ( new_AGEMA_signal_17512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6018 ( .C ( clk ), .D ( new_AGEMA_signal_17517 ), .Q ( new_AGEMA_signal_17518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6024 ( .C ( clk ), .D ( new_AGEMA_signal_17523 ), .Q ( new_AGEMA_signal_17524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6030 ( .C ( clk ), .D ( new_AGEMA_signal_17529 ), .Q ( new_AGEMA_signal_17530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6036 ( .C ( clk ), .D ( new_AGEMA_signal_17535 ), .Q ( new_AGEMA_signal_17536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6042 ( .C ( clk ), .D ( new_AGEMA_signal_17541 ), .Q ( new_AGEMA_signal_17542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6048 ( .C ( clk ), .D ( new_AGEMA_signal_17547 ), .Q ( new_AGEMA_signal_17548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6054 ( .C ( clk ), .D ( new_AGEMA_signal_17553 ), .Q ( new_AGEMA_signal_17554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6058 ( .C ( clk ), .D ( new_AGEMA_signal_17557 ), .Q ( new_AGEMA_signal_17558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6062 ( .C ( clk ), .D ( new_AGEMA_signal_17561 ), .Q ( new_AGEMA_signal_17562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6066 ( .C ( clk ), .D ( new_AGEMA_signal_17565 ), .Q ( new_AGEMA_signal_17566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6070 ( .C ( clk ), .D ( new_AGEMA_signal_17569 ), .Q ( new_AGEMA_signal_17570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6074 ( .C ( clk ), .D ( new_AGEMA_signal_17573 ), .Q ( new_AGEMA_signal_17574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6078 ( .C ( clk ), .D ( new_AGEMA_signal_17577 ), .Q ( new_AGEMA_signal_17578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6082 ( .C ( clk ), .D ( new_AGEMA_signal_17581 ), .Q ( new_AGEMA_signal_17582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6086 ( .C ( clk ), .D ( new_AGEMA_signal_17585 ), .Q ( new_AGEMA_signal_17586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6094 ( .C ( clk ), .D ( new_AGEMA_signal_17593 ), .Q ( new_AGEMA_signal_17594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6102 ( .C ( clk ), .D ( new_AGEMA_signal_17601 ), .Q ( new_AGEMA_signal_17602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6110 ( .C ( clk ), .D ( new_AGEMA_signal_17609 ), .Q ( new_AGEMA_signal_17610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6118 ( .C ( clk ), .D ( new_AGEMA_signal_17617 ), .Q ( new_AGEMA_signal_17618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6124 ( .C ( clk ), .D ( new_AGEMA_signal_17623 ), .Q ( new_AGEMA_signal_17624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6130 ( .C ( clk ), .D ( new_AGEMA_signal_17629 ), .Q ( new_AGEMA_signal_17630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6136 ( .C ( clk ), .D ( new_AGEMA_signal_17635 ), .Q ( new_AGEMA_signal_17636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6142 ( .C ( clk ), .D ( new_AGEMA_signal_17641 ), .Q ( new_AGEMA_signal_17642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6150 ( .C ( clk ), .D ( new_AGEMA_signal_17649 ), .Q ( new_AGEMA_signal_17650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6158 ( .C ( clk ), .D ( new_AGEMA_signal_17657 ), .Q ( new_AGEMA_signal_17658 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6166 ( .C ( clk ), .D ( new_AGEMA_signal_17665 ), .Q ( new_AGEMA_signal_17666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6174 ( .C ( clk ), .D ( new_AGEMA_signal_17673 ), .Q ( new_AGEMA_signal_17674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6182 ( .C ( clk ), .D ( new_AGEMA_signal_17681 ), .Q ( new_AGEMA_signal_17682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6190 ( .C ( clk ), .D ( new_AGEMA_signal_17689 ), .Q ( new_AGEMA_signal_17690 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6198 ( .C ( clk ), .D ( new_AGEMA_signal_17697 ), .Q ( new_AGEMA_signal_17698 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6206 ( .C ( clk ), .D ( new_AGEMA_signal_17705 ), .Q ( new_AGEMA_signal_17706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6208 ( .C ( clk ), .D ( new_AGEMA_signal_17707 ), .Q ( new_AGEMA_signal_17708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6210 ( .C ( clk ), .D ( new_AGEMA_signal_17709 ), .Q ( new_AGEMA_signal_17710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6212 ( .C ( clk ), .D ( new_AGEMA_signal_17711 ), .Q ( new_AGEMA_signal_17712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6214 ( .C ( clk ), .D ( new_AGEMA_signal_17713 ), .Q ( new_AGEMA_signal_17714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6218 ( .C ( clk ), .D ( new_AGEMA_signal_17717 ), .Q ( new_AGEMA_signal_17718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6222 ( .C ( clk ), .D ( new_AGEMA_signal_17721 ), .Q ( new_AGEMA_signal_17722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6226 ( .C ( clk ), .D ( new_AGEMA_signal_17725 ), .Q ( new_AGEMA_signal_17726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6230 ( .C ( clk ), .D ( new_AGEMA_signal_17729 ), .Q ( new_AGEMA_signal_17730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6234 ( .C ( clk ), .D ( new_AGEMA_signal_17733 ), .Q ( new_AGEMA_signal_17734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6238 ( .C ( clk ), .D ( new_AGEMA_signal_17737 ), .Q ( new_AGEMA_signal_17738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6242 ( .C ( clk ), .D ( new_AGEMA_signal_17741 ), .Q ( new_AGEMA_signal_17742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6246 ( .C ( clk ), .D ( new_AGEMA_signal_17745 ), .Q ( new_AGEMA_signal_17746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6254 ( .C ( clk ), .D ( new_AGEMA_signal_17753 ), .Q ( new_AGEMA_signal_17754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6262 ( .C ( clk ), .D ( new_AGEMA_signal_17761 ), .Q ( new_AGEMA_signal_17762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6270 ( .C ( clk ), .D ( new_AGEMA_signal_17769 ), .Q ( new_AGEMA_signal_17770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6278 ( .C ( clk ), .D ( new_AGEMA_signal_17777 ), .Q ( new_AGEMA_signal_17778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6282 ( .C ( clk ), .D ( new_AGEMA_signal_17781 ), .Q ( new_AGEMA_signal_17782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6286 ( .C ( clk ), .D ( new_AGEMA_signal_17785 ), .Q ( new_AGEMA_signal_17786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6290 ( .C ( clk ), .D ( new_AGEMA_signal_17789 ), .Q ( new_AGEMA_signal_17790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6294 ( .C ( clk ), .D ( new_AGEMA_signal_17793 ), .Q ( new_AGEMA_signal_17794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6300 ( .C ( clk ), .D ( new_AGEMA_signal_17799 ), .Q ( new_AGEMA_signal_17800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6308 ( .C ( clk ), .D ( new_AGEMA_signal_17807 ), .Q ( new_AGEMA_signal_17808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6316 ( .C ( clk ), .D ( new_AGEMA_signal_17815 ), .Q ( new_AGEMA_signal_17816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6324 ( .C ( clk ), .D ( new_AGEMA_signal_17823 ), .Q ( new_AGEMA_signal_17824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6336 ( .C ( clk ), .D ( new_AGEMA_signal_17835 ), .Q ( new_AGEMA_signal_17836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6348 ( .C ( clk ), .D ( new_AGEMA_signal_17847 ), .Q ( new_AGEMA_signal_17848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6360 ( .C ( clk ), .D ( new_AGEMA_signal_17859 ), .Q ( new_AGEMA_signal_17860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6372 ( .C ( clk ), .D ( new_AGEMA_signal_17871 ), .Q ( new_AGEMA_signal_17872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6386 ( .C ( clk ), .D ( new_AGEMA_signal_17885 ), .Q ( new_AGEMA_signal_17886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6400 ( .C ( clk ), .D ( new_AGEMA_signal_17899 ), .Q ( new_AGEMA_signal_17900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6414 ( .C ( clk ), .D ( new_AGEMA_signal_17913 ), .Q ( new_AGEMA_signal_17914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6428 ( .C ( clk ), .D ( new_AGEMA_signal_17927 ), .Q ( new_AGEMA_signal_17928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6436 ( .C ( clk ), .D ( new_AGEMA_signal_17935 ), .Q ( new_AGEMA_signal_17936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6444 ( .C ( clk ), .D ( new_AGEMA_signal_17943 ), .Q ( new_AGEMA_signal_17944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6452 ( .C ( clk ), .D ( new_AGEMA_signal_17951 ), .Q ( new_AGEMA_signal_17952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6460 ( .C ( clk ), .D ( new_AGEMA_signal_17959 ), .Q ( new_AGEMA_signal_17960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6474 ( .C ( clk ), .D ( new_AGEMA_signal_17973 ), .Q ( new_AGEMA_signal_17974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6488 ( .C ( clk ), .D ( new_AGEMA_signal_17987 ), .Q ( new_AGEMA_signal_17988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6502 ( .C ( clk ), .D ( new_AGEMA_signal_18001 ), .Q ( new_AGEMA_signal_18002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6516 ( .C ( clk ), .D ( new_AGEMA_signal_18015 ), .Q ( new_AGEMA_signal_18016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6524 ( .C ( clk ), .D ( new_AGEMA_signal_18023 ), .Q ( new_AGEMA_signal_18024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6532 ( .C ( clk ), .D ( new_AGEMA_signal_18031 ), .Q ( new_AGEMA_signal_18032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6540 ( .C ( clk ), .D ( new_AGEMA_signal_18039 ), .Q ( new_AGEMA_signal_18040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6548 ( .C ( clk ), .D ( new_AGEMA_signal_18047 ), .Q ( new_AGEMA_signal_18048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6556 ( .C ( clk ), .D ( new_AGEMA_signal_18055 ), .Q ( new_AGEMA_signal_18056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6564 ( .C ( clk ), .D ( new_AGEMA_signal_18063 ), .Q ( new_AGEMA_signal_18064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6572 ( .C ( clk ), .D ( new_AGEMA_signal_18071 ), .Q ( new_AGEMA_signal_18072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6580 ( .C ( clk ), .D ( new_AGEMA_signal_18079 ), .Q ( new_AGEMA_signal_18080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6618 ( .C ( clk ), .D ( new_AGEMA_signal_18117 ), .Q ( new_AGEMA_signal_18118 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6634 ( .C ( clk ), .D ( new_AGEMA_signal_18133 ), .Q ( new_AGEMA_signal_18134 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6650 ( .C ( clk ), .D ( new_AGEMA_signal_18149 ), .Q ( new_AGEMA_signal_18150 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6666 ( .C ( clk ), .D ( new_AGEMA_signal_18165 ), .Q ( new_AGEMA_signal_18166 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6706 ( .C ( clk ), .D ( new_AGEMA_signal_18205 ), .Q ( new_AGEMA_signal_18206 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6722 ( .C ( clk ), .D ( new_AGEMA_signal_18221 ), .Q ( new_AGEMA_signal_18222 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6738 ( .C ( clk ), .D ( new_AGEMA_signal_18237 ), .Q ( new_AGEMA_signal_18238 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6754 ( .C ( clk ), .D ( new_AGEMA_signal_18253 ), .Q ( new_AGEMA_signal_18254 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6764 ( .C ( clk ), .D ( new_AGEMA_signal_18263 ), .Q ( new_AGEMA_signal_18264 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6774 ( .C ( clk ), .D ( new_AGEMA_signal_18273 ), .Q ( new_AGEMA_signal_18274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6784 ( .C ( clk ), .D ( new_AGEMA_signal_18283 ), .Q ( new_AGEMA_signal_18284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6794 ( .C ( clk ), .D ( new_AGEMA_signal_18293 ), .Q ( new_AGEMA_signal_18294 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6818 ( .C ( clk ), .D ( new_AGEMA_signal_18317 ), .Q ( new_AGEMA_signal_18318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6826 ( .C ( clk ), .D ( new_AGEMA_signal_18325 ), .Q ( new_AGEMA_signal_18326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6834 ( .C ( clk ), .D ( new_AGEMA_signal_18333 ), .Q ( new_AGEMA_signal_18334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6842 ( .C ( clk ), .D ( new_AGEMA_signal_18341 ), .Q ( new_AGEMA_signal_18342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6904 ( .C ( clk ), .D ( new_AGEMA_signal_18403 ), .Q ( new_AGEMA_signal_18404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6920 ( .C ( clk ), .D ( new_AGEMA_signal_18419 ), .Q ( new_AGEMA_signal_18420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6936 ( .C ( clk ), .D ( new_AGEMA_signal_18435 ), .Q ( new_AGEMA_signal_18436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6952 ( .C ( clk ), .D ( new_AGEMA_signal_18451 ), .Q ( new_AGEMA_signal_18452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6962 ( .C ( clk ), .D ( new_AGEMA_signal_18461 ), .Q ( new_AGEMA_signal_18462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6972 ( .C ( clk ), .D ( new_AGEMA_signal_18471 ), .Q ( new_AGEMA_signal_18472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6982 ( .C ( clk ), .D ( new_AGEMA_signal_18481 ), .Q ( new_AGEMA_signal_18482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6992 ( .C ( clk ), .D ( new_AGEMA_signal_18491 ), .Q ( new_AGEMA_signal_18492 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7010 ( .C ( clk ), .D ( new_AGEMA_signal_18509 ), .Q ( new_AGEMA_signal_18510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7028 ( .C ( clk ), .D ( new_AGEMA_signal_18527 ), .Q ( new_AGEMA_signal_18528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7046 ( .C ( clk ), .D ( new_AGEMA_signal_18545 ), .Q ( new_AGEMA_signal_18546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7064 ( .C ( clk ), .D ( new_AGEMA_signal_18563 ), .Q ( new_AGEMA_signal_18564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7088 ( .C ( clk ), .D ( new_AGEMA_signal_18587 ), .Q ( new_AGEMA_signal_18588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7096 ( .C ( clk ), .D ( new_AGEMA_signal_18595 ), .Q ( new_AGEMA_signal_18596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7104 ( .C ( clk ), .D ( new_AGEMA_signal_18603 ), .Q ( new_AGEMA_signal_18604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7112 ( .C ( clk ), .D ( new_AGEMA_signal_18611 ), .Q ( new_AGEMA_signal_18612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7210 ( .C ( clk ), .D ( new_AGEMA_signal_18709 ), .Q ( new_AGEMA_signal_18710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7230 ( .C ( clk ), .D ( new_AGEMA_signal_18729 ), .Q ( new_AGEMA_signal_18730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7250 ( .C ( clk ), .D ( new_AGEMA_signal_18749 ), .Q ( new_AGEMA_signal_18750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7270 ( .C ( clk ), .D ( new_AGEMA_signal_18769 ), .Q ( new_AGEMA_signal_18770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7312 ( .C ( clk ), .D ( new_AGEMA_signal_18811 ), .Q ( new_AGEMA_signal_18812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7324 ( .C ( clk ), .D ( new_AGEMA_signal_18823 ), .Q ( new_AGEMA_signal_18824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7336 ( .C ( clk ), .D ( new_AGEMA_signal_18835 ), .Q ( new_AGEMA_signal_18836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7348 ( .C ( clk ), .D ( new_AGEMA_signal_18847 ), .Q ( new_AGEMA_signal_18848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7360 ( .C ( clk ), .D ( new_AGEMA_signal_18859 ), .Q ( new_AGEMA_signal_18860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7374 ( .C ( clk ), .D ( new_AGEMA_signal_18873 ), .Q ( new_AGEMA_signal_18874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7388 ( .C ( clk ), .D ( new_AGEMA_signal_18887 ), .Q ( new_AGEMA_signal_18888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7402 ( .C ( clk ), .D ( new_AGEMA_signal_18901 ), .Q ( new_AGEMA_signal_18902 ) ) ;

    /* cells in depth 19 */
    buf_clk new_AGEMA_reg_buffer_6301 ( .C ( clk ), .D ( new_AGEMA_signal_17800 ), .Q ( new_AGEMA_signal_17801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6309 ( .C ( clk ), .D ( new_AGEMA_signal_17808 ), .Q ( new_AGEMA_signal_17809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6317 ( .C ( clk ), .D ( new_AGEMA_signal_17816 ), .Q ( new_AGEMA_signal_17817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6325 ( .C ( clk ), .D ( new_AGEMA_signal_17824 ), .Q ( new_AGEMA_signal_17825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6337 ( .C ( clk ), .D ( new_AGEMA_signal_17836 ), .Q ( new_AGEMA_signal_17837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6349 ( .C ( clk ), .D ( new_AGEMA_signal_17848 ), .Q ( new_AGEMA_signal_17849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6361 ( .C ( clk ), .D ( new_AGEMA_signal_17860 ), .Q ( new_AGEMA_signal_17861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6373 ( .C ( clk ), .D ( new_AGEMA_signal_17872 ), .Q ( new_AGEMA_signal_17873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6387 ( .C ( clk ), .D ( new_AGEMA_signal_17886 ), .Q ( new_AGEMA_signal_17887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6401 ( .C ( clk ), .D ( new_AGEMA_signal_17900 ), .Q ( new_AGEMA_signal_17901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6415 ( .C ( clk ), .D ( new_AGEMA_signal_17914 ), .Q ( new_AGEMA_signal_17915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6429 ( .C ( clk ), .D ( new_AGEMA_signal_17928 ), .Q ( new_AGEMA_signal_17929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6437 ( .C ( clk ), .D ( new_AGEMA_signal_17936 ), .Q ( new_AGEMA_signal_17937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6445 ( .C ( clk ), .D ( new_AGEMA_signal_17944 ), .Q ( new_AGEMA_signal_17945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6453 ( .C ( clk ), .D ( new_AGEMA_signal_17952 ), .Q ( new_AGEMA_signal_17953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6461 ( .C ( clk ), .D ( new_AGEMA_signal_17960 ), .Q ( new_AGEMA_signal_17961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6475 ( .C ( clk ), .D ( new_AGEMA_signal_17974 ), .Q ( new_AGEMA_signal_17975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6489 ( .C ( clk ), .D ( new_AGEMA_signal_17988 ), .Q ( new_AGEMA_signal_17989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6503 ( .C ( clk ), .D ( new_AGEMA_signal_18002 ), .Q ( new_AGEMA_signal_18003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6517 ( .C ( clk ), .D ( new_AGEMA_signal_18016 ), .Q ( new_AGEMA_signal_18017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6525 ( .C ( clk ), .D ( new_AGEMA_signal_18024 ), .Q ( new_AGEMA_signal_18025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6533 ( .C ( clk ), .D ( new_AGEMA_signal_18032 ), .Q ( new_AGEMA_signal_18033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6541 ( .C ( clk ), .D ( new_AGEMA_signal_18040 ), .Q ( new_AGEMA_signal_18041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6549 ( .C ( clk ), .D ( new_AGEMA_signal_18048 ), .Q ( new_AGEMA_signal_18049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6557 ( .C ( clk ), .D ( new_AGEMA_signal_18056 ), .Q ( new_AGEMA_signal_18057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6565 ( .C ( clk ), .D ( new_AGEMA_signal_18064 ), .Q ( new_AGEMA_signal_18065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6573 ( .C ( clk ), .D ( new_AGEMA_signal_18072 ), .Q ( new_AGEMA_signal_18073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6581 ( .C ( clk ), .D ( new_AGEMA_signal_18080 ), .Q ( new_AGEMA_signal_18081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6583 ( .C ( clk ), .D ( n2002 ), .Q ( new_AGEMA_signal_18083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6587 ( .C ( clk ), .D ( new_AGEMA_signal_3510 ), .Q ( new_AGEMA_signal_18087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6591 ( .C ( clk ), .D ( new_AGEMA_signal_3511 ), .Q ( new_AGEMA_signal_18091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6595 ( .C ( clk ), .D ( new_AGEMA_signal_3512 ), .Q ( new_AGEMA_signal_18095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6619 ( .C ( clk ), .D ( new_AGEMA_signal_18118 ), .Q ( new_AGEMA_signal_18119 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6635 ( .C ( clk ), .D ( new_AGEMA_signal_18134 ), .Q ( new_AGEMA_signal_18135 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6651 ( .C ( clk ), .D ( new_AGEMA_signal_18150 ), .Q ( new_AGEMA_signal_18151 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6667 ( .C ( clk ), .D ( new_AGEMA_signal_18166 ), .Q ( new_AGEMA_signal_18167 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6671 ( .C ( clk ), .D ( n2208 ), .Q ( new_AGEMA_signal_18171 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6675 ( .C ( clk ), .D ( new_AGEMA_signal_3537 ), .Q ( new_AGEMA_signal_18175 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6679 ( .C ( clk ), .D ( new_AGEMA_signal_3538 ), .Q ( new_AGEMA_signal_18179 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6683 ( .C ( clk ), .D ( new_AGEMA_signal_3539 ), .Q ( new_AGEMA_signal_18183 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6707 ( .C ( clk ), .D ( new_AGEMA_signal_18206 ), .Q ( new_AGEMA_signal_18207 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6723 ( .C ( clk ), .D ( new_AGEMA_signal_18222 ), .Q ( new_AGEMA_signal_18223 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6739 ( .C ( clk ), .D ( new_AGEMA_signal_18238 ), .Q ( new_AGEMA_signal_18239 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6755 ( .C ( clk ), .D ( new_AGEMA_signal_18254 ), .Q ( new_AGEMA_signal_18255 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6765 ( .C ( clk ), .D ( new_AGEMA_signal_18264 ), .Q ( new_AGEMA_signal_18265 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6775 ( .C ( clk ), .D ( new_AGEMA_signal_18274 ), .Q ( new_AGEMA_signal_18275 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6785 ( .C ( clk ), .D ( new_AGEMA_signal_18284 ), .Q ( new_AGEMA_signal_18285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6795 ( .C ( clk ), .D ( new_AGEMA_signal_18294 ), .Q ( new_AGEMA_signal_18295 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6799 ( .C ( clk ), .D ( n2668 ), .Q ( new_AGEMA_signal_18299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6803 ( .C ( clk ), .D ( new_AGEMA_signal_3570 ), .Q ( new_AGEMA_signal_18303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6807 ( .C ( clk ), .D ( new_AGEMA_signal_3571 ), .Q ( new_AGEMA_signal_18307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6811 ( .C ( clk ), .D ( new_AGEMA_signal_3572 ), .Q ( new_AGEMA_signal_18311 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6819 ( .C ( clk ), .D ( new_AGEMA_signal_18318 ), .Q ( new_AGEMA_signal_18319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6827 ( .C ( clk ), .D ( new_AGEMA_signal_18326 ), .Q ( new_AGEMA_signal_18327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6835 ( .C ( clk ), .D ( new_AGEMA_signal_18334 ), .Q ( new_AGEMA_signal_18335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6843 ( .C ( clk ), .D ( new_AGEMA_signal_18342 ), .Q ( new_AGEMA_signal_18343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6847 ( .C ( clk ), .D ( n2016 ), .Q ( new_AGEMA_signal_18347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6853 ( .C ( clk ), .D ( new_AGEMA_signal_3516 ), .Q ( new_AGEMA_signal_18353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6859 ( .C ( clk ), .D ( new_AGEMA_signal_3517 ), .Q ( new_AGEMA_signal_18359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6865 ( .C ( clk ), .D ( new_AGEMA_signal_3518 ), .Q ( new_AGEMA_signal_18365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6871 ( .C ( clk ), .D ( n2111 ), .Q ( new_AGEMA_signal_18371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6877 ( .C ( clk ), .D ( new_AGEMA_signal_3522 ), .Q ( new_AGEMA_signal_18377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6883 ( .C ( clk ), .D ( new_AGEMA_signal_3523 ), .Q ( new_AGEMA_signal_18383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6889 ( .C ( clk ), .D ( new_AGEMA_signal_3524 ), .Q ( new_AGEMA_signal_18389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6905 ( .C ( clk ), .D ( new_AGEMA_signal_18404 ), .Q ( new_AGEMA_signal_18405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6921 ( .C ( clk ), .D ( new_AGEMA_signal_18420 ), .Q ( new_AGEMA_signal_18421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6937 ( .C ( clk ), .D ( new_AGEMA_signal_18436 ), .Q ( new_AGEMA_signal_18437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6953 ( .C ( clk ), .D ( new_AGEMA_signal_18452 ), .Q ( new_AGEMA_signal_18453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6963 ( .C ( clk ), .D ( new_AGEMA_signal_18462 ), .Q ( new_AGEMA_signal_18463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6973 ( .C ( clk ), .D ( new_AGEMA_signal_18472 ), .Q ( new_AGEMA_signal_18473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6983 ( .C ( clk ), .D ( new_AGEMA_signal_18482 ), .Q ( new_AGEMA_signal_18483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6993 ( .C ( clk ), .D ( new_AGEMA_signal_18492 ), .Q ( new_AGEMA_signal_18493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7011 ( .C ( clk ), .D ( new_AGEMA_signal_18510 ), .Q ( new_AGEMA_signal_18511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7029 ( .C ( clk ), .D ( new_AGEMA_signal_18528 ), .Q ( new_AGEMA_signal_18529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7047 ( .C ( clk ), .D ( new_AGEMA_signal_18546 ), .Q ( new_AGEMA_signal_18547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7065 ( .C ( clk ), .D ( new_AGEMA_signal_18564 ), .Q ( new_AGEMA_signal_18565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7089 ( .C ( clk ), .D ( new_AGEMA_signal_18588 ), .Q ( new_AGEMA_signal_18589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7097 ( .C ( clk ), .D ( new_AGEMA_signal_18596 ), .Q ( new_AGEMA_signal_18597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7105 ( .C ( clk ), .D ( new_AGEMA_signal_18604 ), .Q ( new_AGEMA_signal_18605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7113 ( .C ( clk ), .D ( new_AGEMA_signal_18612 ), .Q ( new_AGEMA_signal_18613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7135 ( .C ( clk ), .D ( n2019 ), .Q ( new_AGEMA_signal_18635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7143 ( .C ( clk ), .D ( new_AGEMA_signal_3507 ), .Q ( new_AGEMA_signal_18643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7151 ( .C ( clk ), .D ( new_AGEMA_signal_3508 ), .Q ( new_AGEMA_signal_18651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7159 ( .C ( clk ), .D ( new_AGEMA_signal_3509 ), .Q ( new_AGEMA_signal_18659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7211 ( .C ( clk ), .D ( new_AGEMA_signal_18710 ), .Q ( new_AGEMA_signal_18711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7231 ( .C ( clk ), .D ( new_AGEMA_signal_18730 ), .Q ( new_AGEMA_signal_18731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7251 ( .C ( clk ), .D ( new_AGEMA_signal_18750 ), .Q ( new_AGEMA_signal_18751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7271 ( .C ( clk ), .D ( new_AGEMA_signal_18770 ), .Q ( new_AGEMA_signal_18771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7313 ( .C ( clk ), .D ( new_AGEMA_signal_18812 ), .Q ( new_AGEMA_signal_18813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7325 ( .C ( clk ), .D ( new_AGEMA_signal_18824 ), .Q ( new_AGEMA_signal_18825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7337 ( .C ( clk ), .D ( new_AGEMA_signal_18836 ), .Q ( new_AGEMA_signal_18837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7349 ( .C ( clk ), .D ( new_AGEMA_signal_18848 ), .Q ( new_AGEMA_signal_18849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7361 ( .C ( clk ), .D ( new_AGEMA_signal_18860 ), .Q ( new_AGEMA_signal_18861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7375 ( .C ( clk ), .D ( new_AGEMA_signal_18874 ), .Q ( new_AGEMA_signal_18875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7389 ( .C ( clk ), .D ( new_AGEMA_signal_18888 ), .Q ( new_AGEMA_signal_18889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7403 ( .C ( clk ), .D ( new_AGEMA_signal_18902 ), .Q ( new_AGEMA_signal_18903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7415 ( .C ( clk ), .D ( n2426 ), .Q ( new_AGEMA_signal_18915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7429 ( .C ( clk ), .D ( new_AGEMA_signal_3555 ), .Q ( new_AGEMA_signal_18929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7443 ( .C ( clk ), .D ( new_AGEMA_signal_3556 ), .Q ( new_AGEMA_signal_18943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7457 ( .C ( clk ), .D ( new_AGEMA_signal_3557 ), .Q ( new_AGEMA_signal_18957 ) ) ;

    /* cells in depth 20 */
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2117 ( .ina ({new_AGEMA_signal_17426, new_AGEMA_signal_17420, new_AGEMA_signal_17414, new_AGEMA_signal_17408}), .inb ({new_AGEMA_signal_3515, new_AGEMA_signal_3514, new_AGEMA_signal_3513, n1989}), .clk ( clk ), .rnd ({Fresh[8179], Fresh[8178], Fresh[8177], Fresh[8176], Fresh[8175], Fresh[8174], Fresh[8173], Fresh[8172], Fresh[8171], Fresh[8170]}), .outt ({new_AGEMA_signal_3581, new_AGEMA_signal_3580, new_AGEMA_signal_3579, n2000}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2181 ( .ina ({new_AGEMA_signal_3437, new_AGEMA_signal_3436, new_AGEMA_signal_3435, n2038}), .inb ({new_AGEMA_signal_17442, new_AGEMA_signal_17438, new_AGEMA_signal_17434, new_AGEMA_signal_17430}), .clk ( clk ), .rnd ({Fresh[8189], Fresh[8188], Fresh[8187], Fresh[8186], Fresh[8185], Fresh[8184], Fresh[8183], Fresh[8182], Fresh[8181], Fresh[8180]}), .outt ({new_AGEMA_signal_3521, new_AGEMA_signal_3520, new_AGEMA_signal_3519, n2113}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2231 ( .ina ({new_AGEMA_signal_3527, new_AGEMA_signal_3526, new_AGEMA_signal_3525, n2079}), .inb ({new_AGEMA_signal_17466, new_AGEMA_signal_17460, new_AGEMA_signal_17454, new_AGEMA_signal_17448}), .clk ( clk ), .rnd ({Fresh[8199], Fresh[8198], Fresh[8197], Fresh[8196], Fresh[8195], Fresh[8194], Fresh[8193], Fresh[8192], Fresh[8191], Fresh[8190]}), .outt ({new_AGEMA_signal_3584, new_AGEMA_signal_3583, new_AGEMA_signal_3582, n2109}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2264 ( .ina ({new_AGEMA_signal_17506, new_AGEMA_signal_17496, new_AGEMA_signal_17486, new_AGEMA_signal_17476}), .inb ({new_AGEMA_signal_3530, new_AGEMA_signal_3529, new_AGEMA_signal_3528, n2104}), .clk ( clk ), .rnd ({Fresh[8209], Fresh[8208], Fresh[8207], Fresh[8206], Fresh[8205], Fresh[8204], Fresh[8203], Fresh[8202], Fresh[8201], Fresh[8200]}), .outt ({new_AGEMA_signal_3587, new_AGEMA_signal_3586, new_AGEMA_signal_3585, n2107}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2290 ( .ina ({new_AGEMA_signal_17530, new_AGEMA_signal_17524, new_AGEMA_signal_17518, new_AGEMA_signal_17512}), .inb ({new_AGEMA_signal_3533, new_AGEMA_signal_3532, new_AGEMA_signal_3531, n2127}), .clk ( clk ), .rnd ({Fresh[8219], Fresh[8218], Fresh[8217], Fresh[8216], Fresh[8215], Fresh[8214], Fresh[8213], Fresh[8212], Fresh[8211], Fresh[8210]}), .outt ({new_AGEMA_signal_3590, new_AGEMA_signal_3589, new_AGEMA_signal_3588, n2212}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2316 ( .ina ({new_AGEMA_signal_17554, new_AGEMA_signal_17548, new_AGEMA_signal_17542, new_AGEMA_signal_17536}), .inb ({new_AGEMA_signal_3536, new_AGEMA_signal_3535, new_AGEMA_signal_3534, n2147}), .clk ( clk ), .rnd ({Fresh[8229], Fresh[8228], Fresh[8227], Fresh[8226], Fresh[8225], Fresh[8224], Fresh[8223], Fresh[8222], Fresh[8221], Fresh[8220]}), .outt ({new_AGEMA_signal_3593, new_AGEMA_signal_3592, new_AGEMA_signal_3591, n2149}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2366 ( .ina ({new_AGEMA_signal_3542, new_AGEMA_signal_3541, new_AGEMA_signal_3540, n2199}), .inb ({new_AGEMA_signal_17570, new_AGEMA_signal_17566, new_AGEMA_signal_17562, new_AGEMA_signal_17558}), .clk ( clk ), .rnd ({Fresh[8239], Fresh[8238], Fresh[8237], Fresh[8236], Fresh[8235], Fresh[8234], Fresh[8233], Fresh[8232], Fresh[8231], Fresh[8230]}), .outt ({new_AGEMA_signal_3596, new_AGEMA_signal_3595, new_AGEMA_signal_3594, n2206}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2421 ( .ina ({new_AGEMA_signal_17586, new_AGEMA_signal_17582, new_AGEMA_signal_17578, new_AGEMA_signal_17574}), .inb ({new_AGEMA_signal_3545, new_AGEMA_signal_3544, new_AGEMA_signal_3543, n2257}), .clk ( clk ), .rnd ({Fresh[8249], Fresh[8248], Fresh[8247], Fresh[8246], Fresh[8245], Fresh[8244], Fresh[8243], Fresh[8242], Fresh[8241], Fresh[8240]}), .outt ({new_AGEMA_signal_3599, new_AGEMA_signal_3598, new_AGEMA_signal_3597, n2310}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2447 ( .ina ({new_AGEMA_signal_3548, new_AGEMA_signal_3547, new_AGEMA_signal_3546, n2281}), .inb ({new_AGEMA_signal_17618, new_AGEMA_signal_17610, new_AGEMA_signal_17602, new_AGEMA_signal_17594}), .clk ( clk ), .rnd ({Fresh[8259], Fresh[8258], Fresh[8257], Fresh[8256], Fresh[8255], Fresh[8254], Fresh[8253], Fresh[8252], Fresh[8251], Fresh[8250]}), .outt ({new_AGEMA_signal_3602, new_AGEMA_signal_3601, new_AGEMA_signal_3600, n2308}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2476 ( .ina ({new_AGEMA_signal_17642, new_AGEMA_signal_17636, new_AGEMA_signal_17630, new_AGEMA_signal_17624}), .inb ({new_AGEMA_signal_3551, new_AGEMA_signal_3550, new_AGEMA_signal_3549, n2305}), .clk ( clk ), .rnd ({Fresh[8269], Fresh[8268], Fresh[8267], Fresh[8266], Fresh[8265], Fresh[8264], Fresh[8263], Fresh[8262], Fresh[8261], Fresh[8260]}), .outt ({new_AGEMA_signal_3605, new_AGEMA_signal_3604, new_AGEMA_signal_3603, n2307}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2533 ( .ina ({new_AGEMA_signal_17674, new_AGEMA_signal_17666, new_AGEMA_signal_17658, new_AGEMA_signal_17650}), .inb ({new_AGEMA_signal_3554, new_AGEMA_signal_3553, new_AGEMA_signal_3552, n2368}), .clk ( clk ), .rnd ({Fresh[8279], Fresh[8278], Fresh[8277], Fresh[8276], Fresh[8275], Fresh[8274], Fresh[8273], Fresh[8272], Fresh[8271], Fresh[8270]}), .outt ({new_AGEMA_signal_3608, new_AGEMA_signal_3607, new_AGEMA_signal_3606, n2370}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2611 ( .ina ({new_AGEMA_signal_3560, new_AGEMA_signal_3559, new_AGEMA_signal_3558, n2457}), .inb ({new_AGEMA_signal_17706, new_AGEMA_signal_17698, new_AGEMA_signal_17690, new_AGEMA_signal_17682}), .clk ( clk ), .rnd ({Fresh[8289], Fresh[8288], Fresh[8287], Fresh[8286], Fresh[8285], Fresh[8284], Fresh[8283], Fresh[8282], Fresh[8281], Fresh[8280]}), .outt ({new_AGEMA_signal_3611, new_AGEMA_signal_3610, new_AGEMA_signal_3609, n2530}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2660 ( .ina ({new_AGEMA_signal_17714, new_AGEMA_signal_17712, new_AGEMA_signal_17710, new_AGEMA_signal_17708}), .inb ({new_AGEMA_signal_3563, new_AGEMA_signal_3562, new_AGEMA_signal_3561, n2513}), .clk ( clk ), .rnd ({Fresh[8299], Fresh[8298], Fresh[8297], Fresh[8296], Fresh[8295], Fresh[8294], Fresh[8293], Fresh[8292], Fresh[8291], Fresh[8290]}), .outt ({new_AGEMA_signal_3614, new_AGEMA_signal_3613, new_AGEMA_signal_3612, n2515}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2718 ( .ina ({new_AGEMA_signal_17730, new_AGEMA_signal_17726, new_AGEMA_signal_17722, new_AGEMA_signal_17718}), .inb ({new_AGEMA_signal_3566, new_AGEMA_signal_3565, new_AGEMA_signal_3564, n2592}), .clk ( clk ), .rnd ({Fresh[8309], Fresh[8308], Fresh[8307], Fresh[8306], Fresh[8305], Fresh[8304], Fresh[8303], Fresh[8302], Fresh[8301], Fresh[8300]}), .outt ({new_AGEMA_signal_3617, new_AGEMA_signal_3616, new_AGEMA_signal_3615, n2639}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2749 ( .ina ({new_AGEMA_signal_3497, new_AGEMA_signal_3496, new_AGEMA_signal_3495, n2637}), .inb ({new_AGEMA_signal_17746, new_AGEMA_signal_17742, new_AGEMA_signal_17738, new_AGEMA_signal_17734}), .clk ( clk ), .rnd ({Fresh[8319], Fresh[8318], Fresh[8317], Fresh[8316], Fresh[8315], Fresh[8314], Fresh[8313], Fresh[8312], Fresh[8311], Fresh[8310]}), .outt ({new_AGEMA_signal_3569, new_AGEMA_signal_3568, new_AGEMA_signal_3567, n2638}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2788 ( .ina ({new_AGEMA_signal_17778, new_AGEMA_signal_17770, new_AGEMA_signal_17762, new_AGEMA_signal_17754}), .inb ({new_AGEMA_signal_3575, new_AGEMA_signal_3574, new_AGEMA_signal_3573, n2705}), .clk ( clk ), .rnd ({Fresh[8329], Fresh[8328], Fresh[8327], Fresh[8326], Fresh[8325], Fresh[8324], Fresh[8323], Fresh[8322], Fresh[8321], Fresh[8320]}), .outt ({new_AGEMA_signal_3620, new_AGEMA_signal_3619, new_AGEMA_signal_3618, n2832}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2842 ( .ina ({new_AGEMA_signal_17794, new_AGEMA_signal_17790, new_AGEMA_signal_17786, new_AGEMA_signal_17782}), .inb ({new_AGEMA_signal_3506, new_AGEMA_signal_3505, new_AGEMA_signal_3504, n2805}), .clk ( clk ), .rnd ({Fresh[8339], Fresh[8338], Fresh[8337], Fresh[8336], Fresh[8335], Fresh[8334], Fresh[8333], Fresh[8332], Fresh[8331], Fresh[8330]}), .outt ({new_AGEMA_signal_3578, new_AGEMA_signal_3577, new_AGEMA_signal_3576, n2807}) ) ;
    buf_clk new_AGEMA_reg_buffer_6302 ( .C ( clk ), .D ( new_AGEMA_signal_17801 ), .Q ( new_AGEMA_signal_17802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6310 ( .C ( clk ), .D ( new_AGEMA_signal_17809 ), .Q ( new_AGEMA_signal_17810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6318 ( .C ( clk ), .D ( new_AGEMA_signal_17817 ), .Q ( new_AGEMA_signal_17818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6326 ( .C ( clk ), .D ( new_AGEMA_signal_17825 ), .Q ( new_AGEMA_signal_17826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6338 ( .C ( clk ), .D ( new_AGEMA_signal_17837 ), .Q ( new_AGEMA_signal_17838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6350 ( .C ( clk ), .D ( new_AGEMA_signal_17849 ), .Q ( new_AGEMA_signal_17850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6362 ( .C ( clk ), .D ( new_AGEMA_signal_17861 ), .Q ( new_AGEMA_signal_17862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6374 ( .C ( clk ), .D ( new_AGEMA_signal_17873 ), .Q ( new_AGEMA_signal_17874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6388 ( .C ( clk ), .D ( new_AGEMA_signal_17887 ), .Q ( new_AGEMA_signal_17888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6402 ( .C ( clk ), .D ( new_AGEMA_signal_17901 ), .Q ( new_AGEMA_signal_17902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6416 ( .C ( clk ), .D ( new_AGEMA_signal_17915 ), .Q ( new_AGEMA_signal_17916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6430 ( .C ( clk ), .D ( new_AGEMA_signal_17929 ), .Q ( new_AGEMA_signal_17930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6438 ( .C ( clk ), .D ( new_AGEMA_signal_17937 ), .Q ( new_AGEMA_signal_17938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6446 ( .C ( clk ), .D ( new_AGEMA_signal_17945 ), .Q ( new_AGEMA_signal_17946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6454 ( .C ( clk ), .D ( new_AGEMA_signal_17953 ), .Q ( new_AGEMA_signal_17954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6462 ( .C ( clk ), .D ( new_AGEMA_signal_17961 ), .Q ( new_AGEMA_signal_17962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6476 ( .C ( clk ), .D ( new_AGEMA_signal_17975 ), .Q ( new_AGEMA_signal_17976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6490 ( .C ( clk ), .D ( new_AGEMA_signal_17989 ), .Q ( new_AGEMA_signal_17990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6504 ( .C ( clk ), .D ( new_AGEMA_signal_18003 ), .Q ( new_AGEMA_signal_18004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6518 ( .C ( clk ), .D ( new_AGEMA_signal_18017 ), .Q ( new_AGEMA_signal_18018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6526 ( .C ( clk ), .D ( new_AGEMA_signal_18025 ), .Q ( new_AGEMA_signal_18026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6534 ( .C ( clk ), .D ( new_AGEMA_signal_18033 ), .Q ( new_AGEMA_signal_18034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6542 ( .C ( clk ), .D ( new_AGEMA_signal_18041 ), .Q ( new_AGEMA_signal_18042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6550 ( .C ( clk ), .D ( new_AGEMA_signal_18049 ), .Q ( new_AGEMA_signal_18050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6558 ( .C ( clk ), .D ( new_AGEMA_signal_18057 ), .Q ( new_AGEMA_signal_18058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6566 ( .C ( clk ), .D ( new_AGEMA_signal_18065 ), .Q ( new_AGEMA_signal_18066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6574 ( .C ( clk ), .D ( new_AGEMA_signal_18073 ), .Q ( new_AGEMA_signal_18074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6582 ( .C ( clk ), .D ( new_AGEMA_signal_18081 ), .Q ( new_AGEMA_signal_18082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6584 ( .C ( clk ), .D ( new_AGEMA_signal_18083 ), .Q ( new_AGEMA_signal_18084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6588 ( .C ( clk ), .D ( new_AGEMA_signal_18087 ), .Q ( new_AGEMA_signal_18088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6592 ( .C ( clk ), .D ( new_AGEMA_signal_18091 ), .Q ( new_AGEMA_signal_18092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6596 ( .C ( clk ), .D ( new_AGEMA_signal_18095 ), .Q ( new_AGEMA_signal_18096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6620 ( .C ( clk ), .D ( new_AGEMA_signal_18119 ), .Q ( new_AGEMA_signal_18120 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6636 ( .C ( clk ), .D ( new_AGEMA_signal_18135 ), .Q ( new_AGEMA_signal_18136 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6652 ( .C ( clk ), .D ( new_AGEMA_signal_18151 ), .Q ( new_AGEMA_signal_18152 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6668 ( .C ( clk ), .D ( new_AGEMA_signal_18167 ), .Q ( new_AGEMA_signal_18168 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6672 ( .C ( clk ), .D ( new_AGEMA_signal_18171 ), .Q ( new_AGEMA_signal_18172 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6676 ( .C ( clk ), .D ( new_AGEMA_signal_18175 ), .Q ( new_AGEMA_signal_18176 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6680 ( .C ( clk ), .D ( new_AGEMA_signal_18179 ), .Q ( new_AGEMA_signal_18180 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6684 ( .C ( clk ), .D ( new_AGEMA_signal_18183 ), .Q ( new_AGEMA_signal_18184 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6708 ( .C ( clk ), .D ( new_AGEMA_signal_18207 ), .Q ( new_AGEMA_signal_18208 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6724 ( .C ( clk ), .D ( new_AGEMA_signal_18223 ), .Q ( new_AGEMA_signal_18224 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6740 ( .C ( clk ), .D ( new_AGEMA_signal_18239 ), .Q ( new_AGEMA_signal_18240 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6756 ( .C ( clk ), .D ( new_AGEMA_signal_18255 ), .Q ( new_AGEMA_signal_18256 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6766 ( .C ( clk ), .D ( new_AGEMA_signal_18265 ), .Q ( new_AGEMA_signal_18266 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6776 ( .C ( clk ), .D ( new_AGEMA_signal_18275 ), .Q ( new_AGEMA_signal_18276 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6786 ( .C ( clk ), .D ( new_AGEMA_signal_18285 ), .Q ( new_AGEMA_signal_18286 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6796 ( .C ( clk ), .D ( new_AGEMA_signal_18295 ), .Q ( new_AGEMA_signal_18296 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6800 ( .C ( clk ), .D ( new_AGEMA_signal_18299 ), .Q ( new_AGEMA_signal_18300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6804 ( .C ( clk ), .D ( new_AGEMA_signal_18303 ), .Q ( new_AGEMA_signal_18304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6808 ( .C ( clk ), .D ( new_AGEMA_signal_18307 ), .Q ( new_AGEMA_signal_18308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6812 ( .C ( clk ), .D ( new_AGEMA_signal_18311 ), .Q ( new_AGEMA_signal_18312 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6820 ( .C ( clk ), .D ( new_AGEMA_signal_18319 ), .Q ( new_AGEMA_signal_18320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6828 ( .C ( clk ), .D ( new_AGEMA_signal_18327 ), .Q ( new_AGEMA_signal_18328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6836 ( .C ( clk ), .D ( new_AGEMA_signal_18335 ), .Q ( new_AGEMA_signal_18336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6844 ( .C ( clk ), .D ( new_AGEMA_signal_18343 ), .Q ( new_AGEMA_signal_18344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6848 ( .C ( clk ), .D ( new_AGEMA_signal_18347 ), .Q ( new_AGEMA_signal_18348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6854 ( .C ( clk ), .D ( new_AGEMA_signal_18353 ), .Q ( new_AGEMA_signal_18354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6860 ( .C ( clk ), .D ( new_AGEMA_signal_18359 ), .Q ( new_AGEMA_signal_18360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6866 ( .C ( clk ), .D ( new_AGEMA_signal_18365 ), .Q ( new_AGEMA_signal_18366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6872 ( .C ( clk ), .D ( new_AGEMA_signal_18371 ), .Q ( new_AGEMA_signal_18372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6878 ( .C ( clk ), .D ( new_AGEMA_signal_18377 ), .Q ( new_AGEMA_signal_18378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6884 ( .C ( clk ), .D ( new_AGEMA_signal_18383 ), .Q ( new_AGEMA_signal_18384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6890 ( .C ( clk ), .D ( new_AGEMA_signal_18389 ), .Q ( new_AGEMA_signal_18390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6906 ( .C ( clk ), .D ( new_AGEMA_signal_18405 ), .Q ( new_AGEMA_signal_18406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6922 ( .C ( clk ), .D ( new_AGEMA_signal_18421 ), .Q ( new_AGEMA_signal_18422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6938 ( .C ( clk ), .D ( new_AGEMA_signal_18437 ), .Q ( new_AGEMA_signal_18438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6954 ( .C ( clk ), .D ( new_AGEMA_signal_18453 ), .Q ( new_AGEMA_signal_18454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6964 ( .C ( clk ), .D ( new_AGEMA_signal_18463 ), .Q ( new_AGEMA_signal_18464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6974 ( .C ( clk ), .D ( new_AGEMA_signal_18473 ), .Q ( new_AGEMA_signal_18474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6984 ( .C ( clk ), .D ( new_AGEMA_signal_18483 ), .Q ( new_AGEMA_signal_18484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6994 ( .C ( clk ), .D ( new_AGEMA_signal_18493 ), .Q ( new_AGEMA_signal_18494 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7012 ( .C ( clk ), .D ( new_AGEMA_signal_18511 ), .Q ( new_AGEMA_signal_18512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7030 ( .C ( clk ), .D ( new_AGEMA_signal_18529 ), .Q ( new_AGEMA_signal_18530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7048 ( .C ( clk ), .D ( new_AGEMA_signal_18547 ), .Q ( new_AGEMA_signal_18548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7066 ( .C ( clk ), .D ( new_AGEMA_signal_18565 ), .Q ( new_AGEMA_signal_18566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7090 ( .C ( clk ), .D ( new_AGEMA_signal_18589 ), .Q ( new_AGEMA_signal_18590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7098 ( .C ( clk ), .D ( new_AGEMA_signal_18597 ), .Q ( new_AGEMA_signal_18598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7106 ( .C ( clk ), .D ( new_AGEMA_signal_18605 ), .Q ( new_AGEMA_signal_18606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7114 ( .C ( clk ), .D ( new_AGEMA_signal_18613 ), .Q ( new_AGEMA_signal_18614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7136 ( .C ( clk ), .D ( new_AGEMA_signal_18635 ), .Q ( new_AGEMA_signal_18636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7144 ( .C ( clk ), .D ( new_AGEMA_signal_18643 ), .Q ( new_AGEMA_signal_18644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7152 ( .C ( clk ), .D ( new_AGEMA_signal_18651 ), .Q ( new_AGEMA_signal_18652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7160 ( .C ( clk ), .D ( new_AGEMA_signal_18659 ), .Q ( new_AGEMA_signal_18660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7212 ( .C ( clk ), .D ( new_AGEMA_signal_18711 ), .Q ( new_AGEMA_signal_18712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7232 ( .C ( clk ), .D ( new_AGEMA_signal_18731 ), .Q ( new_AGEMA_signal_18732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7252 ( .C ( clk ), .D ( new_AGEMA_signal_18751 ), .Q ( new_AGEMA_signal_18752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7272 ( .C ( clk ), .D ( new_AGEMA_signal_18771 ), .Q ( new_AGEMA_signal_18772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7314 ( .C ( clk ), .D ( new_AGEMA_signal_18813 ), .Q ( new_AGEMA_signal_18814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7326 ( .C ( clk ), .D ( new_AGEMA_signal_18825 ), .Q ( new_AGEMA_signal_18826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7338 ( .C ( clk ), .D ( new_AGEMA_signal_18837 ), .Q ( new_AGEMA_signal_18838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7350 ( .C ( clk ), .D ( new_AGEMA_signal_18849 ), .Q ( new_AGEMA_signal_18850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7362 ( .C ( clk ), .D ( new_AGEMA_signal_18861 ), .Q ( new_AGEMA_signal_18862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7376 ( .C ( clk ), .D ( new_AGEMA_signal_18875 ), .Q ( new_AGEMA_signal_18876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7390 ( .C ( clk ), .D ( new_AGEMA_signal_18889 ), .Q ( new_AGEMA_signal_18890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7404 ( .C ( clk ), .D ( new_AGEMA_signal_18903 ), .Q ( new_AGEMA_signal_18904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7416 ( .C ( clk ), .D ( new_AGEMA_signal_18915 ), .Q ( new_AGEMA_signal_18916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7430 ( .C ( clk ), .D ( new_AGEMA_signal_18929 ), .Q ( new_AGEMA_signal_18930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7444 ( .C ( clk ), .D ( new_AGEMA_signal_18943 ), .Q ( new_AGEMA_signal_18944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7458 ( .C ( clk ), .D ( new_AGEMA_signal_18957 ), .Q ( new_AGEMA_signal_18958 ) ) ;

    /* cells in depth 21 */
    buf_clk new_AGEMA_reg_buffer_6585 ( .C ( clk ), .D ( new_AGEMA_signal_18084 ), .Q ( new_AGEMA_signal_18085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6589 ( .C ( clk ), .D ( new_AGEMA_signal_18088 ), .Q ( new_AGEMA_signal_18089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6593 ( .C ( clk ), .D ( new_AGEMA_signal_18092 ), .Q ( new_AGEMA_signal_18093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6597 ( .C ( clk ), .D ( new_AGEMA_signal_18096 ), .Q ( new_AGEMA_signal_18097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6599 ( .C ( clk ), .D ( n2109 ), .Q ( new_AGEMA_signal_18099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6601 ( .C ( clk ), .D ( new_AGEMA_signal_3582 ), .Q ( new_AGEMA_signal_18101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6603 ( .C ( clk ), .D ( new_AGEMA_signal_3583 ), .Q ( new_AGEMA_signal_18103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6605 ( .C ( clk ), .D ( new_AGEMA_signal_3584 ), .Q ( new_AGEMA_signal_18105 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6621 ( .C ( clk ), .D ( new_AGEMA_signal_18120 ), .Q ( new_AGEMA_signal_18121 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6637 ( .C ( clk ), .D ( new_AGEMA_signal_18136 ), .Q ( new_AGEMA_signal_18137 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6653 ( .C ( clk ), .D ( new_AGEMA_signal_18152 ), .Q ( new_AGEMA_signal_18153 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6669 ( .C ( clk ), .D ( new_AGEMA_signal_18168 ), .Q ( new_AGEMA_signal_18169 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6673 ( .C ( clk ), .D ( new_AGEMA_signal_18172 ), .Q ( new_AGEMA_signal_18173 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6677 ( .C ( clk ), .D ( new_AGEMA_signal_18176 ), .Q ( new_AGEMA_signal_18177 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6681 ( .C ( clk ), .D ( new_AGEMA_signal_18180 ), .Q ( new_AGEMA_signal_18181 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6685 ( .C ( clk ), .D ( new_AGEMA_signal_18184 ), .Q ( new_AGEMA_signal_18185 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6687 ( .C ( clk ), .D ( n2310 ), .Q ( new_AGEMA_signal_18187 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6689 ( .C ( clk ), .D ( new_AGEMA_signal_3597 ), .Q ( new_AGEMA_signal_18189 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6691 ( .C ( clk ), .D ( new_AGEMA_signal_3598 ), .Q ( new_AGEMA_signal_18191 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6693 ( .C ( clk ), .D ( new_AGEMA_signal_3599 ), .Q ( new_AGEMA_signal_18193 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6709 ( .C ( clk ), .D ( new_AGEMA_signal_18208 ), .Q ( new_AGEMA_signal_18209 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6725 ( .C ( clk ), .D ( new_AGEMA_signal_18224 ), .Q ( new_AGEMA_signal_18225 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6741 ( .C ( clk ), .D ( new_AGEMA_signal_18240 ), .Q ( new_AGEMA_signal_18241 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6757 ( .C ( clk ), .D ( new_AGEMA_signal_18256 ), .Q ( new_AGEMA_signal_18257 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6767 ( .C ( clk ), .D ( new_AGEMA_signal_18266 ), .Q ( new_AGEMA_signal_18267 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6777 ( .C ( clk ), .D ( new_AGEMA_signal_18276 ), .Q ( new_AGEMA_signal_18277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6787 ( .C ( clk ), .D ( new_AGEMA_signal_18286 ), .Q ( new_AGEMA_signal_18287 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6797 ( .C ( clk ), .D ( new_AGEMA_signal_18296 ), .Q ( new_AGEMA_signal_18297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6801 ( .C ( clk ), .D ( new_AGEMA_signal_18300 ), .Q ( new_AGEMA_signal_18301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6805 ( .C ( clk ), .D ( new_AGEMA_signal_18304 ), .Q ( new_AGEMA_signal_18305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6809 ( .C ( clk ), .D ( new_AGEMA_signal_18308 ), .Q ( new_AGEMA_signal_18309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6813 ( .C ( clk ), .D ( new_AGEMA_signal_18312 ), .Q ( new_AGEMA_signal_18313 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6821 ( .C ( clk ), .D ( new_AGEMA_signal_18320 ), .Q ( new_AGEMA_signal_18321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6829 ( .C ( clk ), .D ( new_AGEMA_signal_18328 ), .Q ( new_AGEMA_signal_18329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6837 ( .C ( clk ), .D ( new_AGEMA_signal_18336 ), .Q ( new_AGEMA_signal_18337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6845 ( .C ( clk ), .D ( new_AGEMA_signal_18344 ), .Q ( new_AGEMA_signal_18345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6849 ( .C ( clk ), .D ( new_AGEMA_signal_18348 ), .Q ( new_AGEMA_signal_18349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6855 ( .C ( clk ), .D ( new_AGEMA_signal_18354 ), .Q ( new_AGEMA_signal_18355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6861 ( .C ( clk ), .D ( new_AGEMA_signal_18360 ), .Q ( new_AGEMA_signal_18361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6867 ( .C ( clk ), .D ( new_AGEMA_signal_18366 ), .Q ( new_AGEMA_signal_18367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6873 ( .C ( clk ), .D ( new_AGEMA_signal_18372 ), .Q ( new_AGEMA_signal_18373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6879 ( .C ( clk ), .D ( new_AGEMA_signal_18378 ), .Q ( new_AGEMA_signal_18379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6885 ( .C ( clk ), .D ( new_AGEMA_signal_18384 ), .Q ( new_AGEMA_signal_18385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6891 ( .C ( clk ), .D ( new_AGEMA_signal_18390 ), .Q ( new_AGEMA_signal_18391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6907 ( .C ( clk ), .D ( new_AGEMA_signal_18406 ), .Q ( new_AGEMA_signal_18407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6923 ( .C ( clk ), .D ( new_AGEMA_signal_18422 ), .Q ( new_AGEMA_signal_18423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6939 ( .C ( clk ), .D ( new_AGEMA_signal_18438 ), .Q ( new_AGEMA_signal_18439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6955 ( .C ( clk ), .D ( new_AGEMA_signal_18454 ), .Q ( new_AGEMA_signal_18455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6965 ( .C ( clk ), .D ( new_AGEMA_signal_18464 ), .Q ( new_AGEMA_signal_18465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6975 ( .C ( clk ), .D ( new_AGEMA_signal_18474 ), .Q ( new_AGEMA_signal_18475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6985 ( .C ( clk ), .D ( new_AGEMA_signal_18484 ), .Q ( new_AGEMA_signal_18485 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6995 ( .C ( clk ), .D ( new_AGEMA_signal_18494 ), .Q ( new_AGEMA_signal_18495 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7013 ( .C ( clk ), .D ( new_AGEMA_signal_18512 ), .Q ( new_AGEMA_signal_18513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7031 ( .C ( clk ), .D ( new_AGEMA_signal_18530 ), .Q ( new_AGEMA_signal_18531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7049 ( .C ( clk ), .D ( new_AGEMA_signal_18548 ), .Q ( new_AGEMA_signal_18549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7067 ( .C ( clk ), .D ( new_AGEMA_signal_18566 ), .Q ( new_AGEMA_signal_18567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7071 ( .C ( clk ), .D ( n2530 ), .Q ( new_AGEMA_signal_18571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7075 ( .C ( clk ), .D ( new_AGEMA_signal_3609 ), .Q ( new_AGEMA_signal_18575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7079 ( .C ( clk ), .D ( new_AGEMA_signal_3610 ), .Q ( new_AGEMA_signal_18579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7083 ( .C ( clk ), .D ( new_AGEMA_signal_3611 ), .Q ( new_AGEMA_signal_18583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7091 ( .C ( clk ), .D ( new_AGEMA_signal_18590 ), .Q ( new_AGEMA_signal_18591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7099 ( .C ( clk ), .D ( new_AGEMA_signal_18598 ), .Q ( new_AGEMA_signal_18599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7107 ( .C ( clk ), .D ( new_AGEMA_signal_18606 ), .Q ( new_AGEMA_signal_18607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7115 ( .C ( clk ), .D ( new_AGEMA_signal_18614 ), .Q ( new_AGEMA_signal_18615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7119 ( .C ( clk ), .D ( n2832 ), .Q ( new_AGEMA_signal_18619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7123 ( .C ( clk ), .D ( new_AGEMA_signal_3618 ), .Q ( new_AGEMA_signal_18623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7127 ( .C ( clk ), .D ( new_AGEMA_signal_3619 ), .Q ( new_AGEMA_signal_18627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7131 ( .C ( clk ), .D ( new_AGEMA_signal_3620 ), .Q ( new_AGEMA_signal_18631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7137 ( .C ( clk ), .D ( new_AGEMA_signal_18636 ), .Q ( new_AGEMA_signal_18637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7145 ( .C ( clk ), .D ( new_AGEMA_signal_18644 ), .Q ( new_AGEMA_signal_18645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7153 ( .C ( clk ), .D ( new_AGEMA_signal_18652 ), .Q ( new_AGEMA_signal_18653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7161 ( .C ( clk ), .D ( new_AGEMA_signal_18660 ), .Q ( new_AGEMA_signal_18661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7167 ( .C ( clk ), .D ( n2113 ), .Q ( new_AGEMA_signal_18667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7173 ( .C ( clk ), .D ( new_AGEMA_signal_3519 ), .Q ( new_AGEMA_signal_18673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7179 ( .C ( clk ), .D ( new_AGEMA_signal_3520 ), .Q ( new_AGEMA_signal_18679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7185 ( .C ( clk ), .D ( new_AGEMA_signal_3521 ), .Q ( new_AGEMA_signal_18685 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7213 ( .C ( clk ), .D ( new_AGEMA_signal_18712 ), .Q ( new_AGEMA_signal_18713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7233 ( .C ( clk ), .D ( new_AGEMA_signal_18732 ), .Q ( new_AGEMA_signal_18733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7253 ( .C ( clk ), .D ( new_AGEMA_signal_18752 ), .Q ( new_AGEMA_signal_18753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7273 ( .C ( clk ), .D ( new_AGEMA_signal_18772 ), .Q ( new_AGEMA_signal_18773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7279 ( .C ( clk ), .D ( n2212 ), .Q ( new_AGEMA_signal_18779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7287 ( .C ( clk ), .D ( new_AGEMA_signal_3588 ), .Q ( new_AGEMA_signal_18787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7295 ( .C ( clk ), .D ( new_AGEMA_signal_3589 ), .Q ( new_AGEMA_signal_18795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7303 ( .C ( clk ), .D ( new_AGEMA_signal_3590 ), .Q ( new_AGEMA_signal_18803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7315 ( .C ( clk ), .D ( new_AGEMA_signal_18814 ), .Q ( new_AGEMA_signal_18815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7327 ( .C ( clk ), .D ( new_AGEMA_signal_18826 ), .Q ( new_AGEMA_signal_18827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7339 ( .C ( clk ), .D ( new_AGEMA_signal_18838 ), .Q ( new_AGEMA_signal_18839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7351 ( .C ( clk ), .D ( new_AGEMA_signal_18850 ), .Q ( new_AGEMA_signal_18851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7363 ( .C ( clk ), .D ( new_AGEMA_signal_18862 ), .Q ( new_AGEMA_signal_18863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7377 ( .C ( clk ), .D ( new_AGEMA_signal_18876 ), .Q ( new_AGEMA_signal_18877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7391 ( .C ( clk ), .D ( new_AGEMA_signal_18890 ), .Q ( new_AGEMA_signal_18891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7405 ( .C ( clk ), .D ( new_AGEMA_signal_18904 ), .Q ( new_AGEMA_signal_18905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7417 ( .C ( clk ), .D ( new_AGEMA_signal_18916 ), .Q ( new_AGEMA_signal_18917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7431 ( .C ( clk ), .D ( new_AGEMA_signal_18930 ), .Q ( new_AGEMA_signal_18931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7445 ( .C ( clk ), .D ( new_AGEMA_signal_18944 ), .Q ( new_AGEMA_signal_18945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7459 ( .C ( clk ), .D ( new_AGEMA_signal_18958 ), .Q ( new_AGEMA_signal_18959 ) ) ;

    /* cells in depth 22 */
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2129 ( .ina ({new_AGEMA_signal_3581, new_AGEMA_signal_3580, new_AGEMA_signal_3579, n2000}), .inb ({new_AGEMA_signal_17826, new_AGEMA_signal_17818, new_AGEMA_signal_17810, new_AGEMA_signal_17802}), .clk ( clk ), .rnd ({Fresh[8349], Fresh[8348], Fresh[8347], Fresh[8346], Fresh[8345], Fresh[8344], Fresh[8343], Fresh[8342], Fresh[8341], Fresh[8340]}), .outt ({new_AGEMA_signal_3626, new_AGEMA_signal_3625, new_AGEMA_signal_3624, n2001}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2267 ( .ina ({new_AGEMA_signal_3587, new_AGEMA_signal_3586, new_AGEMA_signal_3585, n2107}), .inb ({new_AGEMA_signal_17874, new_AGEMA_signal_17862, new_AGEMA_signal_17850, new_AGEMA_signal_17838}), .clk ( clk ), .rnd ({Fresh[8359], Fresh[8358], Fresh[8357], Fresh[8356], Fresh[8355], Fresh[8354], Fresh[8353], Fresh[8352], Fresh[8351], Fresh[8350]}), .outt ({new_AGEMA_signal_3629, new_AGEMA_signal_3628, new_AGEMA_signal_3627, n2108}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2317 ( .ina ({new_AGEMA_signal_17930, new_AGEMA_signal_17916, new_AGEMA_signal_17902, new_AGEMA_signal_17888}), .inb ({new_AGEMA_signal_3593, new_AGEMA_signal_3592, new_AGEMA_signal_3591, n2149}), .clk ( clk ), .rnd ({Fresh[8369], Fresh[8368], Fresh[8367], Fresh[8366], Fresh[8365], Fresh[8364], Fresh[8363], Fresh[8362], Fresh[8361], Fresh[8360]}), .outt ({new_AGEMA_signal_3632, new_AGEMA_signal_3631, new_AGEMA_signal_3630, n2153}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2374 ( .ina ({new_AGEMA_signal_3596, new_AGEMA_signal_3595, new_AGEMA_signal_3594, n2206}), .inb ({new_AGEMA_signal_17962, new_AGEMA_signal_17954, new_AGEMA_signal_17946, new_AGEMA_signal_17938}), .clk ( clk ), .rnd ({Fresh[8379], Fresh[8378], Fresh[8377], Fresh[8376], Fresh[8375], Fresh[8374], Fresh[8373], Fresh[8372], Fresh[8371], Fresh[8370]}), .outt ({new_AGEMA_signal_3635, new_AGEMA_signal_3634, new_AGEMA_signal_3633, n2207}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2477 ( .ina ({new_AGEMA_signal_3602, new_AGEMA_signal_3601, new_AGEMA_signal_3600, n2308}), .inb ({new_AGEMA_signal_3605, new_AGEMA_signal_3604, new_AGEMA_signal_3603, n2307}), .clk ( clk ), .rnd ({Fresh[8389], Fresh[8388], Fresh[8387], Fresh[8386], Fresh[8385], Fresh[8384], Fresh[8383], Fresh[8382], Fresh[8381], Fresh[8380]}), .outt ({new_AGEMA_signal_3638, new_AGEMA_signal_3637, new_AGEMA_signal_3636, n2309}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2535 ( .ina ({new_AGEMA_signal_3608, new_AGEMA_signal_3607, new_AGEMA_signal_3606, n2370}), .inb ({new_AGEMA_signal_18018, new_AGEMA_signal_18004, new_AGEMA_signal_17990, new_AGEMA_signal_17976}), .clk ( clk ), .rnd ({Fresh[8399], Fresh[8398], Fresh[8397], Fresh[8396], Fresh[8395], Fresh[8394], Fresh[8393], Fresh[8392], Fresh[8391], Fresh[8390]}), .outt ({new_AGEMA_signal_3641, new_AGEMA_signal_3640, new_AGEMA_signal_3639, n2373}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2661 ( .ina ({new_AGEMA_signal_18050, new_AGEMA_signal_18042, new_AGEMA_signal_18034, new_AGEMA_signal_18026}), .inb ({new_AGEMA_signal_3614, new_AGEMA_signal_3613, new_AGEMA_signal_3612, n2515}), .clk ( clk ), .rnd ({Fresh[8409], Fresh[8408], Fresh[8407], Fresh[8406], Fresh[8405], Fresh[8404], Fresh[8403], Fresh[8402], Fresh[8401], Fresh[8400]}), .outt ({new_AGEMA_signal_3644, new_AGEMA_signal_3643, new_AGEMA_signal_3642, n2528}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2750 ( .ina ({new_AGEMA_signal_3617, new_AGEMA_signal_3616, new_AGEMA_signal_3615, n2639}), .inb ({new_AGEMA_signal_3569, new_AGEMA_signal_3568, new_AGEMA_signal_3567, n2638}), .clk ( clk ), .rnd ({Fresh[8419], Fresh[8418], Fresh[8417], Fresh[8416], Fresh[8415], Fresh[8414], Fresh[8413], Fresh[8412], Fresh[8411], Fresh[8410]}), .outt ({new_AGEMA_signal_3647, new_AGEMA_signal_3646, new_AGEMA_signal_3645, n2669}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2843 ( .ina ({new_AGEMA_signal_18082, new_AGEMA_signal_18074, new_AGEMA_signal_18066, new_AGEMA_signal_18058}), .inb ({new_AGEMA_signal_3578, new_AGEMA_signal_3577, new_AGEMA_signal_3576, n2807}), .clk ( clk ), .rnd ({Fresh[8429], Fresh[8428], Fresh[8427], Fresh[8426], Fresh[8425], Fresh[8424], Fresh[8423], Fresh[8422], Fresh[8421], Fresh[8420]}), .outt ({new_AGEMA_signal_3623, new_AGEMA_signal_3622, new_AGEMA_signal_3621, n2830}) ) ;
    buf_clk new_AGEMA_reg_buffer_6586 ( .C ( clk ), .D ( new_AGEMA_signal_18085 ), .Q ( new_AGEMA_signal_18086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6590 ( .C ( clk ), .D ( new_AGEMA_signal_18089 ), .Q ( new_AGEMA_signal_18090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6594 ( .C ( clk ), .D ( new_AGEMA_signal_18093 ), .Q ( new_AGEMA_signal_18094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6598 ( .C ( clk ), .D ( new_AGEMA_signal_18097 ), .Q ( new_AGEMA_signal_18098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6600 ( .C ( clk ), .D ( new_AGEMA_signal_18099 ), .Q ( new_AGEMA_signal_18100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6602 ( .C ( clk ), .D ( new_AGEMA_signal_18101 ), .Q ( new_AGEMA_signal_18102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6604 ( .C ( clk ), .D ( new_AGEMA_signal_18103 ), .Q ( new_AGEMA_signal_18104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6606 ( .C ( clk ), .D ( new_AGEMA_signal_18105 ), .Q ( new_AGEMA_signal_18106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6622 ( .C ( clk ), .D ( new_AGEMA_signal_18121 ), .Q ( new_AGEMA_signal_18122 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6638 ( .C ( clk ), .D ( new_AGEMA_signal_18137 ), .Q ( new_AGEMA_signal_18138 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6654 ( .C ( clk ), .D ( new_AGEMA_signal_18153 ), .Q ( new_AGEMA_signal_18154 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6670 ( .C ( clk ), .D ( new_AGEMA_signal_18169 ), .Q ( new_AGEMA_signal_18170 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6674 ( .C ( clk ), .D ( new_AGEMA_signal_18173 ), .Q ( new_AGEMA_signal_18174 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6678 ( .C ( clk ), .D ( new_AGEMA_signal_18177 ), .Q ( new_AGEMA_signal_18178 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6682 ( .C ( clk ), .D ( new_AGEMA_signal_18181 ), .Q ( new_AGEMA_signal_18182 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6686 ( .C ( clk ), .D ( new_AGEMA_signal_18185 ), .Q ( new_AGEMA_signal_18186 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6688 ( .C ( clk ), .D ( new_AGEMA_signal_18187 ), .Q ( new_AGEMA_signal_18188 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6690 ( .C ( clk ), .D ( new_AGEMA_signal_18189 ), .Q ( new_AGEMA_signal_18190 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6692 ( .C ( clk ), .D ( new_AGEMA_signal_18191 ), .Q ( new_AGEMA_signal_18192 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6694 ( .C ( clk ), .D ( new_AGEMA_signal_18193 ), .Q ( new_AGEMA_signal_18194 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6710 ( .C ( clk ), .D ( new_AGEMA_signal_18209 ), .Q ( new_AGEMA_signal_18210 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6726 ( .C ( clk ), .D ( new_AGEMA_signal_18225 ), .Q ( new_AGEMA_signal_18226 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6742 ( .C ( clk ), .D ( new_AGEMA_signal_18241 ), .Q ( new_AGEMA_signal_18242 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6758 ( .C ( clk ), .D ( new_AGEMA_signal_18257 ), .Q ( new_AGEMA_signal_18258 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6768 ( .C ( clk ), .D ( new_AGEMA_signal_18267 ), .Q ( new_AGEMA_signal_18268 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6778 ( .C ( clk ), .D ( new_AGEMA_signal_18277 ), .Q ( new_AGEMA_signal_18278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6788 ( .C ( clk ), .D ( new_AGEMA_signal_18287 ), .Q ( new_AGEMA_signal_18288 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6798 ( .C ( clk ), .D ( new_AGEMA_signal_18297 ), .Q ( new_AGEMA_signal_18298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6802 ( .C ( clk ), .D ( new_AGEMA_signal_18301 ), .Q ( new_AGEMA_signal_18302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6806 ( .C ( clk ), .D ( new_AGEMA_signal_18305 ), .Q ( new_AGEMA_signal_18306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6810 ( .C ( clk ), .D ( new_AGEMA_signal_18309 ), .Q ( new_AGEMA_signal_18310 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6814 ( .C ( clk ), .D ( new_AGEMA_signal_18313 ), .Q ( new_AGEMA_signal_18314 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6822 ( .C ( clk ), .D ( new_AGEMA_signal_18321 ), .Q ( new_AGEMA_signal_18322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6830 ( .C ( clk ), .D ( new_AGEMA_signal_18329 ), .Q ( new_AGEMA_signal_18330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6838 ( .C ( clk ), .D ( new_AGEMA_signal_18337 ), .Q ( new_AGEMA_signal_18338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6846 ( .C ( clk ), .D ( new_AGEMA_signal_18345 ), .Q ( new_AGEMA_signal_18346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6850 ( .C ( clk ), .D ( new_AGEMA_signal_18349 ), .Q ( new_AGEMA_signal_18350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6856 ( .C ( clk ), .D ( new_AGEMA_signal_18355 ), .Q ( new_AGEMA_signal_18356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6862 ( .C ( clk ), .D ( new_AGEMA_signal_18361 ), .Q ( new_AGEMA_signal_18362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6868 ( .C ( clk ), .D ( new_AGEMA_signal_18367 ), .Q ( new_AGEMA_signal_18368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6874 ( .C ( clk ), .D ( new_AGEMA_signal_18373 ), .Q ( new_AGEMA_signal_18374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6880 ( .C ( clk ), .D ( new_AGEMA_signal_18379 ), .Q ( new_AGEMA_signal_18380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6886 ( .C ( clk ), .D ( new_AGEMA_signal_18385 ), .Q ( new_AGEMA_signal_18386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6892 ( .C ( clk ), .D ( new_AGEMA_signal_18391 ), .Q ( new_AGEMA_signal_18392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6908 ( .C ( clk ), .D ( new_AGEMA_signal_18407 ), .Q ( new_AGEMA_signal_18408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6924 ( .C ( clk ), .D ( new_AGEMA_signal_18423 ), .Q ( new_AGEMA_signal_18424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6940 ( .C ( clk ), .D ( new_AGEMA_signal_18439 ), .Q ( new_AGEMA_signal_18440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6956 ( .C ( clk ), .D ( new_AGEMA_signal_18455 ), .Q ( new_AGEMA_signal_18456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6966 ( .C ( clk ), .D ( new_AGEMA_signal_18465 ), .Q ( new_AGEMA_signal_18466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6976 ( .C ( clk ), .D ( new_AGEMA_signal_18475 ), .Q ( new_AGEMA_signal_18476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6986 ( .C ( clk ), .D ( new_AGEMA_signal_18485 ), .Q ( new_AGEMA_signal_18486 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6996 ( .C ( clk ), .D ( new_AGEMA_signal_18495 ), .Q ( new_AGEMA_signal_18496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7014 ( .C ( clk ), .D ( new_AGEMA_signal_18513 ), .Q ( new_AGEMA_signal_18514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7032 ( .C ( clk ), .D ( new_AGEMA_signal_18531 ), .Q ( new_AGEMA_signal_18532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7050 ( .C ( clk ), .D ( new_AGEMA_signal_18549 ), .Q ( new_AGEMA_signal_18550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7068 ( .C ( clk ), .D ( new_AGEMA_signal_18567 ), .Q ( new_AGEMA_signal_18568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7072 ( .C ( clk ), .D ( new_AGEMA_signal_18571 ), .Q ( new_AGEMA_signal_18572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7076 ( .C ( clk ), .D ( new_AGEMA_signal_18575 ), .Q ( new_AGEMA_signal_18576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7080 ( .C ( clk ), .D ( new_AGEMA_signal_18579 ), .Q ( new_AGEMA_signal_18580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7084 ( .C ( clk ), .D ( new_AGEMA_signal_18583 ), .Q ( new_AGEMA_signal_18584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7092 ( .C ( clk ), .D ( new_AGEMA_signal_18591 ), .Q ( new_AGEMA_signal_18592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7100 ( .C ( clk ), .D ( new_AGEMA_signal_18599 ), .Q ( new_AGEMA_signal_18600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7108 ( .C ( clk ), .D ( new_AGEMA_signal_18607 ), .Q ( new_AGEMA_signal_18608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7116 ( .C ( clk ), .D ( new_AGEMA_signal_18615 ), .Q ( new_AGEMA_signal_18616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7120 ( .C ( clk ), .D ( new_AGEMA_signal_18619 ), .Q ( new_AGEMA_signal_18620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7124 ( .C ( clk ), .D ( new_AGEMA_signal_18623 ), .Q ( new_AGEMA_signal_18624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7128 ( .C ( clk ), .D ( new_AGEMA_signal_18627 ), .Q ( new_AGEMA_signal_18628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7132 ( .C ( clk ), .D ( new_AGEMA_signal_18631 ), .Q ( new_AGEMA_signal_18632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7138 ( .C ( clk ), .D ( new_AGEMA_signal_18637 ), .Q ( new_AGEMA_signal_18638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7146 ( .C ( clk ), .D ( new_AGEMA_signal_18645 ), .Q ( new_AGEMA_signal_18646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7154 ( .C ( clk ), .D ( new_AGEMA_signal_18653 ), .Q ( new_AGEMA_signal_18654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7162 ( .C ( clk ), .D ( new_AGEMA_signal_18661 ), .Q ( new_AGEMA_signal_18662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7168 ( .C ( clk ), .D ( new_AGEMA_signal_18667 ), .Q ( new_AGEMA_signal_18668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7174 ( .C ( clk ), .D ( new_AGEMA_signal_18673 ), .Q ( new_AGEMA_signal_18674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7180 ( .C ( clk ), .D ( new_AGEMA_signal_18679 ), .Q ( new_AGEMA_signal_18680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7186 ( .C ( clk ), .D ( new_AGEMA_signal_18685 ), .Q ( new_AGEMA_signal_18686 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7214 ( .C ( clk ), .D ( new_AGEMA_signal_18713 ), .Q ( new_AGEMA_signal_18714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7234 ( .C ( clk ), .D ( new_AGEMA_signal_18733 ), .Q ( new_AGEMA_signal_18734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7254 ( .C ( clk ), .D ( new_AGEMA_signal_18753 ), .Q ( new_AGEMA_signal_18754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7274 ( .C ( clk ), .D ( new_AGEMA_signal_18773 ), .Q ( new_AGEMA_signal_18774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7280 ( .C ( clk ), .D ( new_AGEMA_signal_18779 ), .Q ( new_AGEMA_signal_18780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7288 ( .C ( clk ), .D ( new_AGEMA_signal_18787 ), .Q ( new_AGEMA_signal_18788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7296 ( .C ( clk ), .D ( new_AGEMA_signal_18795 ), .Q ( new_AGEMA_signal_18796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7304 ( .C ( clk ), .D ( new_AGEMA_signal_18803 ), .Q ( new_AGEMA_signal_18804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7316 ( .C ( clk ), .D ( new_AGEMA_signal_18815 ), .Q ( new_AGEMA_signal_18816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7328 ( .C ( clk ), .D ( new_AGEMA_signal_18827 ), .Q ( new_AGEMA_signal_18828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7340 ( .C ( clk ), .D ( new_AGEMA_signal_18839 ), .Q ( new_AGEMA_signal_18840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7352 ( .C ( clk ), .D ( new_AGEMA_signal_18851 ), .Q ( new_AGEMA_signal_18852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7364 ( .C ( clk ), .D ( new_AGEMA_signal_18863 ), .Q ( new_AGEMA_signal_18864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7378 ( .C ( clk ), .D ( new_AGEMA_signal_18877 ), .Q ( new_AGEMA_signal_18878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7392 ( .C ( clk ), .D ( new_AGEMA_signal_18891 ), .Q ( new_AGEMA_signal_18892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7406 ( .C ( clk ), .D ( new_AGEMA_signal_18905 ), .Q ( new_AGEMA_signal_18906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7418 ( .C ( clk ), .D ( new_AGEMA_signal_18917 ), .Q ( new_AGEMA_signal_18918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7432 ( .C ( clk ), .D ( new_AGEMA_signal_18931 ), .Q ( new_AGEMA_signal_18932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7446 ( .C ( clk ), .D ( new_AGEMA_signal_18945 ), .Q ( new_AGEMA_signal_18946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7460 ( .C ( clk ), .D ( new_AGEMA_signal_18959 ), .Q ( new_AGEMA_signal_18960 ) ) ;

    /* cells in depth 23 */
    buf_clk new_AGEMA_reg_buffer_6851 ( .C ( clk ), .D ( new_AGEMA_signal_18350 ), .Q ( new_AGEMA_signal_18351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6857 ( .C ( clk ), .D ( new_AGEMA_signal_18356 ), .Q ( new_AGEMA_signal_18357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6863 ( .C ( clk ), .D ( new_AGEMA_signal_18362 ), .Q ( new_AGEMA_signal_18363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6869 ( .C ( clk ), .D ( new_AGEMA_signal_18368 ), .Q ( new_AGEMA_signal_18369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6875 ( .C ( clk ), .D ( new_AGEMA_signal_18374 ), .Q ( new_AGEMA_signal_18375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6881 ( .C ( clk ), .D ( new_AGEMA_signal_18380 ), .Q ( new_AGEMA_signal_18381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6887 ( .C ( clk ), .D ( new_AGEMA_signal_18386 ), .Q ( new_AGEMA_signal_18387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6893 ( .C ( clk ), .D ( new_AGEMA_signal_18392 ), .Q ( new_AGEMA_signal_18393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6909 ( .C ( clk ), .D ( new_AGEMA_signal_18408 ), .Q ( new_AGEMA_signal_18409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6925 ( .C ( clk ), .D ( new_AGEMA_signal_18424 ), .Q ( new_AGEMA_signal_18425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6941 ( .C ( clk ), .D ( new_AGEMA_signal_18440 ), .Q ( new_AGEMA_signal_18441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6957 ( .C ( clk ), .D ( new_AGEMA_signal_18456 ), .Q ( new_AGEMA_signal_18457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6967 ( .C ( clk ), .D ( new_AGEMA_signal_18466 ), .Q ( new_AGEMA_signal_18467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6977 ( .C ( clk ), .D ( new_AGEMA_signal_18476 ), .Q ( new_AGEMA_signal_18477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6987 ( .C ( clk ), .D ( new_AGEMA_signal_18486 ), .Q ( new_AGEMA_signal_18487 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6997 ( .C ( clk ), .D ( new_AGEMA_signal_18496 ), .Q ( new_AGEMA_signal_18497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7015 ( .C ( clk ), .D ( new_AGEMA_signal_18514 ), .Q ( new_AGEMA_signal_18515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7033 ( .C ( clk ), .D ( new_AGEMA_signal_18532 ), .Q ( new_AGEMA_signal_18533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7051 ( .C ( clk ), .D ( new_AGEMA_signal_18550 ), .Q ( new_AGEMA_signal_18551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7069 ( .C ( clk ), .D ( new_AGEMA_signal_18568 ), .Q ( new_AGEMA_signal_18569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7073 ( .C ( clk ), .D ( new_AGEMA_signal_18572 ), .Q ( new_AGEMA_signal_18573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7077 ( .C ( clk ), .D ( new_AGEMA_signal_18576 ), .Q ( new_AGEMA_signal_18577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7081 ( .C ( clk ), .D ( new_AGEMA_signal_18580 ), .Q ( new_AGEMA_signal_18581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7085 ( .C ( clk ), .D ( new_AGEMA_signal_18584 ), .Q ( new_AGEMA_signal_18585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7093 ( .C ( clk ), .D ( new_AGEMA_signal_18592 ), .Q ( new_AGEMA_signal_18593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7101 ( .C ( clk ), .D ( new_AGEMA_signal_18600 ), .Q ( new_AGEMA_signal_18601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7109 ( .C ( clk ), .D ( new_AGEMA_signal_18608 ), .Q ( new_AGEMA_signal_18609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7117 ( .C ( clk ), .D ( new_AGEMA_signal_18616 ), .Q ( new_AGEMA_signal_18617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7121 ( .C ( clk ), .D ( new_AGEMA_signal_18620 ), .Q ( new_AGEMA_signal_18621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7125 ( .C ( clk ), .D ( new_AGEMA_signal_18624 ), .Q ( new_AGEMA_signal_18625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7129 ( .C ( clk ), .D ( new_AGEMA_signal_18628 ), .Q ( new_AGEMA_signal_18629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7133 ( .C ( clk ), .D ( new_AGEMA_signal_18632 ), .Q ( new_AGEMA_signal_18633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7139 ( .C ( clk ), .D ( new_AGEMA_signal_18638 ), .Q ( new_AGEMA_signal_18639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7147 ( .C ( clk ), .D ( new_AGEMA_signal_18646 ), .Q ( new_AGEMA_signal_18647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7155 ( .C ( clk ), .D ( new_AGEMA_signal_18654 ), .Q ( new_AGEMA_signal_18655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7163 ( .C ( clk ), .D ( new_AGEMA_signal_18662 ), .Q ( new_AGEMA_signal_18663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7169 ( .C ( clk ), .D ( new_AGEMA_signal_18668 ), .Q ( new_AGEMA_signal_18669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7175 ( .C ( clk ), .D ( new_AGEMA_signal_18674 ), .Q ( new_AGEMA_signal_18675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7181 ( .C ( clk ), .D ( new_AGEMA_signal_18680 ), .Q ( new_AGEMA_signal_18681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7187 ( .C ( clk ), .D ( new_AGEMA_signal_18686 ), .Q ( new_AGEMA_signal_18687 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7215 ( .C ( clk ), .D ( new_AGEMA_signal_18714 ), .Q ( new_AGEMA_signal_18715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7235 ( .C ( clk ), .D ( new_AGEMA_signal_18734 ), .Q ( new_AGEMA_signal_18735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7255 ( .C ( clk ), .D ( new_AGEMA_signal_18754 ), .Q ( new_AGEMA_signal_18755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7275 ( .C ( clk ), .D ( new_AGEMA_signal_18774 ), .Q ( new_AGEMA_signal_18775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7281 ( .C ( clk ), .D ( new_AGEMA_signal_18780 ), .Q ( new_AGEMA_signal_18781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7289 ( .C ( clk ), .D ( new_AGEMA_signal_18788 ), .Q ( new_AGEMA_signal_18789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7297 ( .C ( clk ), .D ( new_AGEMA_signal_18796 ), .Q ( new_AGEMA_signal_18797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7305 ( .C ( clk ), .D ( new_AGEMA_signal_18804 ), .Q ( new_AGEMA_signal_18805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7317 ( .C ( clk ), .D ( new_AGEMA_signal_18816 ), .Q ( new_AGEMA_signal_18817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7329 ( .C ( clk ), .D ( new_AGEMA_signal_18828 ), .Q ( new_AGEMA_signal_18829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7341 ( .C ( clk ), .D ( new_AGEMA_signal_18840 ), .Q ( new_AGEMA_signal_18841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7353 ( .C ( clk ), .D ( new_AGEMA_signal_18852 ), .Q ( new_AGEMA_signal_18853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7365 ( .C ( clk ), .D ( new_AGEMA_signal_18864 ), .Q ( new_AGEMA_signal_18865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7379 ( .C ( clk ), .D ( new_AGEMA_signal_18878 ), .Q ( new_AGEMA_signal_18879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7393 ( .C ( clk ), .D ( new_AGEMA_signal_18892 ), .Q ( new_AGEMA_signal_18893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7407 ( .C ( clk ), .D ( new_AGEMA_signal_18906 ), .Q ( new_AGEMA_signal_18907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7419 ( .C ( clk ), .D ( new_AGEMA_signal_18918 ), .Q ( new_AGEMA_signal_18919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7433 ( .C ( clk ), .D ( new_AGEMA_signal_18932 ), .Q ( new_AGEMA_signal_18933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7447 ( .C ( clk ), .D ( new_AGEMA_signal_18946 ), .Q ( new_AGEMA_signal_18947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7461 ( .C ( clk ), .D ( new_AGEMA_signal_18960 ), .Q ( new_AGEMA_signal_18961 ) ) ;

    /* cells in depth 24 */
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2130 ( .ina ({new_AGEMA_signal_18098, new_AGEMA_signal_18094, new_AGEMA_signal_18090, new_AGEMA_signal_18086}), .inb ({new_AGEMA_signal_3626, new_AGEMA_signal_3625, new_AGEMA_signal_3624, n2001}), .clk ( clk ), .rnd ({Fresh[8439], Fresh[8438], Fresh[8437], Fresh[8436], Fresh[8435], Fresh[8434], Fresh[8433], Fresh[8432], Fresh[8431], Fresh[8430]}), .outt ({new_AGEMA_signal_3653, new_AGEMA_signal_3652, new_AGEMA_signal_3651, n2017}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2268 ( .ina ({new_AGEMA_signal_18106, new_AGEMA_signal_18104, new_AGEMA_signal_18102, new_AGEMA_signal_18100}), .inb ({new_AGEMA_signal_3629, new_AGEMA_signal_3628, new_AGEMA_signal_3627, n2108}), .clk ( clk ), .rnd ({Fresh[8449], Fresh[8448], Fresh[8447], Fresh[8446], Fresh[8445], Fresh[8444], Fresh[8443], Fresh[8442], Fresh[8441], Fresh[8440]}), .outt ({new_AGEMA_signal_3656, new_AGEMA_signal_3655, new_AGEMA_signal_3654, n2110}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2319 ( .ina ({new_AGEMA_signal_3632, new_AGEMA_signal_3631, new_AGEMA_signal_3630, n2153}), .inb ({new_AGEMA_signal_18170, new_AGEMA_signal_18154, new_AGEMA_signal_18138, new_AGEMA_signal_18122}), .clk ( clk ), .rnd ({Fresh[8459], Fresh[8458], Fresh[8457], Fresh[8456], Fresh[8455], Fresh[8454], Fresh[8453], Fresh[8452], Fresh[8451], Fresh[8450]}), .outt ({new_AGEMA_signal_3659, new_AGEMA_signal_3658, new_AGEMA_signal_3657, n2154}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2375 ( .ina ({new_AGEMA_signal_18186, new_AGEMA_signal_18182, new_AGEMA_signal_18178, new_AGEMA_signal_18174}), .inb ({new_AGEMA_signal_3635, new_AGEMA_signal_3634, new_AGEMA_signal_3633, n2207}), .clk ( clk ), .rnd ({Fresh[8469], Fresh[8468], Fresh[8467], Fresh[8466], Fresh[8465], Fresh[8464], Fresh[8463], Fresh[8462], Fresh[8461], Fresh[8460]}), .outt ({new_AGEMA_signal_3662, new_AGEMA_signal_3661, new_AGEMA_signal_3660, n2209}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2478 ( .ina ({new_AGEMA_signal_18194, new_AGEMA_signal_18192, new_AGEMA_signal_18190, new_AGEMA_signal_18188}), .inb ({new_AGEMA_signal_3638, new_AGEMA_signal_3637, new_AGEMA_signal_3636, n2309}), .clk ( clk ), .rnd ({Fresh[8479], Fresh[8478], Fresh[8477], Fresh[8476], Fresh[8475], Fresh[8474], Fresh[8473], Fresh[8472], Fresh[8471], Fresh[8470]}), .outt ({new_AGEMA_signal_3665, new_AGEMA_signal_3664, new_AGEMA_signal_3663, n2311}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2537 ( .ina ({new_AGEMA_signal_3641, new_AGEMA_signal_3640, new_AGEMA_signal_3639, n2373}), .inb ({new_AGEMA_signal_18258, new_AGEMA_signal_18242, new_AGEMA_signal_18226, new_AGEMA_signal_18210}), .clk ( clk ), .rnd ({Fresh[8489], Fresh[8488], Fresh[8487], Fresh[8486], Fresh[8485], Fresh[8484], Fresh[8483], Fresh[8482], Fresh[8481], Fresh[8480]}), .outt ({new_AGEMA_signal_3668, new_AGEMA_signal_3667, new_AGEMA_signal_3666, n2374}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2672 ( .ina ({new_AGEMA_signal_3644, new_AGEMA_signal_3643, new_AGEMA_signal_3642, n2528}), .inb ({new_AGEMA_signal_18298, new_AGEMA_signal_18288, new_AGEMA_signal_18278, new_AGEMA_signal_18268}), .clk ( clk ), .rnd ({Fresh[8499], Fresh[8498], Fresh[8497], Fresh[8496], Fresh[8495], Fresh[8494], Fresh[8493], Fresh[8492], Fresh[8491], Fresh[8490]}), .outt ({new_AGEMA_signal_3671, new_AGEMA_signal_3670, new_AGEMA_signal_3669, n2529}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2768 ( .ina ({new_AGEMA_signal_3647, new_AGEMA_signal_3646, new_AGEMA_signal_3645, n2669}), .inb ({new_AGEMA_signal_18314, new_AGEMA_signal_18310, new_AGEMA_signal_18306, new_AGEMA_signal_18302}), .clk ( clk ), .rnd ({Fresh[8509], Fresh[8508], Fresh[8507], Fresh[8506], Fresh[8505], Fresh[8504], Fresh[8503], Fresh[8502], Fresh[8501], Fresh[8500]}), .outt ({new_AGEMA_signal_3674, new_AGEMA_signal_3673, new_AGEMA_signal_3672, n2670}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2854 ( .ina ({new_AGEMA_signal_3623, new_AGEMA_signal_3622, new_AGEMA_signal_3621, n2830}), .inb ({new_AGEMA_signal_18346, new_AGEMA_signal_18338, new_AGEMA_signal_18330, new_AGEMA_signal_18322}), .clk ( clk ), .rnd ({Fresh[8519], Fresh[8518], Fresh[8517], Fresh[8516], Fresh[8515], Fresh[8514], Fresh[8513], Fresh[8512], Fresh[8511], Fresh[8510]}), .outt ({new_AGEMA_signal_3650, new_AGEMA_signal_3649, new_AGEMA_signal_3648, n2831}) ) ;
    buf_clk new_AGEMA_reg_buffer_6852 ( .C ( clk ), .D ( new_AGEMA_signal_18351 ), .Q ( new_AGEMA_signal_18352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6858 ( .C ( clk ), .D ( new_AGEMA_signal_18357 ), .Q ( new_AGEMA_signal_18358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6864 ( .C ( clk ), .D ( new_AGEMA_signal_18363 ), .Q ( new_AGEMA_signal_18364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6870 ( .C ( clk ), .D ( new_AGEMA_signal_18369 ), .Q ( new_AGEMA_signal_18370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6876 ( .C ( clk ), .D ( new_AGEMA_signal_18375 ), .Q ( new_AGEMA_signal_18376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6882 ( .C ( clk ), .D ( new_AGEMA_signal_18381 ), .Q ( new_AGEMA_signal_18382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6888 ( .C ( clk ), .D ( new_AGEMA_signal_18387 ), .Q ( new_AGEMA_signal_18388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6894 ( .C ( clk ), .D ( new_AGEMA_signal_18393 ), .Q ( new_AGEMA_signal_18394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6910 ( .C ( clk ), .D ( new_AGEMA_signal_18409 ), .Q ( new_AGEMA_signal_18410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6926 ( .C ( clk ), .D ( new_AGEMA_signal_18425 ), .Q ( new_AGEMA_signal_18426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6942 ( .C ( clk ), .D ( new_AGEMA_signal_18441 ), .Q ( new_AGEMA_signal_18442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6958 ( .C ( clk ), .D ( new_AGEMA_signal_18457 ), .Q ( new_AGEMA_signal_18458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6968 ( .C ( clk ), .D ( new_AGEMA_signal_18467 ), .Q ( new_AGEMA_signal_18468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6978 ( .C ( clk ), .D ( new_AGEMA_signal_18477 ), .Q ( new_AGEMA_signal_18478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6988 ( .C ( clk ), .D ( new_AGEMA_signal_18487 ), .Q ( new_AGEMA_signal_18488 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6998 ( .C ( clk ), .D ( new_AGEMA_signal_18497 ), .Q ( new_AGEMA_signal_18498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7016 ( .C ( clk ), .D ( new_AGEMA_signal_18515 ), .Q ( new_AGEMA_signal_18516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7034 ( .C ( clk ), .D ( new_AGEMA_signal_18533 ), .Q ( new_AGEMA_signal_18534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7052 ( .C ( clk ), .D ( new_AGEMA_signal_18551 ), .Q ( new_AGEMA_signal_18552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7070 ( .C ( clk ), .D ( new_AGEMA_signal_18569 ), .Q ( new_AGEMA_signal_18570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7074 ( .C ( clk ), .D ( new_AGEMA_signal_18573 ), .Q ( new_AGEMA_signal_18574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7078 ( .C ( clk ), .D ( new_AGEMA_signal_18577 ), .Q ( new_AGEMA_signal_18578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7082 ( .C ( clk ), .D ( new_AGEMA_signal_18581 ), .Q ( new_AGEMA_signal_18582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7086 ( .C ( clk ), .D ( new_AGEMA_signal_18585 ), .Q ( new_AGEMA_signal_18586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7094 ( .C ( clk ), .D ( new_AGEMA_signal_18593 ), .Q ( new_AGEMA_signal_18594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7102 ( .C ( clk ), .D ( new_AGEMA_signal_18601 ), .Q ( new_AGEMA_signal_18602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7110 ( .C ( clk ), .D ( new_AGEMA_signal_18609 ), .Q ( new_AGEMA_signal_18610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7118 ( .C ( clk ), .D ( new_AGEMA_signal_18617 ), .Q ( new_AGEMA_signal_18618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7122 ( .C ( clk ), .D ( new_AGEMA_signal_18621 ), .Q ( new_AGEMA_signal_18622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7126 ( .C ( clk ), .D ( new_AGEMA_signal_18625 ), .Q ( new_AGEMA_signal_18626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7130 ( .C ( clk ), .D ( new_AGEMA_signal_18629 ), .Q ( new_AGEMA_signal_18630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7134 ( .C ( clk ), .D ( new_AGEMA_signal_18633 ), .Q ( new_AGEMA_signal_18634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7140 ( .C ( clk ), .D ( new_AGEMA_signal_18639 ), .Q ( new_AGEMA_signal_18640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7148 ( .C ( clk ), .D ( new_AGEMA_signal_18647 ), .Q ( new_AGEMA_signal_18648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7156 ( .C ( clk ), .D ( new_AGEMA_signal_18655 ), .Q ( new_AGEMA_signal_18656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7164 ( .C ( clk ), .D ( new_AGEMA_signal_18663 ), .Q ( new_AGEMA_signal_18664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7170 ( .C ( clk ), .D ( new_AGEMA_signal_18669 ), .Q ( new_AGEMA_signal_18670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7176 ( .C ( clk ), .D ( new_AGEMA_signal_18675 ), .Q ( new_AGEMA_signal_18676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7182 ( .C ( clk ), .D ( new_AGEMA_signal_18681 ), .Q ( new_AGEMA_signal_18682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7188 ( .C ( clk ), .D ( new_AGEMA_signal_18687 ), .Q ( new_AGEMA_signal_18688 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7216 ( .C ( clk ), .D ( new_AGEMA_signal_18715 ), .Q ( new_AGEMA_signal_18716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7236 ( .C ( clk ), .D ( new_AGEMA_signal_18735 ), .Q ( new_AGEMA_signal_18736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7256 ( .C ( clk ), .D ( new_AGEMA_signal_18755 ), .Q ( new_AGEMA_signal_18756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7276 ( .C ( clk ), .D ( new_AGEMA_signal_18775 ), .Q ( new_AGEMA_signal_18776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7282 ( .C ( clk ), .D ( new_AGEMA_signal_18781 ), .Q ( new_AGEMA_signal_18782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7290 ( .C ( clk ), .D ( new_AGEMA_signal_18789 ), .Q ( new_AGEMA_signal_18790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7298 ( .C ( clk ), .D ( new_AGEMA_signal_18797 ), .Q ( new_AGEMA_signal_18798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7306 ( .C ( clk ), .D ( new_AGEMA_signal_18805 ), .Q ( new_AGEMA_signal_18806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7318 ( .C ( clk ), .D ( new_AGEMA_signal_18817 ), .Q ( new_AGEMA_signal_18818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7330 ( .C ( clk ), .D ( new_AGEMA_signal_18829 ), .Q ( new_AGEMA_signal_18830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7342 ( .C ( clk ), .D ( new_AGEMA_signal_18841 ), .Q ( new_AGEMA_signal_18842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7354 ( .C ( clk ), .D ( new_AGEMA_signal_18853 ), .Q ( new_AGEMA_signal_18854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7366 ( .C ( clk ), .D ( new_AGEMA_signal_18865 ), .Q ( new_AGEMA_signal_18866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7380 ( .C ( clk ), .D ( new_AGEMA_signal_18879 ), .Q ( new_AGEMA_signal_18880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7394 ( .C ( clk ), .D ( new_AGEMA_signal_18893 ), .Q ( new_AGEMA_signal_18894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7408 ( .C ( clk ), .D ( new_AGEMA_signal_18907 ), .Q ( new_AGEMA_signal_18908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7420 ( .C ( clk ), .D ( new_AGEMA_signal_18919 ), .Q ( new_AGEMA_signal_18920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7434 ( .C ( clk ), .D ( new_AGEMA_signal_18933 ), .Q ( new_AGEMA_signal_18934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7448 ( .C ( clk ), .D ( new_AGEMA_signal_18947 ), .Q ( new_AGEMA_signal_18948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7462 ( .C ( clk ), .D ( new_AGEMA_signal_18961 ), .Q ( new_AGEMA_signal_18962 ) ) ;

    /* cells in depth 25 */
    buf_clk new_AGEMA_reg_buffer_7141 ( .C ( clk ), .D ( new_AGEMA_signal_18640 ), .Q ( new_AGEMA_signal_18641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7149 ( .C ( clk ), .D ( new_AGEMA_signal_18648 ), .Q ( new_AGEMA_signal_18649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7157 ( .C ( clk ), .D ( new_AGEMA_signal_18656 ), .Q ( new_AGEMA_signal_18657 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7165 ( .C ( clk ), .D ( new_AGEMA_signal_18664 ), .Q ( new_AGEMA_signal_18665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7171 ( .C ( clk ), .D ( new_AGEMA_signal_18670 ), .Q ( new_AGEMA_signal_18671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7177 ( .C ( clk ), .D ( new_AGEMA_signal_18676 ), .Q ( new_AGEMA_signal_18677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7183 ( .C ( clk ), .D ( new_AGEMA_signal_18682 ), .Q ( new_AGEMA_signal_18683 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7189 ( .C ( clk ), .D ( new_AGEMA_signal_18688 ), .Q ( new_AGEMA_signal_18689 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7191 ( .C ( clk ), .D ( n2209 ), .Q ( new_AGEMA_signal_18691 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7193 ( .C ( clk ), .D ( new_AGEMA_signal_3660 ), .Q ( new_AGEMA_signal_18693 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7195 ( .C ( clk ), .D ( new_AGEMA_signal_3661 ), .Q ( new_AGEMA_signal_18695 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7197 ( .C ( clk ), .D ( new_AGEMA_signal_3662 ), .Q ( new_AGEMA_signal_18697 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7217 ( .C ( clk ), .D ( new_AGEMA_signal_18716 ), .Q ( new_AGEMA_signal_18717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7237 ( .C ( clk ), .D ( new_AGEMA_signal_18736 ), .Q ( new_AGEMA_signal_18737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7257 ( .C ( clk ), .D ( new_AGEMA_signal_18756 ), .Q ( new_AGEMA_signal_18757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7277 ( .C ( clk ), .D ( new_AGEMA_signal_18776 ), .Q ( new_AGEMA_signal_18777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7283 ( .C ( clk ), .D ( new_AGEMA_signal_18782 ), .Q ( new_AGEMA_signal_18783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7291 ( .C ( clk ), .D ( new_AGEMA_signal_18790 ), .Q ( new_AGEMA_signal_18791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7299 ( .C ( clk ), .D ( new_AGEMA_signal_18798 ), .Q ( new_AGEMA_signal_18799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7307 ( .C ( clk ), .D ( new_AGEMA_signal_18806 ), .Q ( new_AGEMA_signal_18807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7319 ( .C ( clk ), .D ( new_AGEMA_signal_18818 ), .Q ( new_AGEMA_signal_18819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7331 ( .C ( clk ), .D ( new_AGEMA_signal_18830 ), .Q ( new_AGEMA_signal_18831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7343 ( .C ( clk ), .D ( new_AGEMA_signal_18842 ), .Q ( new_AGEMA_signal_18843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7355 ( .C ( clk ), .D ( new_AGEMA_signal_18854 ), .Q ( new_AGEMA_signal_18855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7367 ( .C ( clk ), .D ( new_AGEMA_signal_18866 ), .Q ( new_AGEMA_signal_18867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7381 ( .C ( clk ), .D ( new_AGEMA_signal_18880 ), .Q ( new_AGEMA_signal_18881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7395 ( .C ( clk ), .D ( new_AGEMA_signal_18894 ), .Q ( new_AGEMA_signal_18895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7409 ( .C ( clk ), .D ( new_AGEMA_signal_18908 ), .Q ( new_AGEMA_signal_18909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7421 ( .C ( clk ), .D ( new_AGEMA_signal_18920 ), .Q ( new_AGEMA_signal_18921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7435 ( .C ( clk ), .D ( new_AGEMA_signal_18934 ), .Q ( new_AGEMA_signal_18935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7449 ( .C ( clk ), .D ( new_AGEMA_signal_18948 ), .Q ( new_AGEMA_signal_18949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7463 ( .C ( clk ), .D ( new_AGEMA_signal_18962 ), .Q ( new_AGEMA_signal_18963 ) ) ;

    /* cells in depth 26 */
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2155 ( .ina ({new_AGEMA_signal_3653, new_AGEMA_signal_3652, new_AGEMA_signal_3651, n2017}), .inb ({new_AGEMA_signal_18370, new_AGEMA_signal_18364, new_AGEMA_signal_18358, new_AGEMA_signal_18352}), .clk ( clk ), .rnd ({Fresh[8529], Fresh[8528], Fresh[8527], Fresh[8526], Fresh[8525], Fresh[8524], Fresh[8523], Fresh[8522], Fresh[8521], Fresh[8520]}), .outt ({new_AGEMA_signal_3680, new_AGEMA_signal_3679, new_AGEMA_signal_3678, n2018}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2269 ( .ina ({new_AGEMA_signal_18394, new_AGEMA_signal_18388, new_AGEMA_signal_18382, new_AGEMA_signal_18376}), .inb ({new_AGEMA_signal_3656, new_AGEMA_signal_3655, new_AGEMA_signal_3654, n2110}), .clk ( clk ), .rnd ({Fresh[8539], Fresh[8538], Fresh[8537], Fresh[8536], Fresh[8535], Fresh[8534], Fresh[8533], Fresh[8532], Fresh[8531], Fresh[8530]}), .outt ({new_AGEMA_signal_3683, new_AGEMA_signal_3682, new_AGEMA_signal_3681, n2112}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2320 ( .ina ({new_AGEMA_signal_18458, new_AGEMA_signal_18442, new_AGEMA_signal_18426, new_AGEMA_signal_18410}), .inb ({new_AGEMA_signal_3659, new_AGEMA_signal_3658, new_AGEMA_signal_3657, n2154}), .clk ( clk ), .rnd ({Fresh[8549], Fresh[8548], Fresh[8547], Fresh[8546], Fresh[8545], Fresh[8544], Fresh[8543], Fresh[8542], Fresh[8541], Fresh[8540]}), .outt ({new_AGEMA_signal_3686, new_AGEMA_signal_3685, new_AGEMA_signal_3684, n2210}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2479 ( .ina ({new_AGEMA_signal_18498, new_AGEMA_signal_18488, new_AGEMA_signal_18478, new_AGEMA_signal_18468}), .inb ({new_AGEMA_signal_3665, new_AGEMA_signal_3664, new_AGEMA_signal_3663, n2311}), .clk ( clk ), .rnd ({Fresh[8559], Fresh[8558], Fresh[8557], Fresh[8556], Fresh[8555], Fresh[8554], Fresh[8553], Fresh[8552], Fresh[8551], Fresh[8550]}), .outt ({new_AGEMA_signal_3689, new_AGEMA_signal_3688, new_AGEMA_signal_3687, N470}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2538 ( .ina ({new_AGEMA_signal_18570, new_AGEMA_signal_18552, new_AGEMA_signal_18534, new_AGEMA_signal_18516}), .inb ({new_AGEMA_signal_3668, new_AGEMA_signal_3667, new_AGEMA_signal_3666, n2374}), .clk ( clk ), .rnd ({Fresh[8569], Fresh[8568], Fresh[8567], Fresh[8566], Fresh[8565], Fresh[8564], Fresh[8563], Fresh[8562], Fresh[8561], Fresh[8560]}), .outt ({new_AGEMA_signal_3692, new_AGEMA_signal_3691, new_AGEMA_signal_3690, n2378}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2673 ( .ina ({new_AGEMA_signal_18586, new_AGEMA_signal_18582, new_AGEMA_signal_18578, new_AGEMA_signal_18574}), .inb ({new_AGEMA_signal_3671, new_AGEMA_signal_3670, new_AGEMA_signal_3669, n2529}), .clk ( clk ), .rnd ({Fresh[8579], Fresh[8578], Fresh[8577], Fresh[8576], Fresh[8575], Fresh[8574], Fresh[8573], Fresh[8572], Fresh[8571], Fresh[8570]}), .outt ({new_AGEMA_signal_3695, new_AGEMA_signal_3694, new_AGEMA_signal_3693, N639}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2769 ( .ina ({new_AGEMA_signal_18618, new_AGEMA_signal_18610, new_AGEMA_signal_18602, new_AGEMA_signal_18594}), .inb ({new_AGEMA_signal_3674, new_AGEMA_signal_3673, new_AGEMA_signal_3672, n2670}), .clk ( clk ), .rnd ({Fresh[8589], Fresh[8588], Fresh[8587], Fresh[8586], Fresh[8585], Fresh[8584], Fresh[8583], Fresh[8582], Fresh[8581], Fresh[8580]}), .outt ({new_AGEMA_signal_3698, new_AGEMA_signal_3697, new_AGEMA_signal_3696, N723}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2855 ( .ina ({new_AGEMA_signal_18634, new_AGEMA_signal_18630, new_AGEMA_signal_18626, new_AGEMA_signal_18622}), .inb ({new_AGEMA_signal_3650, new_AGEMA_signal_3649, new_AGEMA_signal_3648, n2831}), .clk ( clk ), .rnd ({Fresh[8599], Fresh[8598], Fresh[8597], Fresh[8596], Fresh[8595], Fresh[8594], Fresh[8593], Fresh[8592], Fresh[8591], Fresh[8590]}), .outt ({new_AGEMA_signal_3677, new_AGEMA_signal_3676, new_AGEMA_signal_3675, N789}) ) ;
    buf_clk new_AGEMA_reg_buffer_7142 ( .C ( clk ), .D ( new_AGEMA_signal_18641 ), .Q ( new_AGEMA_signal_18642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7150 ( .C ( clk ), .D ( new_AGEMA_signal_18649 ), .Q ( new_AGEMA_signal_18650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7158 ( .C ( clk ), .D ( new_AGEMA_signal_18657 ), .Q ( new_AGEMA_signal_18658 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7166 ( .C ( clk ), .D ( new_AGEMA_signal_18665 ), .Q ( new_AGEMA_signal_18666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7172 ( .C ( clk ), .D ( new_AGEMA_signal_18671 ), .Q ( new_AGEMA_signal_18672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7178 ( .C ( clk ), .D ( new_AGEMA_signal_18677 ), .Q ( new_AGEMA_signal_18678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7184 ( .C ( clk ), .D ( new_AGEMA_signal_18683 ), .Q ( new_AGEMA_signal_18684 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7190 ( .C ( clk ), .D ( new_AGEMA_signal_18689 ), .Q ( new_AGEMA_signal_18690 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7192 ( .C ( clk ), .D ( new_AGEMA_signal_18691 ), .Q ( new_AGEMA_signal_18692 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7194 ( .C ( clk ), .D ( new_AGEMA_signal_18693 ), .Q ( new_AGEMA_signal_18694 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7196 ( .C ( clk ), .D ( new_AGEMA_signal_18695 ), .Q ( new_AGEMA_signal_18696 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7198 ( .C ( clk ), .D ( new_AGEMA_signal_18697 ), .Q ( new_AGEMA_signal_18698 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7218 ( .C ( clk ), .D ( new_AGEMA_signal_18717 ), .Q ( new_AGEMA_signal_18718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7238 ( .C ( clk ), .D ( new_AGEMA_signal_18737 ), .Q ( new_AGEMA_signal_18738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7258 ( .C ( clk ), .D ( new_AGEMA_signal_18757 ), .Q ( new_AGEMA_signal_18758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7278 ( .C ( clk ), .D ( new_AGEMA_signal_18777 ), .Q ( new_AGEMA_signal_18778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7284 ( .C ( clk ), .D ( new_AGEMA_signal_18783 ), .Q ( new_AGEMA_signal_18784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7292 ( .C ( clk ), .D ( new_AGEMA_signal_18791 ), .Q ( new_AGEMA_signal_18792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7300 ( .C ( clk ), .D ( new_AGEMA_signal_18799 ), .Q ( new_AGEMA_signal_18800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7308 ( .C ( clk ), .D ( new_AGEMA_signal_18807 ), .Q ( new_AGEMA_signal_18808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7320 ( .C ( clk ), .D ( new_AGEMA_signal_18819 ), .Q ( new_AGEMA_signal_18820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7332 ( .C ( clk ), .D ( new_AGEMA_signal_18831 ), .Q ( new_AGEMA_signal_18832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7344 ( .C ( clk ), .D ( new_AGEMA_signal_18843 ), .Q ( new_AGEMA_signal_18844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7356 ( .C ( clk ), .D ( new_AGEMA_signal_18855 ), .Q ( new_AGEMA_signal_18856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7368 ( .C ( clk ), .D ( new_AGEMA_signal_18867 ), .Q ( new_AGEMA_signal_18868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7382 ( .C ( clk ), .D ( new_AGEMA_signal_18881 ), .Q ( new_AGEMA_signal_18882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7396 ( .C ( clk ), .D ( new_AGEMA_signal_18895 ), .Q ( new_AGEMA_signal_18896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7410 ( .C ( clk ), .D ( new_AGEMA_signal_18909 ), .Q ( new_AGEMA_signal_18910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7422 ( .C ( clk ), .D ( new_AGEMA_signal_18921 ), .Q ( new_AGEMA_signal_18922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7436 ( .C ( clk ), .D ( new_AGEMA_signal_18935 ), .Q ( new_AGEMA_signal_18936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7450 ( .C ( clk ), .D ( new_AGEMA_signal_18949 ), .Q ( new_AGEMA_signal_18950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7464 ( .C ( clk ), .D ( new_AGEMA_signal_18963 ), .Q ( new_AGEMA_signal_18964 ) ) ;

    /* cells in depth 27 */
    buf_clk new_AGEMA_reg_buffer_7285 ( .C ( clk ), .D ( new_AGEMA_signal_18784 ), .Q ( new_AGEMA_signal_18785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7293 ( .C ( clk ), .D ( new_AGEMA_signal_18792 ), .Q ( new_AGEMA_signal_18793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7301 ( .C ( clk ), .D ( new_AGEMA_signal_18800 ), .Q ( new_AGEMA_signal_18801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7309 ( .C ( clk ), .D ( new_AGEMA_signal_18808 ), .Q ( new_AGEMA_signal_18809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7321 ( .C ( clk ), .D ( new_AGEMA_signal_18820 ), .Q ( new_AGEMA_signal_18821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7333 ( .C ( clk ), .D ( new_AGEMA_signal_18832 ), .Q ( new_AGEMA_signal_18833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7345 ( .C ( clk ), .D ( new_AGEMA_signal_18844 ), .Q ( new_AGEMA_signal_18845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7357 ( .C ( clk ), .D ( new_AGEMA_signal_18856 ), .Q ( new_AGEMA_signal_18857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7369 ( .C ( clk ), .D ( new_AGEMA_signal_18868 ), .Q ( new_AGEMA_signal_18869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7383 ( .C ( clk ), .D ( new_AGEMA_signal_18882 ), .Q ( new_AGEMA_signal_18883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7397 ( .C ( clk ), .D ( new_AGEMA_signal_18896 ), .Q ( new_AGEMA_signal_18897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7411 ( .C ( clk ), .D ( new_AGEMA_signal_18910 ), .Q ( new_AGEMA_signal_18911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7423 ( .C ( clk ), .D ( new_AGEMA_signal_18922 ), .Q ( new_AGEMA_signal_18923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7437 ( .C ( clk ), .D ( new_AGEMA_signal_18936 ), .Q ( new_AGEMA_signal_18937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7451 ( .C ( clk ), .D ( new_AGEMA_signal_18950 ), .Q ( new_AGEMA_signal_18951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7465 ( .C ( clk ), .D ( new_AGEMA_signal_18964 ), .Q ( new_AGEMA_signal_18965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7535 ( .C ( clk ), .D ( N470 ), .Q ( new_AGEMA_signal_19035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7543 ( .C ( clk ), .D ( new_AGEMA_signal_3687 ), .Q ( new_AGEMA_signal_19043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7551 ( .C ( clk ), .D ( new_AGEMA_signal_3688 ), .Q ( new_AGEMA_signal_19051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7559 ( .C ( clk ), .D ( new_AGEMA_signal_3689 ), .Q ( new_AGEMA_signal_19059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7567 ( .C ( clk ), .D ( N639 ), .Q ( new_AGEMA_signal_19067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7575 ( .C ( clk ), .D ( new_AGEMA_signal_3693 ), .Q ( new_AGEMA_signal_19075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7583 ( .C ( clk ), .D ( new_AGEMA_signal_3694 ), .Q ( new_AGEMA_signal_19083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7591 ( .C ( clk ), .D ( new_AGEMA_signal_3695 ), .Q ( new_AGEMA_signal_19091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7599 ( .C ( clk ), .D ( N723 ), .Q ( new_AGEMA_signal_19099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7607 ( .C ( clk ), .D ( new_AGEMA_signal_3696 ), .Q ( new_AGEMA_signal_19107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7615 ( .C ( clk ), .D ( new_AGEMA_signal_3697 ), .Q ( new_AGEMA_signal_19115 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7623 ( .C ( clk ), .D ( new_AGEMA_signal_3698 ), .Q ( new_AGEMA_signal_19123 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7631 ( .C ( clk ), .D ( N789 ), .Q ( new_AGEMA_signal_19131 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7639 ( .C ( clk ), .D ( new_AGEMA_signal_3675 ), .Q ( new_AGEMA_signal_19139 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7647 ( .C ( clk ), .D ( new_AGEMA_signal_3676 ), .Q ( new_AGEMA_signal_19147 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7655 ( .C ( clk ), .D ( new_AGEMA_signal_3677 ), .Q ( new_AGEMA_signal_19155 ) ) ;

    /* cells in depth 28 */
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2156 ( .ina ({new_AGEMA_signal_18666, new_AGEMA_signal_18658, new_AGEMA_signal_18650, new_AGEMA_signal_18642}), .inb ({new_AGEMA_signal_3680, new_AGEMA_signal_3679, new_AGEMA_signal_3678, n2018}), .clk ( clk ), .rnd ({Fresh[8609], Fresh[8608], Fresh[8607], Fresh[8606], Fresh[8605], Fresh[8604], Fresh[8603], Fresh[8602], Fresh[8601], Fresh[8600]}), .outt ({new_AGEMA_signal_3701, new_AGEMA_signal_3700, new_AGEMA_signal_3699, N169}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2270 ( .ina ({new_AGEMA_signal_18690, new_AGEMA_signal_18684, new_AGEMA_signal_18678, new_AGEMA_signal_18672}), .inb ({new_AGEMA_signal_3683, new_AGEMA_signal_3682, new_AGEMA_signal_3681, n2112}), .clk ( clk ), .rnd ({Fresh[8619], Fresh[8618], Fresh[8617], Fresh[8616], Fresh[8615], Fresh[8614], Fresh[8613], Fresh[8612], Fresh[8611], Fresh[8610]}), .outt ({new_AGEMA_signal_3704, new_AGEMA_signal_3703, new_AGEMA_signal_3702, N277}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2376 ( .ina ({new_AGEMA_signal_3686, new_AGEMA_signal_3685, new_AGEMA_signal_3684, n2210}), .inb ({new_AGEMA_signal_18698, new_AGEMA_signal_18696, new_AGEMA_signal_18694, new_AGEMA_signal_18692}), .clk ( clk ), .rnd ({Fresh[8629], Fresh[8628], Fresh[8627], Fresh[8626], Fresh[8625], Fresh[8624], Fresh[8623], Fresh[8622], Fresh[8621], Fresh[8620]}), .outt ({new_AGEMA_signal_3707, new_AGEMA_signal_3706, new_AGEMA_signal_3705, n2211}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2540 ( .ina ({new_AGEMA_signal_3692, new_AGEMA_signal_3691, new_AGEMA_signal_3690, n2378}), .inb ({new_AGEMA_signal_18778, new_AGEMA_signal_18758, new_AGEMA_signal_18738, new_AGEMA_signal_18718}), .clk ( clk ), .rnd ({Fresh[8639], Fresh[8638], Fresh[8637], Fresh[8636], Fresh[8635], Fresh[8634], Fresh[8633], Fresh[8632], Fresh[8631], Fresh[8630]}), .outt ({new_AGEMA_signal_3710, new_AGEMA_signal_3709, new_AGEMA_signal_3708, n2379}) ) ;
    buf_clk new_AGEMA_reg_buffer_7286 ( .C ( clk ), .D ( new_AGEMA_signal_18785 ), .Q ( new_AGEMA_signal_18786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7294 ( .C ( clk ), .D ( new_AGEMA_signal_18793 ), .Q ( new_AGEMA_signal_18794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7302 ( .C ( clk ), .D ( new_AGEMA_signal_18801 ), .Q ( new_AGEMA_signal_18802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7310 ( .C ( clk ), .D ( new_AGEMA_signal_18809 ), .Q ( new_AGEMA_signal_18810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7322 ( .C ( clk ), .D ( new_AGEMA_signal_18821 ), .Q ( new_AGEMA_signal_18822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7334 ( .C ( clk ), .D ( new_AGEMA_signal_18833 ), .Q ( new_AGEMA_signal_18834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7346 ( .C ( clk ), .D ( new_AGEMA_signal_18845 ), .Q ( new_AGEMA_signal_18846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7358 ( .C ( clk ), .D ( new_AGEMA_signal_18857 ), .Q ( new_AGEMA_signal_18858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7370 ( .C ( clk ), .D ( new_AGEMA_signal_18869 ), .Q ( new_AGEMA_signal_18870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7384 ( .C ( clk ), .D ( new_AGEMA_signal_18883 ), .Q ( new_AGEMA_signal_18884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7398 ( .C ( clk ), .D ( new_AGEMA_signal_18897 ), .Q ( new_AGEMA_signal_18898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7412 ( .C ( clk ), .D ( new_AGEMA_signal_18911 ), .Q ( new_AGEMA_signal_18912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7424 ( .C ( clk ), .D ( new_AGEMA_signal_18923 ), .Q ( new_AGEMA_signal_18924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7438 ( .C ( clk ), .D ( new_AGEMA_signal_18937 ), .Q ( new_AGEMA_signal_18938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7452 ( .C ( clk ), .D ( new_AGEMA_signal_18951 ), .Q ( new_AGEMA_signal_18952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7466 ( .C ( clk ), .D ( new_AGEMA_signal_18965 ), .Q ( new_AGEMA_signal_18966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7536 ( .C ( clk ), .D ( new_AGEMA_signal_19035 ), .Q ( new_AGEMA_signal_19036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7544 ( .C ( clk ), .D ( new_AGEMA_signal_19043 ), .Q ( new_AGEMA_signal_19044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7552 ( .C ( clk ), .D ( new_AGEMA_signal_19051 ), .Q ( new_AGEMA_signal_19052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7560 ( .C ( clk ), .D ( new_AGEMA_signal_19059 ), .Q ( new_AGEMA_signal_19060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7568 ( .C ( clk ), .D ( new_AGEMA_signal_19067 ), .Q ( new_AGEMA_signal_19068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7576 ( .C ( clk ), .D ( new_AGEMA_signal_19075 ), .Q ( new_AGEMA_signal_19076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7584 ( .C ( clk ), .D ( new_AGEMA_signal_19083 ), .Q ( new_AGEMA_signal_19084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7592 ( .C ( clk ), .D ( new_AGEMA_signal_19091 ), .Q ( new_AGEMA_signal_19092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7600 ( .C ( clk ), .D ( new_AGEMA_signal_19099 ), .Q ( new_AGEMA_signal_19100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7608 ( .C ( clk ), .D ( new_AGEMA_signal_19107 ), .Q ( new_AGEMA_signal_19108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7616 ( .C ( clk ), .D ( new_AGEMA_signal_19115 ), .Q ( new_AGEMA_signal_19116 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7624 ( .C ( clk ), .D ( new_AGEMA_signal_19123 ), .Q ( new_AGEMA_signal_19124 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7632 ( .C ( clk ), .D ( new_AGEMA_signal_19131 ), .Q ( new_AGEMA_signal_19132 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7640 ( .C ( clk ), .D ( new_AGEMA_signal_19139 ), .Q ( new_AGEMA_signal_19140 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7648 ( .C ( clk ), .D ( new_AGEMA_signal_19147 ), .Q ( new_AGEMA_signal_19148 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7656 ( .C ( clk ), .D ( new_AGEMA_signal_19155 ), .Q ( new_AGEMA_signal_19156 ) ) ;

    /* cells in depth 29 */
    buf_clk new_AGEMA_reg_buffer_7371 ( .C ( clk ), .D ( new_AGEMA_signal_18870 ), .Q ( new_AGEMA_signal_18871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7385 ( .C ( clk ), .D ( new_AGEMA_signal_18884 ), .Q ( new_AGEMA_signal_18885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7399 ( .C ( clk ), .D ( new_AGEMA_signal_18898 ), .Q ( new_AGEMA_signal_18899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7413 ( .C ( clk ), .D ( new_AGEMA_signal_18912 ), .Q ( new_AGEMA_signal_18913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7425 ( .C ( clk ), .D ( new_AGEMA_signal_18924 ), .Q ( new_AGEMA_signal_18925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7439 ( .C ( clk ), .D ( new_AGEMA_signal_18938 ), .Q ( new_AGEMA_signal_18939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7453 ( .C ( clk ), .D ( new_AGEMA_signal_18952 ), .Q ( new_AGEMA_signal_18953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7467 ( .C ( clk ), .D ( new_AGEMA_signal_18966 ), .Q ( new_AGEMA_signal_18967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7471 ( .C ( clk ), .D ( N169 ), .Q ( new_AGEMA_signal_18971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7477 ( .C ( clk ), .D ( new_AGEMA_signal_3699 ), .Q ( new_AGEMA_signal_18977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7483 ( .C ( clk ), .D ( new_AGEMA_signal_3700 ), .Q ( new_AGEMA_signal_18983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7489 ( .C ( clk ), .D ( new_AGEMA_signal_3701 ), .Q ( new_AGEMA_signal_18989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7495 ( .C ( clk ), .D ( N277 ), .Q ( new_AGEMA_signal_18995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7501 ( .C ( clk ), .D ( new_AGEMA_signal_3702 ), .Q ( new_AGEMA_signal_19001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7507 ( .C ( clk ), .D ( new_AGEMA_signal_3703 ), .Q ( new_AGEMA_signal_19007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7513 ( .C ( clk ), .D ( new_AGEMA_signal_3704 ), .Q ( new_AGEMA_signal_19013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7537 ( .C ( clk ), .D ( new_AGEMA_signal_19036 ), .Q ( new_AGEMA_signal_19037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7545 ( .C ( clk ), .D ( new_AGEMA_signal_19044 ), .Q ( new_AGEMA_signal_19045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7553 ( .C ( clk ), .D ( new_AGEMA_signal_19052 ), .Q ( new_AGEMA_signal_19053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7561 ( .C ( clk ), .D ( new_AGEMA_signal_19060 ), .Q ( new_AGEMA_signal_19061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7569 ( .C ( clk ), .D ( new_AGEMA_signal_19068 ), .Q ( new_AGEMA_signal_19069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7577 ( .C ( clk ), .D ( new_AGEMA_signal_19076 ), .Q ( new_AGEMA_signal_19077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7585 ( .C ( clk ), .D ( new_AGEMA_signal_19084 ), .Q ( new_AGEMA_signal_19085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7593 ( .C ( clk ), .D ( new_AGEMA_signal_19092 ), .Q ( new_AGEMA_signal_19093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7601 ( .C ( clk ), .D ( new_AGEMA_signal_19100 ), .Q ( new_AGEMA_signal_19101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7609 ( .C ( clk ), .D ( new_AGEMA_signal_19108 ), .Q ( new_AGEMA_signal_19109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7617 ( .C ( clk ), .D ( new_AGEMA_signal_19116 ), .Q ( new_AGEMA_signal_19117 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7625 ( .C ( clk ), .D ( new_AGEMA_signal_19124 ), .Q ( new_AGEMA_signal_19125 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7633 ( .C ( clk ), .D ( new_AGEMA_signal_19132 ), .Q ( new_AGEMA_signal_19133 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7641 ( .C ( clk ), .D ( new_AGEMA_signal_19140 ), .Q ( new_AGEMA_signal_19141 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7649 ( .C ( clk ), .D ( new_AGEMA_signal_19148 ), .Q ( new_AGEMA_signal_19149 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7657 ( .C ( clk ), .D ( new_AGEMA_signal_19156 ), .Q ( new_AGEMA_signal_19157 ) ) ;

    /* cells in depth 30 */
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2377 ( .ina ({new_AGEMA_signal_18810, new_AGEMA_signal_18802, new_AGEMA_signal_18794, new_AGEMA_signal_18786}), .inb ({new_AGEMA_signal_3707, new_AGEMA_signal_3706, new_AGEMA_signal_3705, n2211}), .clk ( clk ), .rnd ({Fresh[8649], Fresh[8648], Fresh[8647], Fresh[8646], Fresh[8645], Fresh[8644], Fresh[8643], Fresh[8642], Fresh[8641], Fresh[8640]}), .outt ({new_AGEMA_signal_3713, new_AGEMA_signal_3712, new_AGEMA_signal_3711, N379}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2541 ( .ina ({new_AGEMA_signal_18858, new_AGEMA_signal_18846, new_AGEMA_signal_18834, new_AGEMA_signal_18822}), .inb ({new_AGEMA_signal_3710, new_AGEMA_signal_3709, new_AGEMA_signal_3708, n2379}), .clk ( clk ), .rnd ({Fresh[8659], Fresh[8658], Fresh[8657], Fresh[8656], Fresh[8655], Fresh[8654], Fresh[8653], Fresh[8652], Fresh[8651], Fresh[8650]}), .outt ({new_AGEMA_signal_3716, new_AGEMA_signal_3715, new_AGEMA_signal_3714, n2381}) ) ;
    buf_clk new_AGEMA_reg_buffer_7372 ( .C ( clk ), .D ( new_AGEMA_signal_18871 ), .Q ( new_AGEMA_signal_18872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7386 ( .C ( clk ), .D ( new_AGEMA_signal_18885 ), .Q ( new_AGEMA_signal_18886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7400 ( .C ( clk ), .D ( new_AGEMA_signal_18899 ), .Q ( new_AGEMA_signal_18900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7414 ( .C ( clk ), .D ( new_AGEMA_signal_18913 ), .Q ( new_AGEMA_signal_18914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7426 ( .C ( clk ), .D ( new_AGEMA_signal_18925 ), .Q ( new_AGEMA_signal_18926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7440 ( .C ( clk ), .D ( new_AGEMA_signal_18939 ), .Q ( new_AGEMA_signal_18940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7454 ( .C ( clk ), .D ( new_AGEMA_signal_18953 ), .Q ( new_AGEMA_signal_18954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7468 ( .C ( clk ), .D ( new_AGEMA_signal_18967 ), .Q ( new_AGEMA_signal_18968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7472 ( .C ( clk ), .D ( new_AGEMA_signal_18971 ), .Q ( new_AGEMA_signal_18972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7478 ( .C ( clk ), .D ( new_AGEMA_signal_18977 ), .Q ( new_AGEMA_signal_18978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7484 ( .C ( clk ), .D ( new_AGEMA_signal_18983 ), .Q ( new_AGEMA_signal_18984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7490 ( .C ( clk ), .D ( new_AGEMA_signal_18989 ), .Q ( new_AGEMA_signal_18990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7496 ( .C ( clk ), .D ( new_AGEMA_signal_18995 ), .Q ( new_AGEMA_signal_18996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7502 ( .C ( clk ), .D ( new_AGEMA_signal_19001 ), .Q ( new_AGEMA_signal_19002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7508 ( .C ( clk ), .D ( new_AGEMA_signal_19007 ), .Q ( new_AGEMA_signal_19008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7514 ( .C ( clk ), .D ( new_AGEMA_signal_19013 ), .Q ( new_AGEMA_signal_19014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7538 ( .C ( clk ), .D ( new_AGEMA_signal_19037 ), .Q ( new_AGEMA_signal_19038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7546 ( .C ( clk ), .D ( new_AGEMA_signal_19045 ), .Q ( new_AGEMA_signal_19046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7554 ( .C ( clk ), .D ( new_AGEMA_signal_19053 ), .Q ( new_AGEMA_signal_19054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7562 ( .C ( clk ), .D ( new_AGEMA_signal_19061 ), .Q ( new_AGEMA_signal_19062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7570 ( .C ( clk ), .D ( new_AGEMA_signal_19069 ), .Q ( new_AGEMA_signal_19070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7578 ( .C ( clk ), .D ( new_AGEMA_signal_19077 ), .Q ( new_AGEMA_signal_19078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7586 ( .C ( clk ), .D ( new_AGEMA_signal_19085 ), .Q ( new_AGEMA_signal_19086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7594 ( .C ( clk ), .D ( new_AGEMA_signal_19093 ), .Q ( new_AGEMA_signal_19094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7602 ( .C ( clk ), .D ( new_AGEMA_signal_19101 ), .Q ( new_AGEMA_signal_19102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7610 ( .C ( clk ), .D ( new_AGEMA_signal_19109 ), .Q ( new_AGEMA_signal_19110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7618 ( .C ( clk ), .D ( new_AGEMA_signal_19117 ), .Q ( new_AGEMA_signal_19118 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7626 ( .C ( clk ), .D ( new_AGEMA_signal_19125 ), .Q ( new_AGEMA_signal_19126 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7634 ( .C ( clk ), .D ( new_AGEMA_signal_19133 ), .Q ( new_AGEMA_signal_19134 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7642 ( .C ( clk ), .D ( new_AGEMA_signal_19141 ), .Q ( new_AGEMA_signal_19142 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7650 ( .C ( clk ), .D ( new_AGEMA_signal_19149 ), .Q ( new_AGEMA_signal_19150 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7658 ( .C ( clk ), .D ( new_AGEMA_signal_19157 ), .Q ( new_AGEMA_signal_19158 ) ) ;

    /* cells in depth 31 */
    buf_clk new_AGEMA_reg_buffer_7427 ( .C ( clk ), .D ( new_AGEMA_signal_18926 ), .Q ( new_AGEMA_signal_18927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7441 ( .C ( clk ), .D ( new_AGEMA_signal_18940 ), .Q ( new_AGEMA_signal_18941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7455 ( .C ( clk ), .D ( new_AGEMA_signal_18954 ), .Q ( new_AGEMA_signal_18955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7469 ( .C ( clk ), .D ( new_AGEMA_signal_18968 ), .Q ( new_AGEMA_signal_18969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7473 ( .C ( clk ), .D ( new_AGEMA_signal_18972 ), .Q ( new_AGEMA_signal_18973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7479 ( .C ( clk ), .D ( new_AGEMA_signal_18978 ), .Q ( new_AGEMA_signal_18979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7485 ( .C ( clk ), .D ( new_AGEMA_signal_18984 ), .Q ( new_AGEMA_signal_18985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7491 ( .C ( clk ), .D ( new_AGEMA_signal_18990 ), .Q ( new_AGEMA_signal_18991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7497 ( .C ( clk ), .D ( new_AGEMA_signal_18996 ), .Q ( new_AGEMA_signal_18997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7503 ( .C ( clk ), .D ( new_AGEMA_signal_19002 ), .Q ( new_AGEMA_signal_19003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7509 ( .C ( clk ), .D ( new_AGEMA_signal_19008 ), .Q ( new_AGEMA_signal_19009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7515 ( .C ( clk ), .D ( new_AGEMA_signal_19014 ), .Q ( new_AGEMA_signal_19015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7519 ( .C ( clk ), .D ( N379 ), .Q ( new_AGEMA_signal_19019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7523 ( .C ( clk ), .D ( new_AGEMA_signal_3711 ), .Q ( new_AGEMA_signal_19023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7527 ( .C ( clk ), .D ( new_AGEMA_signal_3712 ), .Q ( new_AGEMA_signal_19027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7531 ( .C ( clk ), .D ( new_AGEMA_signal_3713 ), .Q ( new_AGEMA_signal_19031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7539 ( .C ( clk ), .D ( new_AGEMA_signal_19038 ), .Q ( new_AGEMA_signal_19039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7547 ( .C ( clk ), .D ( new_AGEMA_signal_19046 ), .Q ( new_AGEMA_signal_19047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7555 ( .C ( clk ), .D ( new_AGEMA_signal_19054 ), .Q ( new_AGEMA_signal_19055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7563 ( .C ( clk ), .D ( new_AGEMA_signal_19062 ), .Q ( new_AGEMA_signal_19063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7571 ( .C ( clk ), .D ( new_AGEMA_signal_19070 ), .Q ( new_AGEMA_signal_19071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7579 ( .C ( clk ), .D ( new_AGEMA_signal_19078 ), .Q ( new_AGEMA_signal_19079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7587 ( .C ( clk ), .D ( new_AGEMA_signal_19086 ), .Q ( new_AGEMA_signal_19087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7595 ( .C ( clk ), .D ( new_AGEMA_signal_19094 ), .Q ( new_AGEMA_signal_19095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7603 ( .C ( clk ), .D ( new_AGEMA_signal_19102 ), .Q ( new_AGEMA_signal_19103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7611 ( .C ( clk ), .D ( new_AGEMA_signal_19110 ), .Q ( new_AGEMA_signal_19111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7619 ( .C ( clk ), .D ( new_AGEMA_signal_19118 ), .Q ( new_AGEMA_signal_19119 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7627 ( .C ( clk ), .D ( new_AGEMA_signal_19126 ), .Q ( new_AGEMA_signal_19127 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7635 ( .C ( clk ), .D ( new_AGEMA_signal_19134 ), .Q ( new_AGEMA_signal_19135 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7643 ( .C ( clk ), .D ( new_AGEMA_signal_19142 ), .Q ( new_AGEMA_signal_19143 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7651 ( .C ( clk ), .D ( new_AGEMA_signal_19150 ), .Q ( new_AGEMA_signal_19151 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7659 ( .C ( clk ), .D ( new_AGEMA_signal_19158 ), .Q ( new_AGEMA_signal_19159 ) ) ;

    /* cells in depth 32 */
    nor_HPC1 #(.security_order(3), .pipeline(1)) U2542 ( .ina ({new_AGEMA_signal_18914, new_AGEMA_signal_18900, new_AGEMA_signal_18886, new_AGEMA_signal_18872}), .inb ({new_AGEMA_signal_3716, new_AGEMA_signal_3715, new_AGEMA_signal_3714, n2381}), .clk ( clk ), .rnd ({Fresh[8669], Fresh[8668], Fresh[8667], Fresh[8666], Fresh[8665], Fresh[8664], Fresh[8663], Fresh[8662], Fresh[8661], Fresh[8660]}), .outt ({new_AGEMA_signal_3719, new_AGEMA_signal_3718, new_AGEMA_signal_3717, n2427}) ) ;
    buf_clk new_AGEMA_reg_buffer_7428 ( .C ( clk ), .D ( new_AGEMA_signal_18927 ), .Q ( new_AGEMA_signal_18928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7442 ( .C ( clk ), .D ( new_AGEMA_signal_18941 ), .Q ( new_AGEMA_signal_18942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7456 ( .C ( clk ), .D ( new_AGEMA_signal_18955 ), .Q ( new_AGEMA_signal_18956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7470 ( .C ( clk ), .D ( new_AGEMA_signal_18969 ), .Q ( new_AGEMA_signal_18970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7474 ( .C ( clk ), .D ( new_AGEMA_signal_18973 ), .Q ( new_AGEMA_signal_18974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7480 ( .C ( clk ), .D ( new_AGEMA_signal_18979 ), .Q ( new_AGEMA_signal_18980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7486 ( .C ( clk ), .D ( new_AGEMA_signal_18985 ), .Q ( new_AGEMA_signal_18986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7492 ( .C ( clk ), .D ( new_AGEMA_signal_18991 ), .Q ( new_AGEMA_signal_18992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7498 ( .C ( clk ), .D ( new_AGEMA_signal_18997 ), .Q ( new_AGEMA_signal_18998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7504 ( .C ( clk ), .D ( new_AGEMA_signal_19003 ), .Q ( new_AGEMA_signal_19004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7510 ( .C ( clk ), .D ( new_AGEMA_signal_19009 ), .Q ( new_AGEMA_signal_19010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7516 ( .C ( clk ), .D ( new_AGEMA_signal_19015 ), .Q ( new_AGEMA_signal_19016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7520 ( .C ( clk ), .D ( new_AGEMA_signal_19019 ), .Q ( new_AGEMA_signal_19020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7524 ( .C ( clk ), .D ( new_AGEMA_signal_19023 ), .Q ( new_AGEMA_signal_19024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7528 ( .C ( clk ), .D ( new_AGEMA_signal_19027 ), .Q ( new_AGEMA_signal_19028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7532 ( .C ( clk ), .D ( new_AGEMA_signal_19031 ), .Q ( new_AGEMA_signal_19032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7540 ( .C ( clk ), .D ( new_AGEMA_signal_19039 ), .Q ( new_AGEMA_signal_19040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7548 ( .C ( clk ), .D ( new_AGEMA_signal_19047 ), .Q ( new_AGEMA_signal_19048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7556 ( .C ( clk ), .D ( new_AGEMA_signal_19055 ), .Q ( new_AGEMA_signal_19056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7564 ( .C ( clk ), .D ( new_AGEMA_signal_19063 ), .Q ( new_AGEMA_signal_19064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7572 ( .C ( clk ), .D ( new_AGEMA_signal_19071 ), .Q ( new_AGEMA_signal_19072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7580 ( .C ( clk ), .D ( new_AGEMA_signal_19079 ), .Q ( new_AGEMA_signal_19080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7588 ( .C ( clk ), .D ( new_AGEMA_signal_19087 ), .Q ( new_AGEMA_signal_19088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7596 ( .C ( clk ), .D ( new_AGEMA_signal_19095 ), .Q ( new_AGEMA_signal_19096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7604 ( .C ( clk ), .D ( new_AGEMA_signal_19103 ), .Q ( new_AGEMA_signal_19104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7612 ( .C ( clk ), .D ( new_AGEMA_signal_19111 ), .Q ( new_AGEMA_signal_19112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7620 ( .C ( clk ), .D ( new_AGEMA_signal_19119 ), .Q ( new_AGEMA_signal_19120 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7628 ( .C ( clk ), .D ( new_AGEMA_signal_19127 ), .Q ( new_AGEMA_signal_19128 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7636 ( .C ( clk ), .D ( new_AGEMA_signal_19135 ), .Q ( new_AGEMA_signal_19136 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7644 ( .C ( clk ), .D ( new_AGEMA_signal_19143 ), .Q ( new_AGEMA_signal_19144 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7652 ( .C ( clk ), .D ( new_AGEMA_signal_19151 ), .Q ( new_AGEMA_signal_19152 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7660 ( .C ( clk ), .D ( new_AGEMA_signal_19159 ), .Q ( new_AGEMA_signal_19160 ) ) ;

    /* cells in depth 33 */
    buf_clk new_AGEMA_reg_buffer_7475 ( .C ( clk ), .D ( new_AGEMA_signal_18974 ), .Q ( new_AGEMA_signal_18975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7481 ( .C ( clk ), .D ( new_AGEMA_signal_18980 ), .Q ( new_AGEMA_signal_18981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7487 ( .C ( clk ), .D ( new_AGEMA_signal_18986 ), .Q ( new_AGEMA_signal_18987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7493 ( .C ( clk ), .D ( new_AGEMA_signal_18992 ), .Q ( new_AGEMA_signal_18993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7499 ( .C ( clk ), .D ( new_AGEMA_signal_18998 ), .Q ( new_AGEMA_signal_18999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7505 ( .C ( clk ), .D ( new_AGEMA_signal_19004 ), .Q ( new_AGEMA_signal_19005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7511 ( .C ( clk ), .D ( new_AGEMA_signal_19010 ), .Q ( new_AGEMA_signal_19011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7517 ( .C ( clk ), .D ( new_AGEMA_signal_19016 ), .Q ( new_AGEMA_signal_19017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7521 ( .C ( clk ), .D ( new_AGEMA_signal_19020 ), .Q ( new_AGEMA_signal_19021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7525 ( .C ( clk ), .D ( new_AGEMA_signal_19024 ), .Q ( new_AGEMA_signal_19025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7529 ( .C ( clk ), .D ( new_AGEMA_signal_19028 ), .Q ( new_AGEMA_signal_19029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7533 ( .C ( clk ), .D ( new_AGEMA_signal_19032 ), .Q ( new_AGEMA_signal_19033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7541 ( .C ( clk ), .D ( new_AGEMA_signal_19040 ), .Q ( new_AGEMA_signal_19041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7549 ( .C ( clk ), .D ( new_AGEMA_signal_19048 ), .Q ( new_AGEMA_signal_19049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7557 ( .C ( clk ), .D ( new_AGEMA_signal_19056 ), .Q ( new_AGEMA_signal_19057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7565 ( .C ( clk ), .D ( new_AGEMA_signal_19064 ), .Q ( new_AGEMA_signal_19065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7573 ( .C ( clk ), .D ( new_AGEMA_signal_19072 ), .Q ( new_AGEMA_signal_19073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7581 ( .C ( clk ), .D ( new_AGEMA_signal_19080 ), .Q ( new_AGEMA_signal_19081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7589 ( .C ( clk ), .D ( new_AGEMA_signal_19088 ), .Q ( new_AGEMA_signal_19089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7597 ( .C ( clk ), .D ( new_AGEMA_signal_19096 ), .Q ( new_AGEMA_signal_19097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7605 ( .C ( clk ), .D ( new_AGEMA_signal_19104 ), .Q ( new_AGEMA_signal_19105 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7613 ( .C ( clk ), .D ( new_AGEMA_signal_19112 ), .Q ( new_AGEMA_signal_19113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7621 ( .C ( clk ), .D ( new_AGEMA_signal_19120 ), .Q ( new_AGEMA_signal_19121 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7629 ( .C ( clk ), .D ( new_AGEMA_signal_19128 ), .Q ( new_AGEMA_signal_19129 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7637 ( .C ( clk ), .D ( new_AGEMA_signal_19136 ), .Q ( new_AGEMA_signal_19137 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7645 ( .C ( clk ), .D ( new_AGEMA_signal_19144 ), .Q ( new_AGEMA_signal_19145 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7653 ( .C ( clk ), .D ( new_AGEMA_signal_19152 ), .Q ( new_AGEMA_signal_19153 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7661 ( .C ( clk ), .D ( new_AGEMA_signal_19160 ), .Q ( new_AGEMA_signal_19161 ) ) ;

    /* cells in depth 34 */
    nand_HPC1 #(.security_order(3), .pipeline(1)) U2584 ( .ina ({new_AGEMA_signal_3719, new_AGEMA_signal_3718, new_AGEMA_signal_3717, n2427}), .inb ({new_AGEMA_signal_18970, new_AGEMA_signal_18956, new_AGEMA_signal_18942, new_AGEMA_signal_18928}), .clk ( clk ), .rnd ({Fresh[8679], Fresh[8678], Fresh[8677], Fresh[8676], Fresh[8675], Fresh[8674], Fresh[8673], Fresh[8672], Fresh[8671], Fresh[8670]}), .outt ({new_AGEMA_signal_3722, new_AGEMA_signal_3721, new_AGEMA_signal_3720, N563}) ) ;
    buf_clk new_AGEMA_reg_buffer_7476 ( .C ( clk ), .D ( new_AGEMA_signal_18975 ), .Q ( new_AGEMA_signal_18976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7482 ( .C ( clk ), .D ( new_AGEMA_signal_18981 ), .Q ( new_AGEMA_signal_18982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7488 ( .C ( clk ), .D ( new_AGEMA_signal_18987 ), .Q ( new_AGEMA_signal_18988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7494 ( .C ( clk ), .D ( new_AGEMA_signal_18993 ), .Q ( new_AGEMA_signal_18994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7500 ( .C ( clk ), .D ( new_AGEMA_signal_18999 ), .Q ( new_AGEMA_signal_19000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7506 ( .C ( clk ), .D ( new_AGEMA_signal_19005 ), .Q ( new_AGEMA_signal_19006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7512 ( .C ( clk ), .D ( new_AGEMA_signal_19011 ), .Q ( new_AGEMA_signal_19012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7518 ( .C ( clk ), .D ( new_AGEMA_signal_19017 ), .Q ( new_AGEMA_signal_19018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7522 ( .C ( clk ), .D ( new_AGEMA_signal_19021 ), .Q ( new_AGEMA_signal_19022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7526 ( .C ( clk ), .D ( new_AGEMA_signal_19025 ), .Q ( new_AGEMA_signal_19026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7530 ( .C ( clk ), .D ( new_AGEMA_signal_19029 ), .Q ( new_AGEMA_signal_19030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7534 ( .C ( clk ), .D ( new_AGEMA_signal_19033 ), .Q ( new_AGEMA_signal_19034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7542 ( .C ( clk ), .D ( new_AGEMA_signal_19041 ), .Q ( new_AGEMA_signal_19042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7550 ( .C ( clk ), .D ( new_AGEMA_signal_19049 ), .Q ( new_AGEMA_signal_19050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7558 ( .C ( clk ), .D ( new_AGEMA_signal_19057 ), .Q ( new_AGEMA_signal_19058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7566 ( .C ( clk ), .D ( new_AGEMA_signal_19065 ), .Q ( new_AGEMA_signal_19066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7574 ( .C ( clk ), .D ( new_AGEMA_signal_19073 ), .Q ( new_AGEMA_signal_19074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7582 ( .C ( clk ), .D ( new_AGEMA_signal_19081 ), .Q ( new_AGEMA_signal_19082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7590 ( .C ( clk ), .D ( new_AGEMA_signal_19089 ), .Q ( new_AGEMA_signal_19090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7598 ( .C ( clk ), .D ( new_AGEMA_signal_19097 ), .Q ( new_AGEMA_signal_19098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7606 ( .C ( clk ), .D ( new_AGEMA_signal_19105 ), .Q ( new_AGEMA_signal_19106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7614 ( .C ( clk ), .D ( new_AGEMA_signal_19113 ), .Q ( new_AGEMA_signal_19114 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7622 ( .C ( clk ), .D ( new_AGEMA_signal_19121 ), .Q ( new_AGEMA_signal_19122 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7630 ( .C ( clk ), .D ( new_AGEMA_signal_19129 ), .Q ( new_AGEMA_signal_19130 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7638 ( .C ( clk ), .D ( new_AGEMA_signal_19137 ), .Q ( new_AGEMA_signal_19138 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7646 ( .C ( clk ), .D ( new_AGEMA_signal_19145 ), .Q ( new_AGEMA_signal_19146 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7654 ( .C ( clk ), .D ( new_AGEMA_signal_19153 ), .Q ( new_AGEMA_signal_19154 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7662 ( .C ( clk ), .D ( new_AGEMA_signal_19161 ), .Q ( new_AGEMA_signal_19162 ) ) ;

    /* register cells */
    reg_masked #(.security_order(3), .pipeline(1)) SO_reg_7_ ( .clk ( clk ), .D ({new_AGEMA_signal_18994, new_AGEMA_signal_18988, new_AGEMA_signal_18982, new_AGEMA_signal_18976}), .Q ({SO_s3[7], SO_s2[7], SO_s1[7], SO_s0[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) SO_reg_6_ ( .clk ( clk ), .D ({new_AGEMA_signal_19018, new_AGEMA_signal_19012, new_AGEMA_signal_19006, new_AGEMA_signal_19000}), .Q ({SO_s3[6], SO_s2[6], SO_s1[6], SO_s0[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) SO_reg_5_ ( .clk ( clk ), .D ({new_AGEMA_signal_19034, new_AGEMA_signal_19030, new_AGEMA_signal_19026, new_AGEMA_signal_19022}), .Q ({SO_s3[5], SO_s2[5], SO_s1[5], SO_s0[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) SO_reg_4_ ( .clk ( clk ), .D ({new_AGEMA_signal_19066, new_AGEMA_signal_19058, new_AGEMA_signal_19050, new_AGEMA_signal_19042}), .Q ({SO_s3[4], SO_s2[4], SO_s1[4], SO_s0[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) SO_reg_3_ ( .clk ( clk ), .D ({new_AGEMA_signal_3722, new_AGEMA_signal_3721, new_AGEMA_signal_3720, N563}), .Q ({SO_s3[3], SO_s2[3], SO_s1[3], SO_s0[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) SO_reg_2_ ( .clk ( clk ), .D ({new_AGEMA_signal_19098, new_AGEMA_signal_19090, new_AGEMA_signal_19082, new_AGEMA_signal_19074}), .Q ({SO_s3[2], SO_s2[2], SO_s1[2], SO_s0[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) SO_reg_1_ ( .clk ( clk ), .D ({new_AGEMA_signal_19130, new_AGEMA_signal_19122, new_AGEMA_signal_19114, new_AGEMA_signal_19106}), .Q ({SO_s3[1], SO_s2[1], SO_s1[1], SO_s0[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) SO_reg_0_ ( .clk ( clk ), .D ({new_AGEMA_signal_19162, new_AGEMA_signal_19154, new_AGEMA_signal_19146, new_AGEMA_signal_19138}), .Q ({SO_s3[0], SO_s2[0], SO_s1[0], SO_s0[0]}) ) ;
endmodule
