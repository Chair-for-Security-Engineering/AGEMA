/* modified netlist. Source: module sbox in file Designs/AESSbox//Canright/AGEMA/sbox.v */
/* clock gating is added to the circuit, the latency increased 16 time(s)  */

module sbox_HPC2_AIG_ClockGating_d2 (X_s0, clk, X_s1, X_s2, Fresh, rst, Y_s0, Y_s1, Y_s2, Synch);
    input [7:0] X_s0 ;
    input clk ;
    input [7:0] X_s1 ;
    input [7:0] X_s2 ;
    input rst ;
    input [263:0] Fresh ;
    output [7:0] Y_s0 ;
    output [7:0] Y_s1 ;
    output [7:0] Y_s2 ;
    output Synch ;
    wire signal_160 ;
    wire signal_161 ;
    wire signal_162 ;
    wire signal_163 ;
    wire signal_164 ;
    wire signal_165 ;
    wire signal_166 ;
    wire signal_167 ;
    wire signal_192 ;
    wire signal_193 ;
    wire signal_194 ;
    wire signal_195 ;
    wire signal_196 ;
    wire signal_197 ;
    wire signal_198 ;
    wire signal_199 ;
    wire signal_200 ;
    wire signal_201 ;
    wire signal_202 ;
    wire signal_203 ;
    wire signal_204 ;
    wire signal_205 ;
    wire signal_206 ;
    wire signal_207 ;
    wire signal_208 ;
    wire signal_209 ;
    wire signal_210 ;
    wire signal_211 ;
    wire signal_212 ;
    wire signal_213 ;
    wire signal_214 ;
    wire signal_215 ;
    wire signal_216 ;
    wire signal_217 ;
    wire signal_218 ;
    wire signal_219 ;
    wire signal_220 ;
    wire signal_221 ;
    wire signal_222 ;
    wire signal_223 ;
    wire signal_224 ;
    wire signal_225 ;
    wire signal_226 ;
    wire signal_227 ;
    wire signal_228 ;
    wire signal_229 ;
    wire signal_230 ;
    wire signal_231 ;
    wire signal_232 ;
    wire signal_233 ;
    wire signal_234 ;
    wire signal_235 ;
    wire signal_236 ;
    wire signal_237 ;
    wire signal_238 ;
    wire signal_239 ;
    wire signal_240 ;
    wire signal_241 ;
    wire signal_242 ;
    wire signal_243 ;
    wire signal_244 ;
    wire signal_245 ;
    wire signal_246 ;
    wire signal_247 ;
    wire signal_248 ;
    wire signal_249 ;
    wire signal_250 ;
    wire signal_251 ;
    wire signal_252 ;
    wire signal_253 ;
    wire signal_254 ;
    wire signal_255 ;
    wire signal_256 ;
    wire signal_257 ;
    wire signal_258 ;
    wire signal_259 ;
    wire signal_260 ;
    wire signal_261 ;
    wire signal_262 ;
    wire signal_263 ;
    wire signal_264 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_285 ;
    wire signal_286 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_295 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_352 ;
    wire signal_353 ;
    wire signal_354 ;
    wire signal_355 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_359 ;
    wire signal_360 ;
    wire signal_361 ;
    wire signal_362 ;
    wire signal_363 ;
    wire signal_364 ;
    wire signal_365 ;
    wire signal_366 ;
    wire signal_367 ;
    wire signal_368 ;
    wire signal_369 ;
    wire signal_370 ;
    wire signal_371 ;
    wire signal_372 ;
    wire signal_373 ;
    wire signal_374 ;
    wire signal_375 ;
    wire signal_376 ;
    wire signal_377 ;
    wire signal_378 ;
    wire signal_379 ;
    wire signal_380 ;
    wire signal_381 ;
    wire signal_382 ;
    wire signal_383 ;
    wire signal_384 ;
    wire signal_385 ;
    wire signal_386 ;
    wire signal_387 ;
    wire signal_388 ;
    wire signal_389 ;
    wire signal_390 ;
    wire signal_391 ;
    wire signal_392 ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_415 ;
    wire signal_416 ;
    wire signal_417 ;
    wire signal_418 ;
    wire signal_419 ;
    wire signal_420 ;
    wire signal_421 ;
    wire signal_422 ;
    wire signal_423 ;
    wire signal_424 ;
    wire signal_425 ;
    wire signal_426 ;
    wire signal_427 ;
    wire signal_428 ;
    wire signal_429 ;
    wire signal_430 ;
    wire signal_431 ;
    wire signal_432 ;
    wire signal_433 ;
    wire signal_434 ;
    wire signal_435 ;
    wire signal_436 ;
    wire signal_439 ;
    wire signal_440 ;
    wire signal_445 ;
    wire signal_446 ;
    wire signal_451 ;
    wire signal_452 ;
    wire signal_453 ;
    wire signal_454 ;
    wire signal_455 ;
    wire signal_456 ;
    wire signal_459 ;
    wire signal_460 ;
    wire signal_461 ;
    wire signal_462 ;
    wire signal_463 ;
    wire signal_464 ;
    wire signal_465 ;
    wire signal_466 ;
    wire signal_467 ;
    wire signal_468 ;
    wire signal_471 ;
    wire signal_472 ;
    wire signal_473 ;
    wire signal_474 ;
    wire signal_477 ;
    wire signal_478 ;
    wire signal_479 ;
    wire signal_480 ;
    wire signal_481 ;
    wire signal_482 ;
    wire signal_483 ;
    wire signal_484 ;
    wire signal_485 ;
    wire signal_486 ;
    wire signal_487 ;
    wire signal_488 ;
    wire signal_489 ;
    wire signal_490 ;
    wire signal_491 ;
    wire signal_492 ;
    wire signal_493 ;
    wire signal_494 ;
    wire signal_495 ;
    wire signal_496 ;
    wire signal_497 ;
    wire signal_498 ;
    wire signal_499 ;
    wire signal_500 ;
    wire signal_501 ;
    wire signal_502 ;
    wire signal_503 ;
    wire signal_504 ;
    wire signal_505 ;
    wire signal_506 ;
    wire signal_507 ;
    wire signal_508 ;
    wire signal_509 ;
    wire signal_510 ;
    wire signal_511 ;
    wire signal_512 ;
    wire signal_513 ;
    wire signal_514 ;
    wire signal_515 ;
    wire signal_516 ;
    wire signal_517 ;
    wire signal_518 ;
    wire signal_519 ;
    wire signal_520 ;
    wire signal_521 ;
    wire signal_522 ;
    wire signal_523 ;
    wire signal_524 ;
    wire signal_525 ;
    wire signal_526 ;
    wire signal_527 ;
    wire signal_528 ;
    wire signal_529 ;
    wire signal_530 ;
    wire signal_531 ;
    wire signal_532 ;
    wire signal_533 ;
    wire signal_534 ;
    wire signal_535 ;
    wire signal_536 ;
    wire signal_537 ;
    wire signal_538 ;
    wire signal_539 ;
    wire signal_540 ;
    wire signal_541 ;
    wire signal_542 ;
    wire signal_543 ;
    wire signal_544 ;
    wire signal_545 ;
    wire signal_546 ;
    wire signal_547 ;
    wire signal_548 ;
    wire signal_549 ;
    wire signal_550 ;
    wire signal_551 ;
    wire signal_552 ;
    wire signal_553 ;
    wire signal_554 ;
    wire signal_555 ;
    wire signal_556 ;
    wire signal_557 ;
    wire signal_558 ;
    wire signal_559 ;
    wire signal_560 ;
    wire signal_561 ;
    wire signal_562 ;
    wire signal_563 ;
    wire signal_564 ;
    wire signal_565 ;
    wire signal_566 ;
    wire signal_567 ;
    wire signal_568 ;
    wire signal_569 ;
    wire signal_570 ;
    wire signal_571 ;
    wire signal_572 ;
    wire signal_573 ;
    wire signal_574 ;
    wire signal_575 ;
    wire signal_576 ;
    wire signal_577 ;
    wire signal_578 ;
    wire signal_579 ;
    wire signal_580 ;
    wire signal_581 ;
    wire signal_582 ;
    wire signal_583 ;
    wire signal_584 ;
    wire signal_585 ;
    wire signal_586 ;
    wire signal_587 ;
    wire signal_588 ;
    wire signal_589 ;
    wire signal_590 ;
    wire signal_591 ;
    wire signal_592 ;
    wire signal_593 ;
    wire signal_594 ;
    wire signal_595 ;
    wire signal_596 ;
    wire signal_597 ;
    wire signal_598 ;
    wire signal_599 ;
    wire signal_600 ;
    wire signal_601 ;
    wire signal_602 ;
    wire signal_603 ;
    wire signal_604 ;
    wire signal_605 ;
    wire signal_606 ;
    wire signal_607 ;
    wire signal_608 ;
    wire signal_609 ;
    wire signal_610 ;
    wire signal_611 ;
    wire signal_612 ;
    wire signal_613 ;
    wire signal_614 ;
    wire signal_615 ;
    wire signal_616 ;
    wire signal_617 ;
    wire signal_618 ;
    wire signal_619 ;
    wire signal_620 ;
    wire signal_621 ;
    wire signal_622 ;
    wire signal_623 ;
    wire signal_624 ;
    wire signal_625 ;
    wire signal_626 ;
    wire signal_627 ;
    wire signal_628 ;
    wire signal_629 ;
    wire signal_630 ;
    wire signal_631 ;
    wire signal_632 ;
    wire signal_633 ;
    wire signal_634 ;
    wire signal_635 ;
    wire signal_636 ;
    wire signal_637 ;
    wire signal_638 ;
    wire signal_639 ;
    wire signal_640 ;
    wire signal_641 ;
    wire signal_642 ;
    wire signal_643 ;
    wire signal_644 ;
    wire signal_645 ;
    wire signal_646 ;
    wire signal_647 ;
    wire signal_648 ;
    wire signal_649 ;
    wire signal_650 ;
    wire signal_651 ;
    wire signal_652 ;
    wire signal_653 ;
    wire signal_654 ;
    wire signal_655 ;
    wire signal_656 ;
    wire signal_657 ;
    wire signal_658 ;
    wire signal_659 ;
    wire signal_660 ;
    wire signal_661 ;
    wire signal_662 ;
    wire signal_663 ;
    wire signal_664 ;
    wire signal_665 ;
    wire signal_666 ;
    wire signal_667 ;
    wire signal_668 ;
    wire signal_669 ;
    wire signal_670 ;
    wire signal_671 ;
    wire signal_672 ;
    wire signal_673 ;
    wire signal_674 ;
    wire signal_675 ;
    wire signal_676 ;
    wire signal_677 ;
    wire signal_678 ;
    wire signal_679 ;
    wire signal_680 ;
    wire signal_681 ;
    wire signal_682 ;
    wire signal_683 ;
    wire signal_684 ;
    wire signal_685 ;
    wire signal_686 ;
    wire signal_687 ;
    wire signal_688 ;
    wire signal_689 ;
    wire signal_690 ;
    wire signal_691 ;
    wire signal_692 ;
    wire signal_693 ;
    wire signal_694 ;
    wire signal_695 ;
    wire signal_696 ;
    wire signal_697 ;
    wire signal_698 ;
    wire signal_699 ;
    wire signal_700 ;
    wire signal_701 ;
    wire signal_702 ;
    wire signal_703 ;
    wire signal_704 ;
    wire signal_705 ;
    wire signal_706 ;
    wire signal_707 ;
    wire signal_708 ;
    wire signal_709 ;
    wire signal_710 ;
    wire signal_711 ;
    wire signal_712 ;
    wire signal_713 ;
    wire signal_714 ;
    wire signal_715 ;
    wire signal_716 ;
    wire signal_717 ;
    wire signal_718 ;
    wire signal_719 ;
    wire signal_720 ;
    wire signal_721 ;
    wire signal_722 ;
    wire signal_723 ;
    wire signal_724 ;
    wire signal_725 ;
    wire signal_726 ;
    wire signal_727 ;
    wire signal_728 ;
    wire signal_729 ;
    wire signal_730 ;
    wire signal_731 ;
    wire signal_732 ;
    wire signal_733 ;
    wire signal_734 ;
    wire signal_735 ;
    wire signal_736 ;
    wire signal_737 ;
    wire signal_738 ;
    wire signal_739 ;
    wire signal_740 ;
    wire signal_741 ;
    wire signal_742 ;
    wire signal_743 ;
    wire signal_744 ;
    wire signal_745 ;
    wire signal_746 ;
    wire signal_747 ;
    wire signal_748 ;
    wire signal_749 ;
    wire signal_750 ;
    wire signal_751 ;
    wire signal_752 ;
    wire signal_753 ;
    wire signal_754 ;
    wire signal_755 ;
    wire signal_756 ;
    wire signal_757 ;
    wire signal_758 ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_768 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_771 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_774 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_777 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_780 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_783 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_786 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_789 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_792 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_809 ;
    wire signal_810 ;
    wire signal_811 ;
    wire signal_812 ;
    wire signal_813 ;
    wire signal_814 ;
    wire signal_815 ;
    wire signal_816 ;
    wire signal_817 ;
    wire signal_818 ;
    wire signal_819 ;
    wire signal_820 ;
    wire signal_821 ;
    wire signal_822 ;
    wire signal_823 ;
    wire signal_824 ;
    wire signal_825 ;
    wire signal_826 ;
    wire signal_827 ;
    wire signal_828 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_831 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_834 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_837 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_840 ;
    wire signal_841 ;
    wire signal_842 ;
    wire signal_843 ;
    wire signal_844 ;
    wire signal_845 ;
    wire signal_846 ;
    wire signal_847 ;
    wire signal_848 ;
    wire signal_849 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_852 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_855 ;
    wire signal_856 ;
    wire signal_857 ;
    wire signal_858 ;
    wire signal_859 ;
    wire signal_860 ;
    wire signal_861 ;
    wire signal_862 ;
    wire signal_863 ;
    wire signal_864 ;
    wire signal_865 ;
    wire signal_866 ;
    wire signal_867 ;
    wire signal_868 ;
    wire signal_869 ;
    wire signal_870 ;
    wire signal_871 ;
    wire signal_872 ;
    wire signal_873 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_879 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_885 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_888 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_891 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_894 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_897 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_900 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_903 ;
    wire signal_904 ;
    wire signal_905 ;
    wire signal_906 ;
    wire signal_907 ;
    wire signal_908 ;
    wire signal_909 ;
    wire signal_910 ;
    wire signal_911 ;
    wire signal_912 ;
    wire signal_913 ;
    wire signal_914 ;
    wire signal_915 ;
    wire signal_916 ;
    wire signal_917 ;
    wire signal_918 ;
    wire signal_919 ;
    wire signal_920 ;
    wire signal_921 ;
    wire signal_922 ;
    wire signal_923 ;
    wire signal_924 ;
    wire signal_925 ;
    wire signal_926 ;
    wire signal_927 ;
    wire signal_928 ;
    wire signal_929 ;
    wire signal_930 ;
    wire signal_931 ;
    wire signal_932 ;
    wire signal_933 ;
    wire signal_934 ;
    wire signal_935 ;
    wire signal_936 ;
    wire signal_937 ;
    wire signal_938 ;
    wire signal_939 ;
    wire signal_940 ;
    wire signal_941 ;
    wire signal_942 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_1238 ;

    /* cells in depth 0 */
    not_masked #(.security_order(2), .pipeline(0)) cell_176 ( .a ({X_s2[0], X_s1[0], X_s0[0]}), .b ({signal_440, signal_439, signal_192}) ) ;
    INV_X1 cell_177 ( .A ( 1'b1 ), .ZN ( signal_193 ) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_178 ( .a ({X_s2[6], X_s1[6], X_s0[6]}), .b ({X_s2[4], X_s1[4], X_s0[4]}), .c ({signal_446, signal_445, signal_194}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_179 ( .a ({X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s2[5], X_s1[5], X_s0[5]}), .c ({signal_452, signal_451, signal_195}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_180 ( .a ({X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s2[4], X_s1[4], X_s0[4]}), .c ({signal_454, signal_453, signal_196}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_181 ( .a ({X_s2[6], X_s1[6], X_s0[6]}), .b ({X_s2[0], X_s1[0], X_s0[0]}), .c ({signal_456, signal_455, signal_197}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_182 ( .a ({X_s2[3], X_s1[3], X_s0[3]}), .b ({X_s2[0], X_s1[0], X_s0[0]}), .c ({signal_460, signal_459, signal_198}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_183 ( .a ({signal_454, signal_453, signal_196}), .b ({signal_462, signal_461, signal_199}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_186 ( .a ({X_s2[6], X_s1[6], X_s0[6]}), .b ({signal_454, signal_453, signal_196}), .c ({signal_468, signal_467, signal_202}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_187 ( .a ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_452, signal_451, signal_195}), .c ({signal_472, signal_471, signal_203}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_188 ( .a ({signal_452, signal_451, signal_195}), .b ({signal_456, signal_455, signal_197}), .c ({signal_474, signal_473, signal_204}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_189 ( .a ({X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_456, signal_455, signal_197}), .c ({signal_478, signal_477, signal_205}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_190 ( .a ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_460, signal_459, signal_198}), .c ({signal_480, signal_479, signal_206}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_191 ( .a ({X_s2[5], X_s1[5], X_s0[5]}), .b ({signal_456, signal_455, signal_197}), .c ({signal_482, signal_481, signal_207}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_192 ( .a ({X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_460, signal_459, signal_198}), .c ({signal_484, signal_483, signal_208}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_193 ( .a ({signal_474, signal_473, signal_204}), .b ({signal_486, signal_485, signal_209}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_194 ( .a ({signal_482, signal_481, signal_207}), .b ({signal_488, signal_487, signal_210}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_201 ( .a ({X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_482, signal_481, signal_207}), .c ({signal_502, signal_501, signal_217}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_202 ( .a ({signal_472, signal_471, signal_203}), .b ({signal_478, signal_477, signal_205}), .c ({signal_504, signal_503, signal_218}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_203 ( .a ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_478, signal_477, signal_205}), .c ({signal_506, signal_505, signal_219}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_204 ( .a ({X_s2[3], X_s1[3], X_s0[3]}), .b ({signal_478, signal_477, signal_205}), .c ({signal_508, signal_507, signal_220}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_205 ( .a ({X_s2[4], X_s1[4], X_s0[4]}), .b ({signal_482, signal_481, signal_207}), .c ({signal_510, signal_509, signal_221}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_206 ( .a ({signal_454, signal_453, signal_196}), .b ({signal_484, signal_483, signal_208}), .c ({signal_512, signal_511, signal_222}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_208 ( .a ({signal_502, signal_501, signal_217}), .b ({signal_516, signal_515, signal_224}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_209 ( .a ({signal_504, signal_503, signal_218}), .b ({signal_518, signal_517, signal_225}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_210 ( .a ({signal_510, signal_509, signal_221}), .b ({signal_520, signal_519, signal_226}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_211 ( .a ({signal_512, signal_511, signal_222}), .b ({signal_522, signal_521, signal_227}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_219 ( .a ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_508, signal_507, signal_220}), .c ({signal_538, signal_537, signal_235}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_220 ( .a ({X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_510, signal_509, signal_221}), .c ({signal_540, signal_539, signal_236}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_222 ( .a ({signal_538, signal_537, signal_235}), .b ({signal_544, signal_543, signal_238}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_223 ( .a ({signal_540, signal_539, signal_236}), .b ({signal_546, signal_545, signal_239}) ) ;
    ClockGatingController #(17) cell_429 ( .clk ( clk ), .rst ( rst ), .GatedClk ( signal_1238 ), .Synch ( Synch ) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_184 ( .a ({signal_440, signal_439, signal_192}), .b ({1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[2], Fresh[1], Fresh[0]}), .c ({signal_464, signal_463, signal_200}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_185 ( .a ({1'b0, 1'b0, signal_193}), .b ({signal_446, signal_445, signal_194}), .clk ( clk ), .r ({Fresh[5], Fresh[4], Fresh[3]}), .c ({signal_466, signal_465, signal_201}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_195 ( .a ({signal_464, signal_463, signal_200}), .b ({signal_490, signal_489, signal_211}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_196 ( .a ({signal_466, signal_465, signal_201}), .b ({signal_492, signal_491, signal_212}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_197 ( .a ({1'b0, 1'b0, signal_193}), .b ({signal_472, signal_471, signal_203}), .clk ( clk ), .r ({Fresh[8], Fresh[7], Fresh[6]}), .c ({signal_494, signal_493, signal_213}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_198 ( .a ({1'b0, 1'b0, signal_193}), .b ({signal_480, signal_479, signal_206}), .clk ( clk ), .r ({Fresh[11], Fresh[10], Fresh[9]}), .c ({signal_496, signal_495, signal_214}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_199 ( .a ({1'b0, 1'b0, signal_193}), .b ({signal_462, signal_461, signal_199}), .clk ( clk ), .r ({Fresh[14], Fresh[13], Fresh[12]}), .c ({signal_498, signal_497, signal_215}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_200 ( .a ({1'b0, 1'b0, signal_193}), .b ({signal_468, signal_467, signal_202}), .clk ( clk ), .r ({Fresh[17], Fresh[16], Fresh[15]}), .c ({signal_500, signal_499, signal_216}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_207 ( .a ({signal_494, signal_493, signal_213}), .b ({signal_514, signal_513, signal_223}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_212 ( .a ({signal_496, signal_495, signal_214}), .b ({signal_524, signal_523, signal_228}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_213 ( .a ({signal_498, signal_497, signal_215}), .b ({signal_526, signal_525, signal_229}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_214 ( .a ({signal_500, signal_499, signal_216}), .b ({signal_528, signal_527, signal_230}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_215 ( .a ({1'b0, 1'b0, 1'b1}), .b ({signal_488, signal_487, signal_210}), .clk ( clk ), .r ({Fresh[20], Fresh[19], Fresh[18]}), .c ({signal_530, signal_529, signal_231}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_216 ( .a ({1'b0, 1'b0, signal_193}), .b ({signal_506, signal_505, signal_219}), .clk ( clk ), .r ({Fresh[23], Fresh[22], Fresh[21]}), .c ({signal_532, signal_531, signal_232}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_217 ( .a ({1'b0, 1'b0, signal_193}), .b ({signal_508, signal_507, signal_220}), .clk ( clk ), .r ({Fresh[26], Fresh[25], Fresh[24]}), .c ({signal_534, signal_533, signal_233}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_218 ( .a ({1'b0, 1'b0, 1'b1}), .b ({signal_486, signal_485, signal_209}), .clk ( clk ), .r ({Fresh[29], Fresh[28], Fresh[27]}), .c ({signal_536, signal_535, signal_234}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_221 ( .a ({signal_530, signal_529, signal_231}), .b ({signal_542, signal_541, signal_237}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_224 ( .a ({signal_532, signal_531, signal_232}), .b ({signal_548, signal_547, signal_240}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_225 ( .a ({signal_534, signal_533, signal_233}), .b ({signal_550, signal_549, signal_241}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_226 ( .a ({signal_536, signal_535, signal_234}), .b ({signal_552, signal_551, signal_242}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_228 ( .a ({1'b0, 1'b0, 1'b1}), .b ({signal_518, signal_517, signal_225}), .clk ( clk ), .r ({Fresh[32], Fresh[31], Fresh[30]}), .c ({signal_556, signal_555, signal_244}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_229 ( .a ({1'b0, 1'b0, 1'b1}), .b ({signal_520, signal_519, signal_226}), .clk ( clk ), .r ({Fresh[35], Fresh[34], Fresh[33]}), .c ({signal_558, signal_557, signal_245}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_230 ( .a ({1'b0, 1'b0, 1'b1}), .b ({signal_516, signal_515, signal_224}), .clk ( clk ), .r ({Fresh[38], Fresh[37], Fresh[36]}), .c ({signal_560, signal_559, signal_246}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_231 ( .a ({1'b0, 1'b0, 1'b1}), .b ({signal_522, signal_521, signal_227}), .clk ( clk ), .r ({Fresh[41], Fresh[40], Fresh[39]}), .c ({signal_562, signal_561, signal_247}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_232 ( .a ({signal_556, signal_555, signal_244}), .b ({signal_564, signal_563, signal_248}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_233 ( .a ({signal_558, signal_557, signal_245}), .b ({signal_566, signal_565, signal_249}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_234 ( .a ({signal_560, signal_559, signal_246}), .b ({signal_568, signal_567, signal_250}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_235 ( .a ({signal_562, signal_561, signal_247}), .b ({signal_570, signal_569, signal_251}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_238 ( .a ({1'b0, 1'b0, signal_193}), .b ({signal_546, signal_545, signal_239}), .clk ( clk ), .r ({Fresh[44], Fresh[43], Fresh[42]}), .c ({signal_576, signal_575, signal_254}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_239 ( .a ({1'b0, 1'b0, 1'b1}), .b ({signal_544, signal_543, signal_238}), .clk ( clk ), .r ({Fresh[47], Fresh[46], Fresh[45]}), .c ({signal_578, signal_577, signal_255}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_241 ( .a ({signal_576, signal_575, signal_254}), .b ({signal_582, signal_581, signal_257}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_242 ( .a ({signal_578, signal_577, signal_255}), .b ({signal_584, signal_583, signal_258}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_227 ( .a ({signal_514, signal_513, signal_223}), .b ({signal_490, signal_489, signal_211}), .clk ( clk ), .r ({Fresh[50], Fresh[49], Fresh[48]}), .c ({signal_554, signal_553, signal_243}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_236 ( .a ({signal_524, signal_523, signal_228}), .b ({signal_542, signal_541, signal_237}), .clk ( clk ), .r ({Fresh[53], Fresh[52], Fresh[51]}), .c ({signal_572, signal_571, signal_252}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_237 ( .a ({signal_550, signal_549, signal_241}), .b ({signal_552, signal_551, signal_242}), .clk ( clk ), .r ({Fresh[56], Fresh[55], Fresh[54]}), .c ({signal_574, signal_573, signal_253}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_240 ( .a ({signal_574, signal_573, signal_253}), .b ({signal_580, signal_579, signal_256}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_243 ( .a ({signal_526, signal_525, signal_229}), .b ({signal_564, signal_563, signal_248}), .clk ( clk ), .r ({Fresh[59], Fresh[58], Fresh[57]}), .c ({signal_586, signal_585, signal_259}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_244 ( .a ({signal_548, signal_547, signal_240}), .b ({signal_566, signal_565, signal_249}), .clk ( clk ), .r ({Fresh[62], Fresh[61], Fresh[60]}), .c ({signal_588, signal_587, signal_260}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_245 ( .a ({signal_492, signal_491, signal_212}), .b ({signal_568, signal_567, signal_250}), .clk ( clk ), .r ({Fresh[65], Fresh[64], Fresh[63]}), .c ({signal_590, signal_589, signal_261}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_246 ( .a ({signal_528, signal_527, signal_230}), .b ({signal_570, signal_569, signal_251}), .clk ( clk ), .r ({Fresh[68], Fresh[67], Fresh[66]}), .c ({signal_592, signal_591, signal_262}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_247 ( .a ({signal_582, signal_581, signal_257}), .b ({signal_584, signal_583, signal_258}), .clk ( clk ), .r ({Fresh[71], Fresh[70], Fresh[69]}), .c ({signal_594, signal_593, signal_263}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_251 ( .a ({signal_554, signal_553, signal_243}), .b ({signal_592, signal_591, signal_262}), .c ({signal_602, signal_601, signal_267}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_252 ( .a ({signal_572, signal_571, signal_252}), .b ({signal_592, signal_591, signal_262}), .c ({signal_604, signal_603, signal_268}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_253 ( .a ({signal_590, signal_589, signal_261}), .b ({signal_574, signal_573, signal_253}), .c ({signal_606, signal_605, signal_269}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_254 ( .a ({signal_586, signal_585, signal_259}), .b ({signal_588, signal_587, signal_260}), .c ({signal_608, signal_607, signal_270}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_255 ( .a ({signal_588, signal_587, signal_260}), .b ({signal_574, signal_573, signal_253}), .c ({signal_610, signal_609, signal_271}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_256 ( .a ({signal_586, signal_585, signal_259}), .b ({signal_590, signal_589, signal_261}), .c ({signal_612, signal_611, signal_272}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_257 ( .a ({signal_594, signal_593, signal_263}), .b ({signal_614, signal_613, signal_273}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_258 ( .a ({signal_604, signal_603, signal_268}), .b ({signal_616, signal_615, signal_274}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_259 ( .a ({signal_606, signal_605, signal_269}), .b ({signal_618, signal_617, signal_275}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_260 ( .a ({signal_610, signal_609, signal_271}), .b ({signal_620, signal_619, signal_276}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_261 ( .a ({signal_612, signal_611, signal_272}), .b ({signal_622, signal_621, signal_277}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_264 ( .a ({signal_572, signal_571, signal_252}), .b ({signal_594, signal_593, signal_263}), .c ({signal_628, signal_627, signal_280}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_265 ( .a ({signal_554, signal_553, signal_243}), .b ({signal_594, signal_593, signal_263}), .c ({signal_630, signal_629, signal_281}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_266 ( .a ({signal_610, signal_609, signal_271}), .b ({signal_612, signal_611, signal_272}), .c ({signal_632, signal_631, signal_282}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_267 ( .a ({signal_628, signal_627, signal_280}), .b ({signal_634, signal_633, signal_283}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_268 ( .a ({signal_630, signal_629, signal_281}), .b ({signal_636, signal_635, signal_284}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_273 ( .a ({signal_604, signal_603, signal_268}), .b ({signal_630, signal_629, signal_281}), .c ({signal_646, signal_645, signal_289}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_248 ( .a ({signal_586, signal_585, signal_259}), .b ({signal_592, signal_591, signal_262}), .clk ( clk ), .r ({Fresh[74], Fresh[73], Fresh[72]}), .c ({signal_596, signal_595, signal_264}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_249 ( .a ({signal_554, signal_553, signal_243}), .b ({signal_588, signal_587, signal_260}), .clk ( clk ), .r ({Fresh[77], Fresh[76], Fresh[75]}), .c ({signal_598, signal_597, signal_265}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_250 ( .a ({signal_572, signal_571, signal_252}), .b ({signal_590, signal_589, signal_261}), .clk ( clk ), .r ({Fresh[80], Fresh[79], Fresh[78]}), .c ({signal_600, signal_599, signal_266}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_262 ( .a ({signal_602, signal_601, signal_267}), .b ({signal_608, signal_607, signal_270}), .clk ( clk ), .r ({Fresh[83], Fresh[82], Fresh[81]}), .c ({signal_624, signal_623, signal_278}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_263 ( .a ({signal_604, signal_603, signal_268}), .b ({signal_612, signal_611, signal_272}), .clk ( clk ), .r ({Fresh[86], Fresh[85], Fresh[84]}), .c ({signal_626, signal_625, signal_279}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_269 ( .a ({signal_616, signal_615, signal_274}), .b ({signal_622, signal_621, signal_277}), .clk ( clk ), .r ({Fresh[89], Fresh[88], Fresh[87]}), .c ({signal_638, signal_637, signal_285}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_270 ( .a ({signal_580, signal_579, signal_256}), .b ({signal_614, signal_613, signal_273}), .clk ( clk ), .r ({Fresh[92], Fresh[91], Fresh[90]}), .c ({signal_640, signal_639, signal_286}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_271 ( .a ({signal_606, signal_605, signal_269}), .b ({signal_628, signal_627, signal_280}), .clk ( clk ), .r ({Fresh[95], Fresh[94], Fresh[93]}), .c ({signal_642, signal_641, signal_287}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_272 ( .a ({signal_610, signal_609, signal_271}), .b ({signal_630, signal_629, signal_281}), .clk ( clk ), .r ({Fresh[98], Fresh[97], Fresh[96]}), .c ({signal_644, signal_643, signal_288}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_274 ( .a ({signal_620, signal_619, signal_276}), .b ({signal_636, signal_635, signal_284}), .clk ( clk ), .r ({Fresh[101], Fresh[100], Fresh[99]}), .c ({signal_648, signal_647, signal_290}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_275 ( .a ({signal_618, signal_617, signal_275}), .b ({signal_634, signal_633, signal_283}), .clk ( clk ), .r ({Fresh[104], Fresh[103], Fresh[102]}), .c ({signal_650, signal_649, signal_291}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_276 ( .a ({signal_632, signal_631, signal_282}), .b ({signal_646, signal_645, signal_289}), .clk ( clk ), .r ({Fresh[107], Fresh[106], Fresh[105]}), .c ({signal_652, signal_651, signal_292}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_277 ( .a ({signal_598, signal_597, signal_265}), .b ({signal_638, signal_637, signal_285}), .c ({signal_654, signal_653, signal_293}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_278 ( .a ({signal_624, signal_623, signal_278}), .b ({signal_644, signal_643, signal_288}), .c ({signal_656, signal_655, signal_294}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_279 ( .a ({signal_640, signal_639, signal_286}), .b ({signal_642, signal_641, signal_287}), .c ({signal_658, signal_657, signal_295}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_280 ( .a ({signal_596, signal_595, signal_264}), .b ({signal_648, signal_647, signal_290}), .c ({signal_660, signal_659, signal_296}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_281 ( .a ({signal_600, signal_599, signal_266}), .b ({signal_650, signal_649, signal_291}), .c ({signal_662, signal_661, signal_297}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_282 ( .a ({signal_624, signal_623, signal_278}), .b ({signal_652, signal_651, signal_292}), .c ({signal_664, signal_663, signal_298}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_283 ( .a ({signal_654, signal_653, signal_293}), .b ({signal_656, signal_655, signal_294}), .c ({signal_666, signal_665, signal_299}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_284 ( .a ({signal_644, signal_643, signal_288}), .b ({signal_652, signal_651, signal_292}), .c ({signal_668, signal_667, signal_300}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_285 ( .a ({signal_626, signal_625, signal_279}), .b ({signal_658, signal_657, signal_295}), .c ({signal_670, signal_669, signal_301}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_286 ( .a ({signal_666, signal_665, signal_299}), .b ({signal_672, signal_671, signal_302}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_287 ( .a ({signal_660, signal_659, signal_296}), .b ({signal_664, signal_663, signal_298}), .c ({signal_674, signal_673, signal_303}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_288 ( .a ({signal_662, signal_661, signal_297}), .b ({signal_668, signal_667, signal_300}), .c ({signal_676, signal_675, signal_304}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_289 ( .a ({signal_644, signal_643, signal_288}), .b ({signal_670, signal_669, signal_301}), .c ({signal_678, signal_677, signal_305}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_290 ( .a ({signal_674, signal_673, signal_303}), .b ({signal_680, signal_679, signal_306}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_291 ( .a ({signal_676, signal_675, signal_304}), .b ({signal_682, signal_681, signal_307}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_292 ( .a ({signal_678, signal_677, signal_305}), .b ({signal_684, signal_683, signal_308}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_294 ( .a ({signal_666, signal_665, signal_299}), .b ({signal_674, signal_673, signal_303}), .c ({signal_688, signal_687, signal_310}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_295 ( .a ({signal_676, signal_675, signal_304}), .b ({signal_678, signal_677, signal_305}), .c ({signal_690, signal_689, signal_311}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_296 ( .a ({signal_688, signal_687, signal_310}), .b ({signal_692, signal_691, signal_312}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_297 ( .a ({signal_690, signal_689, signal_311}), .b ({signal_694, signal_693, signal_313}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_293 ( .a ({signal_674, signal_673, signal_303}), .b ({signal_676, signal_675, signal_304}), .clk ( clk ), .r ({Fresh[110], Fresh[109], Fresh[108]}), .c ({signal_686, signal_685, signal_309}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_298 ( .a ({signal_672, signal_671, signal_302}), .b ({signal_684, signal_683, signal_308}), .clk ( clk ), .r ({Fresh[113], Fresh[112], Fresh[111]}), .c ({signal_696, signal_695, signal_314}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_299 ( .a ({signal_688, signal_687, signal_310}), .b ({signal_690, signal_689, signal_311}), .clk ( clk ), .r ({Fresh[116], Fresh[115], Fresh[114]}), .c ({signal_698, signal_697, signal_315}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_300 ( .a ({signal_692, signal_691, signal_312}), .b ({signal_694, signal_693, signal_313}), .clk ( clk ), .r ({Fresh[119], Fresh[118], Fresh[117]}), .c ({signal_700, signal_699, signal_316}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_301 ( .a ({signal_686, signal_685, signal_309}), .b ({signal_698, signal_697, signal_315}), .c ({signal_702, signal_701, signal_317}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_302 ( .a ({signal_702, signal_701, signal_317}), .b ({signal_704, signal_703, signal_318}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_303 ( .a ({signal_696, signal_695, signal_314}), .b ({signal_700, signal_699, signal_316}), .c ({signal_706, signal_705, signal_319}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_304 ( .a ({signal_706, signal_705, signal_319}), .b ({signal_708, signal_707, signal_320}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_307 ( .a ({signal_702, signal_701, signal_317}), .b ({signal_706, signal_705, signal_319}), .c ({signal_714, signal_713, signal_323}) ) ;

    /* cells in depth 9 */

    /* cells in depth 10 */
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_305 ( .a ({signal_684, signal_683, signal_308}), .b ({signal_704, signal_703, signal_318}), .clk ( clk ), .r ({Fresh[122], Fresh[121], Fresh[120]}), .c ({signal_710, signal_709, signal_321}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_306 ( .a ({signal_672, signal_671, signal_302}), .b ({signal_704, signal_703, signal_318}), .clk ( clk ), .r ({Fresh[125], Fresh[124], Fresh[123]}), .c ({signal_712, signal_711, signal_322}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_308 ( .a ({signal_682, signal_681, signal_307}), .b ({signal_708, signal_707, signal_320}), .clk ( clk ), .r ({Fresh[128], Fresh[127], Fresh[126]}), .c ({signal_716, signal_715, signal_324}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_309 ( .a ({signal_680, signal_679, signal_306}), .b ({signal_708, signal_707, signal_320}), .clk ( clk ), .r ({Fresh[131], Fresh[130], Fresh[129]}), .c ({signal_718, signal_717, signal_325}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_310 ( .a ({signal_690, signal_689, signal_311}), .b ({signal_714, signal_713, signal_323}), .clk ( clk ), .r ({Fresh[134], Fresh[133], Fresh[132]}), .c ({signal_720, signal_719, signal_326}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_311 ( .a ({signal_688, signal_687, signal_310}), .b ({signal_714, signal_713, signal_323}), .clk ( clk ), .r ({Fresh[137], Fresh[136], Fresh[135]}), .c ({signal_722, signal_721, signal_327}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_312 ( .a ({signal_716, signal_715, signal_324}), .b ({signal_720, signal_719, signal_326}), .c ({signal_724, signal_723, signal_328}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_313 ( .a ({signal_710, signal_709, signal_321}), .b ({signal_720, signal_719, signal_326}), .c ({signal_726, signal_725, signal_329}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_314 ( .a ({signal_718, signal_717, signal_325}), .b ({signal_722, signal_721, signal_327}), .c ({signal_728, signal_727, signal_330}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_315 ( .a ({signal_712, signal_711, signal_322}), .b ({signal_722, signal_721, signal_327}), .c ({signal_730, signal_729, signal_331}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_324 ( .a ({signal_728, signal_727, signal_330}), .b ({signal_730, signal_729, signal_331}), .c ({signal_748, signal_747, signal_340}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_325 ( .a ({signal_724, signal_723, signal_328}), .b ({signal_726, signal_725, signal_329}), .c ({signal_750, signal_749, signal_341}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_326 ( .a ({signal_726, signal_725, signal_329}), .b ({signal_730, signal_729, signal_331}), .c ({signal_752, signal_751, signal_342}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_327 ( .a ({signal_724, signal_723, signal_328}), .b ({signal_728, signal_727, signal_330}), .c ({signal_754, signal_753, signal_343}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_336 ( .a ({signal_752, signal_751, signal_342}), .b ({signal_754, signal_753, signal_343}), .c ({signal_772, signal_771, signal_352}) ) ;

    /* cells in depth 11 */

    /* cells in depth 12 */
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_316 ( .a ({signal_592, signal_591, signal_262}), .b ({signal_724, signal_723, signal_328}), .clk ( clk ), .r ({Fresh[140], Fresh[139], Fresh[138]}), .c ({signal_732, signal_731, signal_332}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_317 ( .a ({signal_554, signal_553, signal_243}), .b ({signal_726, signal_725, signal_329}), .clk ( clk ), .r ({Fresh[143], Fresh[142], Fresh[141]}), .c ({signal_734, signal_733, signal_333}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_318 ( .a ({signal_572, signal_571, signal_252}), .b ({signal_728, signal_727, signal_330}), .clk ( clk ), .r ({Fresh[146], Fresh[145], Fresh[144]}), .c ({signal_736, signal_735, signal_334}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_319 ( .a ({signal_594, signal_593, signal_263}), .b ({signal_730, signal_729, signal_331}), .clk ( clk ), .r ({Fresh[149], Fresh[148], Fresh[147]}), .c ({signal_738, signal_737, signal_335}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_320 ( .a ({signal_586, signal_585, signal_259}), .b ({signal_724, signal_723, signal_328}), .clk ( clk ), .r ({Fresh[152], Fresh[151], Fresh[150]}), .c ({signal_740, signal_739, signal_336}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_321 ( .a ({signal_588, signal_587, signal_260}), .b ({signal_726, signal_725, signal_329}), .clk ( clk ), .r ({Fresh[155], Fresh[154], Fresh[153]}), .c ({signal_742, signal_741, signal_337}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_322 ( .a ({signal_590, signal_589, signal_261}), .b ({signal_728, signal_727, signal_330}), .clk ( clk ), .r ({Fresh[158], Fresh[157], Fresh[156]}), .c ({signal_744, signal_743, signal_338}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_323 ( .a ({signal_574, signal_573, signal_253}), .b ({signal_730, signal_729, signal_331}), .clk ( clk ), .r ({Fresh[161], Fresh[160], Fresh[159]}), .c ({signal_746, signal_745, signal_339}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_328 ( .a ({signal_602, signal_601, signal_267}), .b ({signal_750, signal_749, signal_341}), .clk ( clk ), .r ({Fresh[164], Fresh[163], Fresh[162]}), .c ({signal_756, signal_755, signal_344}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_329 ( .a ({signal_628, signal_627, signal_280}), .b ({signal_748, signal_747, signal_340}), .clk ( clk ), .r ({Fresh[167], Fresh[166], Fresh[165]}), .c ({signal_758, signal_757, signal_345}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_330 ( .a ({signal_604, signal_603, signal_268}), .b ({signal_754, signal_753, signal_343}), .clk ( clk ), .r ({Fresh[170], Fresh[169], Fresh[168]}), .c ({signal_760, signal_759, signal_346}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_331 ( .a ({signal_630, signal_629, signal_281}), .b ({signal_752, signal_751, signal_342}), .clk ( clk ), .r ({Fresh[173], Fresh[172], Fresh[171]}), .c ({signal_762, signal_761, signal_347}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_332 ( .a ({signal_608, signal_607, signal_270}), .b ({signal_750, signal_749, signal_341}), .clk ( clk ), .r ({Fresh[176], Fresh[175], Fresh[174]}), .c ({signal_764, signal_763, signal_348}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_333 ( .a ({signal_606, signal_605, signal_269}), .b ({signal_748, signal_747, signal_340}), .clk ( clk ), .r ({Fresh[179], Fresh[178], Fresh[177]}), .c ({signal_766, signal_765, signal_349}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_334 ( .a ({signal_612, signal_611, signal_272}), .b ({signal_754, signal_753, signal_343}), .clk ( clk ), .r ({Fresh[182], Fresh[181], Fresh[180]}), .c ({signal_768, signal_767, signal_350}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_335 ( .a ({signal_610, signal_609, signal_271}), .b ({signal_752, signal_751, signal_342}), .clk ( clk ), .r ({Fresh[185], Fresh[184], Fresh[183]}), .c ({signal_770, signal_769, signal_351}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_337 ( .a ({signal_646, signal_645, signal_289}), .b ({signal_772, signal_771, signal_352}), .clk ( clk ), .r ({Fresh[188], Fresh[187], Fresh[186]}), .c ({signal_774, signal_773, signal_353}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_338 ( .a ({signal_632, signal_631, signal_282}), .b ({signal_772, signal_771, signal_352}), .clk ( clk ), .r ({Fresh[191], Fresh[190], Fresh[189]}), .c ({signal_776, signal_775, signal_354}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_339 ( .a ({signal_732, signal_731, signal_332}), .b ({signal_756, signal_755, signal_344}), .c ({signal_778, signal_777, signal_355}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_340 ( .a ({signal_734, signal_733, signal_333}), .b ({signal_756, signal_755, signal_344}), .c ({signal_780, signal_779, signal_356}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_341 ( .a ({signal_736, signal_735, signal_334}), .b ({signal_758, signal_757, signal_345}), .c ({signal_782, signal_781, signal_357}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_342 ( .a ({signal_738, signal_737, signal_335}), .b ({signal_758, signal_757, signal_345}), .c ({signal_784, signal_783, signal_358}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_343 ( .a ({signal_760, signal_759, signal_346}), .b ({signal_762, signal_761, signal_347}), .c ({signal_786, signal_785, signal_359}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_344 ( .a ({signal_740, signal_739, signal_336}), .b ({signal_764, signal_763, signal_348}), .c ({signal_788, signal_787, signal_360}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_345 ( .a ({signal_742, signal_741, signal_337}), .b ({signal_764, signal_763, signal_348}), .c ({signal_790, signal_789, signal_361}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_346 ( .a ({signal_744, signal_743, signal_338}), .b ({signal_766, signal_765, signal_349}), .c ({signal_792, signal_791, signal_362}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_347 ( .a ({signal_746, signal_745, signal_339}), .b ({signal_766, signal_765, signal_349}), .c ({signal_794, signal_793, signal_363}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_348 ( .a ({signal_768, signal_767, signal_350}), .b ({signal_770, signal_769, signal_351}), .c ({signal_796, signal_795, signal_364}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_349 ( .a ({signal_780, signal_779, signal_356}), .b ({signal_786, signal_785, signal_359}), .c ({signal_798, signal_797, signal_365}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_350 ( .a ({signal_784, signal_783, signal_358}), .b ({signal_786, signal_785, signal_359}), .c ({signal_800, signal_799, signal_366}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_351 ( .a ({signal_762, signal_761, signal_347}), .b ({signal_774, signal_773, signal_353}), .c ({signal_802, signal_801, signal_367}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_352 ( .a ({signal_790, signal_789, signal_361}), .b ({signal_796, signal_795, signal_364}), .c ({signal_804, signal_803, signal_368}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_353 ( .a ({signal_794, signal_793, signal_363}), .b ({signal_796, signal_795, signal_364}), .c ({signal_806, signal_805, signal_369}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_354 ( .a ({signal_770, signal_769, signal_351}), .b ({signal_776, signal_775, signal_354}), .c ({signal_808, signal_807, signal_370}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_355 ( .a ({signal_804, signal_803, signal_368}), .b ({signal_810, signal_809, signal_371}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_356 ( .a ({signal_798, signal_797, signal_365}), .b ({signal_806, signal_805, signal_369}), .c ({signal_812, signal_811, signal_372}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_357 ( .a ({signal_798, signal_797, signal_365}), .b ({signal_800, signal_799, signal_366}), .c ({signal_814, signal_813, signal_373}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_358 ( .a ({signal_778, signal_777, signal_355}), .b ({signal_802, signal_801, signal_367}), .c ({signal_816, signal_815, signal_374}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_359 ( .a ({signal_782, signal_781, signal_357}), .b ({signal_802, signal_801, signal_367}), .c ({signal_818, signal_817, signal_375}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_360 ( .a ({signal_788, signal_787, signal_360}), .b ({signal_808, signal_807, signal_370}), .c ({signal_820, signal_819, signal_376}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_361 ( .a ({signal_792, signal_791, signal_362}), .b ({signal_808, signal_807, signal_370}), .c ({signal_822, signal_821, signal_377}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_364 ( .a ({signal_818, signal_817, signal_375}), .b ({signal_822, signal_821, signal_377}), .c ({signal_828, signal_827, signal_380}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_365 ( .a ({signal_800, signal_799, signal_366}), .b ({signal_822, signal_821, signal_377}), .c ({signal_830, signal_829, signal_381}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_366 ( .a ({signal_798, signal_797, signal_365}), .b ({signal_822, signal_821, signal_377}), .c ({signal_832, signal_831, signal_382}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_367 ( .a ({signal_816, signal_815, signal_374}), .b ({signal_820, signal_819, signal_376}), .c ({signal_834, signal_833, signal_383}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_368 ( .a ({signal_818, signal_817, signal_375}), .b ({signal_820, signal_819, signal_376}), .c ({signal_836, signal_835, signal_384}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_369 ( .a ({signal_814, signal_813, signal_373}), .b ({signal_822, signal_821, signal_377}), .c ({signal_838, signal_837, signal_385}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_370 ( .a ({signal_828, signal_827, signal_380}), .b ({signal_840, signal_839, signal_386}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_371 ( .a ({signal_830, signal_829, signal_381}), .b ({signal_842, signal_841, signal_387}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_372 ( .a ({signal_832, signal_831, signal_382}), .b ({signal_844, signal_843, signal_388}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_373 ( .a ({signal_836, signal_835, signal_384}), .b ({signal_846, signal_845, signal_389}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_378 ( .a ({signal_800, signal_799, signal_366}), .b ({signal_828, signal_827, signal_380}), .c ({signal_856, signal_855, signal_394}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_379 ( .a ({signal_818, signal_817, signal_375}), .b ({signal_834, signal_833, signal_383}), .c ({signal_858, signal_857, signal_395}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_380 ( .a ({signal_804, signal_803, signal_368}), .b ({signal_836, signal_835, signal_384}), .c ({signal_860, signal_859, signal_396}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_381 ( .a ({signal_858, signal_857, signal_395}), .b ({signal_862, signal_861, signal_397}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_389 ( .a ({signal_816, signal_815, signal_374}), .b ({signal_856, signal_855, signal_394}), .c ({signal_878, signal_877, signal_405}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_390 ( .a ({signal_812, signal_811, signal_372}), .b ({signal_858, signal_857, signal_395}), .c ({signal_880, signal_879, signal_406}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_391 ( .a ({signal_838, signal_837, signal_385}), .b ({signal_860, signal_859, signal_396}), .c ({signal_882, signal_881, signal_407}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_392 ( .a ({signal_814, signal_813, signal_373}), .b ({signal_858, signal_857, signal_395}), .c ({signal_884, signal_883, signal_408}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_393 ( .a ({signal_812, signal_811, signal_372}), .b ({signal_860, signal_859, signal_396}), .c ({signal_886, signal_885, signal_409}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_396 ( .a ({signal_878, signal_877, signal_405}), .b ({signal_892, signal_891, signal_412}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_397 ( .a ({signal_882, signal_881, signal_407}), .b ({signal_894, signal_893, signal_413}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_398 ( .a ({signal_884, signal_883, signal_408}), .b ({signal_896, signal_895, signal_414}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_399 ( .a ({signal_886, signal_885, signal_409}), .b ({signal_898, signal_897, signal_415}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_405 ( .a ({signal_822, signal_821, signal_377}), .b ({signal_880, signal_879, signal_406}), .c ({signal_910, signal_909, signal_420}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_406 ( .a ({signal_804, signal_803, signal_368}), .b ({signal_880, signal_879, signal_406}), .c ({signal_912, signal_911, signal_421}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_408 ( .a ({signal_910, signal_909, signal_420}), .b ({signal_916, signal_915, signal_423}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_409 ( .a ({signal_912, signal_911, signal_421}), .b ({signal_918, signal_917, signal_424}) ) ;

    /* cells in depth 13 */

    /* cells in depth 14 */
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_362 ( .a ({1'b0, 1'b0, signal_193}), .b ({signal_810, signal_809, signal_371}), .clk ( clk ), .r ({Fresh[194], Fresh[193], Fresh[192]}), .c ({signal_824, signal_823, signal_378}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_363 ( .a ({1'b0, 1'b0, 1'b1}), .b ({signal_812, signal_811, signal_372}), .clk ( clk ), .r ({Fresh[197], Fresh[196], Fresh[195]}), .c ({signal_826, signal_825, signal_379}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_374 ( .a ({signal_824, signal_823, signal_378}), .b ({signal_848, signal_847, signal_390}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_375 ( .a ({signal_826, signal_825, signal_379}), .b ({signal_850, signal_849, signal_391}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_376 ( .a ({1'b0, 1'b0, 1'b1}), .b ({signal_838, signal_837, signal_385}), .clk ( clk ), .r ({Fresh[200], Fresh[199], Fresh[198]}), .c ({signal_852, signal_851, signal_392}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_377 ( .a ({1'b0, 1'b0, 1'b1}), .b ({signal_834, signal_833, signal_383}), .clk ( clk ), .r ({Fresh[203], Fresh[202], Fresh[201]}), .c ({signal_854, signal_853, signal_393}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_382 ( .a ({signal_852, signal_851, signal_392}), .b ({signal_864, signal_863, signal_398}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_383 ( .a ({signal_854, signal_853, signal_393}), .b ({signal_866, signal_865, signal_399}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_384 ( .a ({1'b0, 1'b0, signal_193}), .b ({signal_842, signal_841, signal_387}), .clk ( clk ), .r ({Fresh[206], Fresh[205], Fresh[204]}), .c ({signal_868, signal_867, signal_400}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_385 ( .a ({1'b0, 1'b0, 1'b1}), .b ({signal_846, signal_845, signal_389}), .clk ( clk ), .r ({Fresh[209], Fresh[208], Fresh[207]}), .c ({signal_870, signal_869, signal_401}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_386 ( .a ({1'b0, 1'b0, signal_193}), .b ({signal_844, signal_843, signal_388}), .clk ( clk ), .r ({Fresh[212], Fresh[211], Fresh[210]}), .c ({signal_872, signal_871, signal_402}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_387 ( .a ({1'b0, 1'b0, signal_193}), .b ({signal_840, signal_839, signal_386}), .clk ( clk ), .r ({Fresh[215], Fresh[214], Fresh[213]}), .c ({signal_874, signal_873, signal_403}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_388 ( .a ({1'b0, 1'b0, 1'b1}), .b ({signal_856, signal_855, signal_394}), .clk ( clk ), .r ({Fresh[218], Fresh[217], Fresh[216]}), .c ({signal_876, signal_875, signal_404}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_394 ( .a ({signal_868, signal_867, signal_400}), .b ({signal_888, signal_887, signal_410}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_395 ( .a ({signal_870, signal_869, signal_401}), .b ({signal_890, signal_889, signal_411}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_400 ( .a ({signal_872, signal_871, signal_402}), .b ({signal_900, signal_899, signal_416}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_401 ( .a ({signal_874, signal_873, signal_403}), .b ({signal_902, signal_901, signal_417}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_402 ( .a ({signal_876, signal_875, signal_404}), .b ({signal_904, signal_903, signal_418}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_404 ( .a ({1'b0, 1'b0, 1'b1}), .b ({signal_862, signal_861, signal_397}), .clk ( clk ), .r ({Fresh[221], Fresh[220], Fresh[219]}), .c ({signal_908, signal_907, signal_419}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_407 ( .a ({signal_908, signal_907, signal_419}), .b ({signal_914, signal_913, signal_422}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_412 ( .a ({1'b0, 1'b0, signal_193}), .b ({signal_894, signal_893, signal_413}), .clk ( clk ), .r ({Fresh[224], Fresh[223], Fresh[222]}), .c ({signal_924, signal_923, signal_425}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_413 ( .a ({1'b0, 1'b0, 1'b1}), .b ({signal_896, signal_895, signal_414}), .clk ( clk ), .r ({Fresh[227], Fresh[226], Fresh[225]}), .c ({signal_926, signal_925, signal_426}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_414 ( .a ({1'b0, 1'b0, signal_193}), .b ({signal_892, signal_891, signal_412}), .clk ( clk ), .r ({Fresh[230], Fresh[229], Fresh[228]}), .c ({signal_928, signal_927, signal_427}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_415 ( .a ({1'b0, 1'b0, 1'b1}), .b ({signal_898, signal_897, signal_415}), .clk ( clk ), .r ({Fresh[233], Fresh[232], Fresh[231]}), .c ({signal_930, signal_929, signal_428}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_416 ( .a ({signal_924, signal_923, signal_425}), .b ({signal_932, signal_931, signal_429}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_417 ( .a ({signal_926, signal_925, signal_426}), .b ({signal_934, signal_933, signal_430}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_418 ( .a ({signal_928, signal_927, signal_427}), .b ({signal_936, signal_935, signal_431}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_419 ( .a ({signal_930, signal_929, signal_428}), .b ({signal_938, signal_937, signal_432}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_421 ( .a ({1'b0, 1'b0, signal_193}), .b ({signal_916, signal_915, signal_423}), .clk ( clk ), .r ({Fresh[236], Fresh[235], Fresh[234]}), .c ({signal_942, signal_941, signal_433}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_422 ( .a ({1'b0, 1'b0, signal_193}), .b ({signal_918, signal_917, signal_424}), .clk ( clk ), .r ({Fresh[239], Fresh[238], Fresh[237]}), .c ({signal_944, signal_943, signal_434}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_423 ( .a ({signal_942, signal_941, signal_433}), .b ({signal_946, signal_945, signal_435}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_424 ( .a ({signal_944, signal_943, signal_434}), .b ({signal_948, signal_947, signal_436}) ) ;

    /* cells in depth 15 */

    /* cells in depth 16 */
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_403 ( .a ({signal_848, signal_847, signal_390}), .b ({signal_864, signal_863, signal_398}), .clk ( clk ), .r ({Fresh[242], Fresh[241], Fresh[240]}), .c ({signal_906, signal_905, signal_167}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_410 ( .a ({signal_888, signal_887, signal_410}), .b ({signal_890, signal_889, signal_411}), .clk ( clk ), .r ({Fresh[245], Fresh[244], Fresh[243]}), .c ({signal_920, signal_919, signal_160}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_411 ( .a ({signal_902, signal_901, signal_417}), .b ({signal_904, signal_903, signal_418}), .clk ( clk ), .r ({Fresh[248], Fresh[247], Fresh[246]}), .c ({signal_922, signal_921, signal_166}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_420 ( .a ({signal_900, signal_899, signal_416}), .b ({signal_914, signal_913, signal_422}), .clk ( clk ), .r ({Fresh[251], Fresh[250], Fresh[249]}), .c ({signal_940, signal_939, signal_163}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_425 ( .a ({signal_932, signal_931, signal_429}), .b ({signal_934, signal_933, signal_430}), .clk ( clk ), .r ({Fresh[254], Fresh[253], Fresh[252]}), .c ({signal_950, signal_949, signal_164}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_426 ( .a ({signal_936, signal_935, signal_431}), .b ({signal_938, signal_937, signal_432}), .clk ( clk ), .r ({Fresh[257], Fresh[256], Fresh[255]}), .c ({signal_952, signal_951, signal_165}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_427 ( .a ({signal_946, signal_945, signal_435}), .b ({signal_866, signal_865, signal_399}), .clk ( clk ), .r ({Fresh[260], Fresh[259], Fresh[258]}), .c ({signal_954, signal_953, signal_161}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_428 ( .a ({signal_948, signal_947, signal_436}), .b ({signal_850, signal_849, signal_391}), .clk ( clk ), .r ({Fresh[263], Fresh[262], Fresh[261]}), .c ({signal_956, signal_955, signal_162}) ) ;

    /* register cells */
    reg_masked #(.security_order(2), .pipeline(0)) cell_0 ( .clk ( signal_1238 ), .D ({signal_920, signal_919, signal_160}), .Q ({Y_s2[7], Y_s1[7], Y_s0[7]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) cell_1 ( .clk ( signal_1238 ), .D ({signal_954, signal_953, signal_161}), .Q ({Y_s2[6], Y_s1[6], Y_s0[6]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) cell_2 ( .clk ( signal_1238 ), .D ({signal_956, signal_955, signal_162}), .Q ({Y_s2[5], Y_s1[5], Y_s0[5]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) cell_3 ( .clk ( signal_1238 ), .D ({signal_940, signal_939, signal_163}), .Q ({Y_s2[4], Y_s1[4], Y_s0[4]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) cell_4 ( .clk ( signal_1238 ), .D ({signal_950, signal_949, signal_164}), .Q ({Y_s2[3], Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) cell_5 ( .clk ( signal_1238 ), .D ({signal_952, signal_951, signal_165}), .Q ({Y_s2[2], Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) cell_6 ( .clk ( signal_1238 ), .D ({signal_922, signal_921, signal_166}), .Q ({Y_s2[1], Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) cell_7 ( .clk ( signal_1238 ), .D ({signal_906, signal_905, signal_167}), .Q ({Y_s2[0], Y_s1[0], Y_s0[0]}) ) ;
endmodule
