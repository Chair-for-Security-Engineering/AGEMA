/* modified netlist. Source: module sbox in file ../sbox_lookup/sbox.v */
/* 12 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 13 register stage(s) in total */

module sbox_HPC2_AIG_Pipeline_d3 (SI_s0, clk, SI_s1, SI_s2, SI_s3, Fresh, SO_s0, SO_s1, SO_s2, SO_s3);
    input [3:0] SI_s0 ;
    input clk ;
    input [3:0] SI_s1 ;
    input [3:0] SI_s2 ;
    input [3:0] SI_s3 ;
    input [101:0] Fresh ;
    output [3:0] SO_s0 ;
    output [3:0] SO_s1 ;
    output [3:0] SO_s2 ;
    output [3:0] SO_s3 ;
    wire signal_15 ;
    wire signal_16 ;
    wire signal_17 ;
    wire signal_18 ;
    wire signal_34 ;
    wire signal_35 ;
    wire signal_36 ;
    wire signal_37 ;
    wire signal_38 ;
    wire signal_39 ;
    wire signal_40 ;
    wire signal_41 ;
    wire signal_42 ;
    wire signal_43 ;
    wire signal_44 ;
    wire signal_45 ;
    wire signal_46 ;
    wire signal_47 ;
    wire signal_48 ;
    wire signal_49 ;
    wire signal_50 ;
    wire signal_51 ;
    wire signal_52 ;
    wire signal_53 ;
    wire signal_54 ;
    wire signal_55 ;
    wire signal_56 ;
    wire signal_57 ;
    wire signal_58 ;
    wire signal_59 ;
    wire signal_60 ;
    wire signal_61 ;
    wire signal_62 ;
    wire signal_63 ;
    wire signal_64 ;
    wire signal_68 ;
    wire signal_69 ;
    wire signal_70 ;
    wire signal_74 ;
    wire signal_75 ;
    wire signal_76 ;
    wire signal_80 ;
    wire signal_81 ;
    wire signal_82 ;
    wire signal_86 ;
    wire signal_87 ;
    wire signal_88 ;
    wire signal_89 ;
    wire signal_90 ;
    wire signal_91 ;
    wire signal_92 ;
    wire signal_93 ;
    wire signal_94 ;
    wire signal_95 ;
    wire signal_96 ;
    wire signal_97 ;
    wire signal_98 ;
    wire signal_99 ;
    wire signal_100 ;
    wire signal_101 ;
    wire signal_102 ;
    wire signal_103 ;
    wire signal_104 ;
    wire signal_105 ;
    wire signal_106 ;
    wire signal_107 ;
    wire signal_108 ;
    wire signal_109 ;
    wire signal_110 ;
    wire signal_111 ;
    wire signal_112 ;
    wire signal_113 ;
    wire signal_114 ;
    wire signal_115 ;
    wire signal_116 ;
    wire signal_117 ;
    wire signal_118 ;
    wire signal_119 ;
    wire signal_120 ;
    wire signal_121 ;
    wire signal_122 ;
    wire signal_123 ;
    wire signal_124 ;
    wire signal_125 ;
    wire signal_126 ;
    wire signal_127 ;
    wire signal_128 ;
    wire signal_129 ;
    wire signal_130 ;
    wire signal_131 ;
    wire signal_132 ;
    wire signal_133 ;
    wire signal_134 ;
    wire signal_135 ;
    wire signal_136 ;
    wire signal_137 ;
    wire signal_138 ;
    wire signal_139 ;
    wire signal_140 ;
    wire signal_141 ;
    wire signal_142 ;
    wire signal_143 ;
    wire signal_144 ;
    wire signal_145 ;
    wire signal_146 ;
    wire signal_147 ;
    wire signal_148 ;
    wire signal_149 ;
    wire signal_150 ;
    wire signal_151 ;
    wire signal_152 ;
    wire signal_153 ;
    wire signal_154 ;
    wire signal_155 ;
    wire signal_156 ;
    wire signal_157 ;
    wire signal_158 ;
    wire signal_159 ;
    wire signal_160 ;
    wire signal_161 ;
    wire signal_162 ;
    wire signal_163 ;
    wire signal_164 ;
    wire signal_165 ;
    wire signal_166 ;
    wire signal_167 ;
    wire signal_168 ;
    wire signal_169 ;
    wire signal_170 ;
    wire signal_171 ;
    wire signal_172 ;
    wire signal_173 ;
    wire signal_174 ;
    wire signal_175 ;
    wire signal_176 ;
    wire signal_177 ;
    wire signal_178 ;
    wire signal_179 ;
    wire signal_180 ;
    wire signal_181 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_352 ;
    wire signal_353 ;
    wire signal_354 ;
    wire signal_355 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_359 ;
    wire signal_360 ;
    wire signal_361 ;
    wire signal_362 ;
    wire signal_363 ;
    wire signal_364 ;
    wire signal_365 ;
    wire signal_366 ;
    wire signal_367 ;
    wire signal_368 ;
    wire signal_369 ;
    wire signal_370 ;
    wire signal_371 ;
    wire signal_372 ;
    wire signal_373 ;
    wire signal_374 ;
    wire signal_375 ;
    wire signal_376 ;
    wire signal_377 ;
    wire signal_378 ;
    wire signal_379 ;
    wire signal_380 ;
    wire signal_381 ;
    wire signal_382 ;
    wire signal_383 ;
    wire signal_384 ;
    wire signal_385 ;
    wire signal_386 ;
    wire signal_387 ;
    wire signal_388 ;
    wire signal_389 ;
    wire signal_390 ;
    wire signal_391 ;
    wire signal_392 ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_415 ;
    wire signal_416 ;
    wire signal_417 ;
    wire signal_418 ;
    wire signal_419 ;
    wire signal_420 ;
    wire signal_421 ;
    wire signal_422 ;
    wire signal_423 ;
    wire signal_424 ;
    wire signal_425 ;
    wire signal_426 ;
    wire signal_427 ;
    wire signal_428 ;
    wire signal_429 ;
    wire signal_430 ;
    wire signal_431 ;
    wire signal_432 ;
    wire signal_433 ;
    wire signal_434 ;
    wire signal_435 ;
    wire signal_436 ;
    wire signal_437 ;
    wire signal_438 ;
    wire signal_439 ;
    wire signal_440 ;
    wire signal_441 ;
    wire signal_442 ;
    wire signal_443 ;
    wire signal_444 ;
    wire signal_445 ;
    wire signal_446 ;
    wire signal_447 ;
    wire signal_448 ;
    wire signal_449 ;
    wire signal_450 ;
    wire signal_451 ;
    wire signal_452 ;
    wire signal_453 ;
    wire signal_454 ;
    wire signal_455 ;
    wire signal_456 ;
    wire signal_457 ;
    wire signal_458 ;
    wire signal_459 ;
    wire signal_460 ;
    wire signal_461 ;
    wire signal_462 ;
    wire signal_463 ;
    wire signal_464 ;
    wire signal_465 ;
    wire signal_466 ;
    wire signal_467 ;
    wire signal_468 ;
    wire signal_469 ;
    wire signal_470 ;
    wire signal_471 ;
    wire signal_472 ;
    wire signal_473 ;
    wire signal_474 ;
    wire signal_475 ;
    wire signal_476 ;
    wire signal_477 ;
    wire signal_478 ;
    wire signal_479 ;
    wire signal_480 ;
    wire signal_481 ;
    wire signal_482 ;
    wire signal_483 ;
    wire signal_484 ;
    wire signal_485 ;
    wire signal_486 ;
    wire signal_487 ;
    wire signal_488 ;
    wire signal_489 ;
    wire signal_490 ;
    wire signal_491 ;
    wire signal_492 ;
    wire signal_493 ;
    wire signal_494 ;
    wire signal_495 ;
    wire signal_496 ;
    wire signal_497 ;
    wire signal_498 ;
    wire signal_499 ;
    wire signal_500 ;
    wire signal_501 ;
    wire signal_502 ;
    wire signal_503 ;
    wire signal_504 ;
    wire signal_505 ;
    wire signal_506 ;
    wire signal_507 ;
    wire signal_508 ;
    wire signal_509 ;
    wire signal_510 ;
    wire signal_511 ;
    wire signal_512 ;
    wire signal_513 ;
    wire signal_514 ;
    wire signal_515 ;
    wire signal_516 ;
    wire signal_517 ;
    wire signal_518 ;
    wire signal_519 ;

    /* cells in depth 0 */
    not_masked #(.security_order(3), .pipeline(1)) cell_23 ( .a ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_70, signal_69, signal_68, signal_34}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_24 ( .a ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_76, signal_75, signal_74, signal_35}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_25 ( .a ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({signal_82, signal_81, signal_80, signal_36}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_26 ( .a ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({signal_88, signal_87, signal_86, signal_37}) ) ;

    /* cells in depth 1 */
    buf_clk cell_58 ( .C ( clk ), .D ( SI_s0[3] ), .Q ( signal_296 ) ) ;
    buf_clk cell_60 ( .C ( clk ), .D ( SI_s1[3] ), .Q ( signal_298 ) ) ;
    buf_clk cell_62 ( .C ( clk ), .D ( SI_s2[3] ), .Q ( signal_300 ) ) ;
    buf_clk cell_64 ( .C ( clk ), .D ( SI_s3[3] ), .Q ( signal_302 ) ) ;
    buf_clk cell_66 ( .C ( clk ), .D ( SI_s0[0] ), .Q ( signal_304 ) ) ;
    buf_clk cell_68 ( .C ( clk ), .D ( SI_s1[0] ), .Q ( signal_306 ) ) ;
    buf_clk cell_70 ( .C ( clk ), .D ( SI_s2[0] ), .Q ( signal_308 ) ) ;
    buf_clk cell_72 ( .C ( clk ), .D ( SI_s3[0] ), .Q ( signal_310 ) ) ;
    buf_clk cell_74 ( .C ( clk ), .D ( SI_s0[2] ), .Q ( signal_312 ) ) ;
    buf_clk cell_76 ( .C ( clk ), .D ( SI_s1[2] ), .Q ( signal_314 ) ) ;
    buf_clk cell_78 ( .C ( clk ), .D ( SI_s2[2] ), .Q ( signal_316 ) ) ;
    buf_clk cell_80 ( .C ( clk ), .D ( SI_s3[2] ), .Q ( signal_318 ) ) ;
    buf_clk cell_82 ( .C ( clk ), .D ( signal_34 ), .Q ( signal_320 ) ) ;
    buf_clk cell_84 ( .C ( clk ), .D ( signal_68 ), .Q ( signal_322 ) ) ;
    buf_clk cell_86 ( .C ( clk ), .D ( signal_69 ), .Q ( signal_324 ) ) ;
    buf_clk cell_88 ( .C ( clk ), .D ( signal_70 ), .Q ( signal_326 ) ) ;
    buf_clk cell_90 ( .C ( clk ), .D ( signal_36 ), .Q ( signal_328 ) ) ;
    buf_clk cell_92 ( .C ( clk ), .D ( signal_80 ), .Q ( signal_330 ) ) ;
    buf_clk cell_94 ( .C ( clk ), .D ( signal_81 ), .Q ( signal_332 ) ) ;
    buf_clk cell_96 ( .C ( clk ), .D ( signal_82 ), .Q ( signal_334 ) ) ;
    buf_clk cell_122 ( .C ( clk ), .D ( SI_s0[1] ), .Q ( signal_360 ) ) ;
    buf_clk cell_128 ( .C ( clk ), .D ( SI_s1[1] ), .Q ( signal_366 ) ) ;
    buf_clk cell_134 ( .C ( clk ), .D ( SI_s2[1] ), .Q ( signal_372 ) ) ;
    buf_clk cell_140 ( .C ( clk ), .D ( SI_s3[1] ), .Q ( signal_378 ) ) ;

    /* cells in depth 2 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_27 ( .a ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({signal_91, signal_90, signal_89, signal_38}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_28 ( .a ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6]}), .c ({signal_94, signal_93, signal_92, signal_39}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_29 ( .a ({signal_91, signal_90, signal_89, signal_38}), .b ({signal_97, signal_96, signal_95, signal_40}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_30 ( .a ({signal_94, signal_93, signal_92, signal_39}), .b ({signal_100, signal_99, signal_98, signal_41}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_31 ( .a ({signal_76, signal_75, signal_74, signal_35}), .b ({signal_82, signal_81, signal_80, signal_36}), .clk ( clk ), .r ({Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({signal_103, signal_102, signal_101, signal_42}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_32 ( .a ({signal_70, signal_69, signal_68, signal_34}), .b ({signal_88, signal_87, signal_86, signal_37}), .clk ( clk ), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18]}), .c ({signal_106, signal_105, signal_104, signal_43}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_33 ( .a ({signal_76, signal_75, signal_74, signal_35}), .b ({signal_88, signal_87, signal_86, signal_37}), .clk ( clk ), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24]}), .c ({signal_109, signal_108, signal_107, signal_44}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_34 ( .a ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_76, signal_75, signal_74, signal_35}), .clk ( clk ), .r ({Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({signal_112, signal_111, signal_110, signal_45}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_35 ( .a ({signal_70, signal_69, signal_68, signal_34}), .b ({signal_76, signal_75, signal_74, signal_35}), .clk ( clk ), .r ({Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36]}), .c ({signal_115, signal_114, signal_113, signal_46}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_36 ( .a ({signal_109, signal_108, signal_107, signal_44}), .b ({signal_118, signal_117, signal_116, signal_47}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_39 ( .a ({signal_303, signal_301, signal_299, signal_297}), .b ({signal_103, signal_102, signal_101, signal_42}), .c ({signal_127, signal_126, signal_125, signal_16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_40 ( .a ({signal_311, signal_309, signal_307, signal_305}), .b ({signal_112, signal_111, signal_110, signal_45}), .c ({signal_130, signal_129, signal_128, signal_50}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_41 ( .a ({signal_311, signal_309, signal_307, signal_305}), .b ({signal_115, signal_114, signal_113, signal_46}), .c ({signal_133, signal_132, signal_131, signal_15}) ) ;
    buf_clk cell_59 ( .C ( clk ), .D ( signal_296 ), .Q ( signal_297 ) ) ;
    buf_clk cell_61 ( .C ( clk ), .D ( signal_298 ), .Q ( signal_299 ) ) ;
    buf_clk cell_63 ( .C ( clk ), .D ( signal_300 ), .Q ( signal_301 ) ) ;
    buf_clk cell_65 ( .C ( clk ), .D ( signal_302 ), .Q ( signal_303 ) ) ;
    buf_clk cell_67 ( .C ( clk ), .D ( signal_304 ), .Q ( signal_305 ) ) ;
    buf_clk cell_69 ( .C ( clk ), .D ( signal_306 ), .Q ( signal_307 ) ) ;
    buf_clk cell_71 ( .C ( clk ), .D ( signal_308 ), .Q ( signal_309 ) ) ;
    buf_clk cell_73 ( .C ( clk ), .D ( signal_310 ), .Q ( signal_311 ) ) ;
    buf_clk cell_75 ( .C ( clk ), .D ( signal_312 ), .Q ( signal_313 ) ) ;
    buf_clk cell_77 ( .C ( clk ), .D ( signal_314 ), .Q ( signal_315 ) ) ;
    buf_clk cell_79 ( .C ( clk ), .D ( signal_316 ), .Q ( signal_317 ) ) ;
    buf_clk cell_81 ( .C ( clk ), .D ( signal_318 ), .Q ( signal_319 ) ) ;
    buf_clk cell_83 ( .C ( clk ), .D ( signal_320 ), .Q ( signal_321 ) ) ;
    buf_clk cell_85 ( .C ( clk ), .D ( signal_322 ), .Q ( signal_323 ) ) ;
    buf_clk cell_87 ( .C ( clk ), .D ( signal_324 ), .Q ( signal_325 ) ) ;
    buf_clk cell_89 ( .C ( clk ), .D ( signal_326 ), .Q ( signal_327 ) ) ;
    buf_clk cell_91 ( .C ( clk ), .D ( signal_328 ), .Q ( signal_329 ) ) ;
    buf_clk cell_93 ( .C ( clk ), .D ( signal_330 ), .Q ( signal_331 ) ) ;
    buf_clk cell_95 ( .C ( clk ), .D ( signal_332 ), .Q ( signal_333 ) ) ;
    buf_clk cell_97 ( .C ( clk ), .D ( signal_334 ), .Q ( signal_335 ) ) ;
    buf_clk cell_123 ( .C ( clk ), .D ( signal_360 ), .Q ( signal_361 ) ) ;
    buf_clk cell_129 ( .C ( clk ), .D ( signal_366 ), .Q ( signal_367 ) ) ;
    buf_clk cell_135 ( .C ( clk ), .D ( signal_372 ), .Q ( signal_373 ) ) ;
    buf_clk cell_141 ( .C ( clk ), .D ( signal_378 ), .Q ( signal_379 ) ) ;

    /* cells in depth 3 */
    buf_clk cell_98 ( .C ( clk ), .D ( signal_40 ), .Q ( signal_336 ) ) ;
    buf_clk cell_100 ( .C ( clk ), .D ( signal_95 ), .Q ( signal_338 ) ) ;
    buf_clk cell_102 ( .C ( clk ), .D ( signal_96 ), .Q ( signal_340 ) ) ;
    buf_clk cell_104 ( .C ( clk ), .D ( signal_97 ), .Q ( signal_342 ) ) ;
    buf_clk cell_106 ( .C ( clk ), .D ( signal_329 ), .Q ( signal_344 ) ) ;
    buf_clk cell_108 ( .C ( clk ), .D ( signal_331 ), .Q ( signal_346 ) ) ;
    buf_clk cell_110 ( .C ( clk ), .D ( signal_333 ), .Q ( signal_348 ) ) ;
    buf_clk cell_112 ( .C ( clk ), .D ( signal_335 ), .Q ( signal_350 ) ) ;
    buf_clk cell_114 ( .C ( clk ), .D ( signal_41 ), .Q ( signal_352 ) ) ;
    buf_clk cell_116 ( .C ( clk ), .D ( signal_98 ), .Q ( signal_354 ) ) ;
    buf_clk cell_118 ( .C ( clk ), .D ( signal_99 ), .Q ( signal_356 ) ) ;
    buf_clk cell_120 ( .C ( clk ), .D ( signal_100 ), .Q ( signal_358 ) ) ;
    buf_clk cell_124 ( .C ( clk ), .D ( signal_361 ), .Q ( signal_362 ) ) ;
    buf_clk cell_130 ( .C ( clk ), .D ( signal_367 ), .Q ( signal_368 ) ) ;
    buf_clk cell_136 ( .C ( clk ), .D ( signal_373 ), .Q ( signal_374 ) ) ;
    buf_clk cell_142 ( .C ( clk ), .D ( signal_379 ), .Q ( signal_380 ) ) ;
    buf_clk cell_178 ( .C ( clk ), .D ( signal_15 ), .Q ( signal_416 ) ) ;
    buf_clk cell_188 ( .C ( clk ), .D ( signal_131 ), .Q ( signal_426 ) ) ;
    buf_clk cell_198 ( .C ( clk ), .D ( signal_132 ), .Q ( signal_436 ) ) ;
    buf_clk cell_208 ( .C ( clk ), .D ( signal_133 ), .Q ( signal_446 ) ) ;
    buf_clk cell_218 ( .C ( clk ), .D ( signal_16 ), .Q ( signal_456 ) ) ;
    buf_clk cell_228 ( .C ( clk ), .D ( signal_125 ), .Q ( signal_466 ) ) ;
    buf_clk cell_238 ( .C ( clk ), .D ( signal_126 ), .Q ( signal_476 ) ) ;
    buf_clk cell_248 ( .C ( clk ), .D ( signal_127 ), .Q ( signal_486 ) ) ;

    /* cells in depth 4 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_37 ( .a ({signal_319, signal_317, signal_315, signal_313}), .b ({signal_106, signal_105, signal_104, signal_43}), .clk ( clk ), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42]}), .c ({signal_121, signal_120, signal_119, signal_48}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_38 ( .a ({signal_303, signal_301, signal_299, signal_297}), .b ({signal_109, signal_108, signal_107, signal_44}), .clk ( clk ), .r ({Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .c ({signal_124, signal_123, signal_122, signal_49}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_42 ( .a ({signal_121, signal_120, signal_119, signal_48}), .b ({signal_136, signal_135, signal_134, signal_51}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_43 ( .a ({signal_124, signal_123, signal_122, signal_49}), .b ({signal_139, signal_138, signal_137, signal_52}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_44 ( .a ({signal_327, signal_325, signal_323, signal_321}), .b ({signal_118, signal_117, signal_116, signal_47}), .clk ( clk ), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54]}), .c ({signal_142, signal_141, signal_140, signal_53}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_45 ( .a ({signal_335, signal_333, signal_331, signal_329}), .b ({signal_130, signal_129, signal_128, signal_50}), .clk ( clk ), .r ({Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({signal_145, signal_144, signal_143, signal_54}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_46 ( .a ({signal_145, signal_144, signal_143, signal_54}), .b ({signal_148, signal_147, signal_146, signal_55}) ) ;
    buf_clk cell_99 ( .C ( clk ), .D ( signal_336 ), .Q ( signal_337 ) ) ;
    buf_clk cell_101 ( .C ( clk ), .D ( signal_338 ), .Q ( signal_339 ) ) ;
    buf_clk cell_103 ( .C ( clk ), .D ( signal_340 ), .Q ( signal_341 ) ) ;
    buf_clk cell_105 ( .C ( clk ), .D ( signal_342 ), .Q ( signal_343 ) ) ;
    buf_clk cell_107 ( .C ( clk ), .D ( signal_344 ), .Q ( signal_345 ) ) ;
    buf_clk cell_109 ( .C ( clk ), .D ( signal_346 ), .Q ( signal_347 ) ) ;
    buf_clk cell_111 ( .C ( clk ), .D ( signal_348 ), .Q ( signal_349 ) ) ;
    buf_clk cell_113 ( .C ( clk ), .D ( signal_350 ), .Q ( signal_351 ) ) ;
    buf_clk cell_115 ( .C ( clk ), .D ( signal_352 ), .Q ( signal_353 ) ) ;
    buf_clk cell_117 ( .C ( clk ), .D ( signal_354 ), .Q ( signal_355 ) ) ;
    buf_clk cell_119 ( .C ( clk ), .D ( signal_356 ), .Q ( signal_357 ) ) ;
    buf_clk cell_121 ( .C ( clk ), .D ( signal_358 ), .Q ( signal_359 ) ) ;
    buf_clk cell_125 ( .C ( clk ), .D ( signal_362 ), .Q ( signal_363 ) ) ;
    buf_clk cell_131 ( .C ( clk ), .D ( signal_368 ), .Q ( signal_369 ) ) ;
    buf_clk cell_137 ( .C ( clk ), .D ( signal_374 ), .Q ( signal_375 ) ) ;
    buf_clk cell_143 ( .C ( clk ), .D ( signal_380 ), .Q ( signal_381 ) ) ;
    buf_clk cell_179 ( .C ( clk ), .D ( signal_416 ), .Q ( signal_417 ) ) ;
    buf_clk cell_189 ( .C ( clk ), .D ( signal_426 ), .Q ( signal_427 ) ) ;
    buf_clk cell_199 ( .C ( clk ), .D ( signal_436 ), .Q ( signal_437 ) ) ;
    buf_clk cell_209 ( .C ( clk ), .D ( signal_446 ), .Q ( signal_447 ) ) ;
    buf_clk cell_219 ( .C ( clk ), .D ( signal_456 ), .Q ( signal_457 ) ) ;
    buf_clk cell_229 ( .C ( clk ), .D ( signal_466 ), .Q ( signal_467 ) ) ;
    buf_clk cell_239 ( .C ( clk ), .D ( signal_476 ), .Q ( signal_477 ) ) ;
    buf_clk cell_249 ( .C ( clk ), .D ( signal_486 ), .Q ( signal_487 ) ) ;

    /* cells in depth 5 */
    buf_clk cell_126 ( .C ( clk ), .D ( signal_363 ), .Q ( signal_364 ) ) ;
    buf_clk cell_132 ( .C ( clk ), .D ( signal_369 ), .Q ( signal_370 ) ) ;
    buf_clk cell_138 ( .C ( clk ), .D ( signal_375 ), .Q ( signal_376 ) ) ;
    buf_clk cell_144 ( .C ( clk ), .D ( signal_381 ), .Q ( signal_382 ) ) ;
    buf_clk cell_154 ( .C ( clk ), .D ( signal_52 ), .Q ( signal_392 ) ) ;
    buf_clk cell_160 ( .C ( clk ), .D ( signal_137 ), .Q ( signal_398 ) ) ;
    buf_clk cell_166 ( .C ( clk ), .D ( signal_138 ), .Q ( signal_404 ) ) ;
    buf_clk cell_172 ( .C ( clk ), .D ( signal_139 ), .Q ( signal_410 ) ) ;
    buf_clk cell_180 ( .C ( clk ), .D ( signal_417 ), .Q ( signal_418 ) ) ;
    buf_clk cell_190 ( .C ( clk ), .D ( signal_427 ), .Q ( signal_428 ) ) ;
    buf_clk cell_200 ( .C ( clk ), .D ( signal_437 ), .Q ( signal_438 ) ) ;
    buf_clk cell_210 ( .C ( clk ), .D ( signal_447 ), .Q ( signal_448 ) ) ;
    buf_clk cell_220 ( .C ( clk ), .D ( signal_457 ), .Q ( signal_458 ) ) ;
    buf_clk cell_230 ( .C ( clk ), .D ( signal_467 ), .Q ( signal_468 ) ) ;
    buf_clk cell_240 ( .C ( clk ), .D ( signal_477 ), .Q ( signal_478 ) ) ;
    buf_clk cell_250 ( .C ( clk ), .D ( signal_487 ), .Q ( signal_488 ) ) ;

    /* cells in depth 6 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_47 ( .a ({signal_343, signal_341, signal_339, signal_337}), .b ({signal_142, signal_141, signal_140, signal_53}), .clk ( clk ), .r ({Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66]}), .c ({signal_151, signal_150, signal_149, signal_56}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_48 ( .a ({signal_351, signal_349, signal_347, signal_345}), .b ({signal_136, signal_135, signal_134, signal_51}), .clk ( clk ), .r ({Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72]}), .c ({signal_154, signal_153, signal_152, signal_57}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_49 ( .a ({signal_154, signal_153, signal_152, signal_57}), .b ({signal_157, signal_156, signal_155, signal_58}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_50 ( .a ({signal_148, signal_147, signal_146, signal_55}), .b ({signal_359, signal_357, signal_355, signal_353}), .clk ( clk ), .r ({Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78]}), .c ({signal_160, signal_159, signal_158, signal_59}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_52 ( .a ({signal_160, signal_159, signal_158, signal_59}), .b ({signal_166, signal_165, signal_164, signal_17}) ) ;
    buf_clk cell_127 ( .C ( clk ), .D ( signal_364 ), .Q ( signal_365 ) ) ;
    buf_clk cell_133 ( .C ( clk ), .D ( signal_370 ), .Q ( signal_371 ) ) ;
    buf_clk cell_139 ( .C ( clk ), .D ( signal_376 ), .Q ( signal_377 ) ) ;
    buf_clk cell_145 ( .C ( clk ), .D ( signal_382 ), .Q ( signal_383 ) ) ;
    buf_clk cell_155 ( .C ( clk ), .D ( signal_392 ), .Q ( signal_393 ) ) ;
    buf_clk cell_161 ( .C ( clk ), .D ( signal_398 ), .Q ( signal_399 ) ) ;
    buf_clk cell_167 ( .C ( clk ), .D ( signal_404 ), .Q ( signal_405 ) ) ;
    buf_clk cell_173 ( .C ( clk ), .D ( signal_410 ), .Q ( signal_411 ) ) ;
    buf_clk cell_181 ( .C ( clk ), .D ( signal_418 ), .Q ( signal_419 ) ) ;
    buf_clk cell_191 ( .C ( clk ), .D ( signal_428 ), .Q ( signal_429 ) ) ;
    buf_clk cell_201 ( .C ( clk ), .D ( signal_438 ), .Q ( signal_439 ) ) ;
    buf_clk cell_211 ( .C ( clk ), .D ( signal_448 ), .Q ( signal_449 ) ) ;
    buf_clk cell_221 ( .C ( clk ), .D ( signal_458 ), .Q ( signal_459 ) ) ;
    buf_clk cell_231 ( .C ( clk ), .D ( signal_468 ), .Q ( signal_469 ) ) ;
    buf_clk cell_241 ( .C ( clk ), .D ( signal_478 ), .Q ( signal_479 ) ) ;
    buf_clk cell_251 ( .C ( clk ), .D ( signal_488 ), .Q ( signal_489 ) ) ;

    /* cells in depth 7 */
    buf_clk cell_146 ( .C ( clk ), .D ( signal_58 ), .Q ( signal_384 ) ) ;
    buf_clk cell_148 ( .C ( clk ), .D ( signal_155 ), .Q ( signal_386 ) ) ;
    buf_clk cell_150 ( .C ( clk ), .D ( signal_156 ), .Q ( signal_388 ) ) ;
    buf_clk cell_152 ( .C ( clk ), .D ( signal_157 ), .Q ( signal_390 ) ) ;
    buf_clk cell_156 ( .C ( clk ), .D ( signal_393 ), .Q ( signal_394 ) ) ;
    buf_clk cell_162 ( .C ( clk ), .D ( signal_399 ), .Q ( signal_400 ) ) ;
    buf_clk cell_168 ( .C ( clk ), .D ( signal_405 ), .Q ( signal_406 ) ) ;
    buf_clk cell_174 ( .C ( clk ), .D ( signal_411 ), .Q ( signal_412 ) ) ;
    buf_clk cell_182 ( .C ( clk ), .D ( signal_419 ), .Q ( signal_420 ) ) ;
    buf_clk cell_192 ( .C ( clk ), .D ( signal_429 ), .Q ( signal_430 ) ) ;
    buf_clk cell_202 ( .C ( clk ), .D ( signal_439 ), .Q ( signal_440 ) ) ;
    buf_clk cell_212 ( .C ( clk ), .D ( signal_449 ), .Q ( signal_450 ) ) ;
    buf_clk cell_222 ( .C ( clk ), .D ( signal_459 ), .Q ( signal_460 ) ) ;
    buf_clk cell_232 ( .C ( clk ), .D ( signal_469 ), .Q ( signal_470 ) ) ;
    buf_clk cell_242 ( .C ( clk ), .D ( signal_479 ), .Q ( signal_480 ) ) ;
    buf_clk cell_252 ( .C ( clk ), .D ( signal_489 ), .Q ( signal_490 ) ) ;
    buf_clk cell_258 ( .C ( clk ), .D ( signal_17 ), .Q ( signal_496 ) ) ;
    buf_clk cell_264 ( .C ( clk ), .D ( signal_164 ), .Q ( signal_502 ) ) ;
    buf_clk cell_270 ( .C ( clk ), .D ( signal_165 ), .Q ( signal_508 ) ) ;
    buf_clk cell_276 ( .C ( clk ), .D ( signal_166 ), .Q ( signal_514 ) ) ;

    /* cells in depth 8 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_51 ( .a ({signal_383, signal_377, signal_371, signal_365}), .b ({signal_151, signal_150, signal_149, signal_56}), .clk ( clk ), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84]}), .c ({signal_163, signal_162, signal_161, signal_60}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_53 ( .a ({signal_163, signal_162, signal_161, signal_60}), .b ({signal_169, signal_168, signal_167, signal_61}) ) ;
    buf_clk cell_147 ( .C ( clk ), .D ( signal_384 ), .Q ( signal_385 ) ) ;
    buf_clk cell_149 ( .C ( clk ), .D ( signal_386 ), .Q ( signal_387 ) ) ;
    buf_clk cell_151 ( .C ( clk ), .D ( signal_388 ), .Q ( signal_389 ) ) ;
    buf_clk cell_153 ( .C ( clk ), .D ( signal_390 ), .Q ( signal_391 ) ) ;
    buf_clk cell_157 ( .C ( clk ), .D ( signal_394 ), .Q ( signal_395 ) ) ;
    buf_clk cell_163 ( .C ( clk ), .D ( signal_400 ), .Q ( signal_401 ) ) ;
    buf_clk cell_169 ( .C ( clk ), .D ( signal_406 ), .Q ( signal_407 ) ) ;
    buf_clk cell_175 ( .C ( clk ), .D ( signal_412 ), .Q ( signal_413 ) ) ;
    buf_clk cell_183 ( .C ( clk ), .D ( signal_420 ), .Q ( signal_421 ) ) ;
    buf_clk cell_193 ( .C ( clk ), .D ( signal_430 ), .Q ( signal_431 ) ) ;
    buf_clk cell_203 ( .C ( clk ), .D ( signal_440 ), .Q ( signal_441 ) ) ;
    buf_clk cell_213 ( .C ( clk ), .D ( signal_450 ), .Q ( signal_451 ) ) ;
    buf_clk cell_223 ( .C ( clk ), .D ( signal_460 ), .Q ( signal_461 ) ) ;
    buf_clk cell_233 ( .C ( clk ), .D ( signal_470 ), .Q ( signal_471 ) ) ;
    buf_clk cell_243 ( .C ( clk ), .D ( signal_480 ), .Q ( signal_481 ) ) ;
    buf_clk cell_253 ( .C ( clk ), .D ( signal_490 ), .Q ( signal_491 ) ) ;
    buf_clk cell_259 ( .C ( clk ), .D ( signal_496 ), .Q ( signal_497 ) ) ;
    buf_clk cell_265 ( .C ( clk ), .D ( signal_502 ), .Q ( signal_503 ) ) ;
    buf_clk cell_271 ( .C ( clk ), .D ( signal_508 ), .Q ( signal_509 ) ) ;
    buf_clk cell_277 ( .C ( clk ), .D ( signal_514 ), .Q ( signal_515 ) ) ;

    /* cells in depth 9 */
    buf_clk cell_158 ( .C ( clk ), .D ( signal_395 ), .Q ( signal_396 ) ) ;
    buf_clk cell_164 ( .C ( clk ), .D ( signal_401 ), .Q ( signal_402 ) ) ;
    buf_clk cell_170 ( .C ( clk ), .D ( signal_407 ), .Q ( signal_408 ) ) ;
    buf_clk cell_176 ( .C ( clk ), .D ( signal_413 ), .Q ( signal_414 ) ) ;
    buf_clk cell_184 ( .C ( clk ), .D ( signal_421 ), .Q ( signal_422 ) ) ;
    buf_clk cell_194 ( .C ( clk ), .D ( signal_431 ), .Q ( signal_432 ) ) ;
    buf_clk cell_204 ( .C ( clk ), .D ( signal_441 ), .Q ( signal_442 ) ) ;
    buf_clk cell_214 ( .C ( clk ), .D ( signal_451 ), .Q ( signal_452 ) ) ;
    buf_clk cell_224 ( .C ( clk ), .D ( signal_461 ), .Q ( signal_462 ) ) ;
    buf_clk cell_234 ( .C ( clk ), .D ( signal_471 ), .Q ( signal_472 ) ) ;
    buf_clk cell_244 ( .C ( clk ), .D ( signal_481 ), .Q ( signal_482 ) ) ;
    buf_clk cell_254 ( .C ( clk ), .D ( signal_491 ), .Q ( signal_492 ) ) ;
    buf_clk cell_260 ( .C ( clk ), .D ( signal_497 ), .Q ( signal_498 ) ) ;
    buf_clk cell_266 ( .C ( clk ), .D ( signal_503 ), .Q ( signal_504 ) ) ;
    buf_clk cell_272 ( .C ( clk ), .D ( signal_509 ), .Q ( signal_510 ) ) ;
    buf_clk cell_278 ( .C ( clk ), .D ( signal_515 ), .Q ( signal_516 ) ) ;

    /* cells in depth 10 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_54 ( .a ({signal_391, signal_389, signal_387, signal_385}), .b ({signal_169, signal_168, signal_167, signal_61}), .clk ( clk ), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({signal_172, signal_171, signal_170, signal_62}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_55 ( .a ({signal_172, signal_171, signal_170, signal_62}), .b ({signal_175, signal_174, signal_173, signal_63}) ) ;
    buf_clk cell_159 ( .C ( clk ), .D ( signal_396 ), .Q ( signal_397 ) ) ;
    buf_clk cell_165 ( .C ( clk ), .D ( signal_402 ), .Q ( signal_403 ) ) ;
    buf_clk cell_171 ( .C ( clk ), .D ( signal_408 ), .Q ( signal_409 ) ) ;
    buf_clk cell_177 ( .C ( clk ), .D ( signal_414 ), .Q ( signal_415 ) ) ;
    buf_clk cell_185 ( .C ( clk ), .D ( signal_422 ), .Q ( signal_423 ) ) ;
    buf_clk cell_195 ( .C ( clk ), .D ( signal_432 ), .Q ( signal_433 ) ) ;
    buf_clk cell_205 ( .C ( clk ), .D ( signal_442 ), .Q ( signal_443 ) ) ;
    buf_clk cell_215 ( .C ( clk ), .D ( signal_452 ), .Q ( signal_453 ) ) ;
    buf_clk cell_225 ( .C ( clk ), .D ( signal_462 ), .Q ( signal_463 ) ) ;
    buf_clk cell_235 ( .C ( clk ), .D ( signal_472 ), .Q ( signal_473 ) ) ;
    buf_clk cell_245 ( .C ( clk ), .D ( signal_482 ), .Q ( signal_483 ) ) ;
    buf_clk cell_255 ( .C ( clk ), .D ( signal_492 ), .Q ( signal_493 ) ) ;
    buf_clk cell_261 ( .C ( clk ), .D ( signal_498 ), .Q ( signal_499 ) ) ;
    buf_clk cell_267 ( .C ( clk ), .D ( signal_504 ), .Q ( signal_505 ) ) ;
    buf_clk cell_273 ( .C ( clk ), .D ( signal_510 ), .Q ( signal_511 ) ) ;
    buf_clk cell_279 ( .C ( clk ), .D ( signal_516 ), .Q ( signal_517 ) ) ;

    /* cells in depth 11 */
    buf_clk cell_186 ( .C ( clk ), .D ( signal_423 ), .Q ( signal_424 ) ) ;
    buf_clk cell_196 ( .C ( clk ), .D ( signal_433 ), .Q ( signal_434 ) ) ;
    buf_clk cell_206 ( .C ( clk ), .D ( signal_443 ), .Q ( signal_444 ) ) ;
    buf_clk cell_216 ( .C ( clk ), .D ( signal_453 ), .Q ( signal_454 ) ) ;
    buf_clk cell_226 ( .C ( clk ), .D ( signal_463 ), .Q ( signal_464 ) ) ;
    buf_clk cell_236 ( .C ( clk ), .D ( signal_473 ), .Q ( signal_474 ) ) ;
    buf_clk cell_246 ( .C ( clk ), .D ( signal_483 ), .Q ( signal_484 ) ) ;
    buf_clk cell_256 ( .C ( clk ), .D ( signal_493 ), .Q ( signal_494 ) ) ;
    buf_clk cell_262 ( .C ( clk ), .D ( signal_499 ), .Q ( signal_500 ) ) ;
    buf_clk cell_268 ( .C ( clk ), .D ( signal_505 ), .Q ( signal_506 ) ) ;
    buf_clk cell_274 ( .C ( clk ), .D ( signal_511 ), .Q ( signal_512 ) ) ;
    buf_clk cell_280 ( .C ( clk ), .D ( signal_517 ), .Q ( signal_518 ) ) ;

    /* cells in depth 12 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_56 ( .a ({signal_415, signal_409, signal_403, signal_397}), .b ({signal_175, signal_174, signal_173, signal_63}), .clk ( clk ), .r ({Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .c ({signal_178, signal_177, signal_176, signal_64}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_57 ( .a ({signal_178, signal_177, signal_176, signal_64}), .b ({signal_181, signal_180, signal_179, signal_18}) ) ;
    buf_clk cell_187 ( .C ( clk ), .D ( signal_424 ), .Q ( signal_425 ) ) ;
    buf_clk cell_197 ( .C ( clk ), .D ( signal_434 ), .Q ( signal_435 ) ) ;
    buf_clk cell_207 ( .C ( clk ), .D ( signal_444 ), .Q ( signal_445 ) ) ;
    buf_clk cell_217 ( .C ( clk ), .D ( signal_454 ), .Q ( signal_455 ) ) ;
    buf_clk cell_227 ( .C ( clk ), .D ( signal_464 ), .Q ( signal_465 ) ) ;
    buf_clk cell_237 ( .C ( clk ), .D ( signal_474 ), .Q ( signal_475 ) ) ;
    buf_clk cell_247 ( .C ( clk ), .D ( signal_484 ), .Q ( signal_485 ) ) ;
    buf_clk cell_257 ( .C ( clk ), .D ( signal_494 ), .Q ( signal_495 ) ) ;
    buf_clk cell_263 ( .C ( clk ), .D ( signal_500 ), .Q ( signal_501 ) ) ;
    buf_clk cell_269 ( .C ( clk ), .D ( signal_506 ), .Q ( signal_507 ) ) ;
    buf_clk cell_275 ( .C ( clk ), .D ( signal_512 ), .Q ( signal_513 ) ) ;
    buf_clk cell_281 ( .C ( clk ), .D ( signal_518 ), .Q ( signal_519 ) ) ;

    /* register cells */
    reg_masked #(.security_order(3), .pipeline(1)) cell_0 ( .clk ( clk ), .D ({signal_455, signal_445, signal_435, signal_425}), .Q ({SO_s3[3], SO_s2[3], SO_s1[3], SO_s0[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_1 ( .clk ( clk ), .D ({signal_495, signal_485, signal_475, signal_465}), .Q ({SO_s3[2], SO_s2[2], SO_s1[2], SO_s0[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_2 ( .clk ( clk ), .D ({signal_519, signal_513, signal_507, signal_501}), .Q ({SO_s3[1], SO_s2[1], SO_s1[1], SO_s0[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_3 ( .clk ( clk ), .D ({signal_181, signal_180, signal_179, signal_18}), .Q ({SO_s3[0], SO_s2[0], SO_s1[0], SO_s0[0]}) ) ;
endmodule
