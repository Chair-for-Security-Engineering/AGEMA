/* modified netlist. Source: module AES in file ../CaseStudies/07_AES128_byte_serial_encryption/FPGA_based/AES_synthesis.v */
/* clock gating is added to the circuit, the latency increased 2 time(s)  */

module AES_GHPCLL_ClockGating_d1 (clk, start, plaintext_s0, key_s0, plaintext_s1, key_s1, Fresh, done, ciphertext_s0, ciphertext_s1, Synch);
    input clk ;
    input start ;
    input [127:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input [127:0] plaintext_s1 ;
    input [127:0] key_s1 ;
    input [2559:0] Fresh ;
    output done ;
    output [127:0] ciphertext_s0 ;
    output [127:0] ciphertext_s1 ;
    output Synch ;
    wire \KeyArray/S13reg/gen_ff[1].gff/GEN[7].SFF/Q_386 ;
    wire \KeyArray/S13reg/gen_ff[1].gff/GEN[6].SFF/Q_387 ;
    wire \KeyArray/S13reg/gen_ff[1].gff/GEN[5].SFF/Q_388 ;
    wire \KeyArray/S13reg/gen_ff[1].gff/GEN[4].SFF/Q_389 ;
    wire \KeyArray/S13reg/gen_ff[1].gff/GEN[3].SFF/Q_390 ;
    wire \KeyArray/S13reg/gen_ff[1].gff/GEN[2].SFF/Q_391 ;
    wire \KeyArray/S13reg/gen_ff[1].gff/GEN[1].SFF/Q_392 ;
    wire \KeyArray/S13reg/gen_ff[1].gff/GEN[0].SFF/Q_393 ;
    wire \KeyArray/S00reg/gen_ff[1].gff/GEN[7].SFF/Q_394 ;
    wire \KeyArray/S00reg/gen_ff[1].gff/GEN[6].SFF/Q_395 ;
    wire \KeyArray/S00reg/gen_ff[1].gff/GEN[5].SFF/Q_396 ;
    wire \KeyArray/S00reg/gen_ff[1].gff/GEN[4].SFF/Q_397 ;
    wire \KeyArray/S00reg/gen_ff[1].gff/GEN[3].SFF/Q_398 ;
    wire \KeyArray/S00reg/gen_ff[1].gff/GEN[2].SFF/Q_399 ;
    wire \KeyArray/S00reg/gen_ff[1].gff/GEN[1].SFF/Q_400 ;
    wire \KeyArray/S00reg/gen_ff[1].gff/GEN[0].SFF/Q_401 ;
    wire selMC ;
    wire selSR ;
    wire selXOR ;
    wire \ctrl/CSenRC_405 ;
    wire intFinal ;
    wire nReset_407 ;
    wire enKS ;
    wire intselXOR_425 ;
    wire \stateArray/S00reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \stateArray/S00reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \stateArray/S00reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \stateArray/S00reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \stateArray/S00reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \stateArray/S00reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \stateArray/S00reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \stateArray/S00reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \stateArray/S01reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \stateArray/S01reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \stateArray/S01reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \stateArray/S01reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \stateArray/S01reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \stateArray/S01reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \stateArray/S01reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \stateArray/S01reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \stateArray/S02reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \stateArray/S02reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \stateArray/S02reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \stateArray/S02reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \stateArray/S02reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \stateArray/S02reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \stateArray/S02reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \stateArray/S02reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \stateArray/S10reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \stateArray/S10reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \stateArray/S10reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \stateArray/S10reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \stateArray/S10reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \stateArray/S10reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \stateArray/S10reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \stateArray/S10reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \stateArray/S11reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \stateArray/S11reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \stateArray/S11reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \stateArray/S11reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \stateArray/S11reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \stateArray/S11reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \stateArray/S11reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \stateArray/S11reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \stateArray/S12reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \stateArray/S12reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \stateArray/S12reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \stateArray/S12reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \stateArray/S12reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \stateArray/S12reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \stateArray/S12reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \stateArray/S12reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \stateArray/S20reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \stateArray/S20reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \stateArray/S20reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \stateArray/S20reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \stateArray/S20reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \stateArray/S20reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \stateArray/S20reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \stateArray/S20reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \stateArray/S21reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \stateArray/S21reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \stateArray/S21reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \stateArray/S21reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \stateArray/S21reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \stateArray/S21reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \stateArray/S21reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \stateArray/S21reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \stateArray/S22reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \stateArray/S22reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \stateArray/S22reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \stateArray/S22reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \stateArray/S22reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \stateArray/S22reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \stateArray/S22reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \stateArray/S22reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \stateArray/S30reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \stateArray/S30reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \stateArray/S30reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \stateArray/S30reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \stateArray/S30reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \stateArray/S30reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \stateArray/S30reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \stateArray/S30reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \stateArray/S31reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \stateArray/S31reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \stateArray/S31reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \stateArray/S31reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \stateArray/S31reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \stateArray/S31reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \stateArray/S31reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \stateArray/S31reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \stateArray/S32reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \stateArray/S32reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \stateArray/S32reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \stateArray/S32reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \stateArray/S32reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \stateArray/S32reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \stateArray/S32reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \stateArray/S32reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \stateArray/S33reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \stateArray/S33reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \stateArray/S33reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \stateArray/S33reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \stateArray/S33reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \stateArray/S33reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \stateArray/S33reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \stateArray/S33reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \KeyArray/S33reg/gen_ff[1].gff/GEN[0].SFF/Q_587 ;
    wire \KeyArray/S33reg/gen_ff[1].gff/GEN[1].SFF/Q_588 ;
    wire \KeyArray/S33reg/gen_ff[1].gff/GEN[2].SFF/Q_589 ;
    wire \KeyArray/S33reg/gen_ff[1].gff/GEN[3].SFF/Q_590 ;
    wire \KeyArray/S33reg/gen_ff[1].gff/GEN[4].SFF/Q_591 ;
    wire \KeyArray/S33reg/gen_ff[1].gff/GEN[5].SFF/Q_592 ;
    wire \KeyArray/S33reg/gen_ff[1].gff/GEN[6].SFF/Q_593 ;
    wire \KeyArray/S33reg/gen_ff[1].gff/GEN[7].SFF/Q_594 ;
    wire \KeyArray/S32reg/gen_ff[1].gff/GEN[0].SFF/Q_595 ;
    wire \KeyArray/S32reg/gen_ff[1].gff/GEN[1].SFF/Q_596 ;
    wire \KeyArray/S32reg/gen_ff[1].gff/GEN[2].SFF/Q_597 ;
    wire \KeyArray/S32reg/gen_ff[1].gff/GEN[3].SFF/Q_598 ;
    wire \KeyArray/S32reg/gen_ff[1].gff/GEN[4].SFF/Q_599 ;
    wire \KeyArray/S32reg/gen_ff[1].gff/GEN[5].SFF/Q_600 ;
    wire \KeyArray/S32reg/gen_ff[1].gff/GEN[6].SFF/Q_601 ;
    wire \KeyArray/S32reg/gen_ff[1].gff/GEN[7].SFF/Q_602 ;
    wire \KeyArray/S31reg/gen_ff[1].gff/GEN[0].SFF/Q_603 ;
    wire \KeyArray/S31reg/gen_ff[1].gff/GEN[1].SFF/Q_604 ;
    wire \KeyArray/S31reg/gen_ff[1].gff/GEN[2].SFF/Q_605 ;
    wire \KeyArray/S31reg/gen_ff[1].gff/GEN[3].SFF/Q_606 ;
    wire \KeyArray/S31reg/gen_ff[1].gff/GEN[4].SFF/Q_607 ;
    wire \KeyArray/S31reg/gen_ff[1].gff/GEN[5].SFF/Q_608 ;
    wire \KeyArray/S31reg/gen_ff[1].gff/GEN[6].SFF/Q_609 ;
    wire \KeyArray/S31reg/gen_ff[1].gff/GEN[7].SFF/Q_610 ;
    wire \KeyArray/S30reg/gen_ff[1].gff/GEN[0].SFF/Q_611 ;
    wire \KeyArray/S30reg/gen_ff[1].gff/GEN[1].SFF/Q_612 ;
    wire \KeyArray/S30reg/gen_ff[1].gff/GEN[2].SFF/Q_613 ;
    wire \KeyArray/S30reg/gen_ff[1].gff/GEN[3].SFF/Q_614 ;
    wire \KeyArray/S30reg/gen_ff[1].gff/GEN[4].SFF/Q_615 ;
    wire \KeyArray/S30reg/gen_ff[1].gff/GEN[5].SFF/Q_616 ;
    wire \KeyArray/S30reg/gen_ff[1].gff/GEN[6].SFF/Q_617 ;
    wire \KeyArray/S30reg/gen_ff[1].gff/GEN[7].SFF/Q_618 ;
    wire \KeyArray/S23reg/gen_ff[1].gff/GEN[0].SFF/Q_619 ;
    wire \KeyArray/S23reg/gen_ff[1].gff/GEN[1].SFF/Q_620 ;
    wire \KeyArray/S23reg/gen_ff[1].gff/GEN[2].SFF/Q_621 ;
    wire \KeyArray/S23reg/gen_ff[1].gff/GEN[3].SFF/Q_622 ;
    wire \KeyArray/S23reg/gen_ff[1].gff/GEN[4].SFF/Q_623 ;
    wire \KeyArray/S23reg/gen_ff[1].gff/GEN[5].SFF/Q_624 ;
    wire \KeyArray/S23reg/gen_ff[1].gff/GEN[6].SFF/Q_625 ;
    wire \KeyArray/S23reg/gen_ff[1].gff/GEN[7].SFF/Q_626 ;
    wire \KeyArray/S22reg/gen_ff[1].gff/GEN[0].SFF/Q_627 ;
    wire \KeyArray/S22reg/gen_ff[1].gff/GEN[1].SFF/Q_628 ;
    wire \KeyArray/S22reg/gen_ff[1].gff/GEN[2].SFF/Q_629 ;
    wire \KeyArray/S22reg/gen_ff[1].gff/GEN[3].SFF/Q_630 ;
    wire \KeyArray/S22reg/gen_ff[1].gff/GEN[4].SFF/Q_631 ;
    wire \KeyArray/S22reg/gen_ff[1].gff/GEN[5].SFF/Q_632 ;
    wire \KeyArray/S22reg/gen_ff[1].gff/GEN[6].SFF/Q_633 ;
    wire \KeyArray/S22reg/gen_ff[1].gff/GEN[7].SFF/Q_634 ;
    wire \KeyArray/S21reg/gen_ff[1].gff/GEN[0].SFF/Q_635 ;
    wire \KeyArray/S21reg/gen_ff[1].gff/GEN[1].SFF/Q_636 ;
    wire \KeyArray/S21reg/gen_ff[1].gff/GEN[2].SFF/Q_637 ;
    wire \KeyArray/S21reg/gen_ff[1].gff/GEN[3].SFF/Q_638 ;
    wire \KeyArray/S21reg/gen_ff[1].gff/GEN[4].SFF/Q_639 ;
    wire \KeyArray/S21reg/gen_ff[1].gff/GEN[5].SFF/Q_640 ;
    wire \KeyArray/S21reg/gen_ff[1].gff/GEN[6].SFF/Q_641 ;
    wire \KeyArray/S21reg/gen_ff[1].gff/GEN[7].SFF/Q_642 ;
    wire \KeyArray/S20reg/gen_ff[1].gff/GEN[0].SFF/Q_643 ;
    wire \KeyArray/S20reg/gen_ff[1].gff/GEN[1].SFF/Q_644 ;
    wire \KeyArray/S20reg/gen_ff[1].gff/GEN[2].SFF/Q_645 ;
    wire \KeyArray/S20reg/gen_ff[1].gff/GEN[3].SFF/Q_646 ;
    wire \KeyArray/S20reg/gen_ff[1].gff/GEN[4].SFF/Q_647 ;
    wire \KeyArray/S20reg/gen_ff[1].gff/GEN[5].SFF/Q_648 ;
    wire \KeyArray/S20reg/gen_ff[1].gff/GEN[6].SFF/Q_649 ;
    wire \KeyArray/S20reg/gen_ff[1].gff/GEN[7].SFF/Q_650 ;
    wire \KeyArray/S12reg/gen_ff[1].gff/GEN[0].SFF/Q_651 ;
    wire \KeyArray/S12reg/gen_ff[1].gff/GEN[1].SFF/Q_652 ;
    wire \KeyArray/S12reg/gen_ff[1].gff/GEN[2].SFF/Q_653 ;
    wire \KeyArray/S12reg/gen_ff[1].gff/GEN[3].SFF/Q_654 ;
    wire \KeyArray/S12reg/gen_ff[1].gff/GEN[4].SFF/Q_655 ;
    wire \KeyArray/S12reg/gen_ff[1].gff/GEN[5].SFF/Q_656 ;
    wire \KeyArray/S12reg/gen_ff[1].gff/GEN[6].SFF/Q_657 ;
    wire \KeyArray/S12reg/gen_ff[1].gff/GEN[7].SFF/Q_658 ;
    wire \KeyArray/S11reg/gen_ff[1].gff/GEN[0].SFF/Q_659 ;
    wire \KeyArray/S11reg/gen_ff[1].gff/GEN[1].SFF/Q_660 ;
    wire \KeyArray/S11reg/gen_ff[1].gff/GEN[2].SFF/Q_661 ;
    wire \KeyArray/S11reg/gen_ff[1].gff/GEN[3].SFF/Q_662 ;
    wire \KeyArray/S11reg/gen_ff[1].gff/GEN[4].SFF/Q_663 ;
    wire \KeyArray/S11reg/gen_ff[1].gff/GEN[5].SFF/Q_664 ;
    wire \KeyArray/S11reg/gen_ff[1].gff/GEN[6].SFF/Q_665 ;
    wire \KeyArray/S11reg/gen_ff[1].gff/GEN[7].SFF/Q_666 ;
    wire \KeyArray/S10reg/gen_ff[1].gff/GEN[0].SFF/Q_667 ;
    wire \KeyArray/S10reg/gen_ff[1].gff/GEN[1].SFF/Q_668 ;
    wire \KeyArray/S10reg/gen_ff[1].gff/GEN[2].SFF/Q_669 ;
    wire \KeyArray/S10reg/gen_ff[1].gff/GEN[3].SFF/Q_670 ;
    wire \KeyArray/S10reg/gen_ff[1].gff/GEN[4].SFF/Q_671 ;
    wire \KeyArray/S10reg/gen_ff[1].gff/GEN[5].SFF/Q_672 ;
    wire \KeyArray/S10reg/gen_ff[1].gff/GEN[6].SFF/Q_673 ;
    wire \KeyArray/S10reg/gen_ff[1].gff/GEN[7].SFF/Q_674 ;
    wire \KeyArray/S03reg/gen_ff[1].gff/GEN[0].SFF/Q_675 ;
    wire \KeyArray/S03reg/gen_ff[1].gff/GEN[1].SFF/Q_676 ;
    wire \KeyArray/S03reg/gen_ff[1].gff/GEN[2].SFF/Q_677 ;
    wire \KeyArray/S03reg/gen_ff[1].gff/GEN[3].SFF/Q_678 ;
    wire \KeyArray/S03reg/gen_ff[1].gff/GEN[4].SFF/Q_679 ;
    wire \KeyArray/S03reg/gen_ff[1].gff/GEN[5].SFF/Q_680 ;
    wire \KeyArray/S03reg/gen_ff[1].gff/GEN[6].SFF/Q_681 ;
    wire \KeyArray/S03reg/gen_ff[1].gff/GEN[7].SFF/Q_682 ;
    wire \KeyArray/S02reg/gen_ff[1].gff/GEN[0].SFF/Q_683 ;
    wire \KeyArray/S02reg/gen_ff[1].gff/GEN[1].SFF/Q_684 ;
    wire \KeyArray/S02reg/gen_ff[1].gff/GEN[2].SFF/Q_685 ;
    wire \KeyArray/S02reg/gen_ff[1].gff/GEN[3].SFF/Q_686 ;
    wire \KeyArray/S02reg/gen_ff[1].gff/GEN[4].SFF/Q_687 ;
    wire \KeyArray/S02reg/gen_ff[1].gff/GEN[5].SFF/Q_688 ;
    wire \KeyArray/S02reg/gen_ff[1].gff/GEN[6].SFF/Q_689 ;
    wire \KeyArray/S02reg/gen_ff[1].gff/GEN[7].SFF/Q_690 ;
    wire \KeyArray/S01reg/gen_ff[1].gff/GEN[0].SFF/Q_691 ;
    wire \KeyArray/S01reg/gen_ff[1].gff/GEN[1].SFF/Q_692 ;
    wire \KeyArray/S01reg/gen_ff[1].gff/GEN[2].SFF/Q_693 ;
    wire \KeyArray/S01reg/gen_ff[1].gff/GEN[3].SFF/Q_694 ;
    wire \KeyArray/S01reg/gen_ff[1].gff/GEN[4].SFF/Q_695 ;
    wire \KeyArray/S01reg/gen_ff[1].gff/GEN[5].SFF/Q_696 ;
    wire \KeyArray/S01reg/gen_ff[1].gff/GEN[6].SFF/Q_697 ;
    wire \KeyArray/S01reg/gen_ff[1].gff/GEN[7].SFF/Q_698 ;
    wire \KeyArray/S00reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \KeyArray/S00reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \KeyArray/S00reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \KeyArray/S00reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \KeyArray/S00reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \KeyArray/S00reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \KeyArray/S00reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \KeyArray/S00reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \KeyArray/S01reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \KeyArray/S01reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \KeyArray/S01reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \KeyArray/S01reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \KeyArray/S01reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \KeyArray/S01reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \KeyArray/S01reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \KeyArray/S01reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \KeyArray/S02reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \KeyArray/S02reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \KeyArray/S02reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \KeyArray/S02reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \KeyArray/S02reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \KeyArray/S02reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \KeyArray/S02reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \KeyArray/S02reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \KeyArray/S03reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \KeyArray/S03reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \KeyArray/S03reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \KeyArray/S03reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \KeyArray/S03reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \KeyArray/S03reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \KeyArray/S03reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \KeyArray/S03reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \KeyArray/S10reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \KeyArray/S10reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \KeyArray/S10reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \KeyArray/S10reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \KeyArray/S10reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \KeyArray/S10reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \KeyArray/S10reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \KeyArray/S10reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \KeyArray/S11reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \KeyArray/S11reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \KeyArray/S11reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \KeyArray/S11reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \KeyArray/S11reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \KeyArray/S11reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \KeyArray/S11reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \KeyArray/S11reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \KeyArray/S12reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \KeyArray/S12reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \KeyArray/S12reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \KeyArray/S12reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \KeyArray/S12reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \KeyArray/S12reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \KeyArray/S12reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \KeyArray/S12reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \KeyArray/S13reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \KeyArray/S13reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \KeyArray/S13reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \KeyArray/S13reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \KeyArray/S13reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \KeyArray/S13reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \KeyArray/S13reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \KeyArray/S13reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \KeyArray/S20reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \KeyArray/S20reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \KeyArray/S20reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \KeyArray/S20reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \KeyArray/S20reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \KeyArray/S20reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \KeyArray/S20reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \KeyArray/S20reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \KeyArray/S21reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \KeyArray/S21reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \KeyArray/S21reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \KeyArray/S21reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \KeyArray/S21reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \KeyArray/S21reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \KeyArray/S21reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \KeyArray/S21reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \KeyArray/S22reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \KeyArray/S22reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \KeyArray/S22reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \KeyArray/S22reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \KeyArray/S22reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \KeyArray/S22reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \KeyArray/S22reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \KeyArray/S22reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \KeyArray/S23reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \KeyArray/S23reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \KeyArray/S23reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \KeyArray/S23reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \KeyArray/S23reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \KeyArray/S23reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \KeyArray/S23reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \KeyArray/S23reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \KeyArray/S30reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \KeyArray/S30reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \KeyArray/S30reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \KeyArray/S30reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \KeyArray/S30reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \KeyArray/S30reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \KeyArray/S30reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \KeyArray/S30reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \KeyArray/S31reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \KeyArray/S31reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \KeyArray/S31reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \KeyArray/S31reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \KeyArray/S31reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \KeyArray/S31reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \KeyArray/S31reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \KeyArray/S31reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \KeyArray/S32reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \KeyArray/S32reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \KeyArray/S32reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \KeyArray/S32reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \KeyArray/S32reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \KeyArray/S32reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \KeyArray/S32reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \KeyArray/S32reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \KeyArray/S33reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \KeyArray/S33reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \KeyArray/S33reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \KeyArray/S33reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \KeyArray/S33reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \KeyArray/S33reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \KeyArray/S33reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \KeyArray/S33reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \ctrl/finalStep1 ;
    wire \ctrl/seq4/GEN[1].SFF/QD ;
    wire \ctrl/seq4/GEN[0].SFF/QD ;
    wire \ctrl/seq6/GEN[4].SFF/QD ;
    wire \ctrl/seq6/GEN[3].SFF/QD ;
    wire \ctrl/seq6/GEN[2].SFF/QD ;
    wire \ctrl/seq6/GEN[1].SFF/QD ;
    wire \ctrl/seq6/GEN[0].SFF/QD ;
    wire \ctrl/CSselMC_835 ;
    wire \ctrl/seq4/GEN[0].SFF/Q_836 ;
    wire \ctrl/seq4/GEN[1].SFF/Q_837 ;
    wire \ctrl/seq6/GEN[1].SFF/Q_838 ;
    wire \ctrl/seq6/GEN[2].SFF/Q_839 ;
    wire \ctrl/seq6/GEN[3].SFF/Q_840 ;
    wire \ctrl/seq6/GEN[0].SFF/Q_841 ;
    wire \ctrl/seq6/GEN[4].SFF/Q_842 ;
    wire \calcRCon/nReset_inv ;
    wire \calcRCon/MSB_s_current_state[0]_XOR_21_o ;
    wire \calcRCon/MSB_s_current_state[2]_XOR_20_o ;
    wire \calcRCon/MSB_s_current_state[3]_XOR_19_o ;
    wire N01 ;
    wire N2 ;
    wire N4 ;
    wire N6 ;
    wire N8 ;
    wire N10 ;
    wire N12 ;
    wire N14 ;
    wire N16 ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q1 ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11_897 ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q12 ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q1 ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11_900 ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q12 ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q12 ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q1 ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11_904 ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q1 ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11_906 ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q1 ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11_908 ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q1 ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11_910 ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q12 ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q1 ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11_913 ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q12 ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q12 ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q1 ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11_917 ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q1 ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11_919 ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q1 ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11_921 ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q1 ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11_923 ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q12 ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q1 ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11_926 ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q12 ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q12 ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q1 ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11_930 ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q1 ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11_932 ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q1 ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11_934 ;
    wire N18 ;
    wire N20 ;
    wire N22 ;
    wire N24 ;
    wire N26 ;
    wire N28 ;
    wire N30 ;
    wire N32 ;
    wire \ctrl/CSselMC_rstpot_1330 ;
    wire nReset_rstpot ;
    wire N34 ;
    wire N36 ;
    wire N38 ;
    wire N40 ;
    wire N42 ;
    wire N44 ;
    wire N46 ;
    wire N48 ;
    wire N50 ;
    wire nReset_1_1341 ;
    wire \ctrl/CSselMC_1_1342 ;
    wire [7:0] StateInMC ;
    wire [7:0] SboxIn ;
    wire [7:0] StateOutXORroundKey ;
    wire [7:0] SboxOut ;
    wire [7:0] \stateArray/input_MC ;
    wire [7:0] \KeyArray/inS00ser ;
    wire [7:0] \calcRCon/s_current_state ;
    wire [3:0] \Inst_bSbox/b7 ;
    wire [3:0] \Inst_bSbox/b6 ;
    wire [3:0] \Inst_bSbox/b5 ;
    wire [3:0] \Inst_bSbox/b4 ;
    wire [3:0] \Inst_bSbox/b3 ;
    wire [3:0] \Inst_bSbox/b2 ;
    wire [3:0] \Inst_bSbox/b1 ;
    wire [3:0] \Inst_bSbox/b0 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1412 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1528 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1564 ;
    wire new_AGEMA_signal_1565 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1573 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1581 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1591 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1609 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1619 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1627 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1645 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1654 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1663 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1699 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1789 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1799 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1870 ;
    wire new_AGEMA_signal_1871 ;
    wire new_AGEMA_signal_1872 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1880 ;
    wire new_AGEMA_signal_1881 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1888 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1896 ;
    wire new_AGEMA_signal_1897 ;
    wire new_AGEMA_signal_1898 ;
    wire new_AGEMA_signal_1899 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1906 ;
    wire new_AGEMA_signal_1907 ;
    wire new_AGEMA_signal_1908 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1914 ;
    wire new_AGEMA_signal_1915 ;
    wire new_AGEMA_signal_1916 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1923 ;
    wire new_AGEMA_signal_1924 ;
    wire new_AGEMA_signal_1927 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1933 ;
    wire new_AGEMA_signal_1936 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1942 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1951 ;
    wire new_AGEMA_signal_1954 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1960 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1969 ;
    wire new_AGEMA_signal_1972 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1978 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1996 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2004 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2016 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2034 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2043 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2052 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2106 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2124 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2130 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2134 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2140 ;
    wire new_AGEMA_signal_2142 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2150 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2154 ;
    wire new_AGEMA_signal_2156 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2158 ;
    wire new_AGEMA_signal_2159 ;
    wire new_AGEMA_signal_2160 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2166 ;
    wire new_AGEMA_signal_2168 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2176 ;
    wire new_AGEMA_signal_2178 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2186 ;
    wire new_AGEMA_signal_2188 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2194 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2212 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2214 ;
    wire new_AGEMA_signal_2215 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2222 ;
    wire new_AGEMA_signal_2224 ;
    wire new_AGEMA_signal_2226 ;
    wire new_AGEMA_signal_2228 ;
    wire new_AGEMA_signal_2230 ;
    wire new_AGEMA_signal_2232 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2236 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2239 ;
    wire new_AGEMA_signal_2240 ;
    wire new_AGEMA_signal_2241 ;
    wire new_AGEMA_signal_2242 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2248 ;
    wire new_AGEMA_signal_2250 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2260 ;
    wire clk_gated ;

    /* cells in depth 0 */
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CCCAAAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CCCAAAA ) ) \KeyArray/gen00ser[7].inS00serInst ( .I0 ({key_s1[127], key_s0[127]}), .I1 ({new_AGEMA_signal_1826, \KeyArray/S01reg/gen_ff[1].gff/GEN[7].SFF/Q_698 }), .I2 ({new_AGEMA_signal_1350, \KeyArray/S00reg/gen_ff[1].gff/GEN[7].SFF/Q_394 }), .I3 ({1'b0, intselXOR_425}), .I4 ({1'b0, nReset_407}), .O ({new_AGEMA_signal_2142, \KeyArray/inS00ser [7]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CCCAAAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CCCAAAA ) ) \KeyArray/gen00ser[6].inS00serInst ( .I0 ({key_s1[126], key_s0[126]}), .I1 ({new_AGEMA_signal_1823, \KeyArray/S01reg/gen_ff[1].gff/GEN[6].SFF/Q_697 }), .I2 ({new_AGEMA_signal_1353, \KeyArray/S00reg/gen_ff[1].gff/GEN[6].SFF/Q_395 }), .I3 ({1'b0, intselXOR_425}), .I4 ({1'b0, nReset_407}), .O ({new_AGEMA_signal_2144, \KeyArray/inS00ser [6]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CCCAAAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CCCAAAA ) ) \KeyArray/gen00ser[5].inS00serInst ( .I0 ({key_s1[125], key_s0[125]}), .I1 ({new_AGEMA_signal_1820, \KeyArray/S01reg/gen_ff[1].gff/GEN[5].SFF/Q_696 }), .I2 ({new_AGEMA_signal_1356, \KeyArray/S00reg/gen_ff[1].gff/GEN[5].SFF/Q_396 }), .I3 ({1'b0, intselXOR_425}), .I4 ({1'b0, nReset_407}), .O ({new_AGEMA_signal_2146, \KeyArray/inS00ser [5]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CCCAAAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CCCAAAA ) ) \KeyArray/gen00ser[4].inS00serInst ( .I0 ({key_s1[124], key_s0[124]}), .I1 ({new_AGEMA_signal_1817, \KeyArray/S01reg/gen_ff[1].gff/GEN[4].SFF/Q_695 }), .I2 ({new_AGEMA_signal_1359, \KeyArray/S00reg/gen_ff[1].gff/GEN[4].SFF/Q_397 }), .I3 ({1'b0, intselXOR_425}), .I4 ({1'b0, nReset_407}), .O ({new_AGEMA_signal_2148, \KeyArray/inS00ser [4]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CCCAAAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CCCAAAA ) ) \KeyArray/gen00ser[3].inS00serInst ( .I0 ({key_s1[123], key_s0[123]}), .I1 ({new_AGEMA_signal_1814, \KeyArray/S01reg/gen_ff[1].gff/GEN[3].SFF/Q_694 }), .I2 ({new_AGEMA_signal_1362, \KeyArray/S00reg/gen_ff[1].gff/GEN[3].SFF/Q_398 }), .I3 ({1'b0, intselXOR_425}), .I4 ({1'b0, nReset_407}), .O ({new_AGEMA_signal_2150, \KeyArray/inS00ser [3]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CCCAAAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CCCAAAA ) ) \KeyArray/gen00ser[2].inS00serInst ( .I0 ({key_s1[122], key_s0[122]}), .I1 ({new_AGEMA_signal_1811, \KeyArray/S01reg/gen_ff[1].gff/GEN[2].SFF/Q_693 }), .I2 ({new_AGEMA_signal_1365, \KeyArray/S00reg/gen_ff[1].gff/GEN[2].SFF/Q_399 }), .I3 ({1'b0, intselXOR_425}), .I4 ({1'b0, nReset_407}), .O ({new_AGEMA_signal_2152, \KeyArray/inS00ser [2]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CCCAAAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CCCAAAA ) ) \KeyArray/gen00ser[1].inS00serInst ( .I0 ({key_s1[121], key_s0[121]}), .I1 ({new_AGEMA_signal_1808, \KeyArray/S01reg/gen_ff[1].gff/GEN[1].SFF/Q_692 }), .I2 ({new_AGEMA_signal_1368, \KeyArray/S00reg/gen_ff[1].gff/GEN[1].SFF/Q_400 }), .I3 ({1'b0, intselXOR_425}), .I4 ({1'b0, nReset_407}), .O ({new_AGEMA_signal_2154, \KeyArray/inS00ser [1]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CCCAAAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CCCAAAA ) ) \KeyArray/gen00ser[0].inS00serInst ( .I0 ({key_s1[120], key_s0[120]}), .I1 ({new_AGEMA_signal_1805, \KeyArray/S01reg/gen_ff[1].gff/GEN[0].SFF/Q_691 }), .I2 ({new_AGEMA_signal_1371, \KeyArray/S00reg/gen_ff[1].gff/GEN[0].SFF/Q_401 }), .I3 ({1'b0, intselXOR_425}), .I4 ({1'b0, nReset_407}), .O ({new_AGEMA_signal_2156, \KeyArray/inS00ser [0]}) ) ;
    LUT5 #( .INIT ( 32'h00800000 ) ) done1 ( .I0 (intFinal), .I1 (nReset_407), .I2 (\ctrl/seq4/GEN[0].SFF/Q_836 ), .I3 (\ctrl/seq4/GEN[1].SFF/Q_837 ), .I4 (\ctrl/finalStep1 ), .O (done) ) ;
    LUT2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \StateOutXORroundKey<7>1 ( .I0 ({ciphertext_s1[127], ciphertext_s0[127]}), .I1 ({new_AGEMA_signal_1350, \KeyArray/S00reg/gen_ff[1].gff/GEN[7].SFF/Q_394 }), .O ({new_AGEMA_signal_1351, StateOutXORroundKey[7]}) ) ;
    LUT2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \StateOutXORroundKey<6>1 ( .I0 ({ciphertext_s1[126], ciphertext_s0[126]}), .I1 ({new_AGEMA_signal_1353, \KeyArray/S00reg/gen_ff[1].gff/GEN[6].SFF/Q_395 }), .O ({new_AGEMA_signal_1354, StateOutXORroundKey[6]}) ) ;
    LUT2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \StateOutXORroundKey<5>1 ( .I0 ({ciphertext_s1[125], ciphertext_s0[125]}), .I1 ({new_AGEMA_signal_1356, \KeyArray/S00reg/gen_ff[1].gff/GEN[5].SFF/Q_396 }), .O ({new_AGEMA_signal_1357, StateOutXORroundKey[5]}) ) ;
    LUT2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \StateOutXORroundKey<4>1 ( .I0 ({ciphertext_s1[124], ciphertext_s0[124]}), .I1 ({new_AGEMA_signal_1359, \KeyArray/S00reg/gen_ff[1].gff/GEN[4].SFF/Q_397 }), .O ({new_AGEMA_signal_1360, StateOutXORroundKey[4]}) ) ;
    LUT2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \StateOutXORroundKey<3>1 ( .I0 ({ciphertext_s1[123], ciphertext_s0[123]}), .I1 ({new_AGEMA_signal_1362, \KeyArray/S00reg/gen_ff[1].gff/GEN[3].SFF/Q_398 }), .O ({new_AGEMA_signal_1363, StateOutXORroundKey[3]}) ) ;
    LUT2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \StateOutXORroundKey<2>1 ( .I0 ({ciphertext_s1[122], ciphertext_s0[122]}), .I1 ({new_AGEMA_signal_1365, \KeyArray/S00reg/gen_ff[1].gff/GEN[2].SFF/Q_399 }), .O ({new_AGEMA_signal_1366, StateOutXORroundKey[2]}) ) ;
    LUT2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \StateOutXORroundKey<1>1 ( .I0 ({ciphertext_s1[121], ciphertext_s0[121]}), .I1 ({new_AGEMA_signal_1368, \KeyArray/S00reg/gen_ff[1].gff/GEN[1].SFF/Q_400 }), .O ({new_AGEMA_signal_1369, StateOutXORroundKey[1]}) ) ;
    LUT2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \StateOutXORroundKey<0>1 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({new_AGEMA_signal_1371, \KeyArray/S00reg/gen_ff[1].gff/GEN[0].SFF/Q_401 }), .O ({new_AGEMA_signal_1372, StateOutXORroundKey[0]}) ) ;
    LUT3 #( .INIT ( 8'hE0 ) ) \ctrl/intSelXOR1 ( .I0 (\ctrl/seq4/GEN[1].SFF/Q_837 ), .I1 (\ctrl/seq4/GEN[0].SFF/Q_836 ), .I2 (nReset_407), .O (selXOR) ) ;
    LUT5 #( .INIT ( 32'h00000001 ) ) \ctrl/finalStep11 ( .I0 (\ctrl/seq6/GEN[0].SFF/Q_841 ), .I1 (\ctrl/seq6/GEN[4].SFF/Q_842 ), .I2 (\ctrl/seq6/GEN[3].SFF/Q_840 ), .I3 (\ctrl/seq6/GEN[1].SFF/Q_838 ), .I4 (\ctrl/seq6/GEN[2].SFF/Q_839 ), .O (\ctrl/finalStep1 ) ) ;
    LUT3 #( .INIT ( 8'h20 ) ) \ctrl/seq4/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 (\ctrl/seq4/GEN[0].SFF/Q_836 ), .I1 (\ctrl/finalStep1 ), .I2 (nReset_407), .O (\ctrl/seq4/GEN[1].SFF/QD ) ) ;
    LUT3 #( .INIT ( 8'hDF ) ) \ctrl/seq4/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 (nReset_407), .I1 (\ctrl/finalStep1 ), .I2 (\ctrl/seq4/GEN[1].SFF/Q_837 ), .O (\ctrl/seq4/GEN[0].SFF/QD ) ) ;
    LUT2 #( .INIT ( 4'hD ) ) \ctrl/seq6/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 (nReset_407), .I1 (\ctrl/seq6/GEN[3].SFF/Q_840 ), .O (\ctrl/seq6/GEN[4].SFF/QD ) ) ;
    LUT2 #( .INIT ( 4'h8 ) ) \ctrl/seq6/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 (\ctrl/seq6/GEN[2].SFF/Q_839 ), .I1 (nReset_407), .O (\ctrl/seq6/GEN[3].SFF/QD ) ) ;
    LUT2 #( .INIT ( 4'hD ) ) \ctrl/seq6/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 (nReset_407), .I1 (\ctrl/seq6/GEN[1].SFF/Q_838 ), .O (\ctrl/seq6/GEN[2].SFF/QD ) ) ;
    LUT2 #( .INIT ( 4'h8 ) ) \ctrl/seq6/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 (\ctrl/seq6/GEN[0].SFF/Q_841 ), .I1 (nReset_407), .O (\ctrl/seq6/GEN[1].SFF/QD ) ) ;
    LUT3 #( .INIT ( 8'h9F ) ) \ctrl/seq6/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 (\ctrl/seq6/GEN[4].SFF/Q_842 ), .I1 (\ctrl/seq6/GEN[0].SFF/Q_841 ), .I2 (nReset_407), .O (\ctrl/seq6/GEN[0].SFF/QD ) ) ;
    LUT2 #( .INIT ( 4'h8 ) ) \ctrl/selMC1 ( .I0 (\ctrl/CSselMC_835 ), .I1 (nReset_407), .O (selMC) ) ;
    LUT2 #( .INIT ( 4'h6 ) ) \calcRCon/Mxor_MSB_s_current_state[0]_XOR_21_o_xo<0>1 ( .I0 (\calcRCon/s_current_state [0]), .I1 (\calcRCon/s_current_state [7]), .O (\calcRCon/MSB_s_current_state[0]_XOR_21_o ) ) ;
    LUT2 #( .INIT ( 4'h6 ) ) \calcRCon/Mxor_MSB_s_current_state[3]_XOR_19_o_xo<0>1 ( .I0 (\calcRCon/s_current_state [3]), .I1 (\calcRCon/s_current_state [7]), .O (\calcRCon/MSB_s_current_state[3]_XOR_19_o ) ) ;
    LUT2 #( .INIT ( 4'h6 ) ) \calcRCon/Mxor_MSB_s_current_state[2]_XOR_20_o_xo<0>1 ( .I0 (\calcRCon/s_current_state [2]), .I1 (\calcRCon/s_current_state [7]), .O (\calcRCon/MSB_s_current_state[2]_XOR_20_o ) ) ;
    LUT4 #( .INIT ( 16'h8000 ) ) \calcRCon/final<1>1 ( .I0 (\calcRCon/s_current_state [1]), .I1 (\calcRCon/s_current_state [2]), .I2 (\calcRCon/s_current_state [4]), .I3 (\calcRCon/s_current_state [5]), .O (intFinal) ) ;
    LUT2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \MUX_StateInMC/gen_mux[0].mux_inst/Mmux_Q1_SW0 ( .I0 ({ciphertext_s1[127], ciphertext_s0[127]}), .I1 ({ciphertext_s1[88], ciphertext_s0[88]}), .O ({new_AGEMA_signal_1374, N01}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \MUX_StateInMC/gen_mux[0].mux_inst/Mmux_Q1 ( .I0 ({1'b0, intFinal}), .I1 ({ciphertext_s1[24], ciphertext_s0[24]}), .I2 ({ciphertext_s1[120], ciphertext_s0[120]}), .I3 ({ciphertext_s1[56], ciphertext_s0[56]}), .I4 ({ciphertext_s1[31], ciphertext_s0[31]}), .I5 ({new_AGEMA_signal_1374, N01}), .O ({new_AGEMA_signal_1893, StateInMC[0]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \MUX_StateInMC/gen_mux[1].mux_inst/Mmux_Q1_SW0 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[31], ciphertext_s0[31]}), .I2 ({ciphertext_s1[127], ciphertext_s0[127]}), .I3 ({ciphertext_s1[24], ciphertext_s0[24]}), .O ({new_AGEMA_signal_1377, N2}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \MUX_StateInMC/gen_mux[1].mux_inst/Mmux_Q1 ( .I0 ({1'b0, intFinal}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[57], ciphertext_s0[57]}), .I3 ({ciphertext_s1[121], ciphertext_s0[121]}), .I4 ({ciphertext_s1[89], ciphertext_s0[89]}), .I5 ({new_AGEMA_signal_1377, N2}), .O ({new_AGEMA_signal_1894, StateInMC[1]}) ) ;
    LUT2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \MUX_StateInMC/gen_mux[2].mux_inst/Mmux_Q1_SW0 ( .I0 ({ciphertext_s1[90], ciphertext_s0[90]}), .I1 ({ciphertext_s1[58], ciphertext_s0[58]}), .O ({new_AGEMA_signal_1380, N4}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \MUX_StateInMC/gen_mux[2].mux_inst/Mmux_Q1 ( .I0 ({1'b0, intFinal}), .I1 ({ciphertext_s1[26], ciphertext_s0[26]}), .I2 ({ciphertext_s1[121], ciphertext_s0[121]}), .I3 ({ciphertext_s1[25], ciphertext_s0[25]}), .I4 ({ciphertext_s1[122], ciphertext_s0[122]}), .I5 ({new_AGEMA_signal_1380, N4}), .O ({new_AGEMA_signal_1895, StateInMC[2]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \MUX_StateInMC/gen_mux[3].mux_inst/Mmux_Q1_SW0 ( .I0 ({ciphertext_s1[122], ciphertext_s0[122]}), .I1 ({ciphertext_s1[31], ciphertext_s0[31]}), .I2 ({ciphertext_s1[127], ciphertext_s0[127]}), .I3 ({ciphertext_s1[26], ciphertext_s0[26]}), .O ({new_AGEMA_signal_1382, N6}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \MUX_StateInMC/gen_mux[3].mux_inst/Mmux_Q1 ( .I0 ({1'b0, intFinal}), .I1 ({ciphertext_s1[27], ciphertext_s0[27]}), .I2 ({ciphertext_s1[123], ciphertext_s0[123]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[59], ciphertext_s0[59]}), .I5 ({new_AGEMA_signal_1382, N6}), .O ({new_AGEMA_signal_1896, StateInMC[3]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \MUX_StateInMC/gen_mux[4].mux_inst/Mmux_Q1_SW0 ( .I0 ({ciphertext_s1[92], ciphertext_s0[92]}), .I1 ({ciphertext_s1[60], ciphertext_s0[60]}), .I2 ({ciphertext_s1[31], ciphertext_s0[31]}), .I3 ({ciphertext_s1[127], ciphertext_s0[127]}), .O ({new_AGEMA_signal_1385, N8}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \MUX_StateInMC/gen_mux[4].mux_inst/Mmux_Q1 ( .I0 ({1'b0, intFinal}), .I1 ({ciphertext_s1[28], ciphertext_s0[28]}), .I2 ({ciphertext_s1[27], ciphertext_s0[27]}), .I3 ({ciphertext_s1[124], ciphertext_s0[124]}), .I4 ({ciphertext_s1[123], ciphertext_s0[123]}), .I5 ({new_AGEMA_signal_1385, N8}), .O ({new_AGEMA_signal_1897, StateInMC[4]}) ) ;
    LUT2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \MUX_StateInMC/gen_mux[5].mux_inst/Mmux_Q1_SW0 ( .I0 ({ciphertext_s1[93], ciphertext_s0[93]}), .I1 ({ciphertext_s1[61], ciphertext_s0[61]}), .O ({new_AGEMA_signal_1388, N10}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \MUX_StateInMC/gen_mux[5].mux_inst/Mmux_Q1 ( .I0 ({1'b0, intFinal}), .I1 ({ciphertext_s1[29], ciphertext_s0[29]}), .I2 ({ciphertext_s1[28], ciphertext_s0[28]}), .I3 ({ciphertext_s1[124], ciphertext_s0[124]}), .I4 ({ciphertext_s1[125], ciphertext_s0[125]}), .I5 ({new_AGEMA_signal_1388, N10}), .O ({new_AGEMA_signal_1898, StateInMC[5]}) ) ;
    LUT2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \MUX_StateInMC/gen_mux[6].mux_inst/Mmux_Q1_SW0 ( .I0 ({ciphertext_s1[94], ciphertext_s0[94]}), .I1 ({ciphertext_s1[62], ciphertext_s0[62]}), .O ({new_AGEMA_signal_1391, N12}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \MUX_StateInMC/gen_mux[6].mux_inst/Mmux_Q1 ( .I0 ({1'b0, intFinal}), .I1 ({ciphertext_s1[30], ciphertext_s0[30]}), .I2 ({ciphertext_s1[125], ciphertext_s0[125]}), .I3 ({ciphertext_s1[29], ciphertext_s0[29]}), .I4 ({ciphertext_s1[126], ciphertext_s0[126]}), .I5 ({new_AGEMA_signal_1391, N12}), .O ({new_AGEMA_signal_1899, StateInMC[6]}) ) ;
    LUT2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \MUX_StateInMC/gen_mux[7].mux_inst/Mmux_Q1_SW0 ( .I0 ({ciphertext_s1[95], ciphertext_s0[95]}), .I1 ({ciphertext_s1[63], ciphertext_s0[63]}), .O ({new_AGEMA_signal_1394, N14}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \MUX_StateInMC/gen_mux[7].mux_inst/Mmux_Q1 ( .I0 ({1'b0, intFinal}), .I1 ({ciphertext_s1[31], ciphertext_s0[31]}), .I2 ({ciphertext_s1[30], ciphertext_s0[30]}), .I3 ({ciphertext_s1[127], ciphertext_s0[127]}), .I4 ({ciphertext_s1[126], ciphertext_s0[126]}), .I5 ({new_AGEMA_signal_1394, N14}), .O ({new_AGEMA_signal_1900, StateInMC[7]}) ) ;
    LUT4 #( .INIT ( 16'h7FFF ) ) intselXOR_SW0 ( .I0 (\calcRCon/s_current_state [2]), .I1 (\calcRCon/s_current_state [7]), .I2 (\calcRCon/s_current_state [3]), .I3 (\calcRCon/s_current_state [0]), .O (N16) ) ;
    LUT6 #( .INIT ( 64'hFFFFFFFE00000000 ) ) intselXOR ( .I0 (\calcRCon/s_current_state [6]), .I1 (\calcRCon/s_current_state [4]), .I2 (\calcRCon/s_current_state [5]), .I3 (\calcRCon/s_current_state [1]), .I4 (N16), .I5 (selXOR), .O (intselXOR_425) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({ciphertext_s1[127], ciphertext_s0[127]}), .I1 ({ciphertext_s1[56], ciphertext_s0[56]}), .I2 ({ciphertext_s1[24], ciphertext_s0[24]}), .O ({new_AGEMA_signal_1396, \stateArray/S03reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q1 }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hFAFAD2785050D278 ) , .MASK ( 6'b010001 ), .INIT2 ( 64'hFAFAD2785050D278 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q12 ( .I0 ({1'b0, selMC}), .I1 ({new_AGEMA_signal_1396, \stateArray/S03reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q1 }), .I2 ({ciphertext_s1[88], ciphertext_s0[88]}), .I3 ({ciphertext_s1[95], ciphertext_s0[95]}), .I4 ({1'b0, intFinal}), .I5 ({ciphertext_s1[120], ciphertext_s0[120]}), .O ({new_AGEMA_signal_1901, \stateArray/S03reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11_897 }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({ciphertext_s1[121], ciphertext_s0[121]}), .I1 ({ciphertext_s1[26], ciphertext_s0[26]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .O ({new_AGEMA_signal_1397, \stateArray/S03reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q1 }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hFAFAD2785050D278 ) , .MASK ( 6'b010001 ), .INIT2 ( 64'hFAFAD2785050D278 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q12 ( .I0 ({1'b0, selMC}), .I1 ({new_AGEMA_signal_1397, \stateArray/S03reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q1 }), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[89], ciphertext_s0[89]}), .I4 ({1'b0, intFinal}), .I5 ({ciphertext_s1[122], ciphertext_s0[122]}), .O ({new_AGEMA_signal_1902, \stateArray/S03reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11_900 }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({ciphertext_s1[124], ciphertext_s0[124]}), .I1 ({ciphertext_s1[29], ciphertext_s0[29]}), .I2 ({ciphertext_s1[61], ciphertext_s0[61]}), .O ({new_AGEMA_signal_1399, \stateArray/S03reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q1 }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hFAFAD2785050D278 ) , .MASK ( 6'b010001 ), .INIT2 ( 64'hFAFAD2785050D278 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q12 ( .I0 ({1'b0, selMC}), .I1 ({new_AGEMA_signal_1399, \stateArray/S03reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q1 }), .I2 ({ciphertext_s1[93], ciphertext_s0[93]}), .I3 ({ciphertext_s1[92], ciphertext_s0[92]}), .I4 ({1'b0, intFinal}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .O ({new_AGEMA_signal_1903, \stateArray/S03reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11_904 }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({ciphertext_s1[125], ciphertext_s0[125]}), .I1 ({ciphertext_s1[30], ciphertext_s0[30]}), .I2 ({ciphertext_s1[62], ciphertext_s0[62]}), .O ({new_AGEMA_signal_1401, \stateArray/S03reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q1 }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hFAFAD2785050D278 ) , .MASK ( 6'b010001 ), .INIT2 ( 64'hFAFAD2785050D278 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q12 ( .I0 ({1'b0, selMC}), .I1 ({new_AGEMA_signal_1401, \stateArray/S03reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q1 }), .I2 ({ciphertext_s1[94], ciphertext_s0[94]}), .I3 ({ciphertext_s1[93], ciphertext_s0[93]}), .I4 ({1'b0, intFinal}), .I5 ({ciphertext_s1[126], ciphertext_s0[126]}), .O ({new_AGEMA_signal_1904, \stateArray/S03reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11_906 }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({ciphertext_s1[126], ciphertext_s0[126]}), .I1 ({ciphertext_s1[31], ciphertext_s0[31]}), .I2 ({ciphertext_s1[63], ciphertext_s0[63]}), .O ({new_AGEMA_signal_1402, \stateArray/S03reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q1 }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hFAFAD2785050D278 ) , .MASK ( 6'b010001 ), .INIT2 ( 64'hFAFAD2785050D278 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q12 ( .I0 ({1'b0, selMC}), .I1 ({new_AGEMA_signal_1402, \stateArray/S03reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q1 }), .I2 ({ciphertext_s1[95], ciphertext_s0[95]}), .I3 ({ciphertext_s1[94], ciphertext_s0[94]}), .I4 ({1'b0, intFinal}), .I5 ({ciphertext_s1[127], ciphertext_s0[127]}), .O ({new_AGEMA_signal_1905, \stateArray/S03reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11_908 }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({ciphertext_s1[95], ciphertext_s0[95]}), .I1 ({ciphertext_s1[120], ciphertext_s0[120]}), .I2 ({ciphertext_s1[24], ciphertext_s0[24]}), .O ({new_AGEMA_signal_1403, \stateArray/S13reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q1 }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hFAFAD2785050D278 ) , .MASK ( 6'b010001 ), .INIT2 ( 64'hFAFAD2785050D278 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q12 ( .I0 ({1'b0, selMC}), .I1 ({new_AGEMA_signal_1403, \stateArray/S13reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q1 }), .I2 ({ciphertext_s1[56], ciphertext_s0[56]}), .I3 ({ciphertext_s1[63], ciphertext_s0[63]}), .I4 ({1'b0, intFinal}), .I5 ({ciphertext_s1[88], ciphertext_s0[88]}), .O ({new_AGEMA_signal_1906, \stateArray/S13reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11_910 }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({ciphertext_s1[122], ciphertext_s0[122]}), .I1 ({ciphertext_s1[26], ciphertext_s0[26]}), .I2 ({ciphertext_s1[89], ciphertext_s0[89]}), .O ({new_AGEMA_signal_1405, \stateArray/S13reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q1 }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hFAFAD2785050D278 ) , .MASK ( 6'b010001 ), .INIT2 ( 64'hFAFAD2785050D278 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q12 ( .I0 ({1'b0, selMC}), .I1 ({new_AGEMA_signal_1405, \stateArray/S13reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q1 }), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[57], ciphertext_s0[57]}), .I4 ({1'b0, intFinal}), .I5 ({ciphertext_s1[90], ciphertext_s0[90]}), .O ({new_AGEMA_signal_1907, \stateArray/S13reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11_913 }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({ciphertext_s1[125], ciphertext_s0[125]}), .I1 ({ciphertext_s1[29], ciphertext_s0[29]}), .I2 ({ciphertext_s1[92], ciphertext_s0[92]}), .O ({new_AGEMA_signal_1406, \stateArray/S13reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q1 }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hFAFAD2785050D278 ) , .MASK ( 6'b010001 ), .INIT2 ( 64'hFAFAD2785050D278 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q12 ( .I0 ({1'b0, selMC}), .I1 ({new_AGEMA_signal_1406, \stateArray/S13reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q1 }), .I2 ({ciphertext_s1[61], ciphertext_s0[61]}), .I3 ({ciphertext_s1[60], ciphertext_s0[60]}), .I4 ({1'b0, intFinal}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .O ({new_AGEMA_signal_1908, \stateArray/S13reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11_917 }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({ciphertext_s1[126], ciphertext_s0[126]}), .I1 ({ciphertext_s1[30], ciphertext_s0[30]}), .I2 ({ciphertext_s1[93], ciphertext_s0[93]}), .O ({new_AGEMA_signal_1407, \stateArray/S13reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q1 }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hFAFAD2785050D278 ) , .MASK ( 6'b010001 ), .INIT2 ( 64'hFAFAD2785050D278 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q12 ( .I0 ({1'b0, selMC}), .I1 ({new_AGEMA_signal_1407, \stateArray/S13reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q1 }), .I2 ({ciphertext_s1[62], ciphertext_s0[62]}), .I3 ({ciphertext_s1[61], ciphertext_s0[61]}), .I4 ({1'b0, intFinal}), .I5 ({ciphertext_s1[94], ciphertext_s0[94]}), .O ({new_AGEMA_signal_1909, \stateArray/S13reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11_919 }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({ciphertext_s1[127], ciphertext_s0[127]}), .I1 ({ciphertext_s1[31], ciphertext_s0[31]}), .I2 ({ciphertext_s1[94], ciphertext_s0[94]}), .O ({new_AGEMA_signal_1408, \stateArray/S13reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q1 }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hFAFAD2785050D278 ) , .MASK ( 6'b010001 ), .INIT2 ( 64'hFAFAD2785050D278 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q12 ( .I0 ({1'b0, selMC}), .I1 ({new_AGEMA_signal_1408, \stateArray/S13reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q1 }), .I2 ({ciphertext_s1[63], ciphertext_s0[63]}), .I3 ({ciphertext_s1[62], ciphertext_s0[62]}), .I4 ({1'b0, intFinal}), .I5 ({ciphertext_s1[95], ciphertext_s0[95]}), .O ({new_AGEMA_signal_1910, \stateArray/S13reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11_921 }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[120], ciphertext_s0[120]}), .I2 ({ciphertext_s1[63], ciphertext_s0[63]}), .O ({new_AGEMA_signal_1409, \stateArray/S23reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q1 }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hFAFAD2785050D278 ) , .MASK ( 6'b010001 ), .INIT2 ( 64'hFAFAD2785050D278 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q12 ( .I0 ({1'b0, selMC}), .I1 ({new_AGEMA_signal_1409, \stateArray/S23reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q1 }), .I2 ({ciphertext_s1[24], ciphertext_s0[24]}), .I3 ({ciphertext_s1[31], ciphertext_s0[31]}), .I4 ({1'b0, intFinal}), .I5 ({ciphertext_s1[56], ciphertext_s0[56]}), .O ({new_AGEMA_signal_1911, \stateArray/S23reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11_923 }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({ciphertext_s1[122], ciphertext_s0[122]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .O ({new_AGEMA_signal_1411, \stateArray/S23reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q1 }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hFAFAD2785050D278 ) , .MASK ( 6'b010001 ), .INIT2 ( 64'hFAFAD2785050D278 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q12 ( .I0 ({1'b0, selMC}), .I1 ({new_AGEMA_signal_1411, \stateArray/S23reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q1 }), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[25], ciphertext_s0[25]}), .I4 ({1'b0, intFinal}), .I5 ({ciphertext_s1[58], ciphertext_s0[58]}), .O ({new_AGEMA_signal_1912, \stateArray/S23reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11_926 }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({ciphertext_s1[93], ciphertext_s0[93]}), .I1 ({ciphertext_s1[125], ciphertext_s0[125]}), .I2 ({ciphertext_s1[60], ciphertext_s0[60]}), .O ({new_AGEMA_signal_1412, \stateArray/S23reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q1 }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hFAFAD2785050D278 ) , .MASK ( 6'b010001 ), .INIT2 ( 64'hFAFAD2785050D278 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q12 ( .I0 ({1'b0, selMC}), .I1 ({new_AGEMA_signal_1412, \stateArray/S23reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q1 }), .I2 ({ciphertext_s1[29], ciphertext_s0[29]}), .I3 ({ciphertext_s1[28], ciphertext_s0[28]}), .I4 ({1'b0, intFinal}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .O ({new_AGEMA_signal_1913, \stateArray/S23reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11_930 }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({ciphertext_s1[94], ciphertext_s0[94]}), .I1 ({ciphertext_s1[126], ciphertext_s0[126]}), .I2 ({ciphertext_s1[61], ciphertext_s0[61]}), .O ({new_AGEMA_signal_1413, \stateArray/S23reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q1 }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hFAFAD2785050D278 ) , .MASK ( 6'b010001 ), .INIT2 ( 64'hFAFAD2785050D278 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q12 ( .I0 ({1'b0, selMC}), .I1 ({new_AGEMA_signal_1413, \stateArray/S23reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q1 }), .I2 ({ciphertext_s1[30], ciphertext_s0[30]}), .I3 ({ciphertext_s1[29], ciphertext_s0[29]}), .I4 ({1'b0, intFinal}), .I5 ({ciphertext_s1[62], ciphertext_s0[62]}), .O ({new_AGEMA_signal_1914, \stateArray/S23reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11_932 }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({ciphertext_s1[95], ciphertext_s0[95]}), .I1 ({ciphertext_s1[127], ciphertext_s0[127]}), .I2 ({ciphertext_s1[62], ciphertext_s0[62]}), .O ({new_AGEMA_signal_1414, \stateArray/S23reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q1 }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hFAFAD2785050D278 ) , .MASK ( 6'b010001 ), .INIT2 ( 64'hFAFAD2785050D278 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q12 ( .I0 ({1'b0, selMC}), .I1 ({new_AGEMA_signal_1414, \stateArray/S23reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q1 }), .I2 ({ciphertext_s1[31], ciphertext_s0[31]}), .I3 ({ciphertext_s1[30], ciphertext_s0[30]}), .I4 ({1'b0, intFinal}), .I5 ({ciphertext_s1[63], ciphertext_s0[63]}), .O ({new_AGEMA_signal_1915, \stateArray/S23reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11_934 }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h95 ) , .MASK ( 3'b110 ), .INIT2 ( 8'hAA ) ) \KeyArray/S30reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_1371, \KeyArray/S00reg/gen_ff[1].gff/GEN[0].SFF/Q_401 }), .I1 ({1'b0, \calcRCon/s_current_state [0]}), .I2 ({1'b0, \ctrl/CSenRC_405 }), .O ({new_AGEMA_signal_1415, N18}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h95 ) , .MASK ( 3'b110 ), .INIT2 ( 8'hAA ) ) \KeyArray/S30reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_1368, \KeyArray/S00reg/gen_ff[1].gff/GEN[1].SFF/Q_400 }), .I1 ({1'b0, \calcRCon/s_current_state [1]}), .I2 ({1'b0, \ctrl/CSenRC_405 }), .O ({new_AGEMA_signal_1416, N20}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h95 ) , .MASK ( 3'b110 ), .INIT2 ( 8'hAA ) ) \KeyArray/S30reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_1365, \KeyArray/S00reg/gen_ff[1].gff/GEN[2].SFF/Q_399 }), .I1 ({1'b0, \calcRCon/s_current_state [2]}), .I2 ({1'b0, \ctrl/CSenRC_405 }), .O ({new_AGEMA_signal_1417, N22}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h95 ) , .MASK ( 3'b110 ), .INIT2 ( 8'hAA ) ) \KeyArray/S30reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_1362, \KeyArray/S00reg/gen_ff[1].gff/GEN[3].SFF/Q_398 }), .I1 ({1'b0, \calcRCon/s_current_state [3]}), .I2 ({1'b0, \ctrl/CSenRC_405 }), .O ({new_AGEMA_signal_1418, N24}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h95 ) , .MASK ( 3'b110 ), .INIT2 ( 8'hAA ) ) \KeyArray/S30reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_1359, \KeyArray/S00reg/gen_ff[1].gff/GEN[4].SFF/Q_397 }), .I1 ({1'b0, \calcRCon/s_current_state [4]}), .I2 ({1'b0, \ctrl/CSenRC_405 }), .O ({new_AGEMA_signal_1419, N26}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h95 ) , .MASK ( 3'b110 ), .INIT2 ( 8'hAA ) ) \KeyArray/S30reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_1356, \KeyArray/S00reg/gen_ff[1].gff/GEN[5].SFF/Q_396 }), .I1 ({1'b0, \calcRCon/s_current_state [5]}), .I2 ({1'b0, \ctrl/CSenRC_405 }), .O ({new_AGEMA_signal_1420, N28}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h95 ) , .MASK ( 3'b110 ), .INIT2 ( 8'hAA ) ) \KeyArray/S30reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_1353, \KeyArray/S00reg/gen_ff[1].gff/GEN[6].SFF/Q_395 }), .I1 ({1'b0, \calcRCon/s_current_state [6]}), .I2 ({1'b0, \ctrl/CSenRC_405 }), .O ({new_AGEMA_signal_1421, N30}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h95 ) , .MASK ( 3'b110 ), .INIT2 ( 8'hAA ) ) \KeyArray/S30reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_1350, \KeyArray/S00reg/gen_ff[1].gff/GEN[7].SFF/Q_394 }), .I1 ({1'b0, \calcRCon/s_current_state [7]}), .I2 ({1'b0, \ctrl/CSenRC_405 }), .O ({new_AGEMA_signal_1422, N32}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hAA3C3C3C ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hAA3C3C3C ) ) \SboxIn<5>1 ( .I0 ({new_AGEMA_signal_1423, \KeyArray/S13reg/gen_ff[1].gff/GEN[5].SFF/Q_388 }), .I1 ({new_AGEMA_signal_1356, \KeyArray/S00reg/gen_ff[1].gff/GEN[5].SFF/Q_396 }), .I2 ({ciphertext_s1[125], ciphertext_s0[125]}), .I3 ({1'b0, \ctrl/CSselMC_1_1342 }), .I4 ({1'b0, nReset_1_1341}), .O ({new_AGEMA_signal_1424, SboxIn[5]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hAA3C3C3C ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hAA3C3C3C ) ) \SboxIn<4>1 ( .I0 ({new_AGEMA_signal_1425, \KeyArray/S13reg/gen_ff[1].gff/GEN[4].SFF/Q_389 }), .I1 ({new_AGEMA_signal_1359, \KeyArray/S00reg/gen_ff[1].gff/GEN[4].SFF/Q_397 }), .I2 ({ciphertext_s1[124], ciphertext_s0[124]}), .I3 ({1'b0, \ctrl/CSselMC_1_1342 }), .I4 ({1'b0, nReset_1_1341}), .O ({new_AGEMA_signal_1426, SboxIn[4]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hAA3C3C3C ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hAA3C3C3C ) ) \SboxIn<3>1 ( .I0 ({new_AGEMA_signal_1427, \KeyArray/S13reg/gen_ff[1].gff/GEN[3].SFF/Q_390 }), .I1 ({new_AGEMA_signal_1362, \KeyArray/S00reg/gen_ff[1].gff/GEN[3].SFF/Q_398 }), .I2 ({ciphertext_s1[123], ciphertext_s0[123]}), .I3 ({1'b0, \ctrl/CSselMC_1_1342 }), .I4 ({1'b0, nReset_1_1341}), .O ({new_AGEMA_signal_1428, SboxIn[3]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hAA3C3C3C ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hAA3C3C3C ) ) \SboxIn<2>1 ( .I0 ({new_AGEMA_signal_1429, \KeyArray/S13reg/gen_ff[1].gff/GEN[2].SFF/Q_391 }), .I1 ({new_AGEMA_signal_1365, \KeyArray/S00reg/gen_ff[1].gff/GEN[2].SFF/Q_399 }), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({1'b0, \ctrl/CSselMC_1_1342 }), .I4 ({1'b0, nReset_1_1341}), .O ({new_AGEMA_signal_1430, SboxIn[2]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hAA3C3C3C ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hAA3C3C3C ) ) \SboxIn<1>1 ( .I0 ({new_AGEMA_signal_1431, \KeyArray/S13reg/gen_ff[1].gff/GEN[1].SFF/Q_392 }), .I1 ({new_AGEMA_signal_1368, \KeyArray/S00reg/gen_ff[1].gff/GEN[1].SFF/Q_400 }), .I2 ({ciphertext_s1[121], ciphertext_s0[121]}), .I3 ({1'b0, \ctrl/CSselMC_1_1342 }), .I4 ({1'b0, nReset_1_1341}), .O ({new_AGEMA_signal_1432, SboxIn[1]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hAA3C3C3C ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hAA3C3C3C ) ) \SboxIn<0>1 ( .I0 ({new_AGEMA_signal_1433, \KeyArray/S13reg/gen_ff[1].gff/GEN[0].SFF/Q_393 }), .I1 ({new_AGEMA_signal_1371, \KeyArray/S00reg/gen_ff[1].gff/GEN[0].SFF/Q_401 }), .I2 ({ciphertext_s1[120], ciphertext_s0[120]}), .I3 ({1'b0, \ctrl/CSselMC_1_1342 }), .I4 ({1'b0, nReset_1_1341}), .O ({new_AGEMA_signal_1434, SboxIn[0]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hAA3C3C3C ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hAA3C3C3C ) ) \SboxIn<7>1 ( .I0 ({new_AGEMA_signal_1435, \KeyArray/S13reg/gen_ff[1].gff/GEN[7].SFF/Q_386 }), .I1 ({new_AGEMA_signal_1350, \KeyArray/S00reg/gen_ff[1].gff/GEN[7].SFF/Q_394 }), .I2 ({ciphertext_s1[127], ciphertext_s0[127]}), .I3 ({1'b0, \ctrl/CSselMC_835 }), .I4 ({1'b0, nReset_407}), .O ({new_AGEMA_signal_1436, SboxIn[7]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hAA3C3C3C ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hAA3C3C3C ) ) \SboxIn<6>1 ( .I0 ({new_AGEMA_signal_1437, \KeyArray/S13reg/gen_ff[1].gff/GEN[6].SFF/Q_387 }), .I1 ({new_AGEMA_signal_1353, \KeyArray/S00reg/gen_ff[1].gff/GEN[6].SFF/Q_395 }), .I2 ({ciphertext_s1[126], ciphertext_s0[126]}), .I3 ({1'b0, \ctrl/CSselMC_835 }), .I4 ({1'b0, nReset_407}), .O ({new_AGEMA_signal_1438, SboxIn[6]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'hBF80 ) , .MASK ( 4'b0110 ), .INIT2 ( 16'hBF80 ) ) \KeyArray/S00reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({new_AGEMA_signal_1589, \KeyArray/S10reg/gen_ff[1].gff/GEN[0].SFF/Q_667 }), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, nReset_407}), .I3 ({new_AGEMA_signal_2156, \KeyArray/inS00ser [0]}), .O ({new_AGEMA_signal_2237, \KeyArray/S00reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'hBF80 ) , .MASK ( 4'b0110 ), .INIT2 ( 16'hBF80 ) ) \KeyArray/S00reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({new_AGEMA_signal_1592, \KeyArray/S10reg/gen_ff[1].gff/GEN[1].SFF/Q_668 }), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, nReset_407}), .I3 ({new_AGEMA_signal_2154, \KeyArray/inS00ser [1]}), .O ({new_AGEMA_signal_2238, \KeyArray/S00reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'hBF80 ) , .MASK ( 4'b0110 ), .INIT2 ( 16'hBF80 ) ) \KeyArray/S00reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({new_AGEMA_signal_1595, \KeyArray/S10reg/gen_ff[1].gff/GEN[2].SFF/Q_669 }), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, nReset_407}), .I3 ({new_AGEMA_signal_2152, \KeyArray/inS00ser [2]}), .O ({new_AGEMA_signal_2239, \KeyArray/S00reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'hBF80 ) , .MASK ( 4'b0110 ), .INIT2 ( 16'hBF80 ) ) \KeyArray/S00reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({new_AGEMA_signal_1598, \KeyArray/S10reg/gen_ff[1].gff/GEN[3].SFF/Q_670 }), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, nReset_407}), .I3 ({new_AGEMA_signal_2150, \KeyArray/inS00ser [3]}), .O ({new_AGEMA_signal_2240, \KeyArray/S00reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'hBF80 ) , .MASK ( 4'b0110 ), .INIT2 ( 16'hBF80 ) ) \KeyArray/S00reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({new_AGEMA_signal_1601, \KeyArray/S10reg/gen_ff[1].gff/GEN[4].SFF/Q_671 }), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, nReset_407}), .I3 ({new_AGEMA_signal_2148, \KeyArray/inS00ser [4]}), .O ({new_AGEMA_signal_2241, \KeyArray/S00reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'hBF80 ) , .MASK ( 4'b0110 ), .INIT2 ( 16'hBF80 ) ) \KeyArray/S00reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({new_AGEMA_signal_1604, \KeyArray/S10reg/gen_ff[1].gff/GEN[5].SFF/Q_672 }), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, nReset_407}), .I3 ({new_AGEMA_signal_2146, \KeyArray/inS00ser [5]}), .O ({new_AGEMA_signal_2242, \KeyArray/S00reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'hBF80 ) , .MASK ( 4'b0110 ), .INIT2 ( 16'hBF80 ) ) \KeyArray/S00reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({new_AGEMA_signal_1607, \KeyArray/S10reg/gen_ff[1].gff/GEN[6].SFF/Q_673 }), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, nReset_407}), .I3 ({new_AGEMA_signal_2144, \KeyArray/inS00ser [6]}), .O ({new_AGEMA_signal_2243, \KeyArray/S00reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'hBF80 ) , .MASK ( 4'b0110 ), .INIT2 ( 16'hBF80 ) ) \KeyArray/S00reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({new_AGEMA_signal_1610, \KeyArray/S10reg/gen_ff[1].gff/GEN[7].SFF/Q_674 }), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, nReset_407}), .I3 ({new_AGEMA_signal_2142, \KeyArray/inS00ser [7]}), .O ({new_AGEMA_signal_2244, \KeyArray/S00reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q13_SW0 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[127], ciphertext_s0[127]}), .I2 ({ciphertext_s1[88], ciphertext_s0[88]}), .I3 ({ciphertext_s1[95], ciphertext_s0[95]}), .I4 ({ciphertext_s1[57], ciphertext_s0[57]}), .I5 ({ciphertext_s1[25], ciphertext_s0[25]}), .O ({new_AGEMA_signal_1440, N34}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hE6EAAAAA262AAAAA ) , .MASK ( 6'b010110 ), .INIT2 ( 64'hE6EAAAAA262AAAAA ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q13 ( .I0 ({ciphertext_s1[89], ciphertext_s0[89]}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, intFinal}), .I3 ({new_AGEMA_signal_1440, N34}), .I4 ({1'b0, nReset_407}), .I5 ({ciphertext_s1[121], ciphertext_s0[121]}), .O ({new_AGEMA_signal_1916, \stateArray/S03reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q12 }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q13_SW0 ( .I0 ({ciphertext_s1[122], ciphertext_s0[122]}), .I1 ({ciphertext_s1[127], ciphertext_s0[127]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[95], ciphertext_s0[95]}), .I4 ({ciphertext_s1[59], ciphertext_s0[59]}), .I5 ({ciphertext_s1[27], ciphertext_s0[27]}), .O ({new_AGEMA_signal_1443, N36}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hE6EAAAAA262AAAAA ) , .MASK ( 6'b010110 ), .INIT2 ( 64'hE6EAAAAA262AAAAA ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q13 ( .I0 ({ciphertext_s1[91], ciphertext_s0[91]}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, intFinal}), .I3 ({new_AGEMA_signal_1443, N36}), .I4 ({1'b0, nReset_407}), .I5 ({ciphertext_s1[123], ciphertext_s0[123]}), .O ({new_AGEMA_signal_1917, \stateArray/S03reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q12 }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q13_SW0 ( .I0 ({ciphertext_s1[123], ciphertext_s0[123]}), .I1 ({ciphertext_s1[127], ciphertext_s0[127]}), .I2 ({ciphertext_s1[91], ciphertext_s0[91]}), .I3 ({ciphertext_s1[95], ciphertext_s0[95]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[28], ciphertext_s0[28]}), .O ({new_AGEMA_signal_1446, N38}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hE6EAAAAA262AAAAA ) , .MASK ( 6'b010110 ), .INIT2 ( 64'hE6EAAAAA262AAAAA ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q13 ( .I0 ({ciphertext_s1[92], ciphertext_s0[92]}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, intFinal}), .I3 ({new_AGEMA_signal_1446, N38}), .I4 ({1'b0, nReset_407}), .I5 ({ciphertext_s1[124], ciphertext_s0[124]}), .O ({new_AGEMA_signal_1918, \stateArray/S03reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q12 }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q13_SW0 ( .I0 ({ciphertext_s1[121], ciphertext_s0[121]}), .I1 ({ciphertext_s1[88], ciphertext_s0[88]}), .I2 ({ciphertext_s1[95], ciphertext_s0[95]}), .I3 ({ciphertext_s1[56], ciphertext_s0[56]}), .I4 ({ciphertext_s1[63], ciphertext_s0[63]}), .I5 ({ciphertext_s1[25], ciphertext_s0[25]}), .O ({new_AGEMA_signal_1447, N40}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hE6EAAAAA262AAAAA ) , .MASK ( 6'b010110 ), .INIT2 ( 64'hE6EAAAAA262AAAAA ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q13 ( .I0 ({ciphertext_s1[57], ciphertext_s0[57]}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, intFinal}), .I3 ({new_AGEMA_signal_1447, N40}), .I4 ({1'b0, nReset_407}), .I5 ({ciphertext_s1[89], ciphertext_s0[89]}), .O ({new_AGEMA_signal_1919, \stateArray/S13reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q12 }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q13_SW0 ( .I0 ({ciphertext_s1[123], ciphertext_s0[123]}), .I1 ({ciphertext_s1[90], ciphertext_s0[90]}), .I2 ({ciphertext_s1[95], ciphertext_s0[95]}), .I3 ({ciphertext_s1[58], ciphertext_s0[58]}), .I4 ({ciphertext_s1[63], ciphertext_s0[63]}), .I5 ({ciphertext_s1[27], ciphertext_s0[27]}), .O ({new_AGEMA_signal_1448, N42}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hE6EAAAAA262AAAAA ) , .MASK ( 6'b010110 ), .INIT2 ( 64'hE6EAAAAA262AAAAA ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q13 ( .I0 ({ciphertext_s1[59], ciphertext_s0[59]}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, intFinal}), .I3 ({new_AGEMA_signal_1448, N42}), .I4 ({1'b0, nReset_407}), .I5 ({ciphertext_s1[91], ciphertext_s0[91]}), .O ({new_AGEMA_signal_1920, \stateArray/S13reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q12 }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q13_SW0 ( .I0 ({ciphertext_s1[124], ciphertext_s0[124]}), .I1 ({ciphertext_s1[91], ciphertext_s0[91]}), .I2 ({ciphertext_s1[95], ciphertext_s0[95]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[63], ciphertext_s0[63]}), .I5 ({ciphertext_s1[28], ciphertext_s0[28]}), .O ({new_AGEMA_signal_1449, N44}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hE6EAAAAA262AAAAA ) , .MASK ( 6'b010110 ), .INIT2 ( 64'hE6EAAAAA262AAAAA ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q13 ( .I0 ({ciphertext_s1[60], ciphertext_s0[60]}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, intFinal}), .I3 ({new_AGEMA_signal_1449, N44}), .I4 ({1'b0, nReset_407}), .I5 ({ciphertext_s1[92], ciphertext_s0[92]}), .O ({new_AGEMA_signal_1921, \stateArray/S13reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q12 }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q13_SW0 ( .I0 ({ciphertext_s1[121], ciphertext_s0[121]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[56], ciphertext_s0[56]}), .I3 ({ciphertext_s1[63], ciphertext_s0[63]}), .I4 ({ciphertext_s1[24], ciphertext_s0[24]}), .I5 ({ciphertext_s1[31], ciphertext_s0[31]}), .O ({new_AGEMA_signal_1450, N46}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hE6EAAAAA262AAAAA ) , .MASK ( 6'b010110 ), .INIT2 ( 64'hE6EAAAAA262AAAAA ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q13 ( .I0 ({ciphertext_s1[25], ciphertext_s0[25]}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, intFinal}), .I3 ({new_AGEMA_signal_1450, N46}), .I4 ({1'b0, nReset_407}), .I5 ({ciphertext_s1[57], ciphertext_s0[57]}), .O ({new_AGEMA_signal_1922, \stateArray/S23reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q12 }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q13_SW0 ( .I0 ({ciphertext_s1[123], ciphertext_s0[123]}), .I1 ({ciphertext_s1[91], ciphertext_s0[91]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[63], ciphertext_s0[63]}), .I4 ({ciphertext_s1[26], ciphertext_s0[26]}), .I5 ({ciphertext_s1[31], ciphertext_s0[31]}), .O ({new_AGEMA_signal_1451, N48}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hE6EAAAAA262AAAAA ) , .MASK ( 6'b010110 ), .INIT2 ( 64'hE6EAAAAA262AAAAA ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q13 ( .I0 ({ciphertext_s1[27], ciphertext_s0[27]}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, intFinal}), .I3 ({new_AGEMA_signal_1451, N48}), .I4 ({1'b0, nReset_407}), .I5 ({ciphertext_s1[59], ciphertext_s0[59]}), .O ({new_AGEMA_signal_1923, \stateArray/S23reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q12 }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q13_SW0 ( .I0 ({ciphertext_s1[124], ciphertext_s0[124]}), .I1 ({ciphertext_s1[92], ciphertext_s0[92]}), .I2 ({ciphertext_s1[59], ciphertext_s0[59]}), .I3 ({ciphertext_s1[63], ciphertext_s0[63]}), .I4 ({ciphertext_s1[27], ciphertext_s0[27]}), .I5 ({ciphertext_s1[31], ciphertext_s0[31]}), .O ({new_AGEMA_signal_1452, N50}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hE6EAAAAA262AAAAA ) , .MASK ( 6'b010110 ), .INIT2 ( 64'hE6EAAAAA262AAAAA ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q13 ( .I0 ({ciphertext_s1[28], ciphertext_s0[28]}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, intFinal}), .I3 ({new_AGEMA_signal_1452, N50}), .I4 ({1'b0, nReset_407}), .I5 ({ciphertext_s1[60], ciphertext_s0[60]}), .O ({new_AGEMA_signal_1924, \stateArray/S23reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q12 }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S10reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[88], plaintext_s0[88]}), .I2 ({ciphertext_s1[80], ciphertext_s0[80]}), .O ({new_AGEMA_signal_1455, \stateArray/S10reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S10reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[89], plaintext_s0[89]}), .I2 ({ciphertext_s1[81], ciphertext_s0[81]}), .O ({new_AGEMA_signal_1458, \stateArray/S10reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S10reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[90], plaintext_s0[90]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .O ({new_AGEMA_signal_1461, \stateArray/S10reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S10reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[91], plaintext_s0[91]}), .I2 ({ciphertext_s1[83], ciphertext_s0[83]}), .O ({new_AGEMA_signal_1464, \stateArray/S10reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S10reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[92], plaintext_s0[92]}), .I2 ({ciphertext_s1[84], ciphertext_s0[84]}), .O ({new_AGEMA_signal_1467, \stateArray/S10reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S10reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[93], plaintext_s0[93]}), .I2 ({ciphertext_s1[85], ciphertext_s0[85]}), .O ({new_AGEMA_signal_1470, \stateArray/S10reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S10reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[94], plaintext_s0[94]}), .I2 ({ciphertext_s1[86], ciphertext_s0[86]}), .O ({new_AGEMA_signal_1473, \stateArray/S10reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S10reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[95], plaintext_s0[95]}), .I2 ({ciphertext_s1[87], ciphertext_s0[87]}), .O ({new_AGEMA_signal_1476, \stateArray/S10reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S11reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[80], plaintext_s0[80]}), .I2 ({ciphertext_s1[72], ciphertext_s0[72]}), .O ({new_AGEMA_signal_1479, \stateArray/S11reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S11reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[81], plaintext_s0[81]}), .I2 ({ciphertext_s1[73], ciphertext_s0[73]}), .O ({new_AGEMA_signal_1482, \stateArray/S11reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S11reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[82], plaintext_s0[82]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .O ({new_AGEMA_signal_1485, \stateArray/S11reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S11reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[83], plaintext_s0[83]}), .I2 ({ciphertext_s1[75], ciphertext_s0[75]}), .O ({new_AGEMA_signal_1488, \stateArray/S11reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S11reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[84], plaintext_s0[84]}), .I2 ({ciphertext_s1[76], ciphertext_s0[76]}), .O ({new_AGEMA_signal_1491, \stateArray/S11reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S11reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[85], plaintext_s0[85]}), .I2 ({ciphertext_s1[77], ciphertext_s0[77]}), .O ({new_AGEMA_signal_1494, \stateArray/S11reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S11reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[86], plaintext_s0[86]}), .I2 ({ciphertext_s1[78], ciphertext_s0[78]}), .O ({new_AGEMA_signal_1497, \stateArray/S11reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S11reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[87], plaintext_s0[87]}), .I2 ({ciphertext_s1[79], ciphertext_s0[79]}), .O ({new_AGEMA_signal_1500, \stateArray/S11reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S12reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[72], plaintext_s0[72]}), .I2 ({ciphertext_s1[64], ciphertext_s0[64]}), .O ({new_AGEMA_signal_1503, \stateArray/S12reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S12reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[73], plaintext_s0[73]}), .I2 ({ciphertext_s1[65], ciphertext_s0[65]}), .O ({new_AGEMA_signal_1506, \stateArray/S12reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S12reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[74], plaintext_s0[74]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .O ({new_AGEMA_signal_1509, \stateArray/S12reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S12reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[75], plaintext_s0[75]}), .I2 ({ciphertext_s1[67], ciphertext_s0[67]}), .O ({new_AGEMA_signal_1512, \stateArray/S12reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S12reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[76], plaintext_s0[76]}), .I2 ({ciphertext_s1[68], ciphertext_s0[68]}), .O ({new_AGEMA_signal_1515, \stateArray/S12reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S12reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[77], plaintext_s0[77]}), .I2 ({ciphertext_s1[69], ciphertext_s0[69]}), .O ({new_AGEMA_signal_1518, \stateArray/S12reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S12reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[78], plaintext_s0[78]}), .I2 ({ciphertext_s1[70], ciphertext_s0[70]}), .O ({new_AGEMA_signal_1521, \stateArray/S12reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S12reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[79], plaintext_s0[79]}), .I2 ({ciphertext_s1[71], ciphertext_s0[71]}), .O ({new_AGEMA_signal_1524, \stateArray/S12reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S00reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[120], ciphertext_s0[120]}), .I3 ({ciphertext_s1[112], ciphertext_s0[112]}), .I4 ({plaintext_s1[120], plaintext_s0[120]}), .O ({new_AGEMA_signal_1927, \stateArray/S00reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S00reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[121], ciphertext_s0[121]}), .I3 ({ciphertext_s1[113], ciphertext_s0[113]}), .I4 ({plaintext_s1[121], plaintext_s0[121]}), .O ({new_AGEMA_signal_1930, \stateArray/S00reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S00reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[114], ciphertext_s0[114]}), .I4 ({plaintext_s1[122], plaintext_s0[122]}), .O ({new_AGEMA_signal_1933, \stateArray/S00reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S00reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[123], ciphertext_s0[123]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({plaintext_s1[123], plaintext_s0[123]}), .O ({new_AGEMA_signal_1936, \stateArray/S00reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S00reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[124], ciphertext_s0[124]}), .I3 ({ciphertext_s1[116], ciphertext_s0[116]}), .I4 ({plaintext_s1[124], plaintext_s0[124]}), .O ({new_AGEMA_signal_1939, \stateArray/S00reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S00reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[125], ciphertext_s0[125]}), .I3 ({ciphertext_s1[117], ciphertext_s0[117]}), .I4 ({plaintext_s1[125], plaintext_s0[125]}), .O ({new_AGEMA_signal_1942, \stateArray/S00reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S00reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[126], ciphertext_s0[126]}), .I3 ({ciphertext_s1[118], ciphertext_s0[118]}), .I4 ({plaintext_s1[126], plaintext_s0[126]}), .O ({new_AGEMA_signal_1945, \stateArray/S00reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S00reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[127], ciphertext_s0[127]}), .I3 ({ciphertext_s1[119], ciphertext_s0[119]}), .I4 ({plaintext_s1[127], plaintext_s0[127]}), .O ({new_AGEMA_signal_1948, \stateArray/S00reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S01reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[112], ciphertext_s0[112]}), .I3 ({ciphertext_s1[104], ciphertext_s0[104]}), .I4 ({plaintext_s1[112], plaintext_s0[112]}), .O ({new_AGEMA_signal_1951, \stateArray/S01reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S01reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[113], ciphertext_s0[113]}), .I3 ({ciphertext_s1[105], ciphertext_s0[105]}), .I4 ({plaintext_s1[113], plaintext_s0[113]}), .O ({new_AGEMA_signal_1954, \stateArray/S01reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S01reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[106], ciphertext_s0[106]}), .I4 ({plaintext_s1[114], plaintext_s0[114]}), .O ({new_AGEMA_signal_1957, \stateArray/S01reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S01reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[115], ciphertext_s0[115]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({plaintext_s1[115], plaintext_s0[115]}), .O ({new_AGEMA_signal_1960, \stateArray/S01reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S01reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[116], ciphertext_s0[116]}), .I3 ({ciphertext_s1[108], ciphertext_s0[108]}), .I4 ({plaintext_s1[116], plaintext_s0[116]}), .O ({new_AGEMA_signal_1963, \stateArray/S01reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S01reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[117], ciphertext_s0[117]}), .I3 ({ciphertext_s1[109], ciphertext_s0[109]}), .I4 ({plaintext_s1[117], plaintext_s0[117]}), .O ({new_AGEMA_signal_1966, \stateArray/S01reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S01reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[118], ciphertext_s0[118]}), .I3 ({ciphertext_s1[110], ciphertext_s0[110]}), .I4 ({plaintext_s1[118], plaintext_s0[118]}), .O ({new_AGEMA_signal_1969, \stateArray/S01reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S01reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[119], ciphertext_s0[119]}), .I3 ({ciphertext_s1[111], ciphertext_s0[111]}), .I4 ({plaintext_s1[119], plaintext_s0[119]}), .O ({new_AGEMA_signal_1972, \stateArray/S01reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S02reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[104], ciphertext_s0[104]}), .I3 ({ciphertext_s1[96], ciphertext_s0[96]}), .I4 ({plaintext_s1[104], plaintext_s0[104]}), .O ({new_AGEMA_signal_1975, \stateArray/S02reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S02reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[105], ciphertext_s0[105]}), .I3 ({ciphertext_s1[97], ciphertext_s0[97]}), .I4 ({plaintext_s1[105], plaintext_s0[105]}), .O ({new_AGEMA_signal_1978, \stateArray/S02reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S02reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[98], ciphertext_s0[98]}), .I4 ({plaintext_s1[106], plaintext_s0[106]}), .O ({new_AGEMA_signal_1981, \stateArray/S02reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S02reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[107], ciphertext_s0[107]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({plaintext_s1[107], plaintext_s0[107]}), .O ({new_AGEMA_signal_1984, \stateArray/S02reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S02reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[108], ciphertext_s0[108]}), .I3 ({ciphertext_s1[100], ciphertext_s0[100]}), .I4 ({plaintext_s1[108], plaintext_s0[108]}), .O ({new_AGEMA_signal_1987, \stateArray/S02reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S02reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[109], ciphertext_s0[109]}), .I3 ({ciphertext_s1[101], ciphertext_s0[101]}), .I4 ({plaintext_s1[109], plaintext_s0[109]}), .O ({new_AGEMA_signal_1990, \stateArray/S02reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S02reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[110], ciphertext_s0[110]}), .I3 ({ciphertext_s1[102], ciphertext_s0[102]}), .I4 ({plaintext_s1[110], plaintext_s0[110]}), .O ({new_AGEMA_signal_1993, \stateArray/S02reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S02reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[111], ciphertext_s0[111]}), .I3 ({ciphertext_s1[103], ciphertext_s0[103]}), .I4 ({plaintext_s1[111], plaintext_s0[111]}), .O ({new_AGEMA_signal_1996, \stateArray/S02reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S20reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[40], ciphertext_s0[40]}), .I3 ({ciphertext_s1[48], ciphertext_s0[48]}), .I4 ({plaintext_s1[56], plaintext_s0[56]}), .O ({new_AGEMA_signal_2000, \stateArray/S20reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S20reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[41], ciphertext_s0[41]}), .I3 ({ciphertext_s1[49], ciphertext_s0[49]}), .I4 ({plaintext_s1[57], plaintext_s0[57]}), .O ({new_AGEMA_signal_2004, \stateArray/S20reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S20reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[50], ciphertext_s0[50]}), .I4 ({plaintext_s1[58], plaintext_s0[58]}), .O ({new_AGEMA_signal_2008, \stateArray/S20reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S20reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[43], ciphertext_s0[43]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({plaintext_s1[59], plaintext_s0[59]}), .O ({new_AGEMA_signal_2012, \stateArray/S20reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S20reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[44], ciphertext_s0[44]}), .I3 ({ciphertext_s1[52], ciphertext_s0[52]}), .I4 ({plaintext_s1[60], plaintext_s0[60]}), .O ({new_AGEMA_signal_2016, \stateArray/S20reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S20reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[45], ciphertext_s0[45]}), .I3 ({ciphertext_s1[53], ciphertext_s0[53]}), .I4 ({plaintext_s1[61], plaintext_s0[61]}), .O ({new_AGEMA_signal_2020, \stateArray/S20reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S20reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[46], ciphertext_s0[46]}), .I3 ({ciphertext_s1[54], ciphertext_s0[54]}), .I4 ({plaintext_s1[62], plaintext_s0[62]}), .O ({new_AGEMA_signal_2024, \stateArray/S20reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S20reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[47], ciphertext_s0[47]}), .I3 ({ciphertext_s1[55], ciphertext_s0[55]}), .I4 ({plaintext_s1[63], plaintext_s0[63]}), .O ({new_AGEMA_signal_2028, \stateArray/S20reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S21reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[32], ciphertext_s0[32]}), .I3 ({ciphertext_s1[40], ciphertext_s0[40]}), .I4 ({plaintext_s1[48], plaintext_s0[48]}), .O ({new_AGEMA_signal_2031, \stateArray/S21reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S21reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[33], ciphertext_s0[33]}), .I3 ({ciphertext_s1[41], ciphertext_s0[41]}), .I4 ({plaintext_s1[49], plaintext_s0[49]}), .O ({new_AGEMA_signal_2034, \stateArray/S21reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S21reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[42], ciphertext_s0[42]}), .I4 ({plaintext_s1[50], plaintext_s0[50]}), .O ({new_AGEMA_signal_2037, \stateArray/S21reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S21reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[35], ciphertext_s0[35]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({plaintext_s1[51], plaintext_s0[51]}), .O ({new_AGEMA_signal_2040, \stateArray/S21reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S21reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[36], ciphertext_s0[36]}), .I3 ({ciphertext_s1[44], ciphertext_s0[44]}), .I4 ({plaintext_s1[52], plaintext_s0[52]}), .O ({new_AGEMA_signal_2043, \stateArray/S21reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S21reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[37], ciphertext_s0[37]}), .I3 ({ciphertext_s1[45], ciphertext_s0[45]}), .I4 ({plaintext_s1[53], plaintext_s0[53]}), .O ({new_AGEMA_signal_2046, \stateArray/S21reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S21reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[38], ciphertext_s0[38]}), .I3 ({ciphertext_s1[46], ciphertext_s0[46]}), .I4 ({plaintext_s1[54], plaintext_s0[54]}), .O ({new_AGEMA_signal_2049, \stateArray/S21reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S21reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[39], ciphertext_s0[39]}), .I3 ({ciphertext_s1[47], ciphertext_s0[47]}), .I4 ({plaintext_s1[55], plaintext_s0[55]}), .O ({new_AGEMA_signal_2052, \stateArray/S21reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S22reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[56], ciphertext_s0[56]}), .I3 ({ciphertext_s1[32], ciphertext_s0[32]}), .I4 ({plaintext_s1[40], plaintext_s0[40]}), .O ({new_AGEMA_signal_2054, \stateArray/S22reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S22reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[57], ciphertext_s0[57]}), .I3 ({ciphertext_s1[33], ciphertext_s0[33]}), .I4 ({plaintext_s1[41], plaintext_s0[41]}), .O ({new_AGEMA_signal_2056, \stateArray/S22reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S22reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[34], ciphertext_s0[34]}), .I4 ({plaintext_s1[42], plaintext_s0[42]}), .O ({new_AGEMA_signal_2058, \stateArray/S22reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S22reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[59], ciphertext_s0[59]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({plaintext_s1[43], plaintext_s0[43]}), .O ({new_AGEMA_signal_2060, \stateArray/S22reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S22reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[60], ciphertext_s0[60]}), .I3 ({ciphertext_s1[36], ciphertext_s0[36]}), .I4 ({plaintext_s1[44], plaintext_s0[44]}), .O ({new_AGEMA_signal_2062, \stateArray/S22reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S22reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[61], ciphertext_s0[61]}), .I3 ({ciphertext_s1[37], ciphertext_s0[37]}), .I4 ({plaintext_s1[45], plaintext_s0[45]}), .O ({new_AGEMA_signal_2064, \stateArray/S22reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S22reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[62], ciphertext_s0[62]}), .I3 ({ciphertext_s1[38], ciphertext_s0[38]}), .I4 ({plaintext_s1[46], plaintext_s0[46]}), .O ({new_AGEMA_signal_2066, \stateArray/S22reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S22reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[63], ciphertext_s0[63]}), .I3 ({ciphertext_s1[39], ciphertext_s0[39]}), .I4 ({plaintext_s1[47], plaintext_s0[47]}), .O ({new_AGEMA_signal_2068, \stateArray/S22reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S30reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[0], ciphertext_s0[0]}), .I3 ({ciphertext_s1[16], ciphertext_s0[16]}), .I4 ({plaintext_s1[24], plaintext_s0[24]}), .O ({new_AGEMA_signal_2072, \stateArray/S30reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S30reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[1], ciphertext_s0[1]}), .I3 ({ciphertext_s1[17], ciphertext_s0[17]}), .I4 ({plaintext_s1[25], plaintext_s0[25]}), .O ({new_AGEMA_signal_2076, \stateArray/S30reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S30reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[18], ciphertext_s0[18]}), .I4 ({plaintext_s1[26], plaintext_s0[26]}), .O ({new_AGEMA_signal_2080, \stateArray/S30reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S30reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[3], ciphertext_s0[3]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({plaintext_s1[27], plaintext_s0[27]}), .O ({new_AGEMA_signal_2084, \stateArray/S30reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S30reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[4], ciphertext_s0[4]}), .I3 ({ciphertext_s1[20], ciphertext_s0[20]}), .I4 ({plaintext_s1[28], plaintext_s0[28]}), .O ({new_AGEMA_signal_2088, \stateArray/S30reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S30reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[5], ciphertext_s0[5]}), .I3 ({ciphertext_s1[21], ciphertext_s0[21]}), .I4 ({plaintext_s1[29], plaintext_s0[29]}), .O ({new_AGEMA_signal_2092, \stateArray/S30reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S30reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[6], ciphertext_s0[6]}), .I3 ({ciphertext_s1[22], ciphertext_s0[22]}), .I4 ({plaintext_s1[30], plaintext_s0[30]}), .O ({new_AGEMA_signal_2096, \stateArray/S30reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S30reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[7], ciphertext_s0[7]}), .I3 ({ciphertext_s1[23], ciphertext_s0[23]}), .I4 ({plaintext_s1[31], plaintext_s0[31]}), .O ({new_AGEMA_signal_2100, \stateArray/S30reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S31reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[24], ciphertext_s0[24]}), .I3 ({ciphertext_s1[8], ciphertext_s0[8]}), .I4 ({plaintext_s1[16], plaintext_s0[16]}), .O ({new_AGEMA_signal_2103, \stateArray/S31reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S31reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[25], ciphertext_s0[25]}), .I3 ({ciphertext_s1[9], ciphertext_s0[9]}), .I4 ({plaintext_s1[17], plaintext_s0[17]}), .O ({new_AGEMA_signal_2106, \stateArray/S31reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S31reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[10], ciphertext_s0[10]}), .I4 ({plaintext_s1[18], plaintext_s0[18]}), .O ({new_AGEMA_signal_2109, \stateArray/S31reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S31reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[27], ciphertext_s0[27]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({plaintext_s1[19], plaintext_s0[19]}), .O ({new_AGEMA_signal_2112, \stateArray/S31reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S31reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[28], ciphertext_s0[28]}), .I3 ({ciphertext_s1[12], ciphertext_s0[12]}), .I4 ({plaintext_s1[20], plaintext_s0[20]}), .O ({new_AGEMA_signal_2115, \stateArray/S31reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S31reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[29], ciphertext_s0[29]}), .I3 ({ciphertext_s1[13], ciphertext_s0[13]}), .I4 ({plaintext_s1[21], plaintext_s0[21]}), .O ({new_AGEMA_signal_2118, \stateArray/S31reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S31reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[30], ciphertext_s0[30]}), .I3 ({ciphertext_s1[14], ciphertext_s0[14]}), .I4 ({plaintext_s1[22], plaintext_s0[22]}), .O ({new_AGEMA_signal_2121, \stateArray/S31reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S31reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[31], ciphertext_s0[31]}), .I3 ({ciphertext_s1[15], ciphertext_s0[15]}), .I4 ({plaintext_s1[23], plaintext_s0[23]}), .O ({new_AGEMA_signal_2124, \stateArray/S31reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S32reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[16], ciphertext_s0[16]}), .I3 ({ciphertext_s1[0], ciphertext_s0[0]}), .I4 ({plaintext_s1[8], plaintext_s0[8]}), .O ({new_AGEMA_signal_2126, \stateArray/S32reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S32reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[17], ciphertext_s0[17]}), .I3 ({ciphertext_s1[1], ciphertext_s0[1]}), .I4 ({plaintext_s1[9], plaintext_s0[9]}), .O ({new_AGEMA_signal_2128, \stateArray/S32reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S32reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[2], ciphertext_s0[2]}), .I4 ({plaintext_s1[10], plaintext_s0[10]}), .O ({new_AGEMA_signal_2130, \stateArray/S32reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S32reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[19], ciphertext_s0[19]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({plaintext_s1[11], plaintext_s0[11]}), .O ({new_AGEMA_signal_2132, \stateArray/S32reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S32reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[20], ciphertext_s0[20]}), .I3 ({ciphertext_s1[4], ciphertext_s0[4]}), .I4 ({plaintext_s1[12], plaintext_s0[12]}), .O ({new_AGEMA_signal_2134, \stateArray/S32reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S32reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[21], ciphertext_s0[21]}), .I3 ({ciphertext_s1[5], ciphertext_s0[5]}), .I4 ({plaintext_s1[13], plaintext_s0[13]}), .O ({new_AGEMA_signal_2136, \stateArray/S32reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S32reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[22], ciphertext_s0[22]}), .I3 ({ciphertext_s1[6], ciphertext_s0[6]}), .I4 ({plaintext_s1[14], plaintext_s0[14]}), .O ({new_AGEMA_signal_2138, \stateArray/S32reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S32reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[23], ciphertext_s0[23]}), .I3 ({ciphertext_s1[7], ciphertext_s0[7]}), .I4 ({plaintext_s1[15], plaintext_s0[15]}), .O ({new_AGEMA_signal_2140, \stateArray/S32reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S01reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1525, \KeyArray/S11reg/gen_ff[1].gff/GEN[0].SFF/Q_659 }), .I3 ({new_AGEMA_signal_1526, \KeyArray/S02reg/gen_ff[1].gff/GEN[0].SFF/Q_683 }), .I4 ({key_s1[112], key_s0[112]}), .O ({new_AGEMA_signal_1528, \KeyArray/S01reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S01reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1529, \KeyArray/S11reg/gen_ff[1].gff/GEN[1].SFF/Q_660 }), .I3 ({new_AGEMA_signal_1530, \KeyArray/S02reg/gen_ff[1].gff/GEN[1].SFF/Q_684 }), .I4 ({key_s1[113], key_s0[113]}), .O ({new_AGEMA_signal_1532, \KeyArray/S01reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S01reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1533, \KeyArray/S11reg/gen_ff[1].gff/GEN[2].SFF/Q_661 }), .I3 ({new_AGEMA_signal_1534, \KeyArray/S02reg/gen_ff[1].gff/GEN[2].SFF/Q_685 }), .I4 ({key_s1[114], key_s0[114]}), .O ({new_AGEMA_signal_1536, \KeyArray/S01reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S01reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1537, \KeyArray/S11reg/gen_ff[1].gff/GEN[3].SFF/Q_662 }), .I3 ({new_AGEMA_signal_1538, \KeyArray/S02reg/gen_ff[1].gff/GEN[3].SFF/Q_686 }), .I4 ({key_s1[115], key_s0[115]}), .O ({new_AGEMA_signal_1540, \KeyArray/S01reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S01reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1541, \KeyArray/S11reg/gen_ff[1].gff/GEN[4].SFF/Q_663 }), .I3 ({new_AGEMA_signal_1542, \KeyArray/S02reg/gen_ff[1].gff/GEN[4].SFF/Q_687 }), .I4 ({key_s1[116], key_s0[116]}), .O ({new_AGEMA_signal_1544, \KeyArray/S01reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S01reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1545, \KeyArray/S11reg/gen_ff[1].gff/GEN[5].SFF/Q_664 }), .I3 ({new_AGEMA_signal_1546, \KeyArray/S02reg/gen_ff[1].gff/GEN[5].SFF/Q_688 }), .I4 ({key_s1[117], key_s0[117]}), .O ({new_AGEMA_signal_1548, \KeyArray/S01reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S01reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1549, \KeyArray/S11reg/gen_ff[1].gff/GEN[6].SFF/Q_665 }), .I3 ({new_AGEMA_signal_1550, \KeyArray/S02reg/gen_ff[1].gff/GEN[6].SFF/Q_689 }), .I4 ({key_s1[118], key_s0[118]}), .O ({new_AGEMA_signal_1552, \KeyArray/S01reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S01reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1553, \KeyArray/S11reg/gen_ff[1].gff/GEN[7].SFF/Q_666 }), .I3 ({new_AGEMA_signal_1554, \KeyArray/S02reg/gen_ff[1].gff/GEN[7].SFF/Q_690 }), .I4 ({key_s1[119], key_s0[119]}), .O ({new_AGEMA_signal_1556, \KeyArray/S01reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S02reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1557, \KeyArray/S12reg/gen_ff[1].gff/GEN[0].SFF/Q_651 }), .I3 ({new_AGEMA_signal_1558, \KeyArray/S03reg/gen_ff[1].gff/GEN[0].SFF/Q_675 }), .I4 ({key_s1[104], key_s0[104]}), .O ({new_AGEMA_signal_1560, \KeyArray/S02reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S02reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1561, \KeyArray/S12reg/gen_ff[1].gff/GEN[1].SFF/Q_652 }), .I3 ({new_AGEMA_signal_1562, \KeyArray/S03reg/gen_ff[1].gff/GEN[1].SFF/Q_676 }), .I4 ({key_s1[105], key_s0[105]}), .O ({new_AGEMA_signal_1564, \KeyArray/S02reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S02reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1565, \KeyArray/S12reg/gen_ff[1].gff/GEN[2].SFF/Q_653 }), .I3 ({new_AGEMA_signal_1566, \KeyArray/S03reg/gen_ff[1].gff/GEN[2].SFF/Q_677 }), .I4 ({key_s1[106], key_s0[106]}), .O ({new_AGEMA_signal_1568, \KeyArray/S02reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S02reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1569, \KeyArray/S12reg/gen_ff[1].gff/GEN[3].SFF/Q_654 }), .I3 ({new_AGEMA_signal_1570, \KeyArray/S03reg/gen_ff[1].gff/GEN[3].SFF/Q_678 }), .I4 ({key_s1[107], key_s0[107]}), .O ({new_AGEMA_signal_1572, \KeyArray/S02reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S02reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1573, \KeyArray/S12reg/gen_ff[1].gff/GEN[4].SFF/Q_655 }), .I3 ({new_AGEMA_signal_1574, \KeyArray/S03reg/gen_ff[1].gff/GEN[4].SFF/Q_679 }), .I4 ({key_s1[108], key_s0[108]}), .O ({new_AGEMA_signal_1576, \KeyArray/S02reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S02reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1577, \KeyArray/S12reg/gen_ff[1].gff/GEN[5].SFF/Q_656 }), .I3 ({new_AGEMA_signal_1578, \KeyArray/S03reg/gen_ff[1].gff/GEN[5].SFF/Q_680 }), .I4 ({key_s1[109], key_s0[109]}), .O ({new_AGEMA_signal_1580, \KeyArray/S02reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S02reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1581, \KeyArray/S12reg/gen_ff[1].gff/GEN[6].SFF/Q_657 }), .I3 ({new_AGEMA_signal_1582, \KeyArray/S03reg/gen_ff[1].gff/GEN[6].SFF/Q_681 }), .I4 ({key_s1[110], key_s0[110]}), .O ({new_AGEMA_signal_1584, \KeyArray/S02reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S02reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1585, \KeyArray/S12reg/gen_ff[1].gff/GEN[7].SFF/Q_658 }), .I3 ({new_AGEMA_signal_1586, \KeyArray/S03reg/gen_ff[1].gff/GEN[7].SFF/Q_682 }), .I4 ({key_s1[111], key_s0[111]}), .O ({new_AGEMA_signal_1588, \KeyArray/S02reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S03reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1433, \KeyArray/S13reg/gen_ff[1].gff/GEN[0].SFF/Q_393 }), .I3 ({new_AGEMA_signal_1589, \KeyArray/S10reg/gen_ff[1].gff/GEN[0].SFF/Q_667 }), .I4 ({key_s1[96], key_s0[96]}), .O ({new_AGEMA_signal_1591, \KeyArray/S03reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S03reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1431, \KeyArray/S13reg/gen_ff[1].gff/GEN[1].SFF/Q_392 }), .I3 ({new_AGEMA_signal_1592, \KeyArray/S10reg/gen_ff[1].gff/GEN[1].SFF/Q_668 }), .I4 ({key_s1[97], key_s0[97]}), .O ({new_AGEMA_signal_1594, \KeyArray/S03reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S03reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1429, \KeyArray/S13reg/gen_ff[1].gff/GEN[2].SFF/Q_391 }), .I3 ({new_AGEMA_signal_1595, \KeyArray/S10reg/gen_ff[1].gff/GEN[2].SFF/Q_669 }), .I4 ({key_s1[98], key_s0[98]}), .O ({new_AGEMA_signal_1597, \KeyArray/S03reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S03reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1427, \KeyArray/S13reg/gen_ff[1].gff/GEN[3].SFF/Q_390 }), .I3 ({new_AGEMA_signal_1598, \KeyArray/S10reg/gen_ff[1].gff/GEN[3].SFF/Q_670 }), .I4 ({key_s1[99], key_s0[99]}), .O ({new_AGEMA_signal_1600, \KeyArray/S03reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S03reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1425, \KeyArray/S13reg/gen_ff[1].gff/GEN[4].SFF/Q_389 }), .I3 ({new_AGEMA_signal_1601, \KeyArray/S10reg/gen_ff[1].gff/GEN[4].SFF/Q_671 }), .I4 ({key_s1[100], key_s0[100]}), .O ({new_AGEMA_signal_1603, \KeyArray/S03reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S03reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1423, \KeyArray/S13reg/gen_ff[1].gff/GEN[5].SFF/Q_388 }), .I3 ({new_AGEMA_signal_1604, \KeyArray/S10reg/gen_ff[1].gff/GEN[5].SFF/Q_672 }), .I4 ({key_s1[101], key_s0[101]}), .O ({new_AGEMA_signal_1606, \KeyArray/S03reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S03reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1437, \KeyArray/S13reg/gen_ff[1].gff/GEN[6].SFF/Q_387 }), .I3 ({new_AGEMA_signal_1607, \KeyArray/S10reg/gen_ff[1].gff/GEN[6].SFF/Q_673 }), .I4 ({key_s1[102], key_s0[102]}), .O ({new_AGEMA_signal_1609, \KeyArray/S03reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S03reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1435, \KeyArray/S13reg/gen_ff[1].gff/GEN[7].SFF/Q_386 }), .I3 ({new_AGEMA_signal_1610, \KeyArray/S10reg/gen_ff[1].gff/GEN[7].SFF/Q_674 }), .I4 ({key_s1[103], key_s0[103]}), .O ({new_AGEMA_signal_1612, \KeyArray/S03reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S10reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1613, \KeyArray/S20reg/gen_ff[1].gff/GEN[0].SFF/Q_643 }), .I3 ({new_AGEMA_signal_1525, \KeyArray/S11reg/gen_ff[1].gff/GEN[0].SFF/Q_659 }), .I4 ({key_s1[88], key_s0[88]}), .O ({new_AGEMA_signal_1615, \KeyArray/S10reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S10reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1616, \KeyArray/S20reg/gen_ff[1].gff/GEN[1].SFF/Q_644 }), .I3 ({new_AGEMA_signal_1529, \KeyArray/S11reg/gen_ff[1].gff/GEN[1].SFF/Q_660 }), .I4 ({key_s1[89], key_s0[89]}), .O ({new_AGEMA_signal_1618, \KeyArray/S10reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S10reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1619, \KeyArray/S20reg/gen_ff[1].gff/GEN[2].SFF/Q_645 }), .I3 ({new_AGEMA_signal_1533, \KeyArray/S11reg/gen_ff[1].gff/GEN[2].SFF/Q_661 }), .I4 ({key_s1[90], key_s0[90]}), .O ({new_AGEMA_signal_1621, \KeyArray/S10reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S10reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1622, \KeyArray/S20reg/gen_ff[1].gff/GEN[3].SFF/Q_646 }), .I3 ({new_AGEMA_signal_1537, \KeyArray/S11reg/gen_ff[1].gff/GEN[3].SFF/Q_662 }), .I4 ({key_s1[91], key_s0[91]}), .O ({new_AGEMA_signal_1624, \KeyArray/S10reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S10reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1625, \KeyArray/S20reg/gen_ff[1].gff/GEN[4].SFF/Q_647 }), .I3 ({new_AGEMA_signal_1541, \KeyArray/S11reg/gen_ff[1].gff/GEN[4].SFF/Q_663 }), .I4 ({key_s1[92], key_s0[92]}), .O ({new_AGEMA_signal_1627, \KeyArray/S10reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S10reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1628, \KeyArray/S20reg/gen_ff[1].gff/GEN[5].SFF/Q_648 }), .I3 ({new_AGEMA_signal_1545, \KeyArray/S11reg/gen_ff[1].gff/GEN[5].SFF/Q_664 }), .I4 ({key_s1[93], key_s0[93]}), .O ({new_AGEMA_signal_1630, \KeyArray/S10reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S10reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1631, \KeyArray/S20reg/gen_ff[1].gff/GEN[6].SFF/Q_649 }), .I3 ({new_AGEMA_signal_1549, \KeyArray/S11reg/gen_ff[1].gff/GEN[6].SFF/Q_665 }), .I4 ({key_s1[94], key_s0[94]}), .O ({new_AGEMA_signal_1633, \KeyArray/S10reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S10reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1634, \KeyArray/S20reg/gen_ff[1].gff/GEN[7].SFF/Q_650 }), .I3 ({new_AGEMA_signal_1553, \KeyArray/S11reg/gen_ff[1].gff/GEN[7].SFF/Q_666 }), .I4 ({key_s1[95], key_s0[95]}), .O ({new_AGEMA_signal_1636, \KeyArray/S10reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S11reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1637, \KeyArray/S21reg/gen_ff[1].gff/GEN[0].SFF/Q_635 }), .I3 ({new_AGEMA_signal_1557, \KeyArray/S12reg/gen_ff[1].gff/GEN[0].SFF/Q_651 }), .I4 ({key_s1[80], key_s0[80]}), .O ({new_AGEMA_signal_1639, \KeyArray/S11reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S11reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1640, \KeyArray/S21reg/gen_ff[1].gff/GEN[1].SFF/Q_636 }), .I3 ({new_AGEMA_signal_1561, \KeyArray/S12reg/gen_ff[1].gff/GEN[1].SFF/Q_652 }), .I4 ({key_s1[81], key_s0[81]}), .O ({new_AGEMA_signal_1642, \KeyArray/S11reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S11reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1643, \KeyArray/S21reg/gen_ff[1].gff/GEN[2].SFF/Q_637 }), .I3 ({new_AGEMA_signal_1565, \KeyArray/S12reg/gen_ff[1].gff/GEN[2].SFF/Q_653 }), .I4 ({key_s1[82], key_s0[82]}), .O ({new_AGEMA_signal_1645, \KeyArray/S11reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S11reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1646, \KeyArray/S21reg/gen_ff[1].gff/GEN[3].SFF/Q_638 }), .I3 ({new_AGEMA_signal_1569, \KeyArray/S12reg/gen_ff[1].gff/GEN[3].SFF/Q_654 }), .I4 ({key_s1[83], key_s0[83]}), .O ({new_AGEMA_signal_1648, \KeyArray/S11reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S11reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1649, \KeyArray/S21reg/gen_ff[1].gff/GEN[4].SFF/Q_639 }), .I3 ({new_AGEMA_signal_1573, \KeyArray/S12reg/gen_ff[1].gff/GEN[4].SFF/Q_655 }), .I4 ({key_s1[84], key_s0[84]}), .O ({new_AGEMA_signal_1651, \KeyArray/S11reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S11reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1652, \KeyArray/S21reg/gen_ff[1].gff/GEN[5].SFF/Q_640 }), .I3 ({new_AGEMA_signal_1577, \KeyArray/S12reg/gen_ff[1].gff/GEN[5].SFF/Q_656 }), .I4 ({key_s1[85], key_s0[85]}), .O ({new_AGEMA_signal_1654, \KeyArray/S11reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S11reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1655, \KeyArray/S21reg/gen_ff[1].gff/GEN[6].SFF/Q_641 }), .I3 ({new_AGEMA_signal_1581, \KeyArray/S12reg/gen_ff[1].gff/GEN[6].SFF/Q_657 }), .I4 ({key_s1[86], key_s0[86]}), .O ({new_AGEMA_signal_1657, \KeyArray/S11reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S11reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1658, \KeyArray/S21reg/gen_ff[1].gff/GEN[7].SFF/Q_642 }), .I3 ({new_AGEMA_signal_1585, \KeyArray/S12reg/gen_ff[1].gff/GEN[7].SFF/Q_658 }), .I4 ({key_s1[87], key_s0[87]}), .O ({new_AGEMA_signal_1660, \KeyArray/S11reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S12reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1661, \KeyArray/S22reg/gen_ff[1].gff/GEN[0].SFF/Q_627 }), .I3 ({new_AGEMA_signal_1433, \KeyArray/S13reg/gen_ff[1].gff/GEN[0].SFF/Q_393 }), .I4 ({key_s1[72], key_s0[72]}), .O ({new_AGEMA_signal_1663, \KeyArray/S12reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S12reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1664, \KeyArray/S22reg/gen_ff[1].gff/GEN[1].SFF/Q_628 }), .I3 ({new_AGEMA_signal_1431, \KeyArray/S13reg/gen_ff[1].gff/GEN[1].SFF/Q_392 }), .I4 ({key_s1[73], key_s0[73]}), .O ({new_AGEMA_signal_1666, \KeyArray/S12reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S12reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1667, \KeyArray/S22reg/gen_ff[1].gff/GEN[2].SFF/Q_629 }), .I3 ({new_AGEMA_signal_1429, \KeyArray/S13reg/gen_ff[1].gff/GEN[2].SFF/Q_391 }), .I4 ({key_s1[74], key_s0[74]}), .O ({new_AGEMA_signal_1669, \KeyArray/S12reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S12reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1670, \KeyArray/S22reg/gen_ff[1].gff/GEN[3].SFF/Q_630 }), .I3 ({new_AGEMA_signal_1427, \KeyArray/S13reg/gen_ff[1].gff/GEN[3].SFF/Q_390 }), .I4 ({key_s1[75], key_s0[75]}), .O ({new_AGEMA_signal_1672, \KeyArray/S12reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S12reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1673, \KeyArray/S22reg/gen_ff[1].gff/GEN[4].SFF/Q_631 }), .I3 ({new_AGEMA_signal_1425, \KeyArray/S13reg/gen_ff[1].gff/GEN[4].SFF/Q_389 }), .I4 ({key_s1[76], key_s0[76]}), .O ({new_AGEMA_signal_1675, \KeyArray/S12reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S12reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1676, \KeyArray/S22reg/gen_ff[1].gff/GEN[5].SFF/Q_632 }), .I3 ({new_AGEMA_signal_1423, \KeyArray/S13reg/gen_ff[1].gff/GEN[5].SFF/Q_388 }), .I4 ({key_s1[77], key_s0[77]}), .O ({new_AGEMA_signal_1678, \KeyArray/S12reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S12reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1679, \KeyArray/S22reg/gen_ff[1].gff/GEN[6].SFF/Q_633 }), .I3 ({new_AGEMA_signal_1437, \KeyArray/S13reg/gen_ff[1].gff/GEN[6].SFF/Q_387 }), .I4 ({key_s1[78], key_s0[78]}), .O ({new_AGEMA_signal_1681, \KeyArray/S12reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S12reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1682, \KeyArray/S22reg/gen_ff[1].gff/GEN[7].SFF/Q_634 }), .I3 ({new_AGEMA_signal_1435, \KeyArray/S13reg/gen_ff[1].gff/GEN[7].SFF/Q_386 }), .I4 ({key_s1[79], key_s0[79]}), .O ({new_AGEMA_signal_1684, \KeyArray/S12reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S13reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1685, \KeyArray/S23reg/gen_ff[1].gff/GEN[0].SFF/Q_619 }), .I3 ({new_AGEMA_signal_1613, \KeyArray/S20reg/gen_ff[1].gff/GEN[0].SFF/Q_643 }), .I4 ({key_s1[64], key_s0[64]}), .O ({new_AGEMA_signal_1687, \KeyArray/S13reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S13reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1688, \KeyArray/S23reg/gen_ff[1].gff/GEN[1].SFF/Q_620 }), .I3 ({new_AGEMA_signal_1616, \KeyArray/S20reg/gen_ff[1].gff/GEN[1].SFF/Q_644 }), .I4 ({key_s1[65], key_s0[65]}), .O ({new_AGEMA_signal_1690, \KeyArray/S13reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S13reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1691, \KeyArray/S23reg/gen_ff[1].gff/GEN[2].SFF/Q_621 }), .I3 ({new_AGEMA_signal_1619, \KeyArray/S20reg/gen_ff[1].gff/GEN[2].SFF/Q_645 }), .I4 ({key_s1[66], key_s0[66]}), .O ({new_AGEMA_signal_1693, \KeyArray/S13reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S13reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1694, \KeyArray/S23reg/gen_ff[1].gff/GEN[3].SFF/Q_622 }), .I3 ({new_AGEMA_signal_1622, \KeyArray/S20reg/gen_ff[1].gff/GEN[3].SFF/Q_646 }), .I4 ({key_s1[67], key_s0[67]}), .O ({new_AGEMA_signal_1696, \KeyArray/S13reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S13reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1697, \KeyArray/S23reg/gen_ff[1].gff/GEN[4].SFF/Q_623 }), .I3 ({new_AGEMA_signal_1625, \KeyArray/S20reg/gen_ff[1].gff/GEN[4].SFF/Q_647 }), .I4 ({key_s1[68], key_s0[68]}), .O ({new_AGEMA_signal_1699, \KeyArray/S13reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S13reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1700, \KeyArray/S23reg/gen_ff[1].gff/GEN[5].SFF/Q_624 }), .I3 ({new_AGEMA_signal_1628, \KeyArray/S20reg/gen_ff[1].gff/GEN[5].SFF/Q_648 }), .I4 ({key_s1[69], key_s0[69]}), .O ({new_AGEMA_signal_1702, \KeyArray/S13reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S13reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1703, \KeyArray/S23reg/gen_ff[1].gff/GEN[6].SFF/Q_625 }), .I3 ({new_AGEMA_signal_1631, \KeyArray/S20reg/gen_ff[1].gff/GEN[6].SFF/Q_649 }), .I4 ({key_s1[70], key_s0[70]}), .O ({new_AGEMA_signal_1705, \KeyArray/S13reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S13reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1706, \KeyArray/S23reg/gen_ff[1].gff/GEN[7].SFF/Q_626 }), .I3 ({new_AGEMA_signal_1634, \KeyArray/S20reg/gen_ff[1].gff/GEN[7].SFF/Q_650 }), .I4 ({key_s1[71], key_s0[71]}), .O ({new_AGEMA_signal_1708, \KeyArray/S13reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S20reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1709, \KeyArray/S30reg/gen_ff[1].gff/GEN[0].SFF/Q_611 }), .I3 ({new_AGEMA_signal_1637, \KeyArray/S21reg/gen_ff[1].gff/GEN[0].SFF/Q_635 }), .I4 ({key_s1[56], key_s0[56]}), .O ({new_AGEMA_signal_1711, \KeyArray/S20reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S20reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1712, \KeyArray/S30reg/gen_ff[1].gff/GEN[1].SFF/Q_612 }), .I3 ({new_AGEMA_signal_1640, \KeyArray/S21reg/gen_ff[1].gff/GEN[1].SFF/Q_636 }), .I4 ({key_s1[57], key_s0[57]}), .O ({new_AGEMA_signal_1714, \KeyArray/S20reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S20reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1715, \KeyArray/S30reg/gen_ff[1].gff/GEN[2].SFF/Q_613 }), .I3 ({new_AGEMA_signal_1643, \KeyArray/S21reg/gen_ff[1].gff/GEN[2].SFF/Q_637 }), .I4 ({key_s1[58], key_s0[58]}), .O ({new_AGEMA_signal_1717, \KeyArray/S20reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S20reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1718, \KeyArray/S30reg/gen_ff[1].gff/GEN[3].SFF/Q_614 }), .I3 ({new_AGEMA_signal_1646, \KeyArray/S21reg/gen_ff[1].gff/GEN[3].SFF/Q_638 }), .I4 ({key_s1[59], key_s0[59]}), .O ({new_AGEMA_signal_1720, \KeyArray/S20reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S20reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1721, \KeyArray/S30reg/gen_ff[1].gff/GEN[4].SFF/Q_615 }), .I3 ({new_AGEMA_signal_1649, \KeyArray/S21reg/gen_ff[1].gff/GEN[4].SFF/Q_639 }), .I4 ({key_s1[60], key_s0[60]}), .O ({new_AGEMA_signal_1723, \KeyArray/S20reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S20reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1724, \KeyArray/S30reg/gen_ff[1].gff/GEN[5].SFF/Q_616 }), .I3 ({new_AGEMA_signal_1652, \KeyArray/S21reg/gen_ff[1].gff/GEN[5].SFF/Q_640 }), .I4 ({key_s1[61], key_s0[61]}), .O ({new_AGEMA_signal_1726, \KeyArray/S20reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S20reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1727, \KeyArray/S30reg/gen_ff[1].gff/GEN[6].SFF/Q_617 }), .I3 ({new_AGEMA_signal_1655, \KeyArray/S21reg/gen_ff[1].gff/GEN[6].SFF/Q_641 }), .I4 ({key_s1[62], key_s0[62]}), .O ({new_AGEMA_signal_1729, \KeyArray/S20reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S20reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1730, \KeyArray/S30reg/gen_ff[1].gff/GEN[7].SFF/Q_618 }), .I3 ({new_AGEMA_signal_1658, \KeyArray/S21reg/gen_ff[1].gff/GEN[7].SFF/Q_642 }), .I4 ({key_s1[63], key_s0[63]}), .O ({new_AGEMA_signal_1732, \KeyArray/S20reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S21reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1733, \KeyArray/S31reg/gen_ff[1].gff/GEN[0].SFF/Q_603 }), .I3 ({new_AGEMA_signal_1661, \KeyArray/S22reg/gen_ff[1].gff/GEN[0].SFF/Q_627 }), .I4 ({key_s1[48], key_s0[48]}), .O ({new_AGEMA_signal_1735, \KeyArray/S21reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S21reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1736, \KeyArray/S31reg/gen_ff[1].gff/GEN[1].SFF/Q_604 }), .I3 ({new_AGEMA_signal_1664, \KeyArray/S22reg/gen_ff[1].gff/GEN[1].SFF/Q_628 }), .I4 ({key_s1[49], key_s0[49]}), .O ({new_AGEMA_signal_1738, \KeyArray/S21reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S21reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1739, \KeyArray/S31reg/gen_ff[1].gff/GEN[2].SFF/Q_605 }), .I3 ({new_AGEMA_signal_1667, \KeyArray/S22reg/gen_ff[1].gff/GEN[2].SFF/Q_629 }), .I4 ({key_s1[50], key_s0[50]}), .O ({new_AGEMA_signal_1741, \KeyArray/S21reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S21reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1742, \KeyArray/S31reg/gen_ff[1].gff/GEN[3].SFF/Q_606 }), .I3 ({new_AGEMA_signal_1670, \KeyArray/S22reg/gen_ff[1].gff/GEN[3].SFF/Q_630 }), .I4 ({key_s1[51], key_s0[51]}), .O ({new_AGEMA_signal_1744, \KeyArray/S21reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S21reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1745, \KeyArray/S31reg/gen_ff[1].gff/GEN[4].SFF/Q_607 }), .I3 ({new_AGEMA_signal_1673, \KeyArray/S22reg/gen_ff[1].gff/GEN[4].SFF/Q_631 }), .I4 ({key_s1[52], key_s0[52]}), .O ({new_AGEMA_signal_1747, \KeyArray/S21reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S21reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1748, \KeyArray/S31reg/gen_ff[1].gff/GEN[5].SFF/Q_608 }), .I3 ({new_AGEMA_signal_1676, \KeyArray/S22reg/gen_ff[1].gff/GEN[5].SFF/Q_632 }), .I4 ({key_s1[53], key_s0[53]}), .O ({new_AGEMA_signal_1750, \KeyArray/S21reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S21reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1751, \KeyArray/S31reg/gen_ff[1].gff/GEN[6].SFF/Q_609 }), .I3 ({new_AGEMA_signal_1679, \KeyArray/S22reg/gen_ff[1].gff/GEN[6].SFF/Q_633 }), .I4 ({key_s1[54], key_s0[54]}), .O ({new_AGEMA_signal_1753, \KeyArray/S21reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S21reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1754, \KeyArray/S31reg/gen_ff[1].gff/GEN[7].SFF/Q_610 }), .I3 ({new_AGEMA_signal_1682, \KeyArray/S22reg/gen_ff[1].gff/GEN[7].SFF/Q_634 }), .I4 ({key_s1[55], key_s0[55]}), .O ({new_AGEMA_signal_1756, \KeyArray/S21reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S22reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1757, \KeyArray/S32reg/gen_ff[1].gff/GEN[0].SFF/Q_595 }), .I3 ({new_AGEMA_signal_1685, \KeyArray/S23reg/gen_ff[1].gff/GEN[0].SFF/Q_619 }), .I4 ({key_s1[40], key_s0[40]}), .O ({new_AGEMA_signal_1759, \KeyArray/S22reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S22reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1760, \KeyArray/S32reg/gen_ff[1].gff/GEN[1].SFF/Q_596 }), .I3 ({new_AGEMA_signal_1688, \KeyArray/S23reg/gen_ff[1].gff/GEN[1].SFF/Q_620 }), .I4 ({key_s1[41], key_s0[41]}), .O ({new_AGEMA_signal_1762, \KeyArray/S22reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S22reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1763, \KeyArray/S32reg/gen_ff[1].gff/GEN[2].SFF/Q_597 }), .I3 ({new_AGEMA_signal_1691, \KeyArray/S23reg/gen_ff[1].gff/GEN[2].SFF/Q_621 }), .I4 ({key_s1[42], key_s0[42]}), .O ({new_AGEMA_signal_1765, \KeyArray/S22reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S22reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1766, \KeyArray/S32reg/gen_ff[1].gff/GEN[3].SFF/Q_598 }), .I3 ({new_AGEMA_signal_1694, \KeyArray/S23reg/gen_ff[1].gff/GEN[3].SFF/Q_622 }), .I4 ({key_s1[43], key_s0[43]}), .O ({new_AGEMA_signal_1768, \KeyArray/S22reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S22reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1769, \KeyArray/S32reg/gen_ff[1].gff/GEN[4].SFF/Q_599 }), .I3 ({new_AGEMA_signal_1697, \KeyArray/S23reg/gen_ff[1].gff/GEN[4].SFF/Q_623 }), .I4 ({key_s1[44], key_s0[44]}), .O ({new_AGEMA_signal_1771, \KeyArray/S22reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S22reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1772, \KeyArray/S32reg/gen_ff[1].gff/GEN[5].SFF/Q_600 }), .I3 ({new_AGEMA_signal_1700, \KeyArray/S23reg/gen_ff[1].gff/GEN[5].SFF/Q_624 }), .I4 ({key_s1[45], key_s0[45]}), .O ({new_AGEMA_signal_1774, \KeyArray/S22reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S22reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1775, \KeyArray/S32reg/gen_ff[1].gff/GEN[6].SFF/Q_601 }), .I3 ({new_AGEMA_signal_1703, \KeyArray/S23reg/gen_ff[1].gff/GEN[6].SFF/Q_625 }), .I4 ({key_s1[46], key_s0[46]}), .O ({new_AGEMA_signal_1777, \KeyArray/S22reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S22reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1778, \KeyArray/S32reg/gen_ff[1].gff/GEN[7].SFF/Q_602 }), .I3 ({new_AGEMA_signal_1706, \KeyArray/S23reg/gen_ff[1].gff/GEN[7].SFF/Q_626 }), .I4 ({key_s1[47], key_s0[47]}), .O ({new_AGEMA_signal_1780, \KeyArray/S22reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S23reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1781, \KeyArray/S33reg/gen_ff[1].gff/GEN[0].SFF/Q_587 }), .I3 ({new_AGEMA_signal_1709, \KeyArray/S30reg/gen_ff[1].gff/GEN[0].SFF/Q_611 }), .I4 ({key_s1[32], key_s0[32]}), .O ({new_AGEMA_signal_1783, \KeyArray/S23reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S23reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1784, \KeyArray/S33reg/gen_ff[1].gff/GEN[1].SFF/Q_588 }), .I3 ({new_AGEMA_signal_1712, \KeyArray/S30reg/gen_ff[1].gff/GEN[1].SFF/Q_612 }), .I4 ({key_s1[33], key_s0[33]}), .O ({new_AGEMA_signal_1786, \KeyArray/S23reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S23reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1787, \KeyArray/S33reg/gen_ff[1].gff/GEN[2].SFF/Q_589 }), .I3 ({new_AGEMA_signal_1715, \KeyArray/S30reg/gen_ff[1].gff/GEN[2].SFF/Q_613 }), .I4 ({key_s1[34], key_s0[34]}), .O ({new_AGEMA_signal_1789, \KeyArray/S23reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S23reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1790, \KeyArray/S33reg/gen_ff[1].gff/GEN[3].SFF/Q_590 }), .I3 ({new_AGEMA_signal_1718, \KeyArray/S30reg/gen_ff[1].gff/GEN[3].SFF/Q_614 }), .I4 ({key_s1[35], key_s0[35]}), .O ({new_AGEMA_signal_1792, \KeyArray/S23reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S23reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1793, \KeyArray/S33reg/gen_ff[1].gff/GEN[4].SFF/Q_591 }), .I3 ({new_AGEMA_signal_1721, \KeyArray/S30reg/gen_ff[1].gff/GEN[4].SFF/Q_615 }), .I4 ({key_s1[36], key_s0[36]}), .O ({new_AGEMA_signal_1795, \KeyArray/S23reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S23reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1796, \KeyArray/S33reg/gen_ff[1].gff/GEN[5].SFF/Q_592 }), .I3 ({new_AGEMA_signal_1724, \KeyArray/S30reg/gen_ff[1].gff/GEN[5].SFF/Q_616 }), .I4 ({key_s1[37], key_s0[37]}), .O ({new_AGEMA_signal_1798, \KeyArray/S23reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S23reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1799, \KeyArray/S33reg/gen_ff[1].gff/GEN[6].SFF/Q_593 }), .I3 ({new_AGEMA_signal_1727, \KeyArray/S30reg/gen_ff[1].gff/GEN[6].SFF/Q_617 }), .I4 ({key_s1[38], key_s0[38]}), .O ({new_AGEMA_signal_1801, \KeyArray/S23reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S23reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1802, \KeyArray/S33reg/gen_ff[1].gff/GEN[7].SFF/Q_594 }), .I3 ({new_AGEMA_signal_1730, \KeyArray/S30reg/gen_ff[1].gff/GEN[7].SFF/Q_618 }), .I4 ({key_s1[39], key_s0[39]}), .O ({new_AGEMA_signal_1804, \KeyArray/S23reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S31reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1805, \KeyArray/S01reg/gen_ff[1].gff/GEN[0].SFF/Q_691 }), .I3 ({new_AGEMA_signal_1757, \KeyArray/S32reg/gen_ff[1].gff/GEN[0].SFF/Q_595 }), .I4 ({key_s1[16], key_s0[16]}), .O ({new_AGEMA_signal_1807, \KeyArray/S31reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S31reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1808, \KeyArray/S01reg/gen_ff[1].gff/GEN[1].SFF/Q_692 }), .I3 ({new_AGEMA_signal_1760, \KeyArray/S32reg/gen_ff[1].gff/GEN[1].SFF/Q_596 }), .I4 ({key_s1[17], key_s0[17]}), .O ({new_AGEMA_signal_1810, \KeyArray/S31reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S31reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1811, \KeyArray/S01reg/gen_ff[1].gff/GEN[2].SFF/Q_693 }), .I3 ({new_AGEMA_signal_1763, \KeyArray/S32reg/gen_ff[1].gff/GEN[2].SFF/Q_597 }), .I4 ({key_s1[18], key_s0[18]}), .O ({new_AGEMA_signal_1813, \KeyArray/S31reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S31reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1814, \KeyArray/S01reg/gen_ff[1].gff/GEN[3].SFF/Q_694 }), .I3 ({new_AGEMA_signal_1766, \KeyArray/S32reg/gen_ff[1].gff/GEN[3].SFF/Q_598 }), .I4 ({key_s1[19], key_s0[19]}), .O ({new_AGEMA_signal_1816, \KeyArray/S31reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S31reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1817, \KeyArray/S01reg/gen_ff[1].gff/GEN[4].SFF/Q_695 }), .I3 ({new_AGEMA_signal_1769, \KeyArray/S32reg/gen_ff[1].gff/GEN[4].SFF/Q_599 }), .I4 ({key_s1[20], key_s0[20]}), .O ({new_AGEMA_signal_1819, \KeyArray/S31reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S31reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1820, \KeyArray/S01reg/gen_ff[1].gff/GEN[5].SFF/Q_696 }), .I3 ({new_AGEMA_signal_1772, \KeyArray/S32reg/gen_ff[1].gff/GEN[5].SFF/Q_600 }), .I4 ({key_s1[21], key_s0[21]}), .O ({new_AGEMA_signal_1822, \KeyArray/S31reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S31reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1823, \KeyArray/S01reg/gen_ff[1].gff/GEN[6].SFF/Q_697 }), .I3 ({new_AGEMA_signal_1775, \KeyArray/S32reg/gen_ff[1].gff/GEN[6].SFF/Q_601 }), .I4 ({key_s1[22], key_s0[22]}), .O ({new_AGEMA_signal_1825, \KeyArray/S31reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S31reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1826, \KeyArray/S01reg/gen_ff[1].gff/GEN[7].SFF/Q_698 }), .I3 ({new_AGEMA_signal_1778, \KeyArray/S32reg/gen_ff[1].gff/GEN[7].SFF/Q_602 }), .I4 ({key_s1[23], key_s0[23]}), .O ({new_AGEMA_signal_1828, \KeyArray/S31reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S32reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1526, \KeyArray/S02reg/gen_ff[1].gff/GEN[0].SFF/Q_683 }), .I3 ({new_AGEMA_signal_1781, \KeyArray/S33reg/gen_ff[1].gff/GEN[0].SFF/Q_587 }), .I4 ({key_s1[8], key_s0[8]}), .O ({new_AGEMA_signal_1830, \KeyArray/S32reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S32reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1530, \KeyArray/S02reg/gen_ff[1].gff/GEN[1].SFF/Q_684 }), .I3 ({new_AGEMA_signal_1784, \KeyArray/S33reg/gen_ff[1].gff/GEN[1].SFF/Q_588 }), .I4 ({key_s1[9], key_s0[9]}), .O ({new_AGEMA_signal_1832, \KeyArray/S32reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S32reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1534, \KeyArray/S02reg/gen_ff[1].gff/GEN[2].SFF/Q_685 }), .I3 ({new_AGEMA_signal_1787, \KeyArray/S33reg/gen_ff[1].gff/GEN[2].SFF/Q_589 }), .I4 ({key_s1[10], key_s0[10]}), .O ({new_AGEMA_signal_1834, \KeyArray/S32reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S32reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1538, \KeyArray/S02reg/gen_ff[1].gff/GEN[3].SFF/Q_686 }), .I3 ({new_AGEMA_signal_1790, \KeyArray/S33reg/gen_ff[1].gff/GEN[3].SFF/Q_590 }), .I4 ({key_s1[11], key_s0[11]}), .O ({new_AGEMA_signal_1836, \KeyArray/S32reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S32reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1542, \KeyArray/S02reg/gen_ff[1].gff/GEN[4].SFF/Q_687 }), .I3 ({new_AGEMA_signal_1793, \KeyArray/S33reg/gen_ff[1].gff/GEN[4].SFF/Q_591 }), .I4 ({key_s1[12], key_s0[12]}), .O ({new_AGEMA_signal_1838, \KeyArray/S32reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S32reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1546, \KeyArray/S02reg/gen_ff[1].gff/GEN[5].SFF/Q_688 }), .I3 ({new_AGEMA_signal_1796, \KeyArray/S33reg/gen_ff[1].gff/GEN[5].SFF/Q_592 }), .I4 ({key_s1[13], key_s0[13]}), .O ({new_AGEMA_signal_1840, \KeyArray/S32reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S32reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1550, \KeyArray/S02reg/gen_ff[1].gff/GEN[6].SFF/Q_689 }), .I3 ({new_AGEMA_signal_1799, \KeyArray/S33reg/gen_ff[1].gff/GEN[6].SFF/Q_593 }), .I4 ({key_s1[14], key_s0[14]}), .O ({new_AGEMA_signal_1842, \KeyArray/S32reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S32reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1554, \KeyArray/S02reg/gen_ff[1].gff/GEN[7].SFF/Q_690 }), .I3 ({new_AGEMA_signal_1802, \KeyArray/S33reg/gen_ff[1].gff/GEN[7].SFF/Q_594 }), .I4 ({key_s1[15], key_s0[15]}), .O ({new_AGEMA_signal_1844, \KeyArray/S32reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S33reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1558, \KeyArray/S03reg/gen_ff[1].gff/GEN[0].SFF/Q_675 }), .I3 ({new_AGEMA_signal_1371, \KeyArray/S00reg/gen_ff[1].gff/GEN[0].SFF/Q_401 }), .I4 ({key_s1[0], key_s0[0]}), .O ({new_AGEMA_signal_1846, \KeyArray/S33reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S33reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1562, \KeyArray/S03reg/gen_ff[1].gff/GEN[1].SFF/Q_676 }), .I3 ({new_AGEMA_signal_1368, \KeyArray/S00reg/gen_ff[1].gff/GEN[1].SFF/Q_400 }), .I4 ({key_s1[1], key_s0[1]}), .O ({new_AGEMA_signal_1848, \KeyArray/S33reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S33reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1566, \KeyArray/S03reg/gen_ff[1].gff/GEN[2].SFF/Q_677 }), .I3 ({new_AGEMA_signal_1365, \KeyArray/S00reg/gen_ff[1].gff/GEN[2].SFF/Q_399 }), .I4 ({key_s1[2], key_s0[2]}), .O ({new_AGEMA_signal_1850, \KeyArray/S33reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S33reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1570, \KeyArray/S03reg/gen_ff[1].gff/GEN[3].SFF/Q_678 }), .I3 ({new_AGEMA_signal_1362, \KeyArray/S00reg/gen_ff[1].gff/GEN[3].SFF/Q_398 }), .I4 ({key_s1[3], key_s0[3]}), .O ({new_AGEMA_signal_1852, \KeyArray/S33reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S33reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1574, \KeyArray/S03reg/gen_ff[1].gff/GEN[4].SFF/Q_679 }), .I3 ({new_AGEMA_signal_1359, \KeyArray/S00reg/gen_ff[1].gff/GEN[4].SFF/Q_397 }), .I4 ({key_s1[4], key_s0[4]}), .O ({new_AGEMA_signal_1854, \KeyArray/S33reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S33reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1578, \KeyArray/S03reg/gen_ff[1].gff/GEN[5].SFF/Q_680 }), .I3 ({new_AGEMA_signal_1356, \KeyArray/S00reg/gen_ff[1].gff/GEN[5].SFF/Q_396 }), .I4 ({key_s1[5], key_s0[5]}), .O ({new_AGEMA_signal_1856, \KeyArray/S33reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S33reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1582, \KeyArray/S03reg/gen_ff[1].gff/GEN[6].SFF/Q_681 }), .I3 ({new_AGEMA_signal_1353, \KeyArray/S00reg/gen_ff[1].gff/GEN[6].SFF/Q_395 }), .I4 ({key_s1[6], key_s0[6]}), .O ({new_AGEMA_signal_1858, \KeyArray/S33reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S33reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1586, \KeyArray/S03reg/gen_ff[1].gff/GEN[7].SFF/Q_682 }), .I3 ({new_AGEMA_signal_1350, \KeyArray/S00reg/gen_ff[1].gff/GEN[7].SFF/Q_394 }), .I4 ({key_s1[7], key_s0[7]}), .O ({new_AGEMA_signal_1860, \KeyArray/S33reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q13 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[96], ciphertext_s0[96]}), .I3 ({new_AGEMA_signal_1901, \stateArray/S03reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11_897 }), .I4 ({plaintext_s1[96], plaintext_s0[96]}), .O ({new_AGEMA_signal_2166, \stateArray/S03reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q14 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[97], ciphertext_s0[97]}), .I3 ({new_AGEMA_signal_1916, \stateArray/S03reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q12 }), .I4 ({plaintext_s1[97], plaintext_s0[97]}), .O ({new_AGEMA_signal_2168, \stateArray/S03reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q13 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({new_AGEMA_signal_1902, \stateArray/S03reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11_900 }), .I4 ({plaintext_s1[98], plaintext_s0[98]}), .O ({new_AGEMA_signal_2170, \stateArray/S03reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q14 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[99], ciphertext_s0[99]}), .I3 ({new_AGEMA_signal_1917, \stateArray/S03reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q12 }), .I4 ({plaintext_s1[99], plaintext_s0[99]}), .O ({new_AGEMA_signal_2172, \stateArray/S03reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q14 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[100], ciphertext_s0[100]}), .I3 ({new_AGEMA_signal_1918, \stateArray/S03reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q12 }), .I4 ({plaintext_s1[100], plaintext_s0[100]}), .O ({new_AGEMA_signal_2174, \stateArray/S03reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q13 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[101], ciphertext_s0[101]}), .I3 ({new_AGEMA_signal_1903, \stateArray/S03reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11_904 }), .I4 ({plaintext_s1[101], plaintext_s0[101]}), .O ({new_AGEMA_signal_2176, \stateArray/S03reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q13 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[102], ciphertext_s0[102]}), .I3 ({new_AGEMA_signal_1904, \stateArray/S03reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11_906 }), .I4 ({plaintext_s1[102], plaintext_s0[102]}), .O ({new_AGEMA_signal_2178, \stateArray/S03reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q13 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[103], ciphertext_s0[103]}), .I3 ({new_AGEMA_signal_1905, \stateArray/S03reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11_908 }), .I4 ({plaintext_s1[103], plaintext_s0[103]}), .O ({new_AGEMA_signal_2180, \stateArray/S03reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q13 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[88], ciphertext_s0[88]}), .I3 ({new_AGEMA_signal_1906, \stateArray/S13reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11_910 }), .I4 ({plaintext_s1[64], plaintext_s0[64]}), .O ({new_AGEMA_signal_2182, \stateArray/S13reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q14 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[89], ciphertext_s0[89]}), .I3 ({new_AGEMA_signal_1919, \stateArray/S13reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q12 }), .I4 ({plaintext_s1[65], plaintext_s0[65]}), .O ({new_AGEMA_signal_2184, \stateArray/S13reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q13 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({new_AGEMA_signal_1907, \stateArray/S13reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11_913 }), .I4 ({plaintext_s1[66], plaintext_s0[66]}), .O ({new_AGEMA_signal_2186, \stateArray/S13reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q14 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[91], ciphertext_s0[91]}), .I3 ({new_AGEMA_signal_1920, \stateArray/S13reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q12 }), .I4 ({plaintext_s1[67], plaintext_s0[67]}), .O ({new_AGEMA_signal_2188, \stateArray/S13reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q14 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[92], ciphertext_s0[92]}), .I3 ({new_AGEMA_signal_1921, \stateArray/S13reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q12 }), .I4 ({plaintext_s1[68], plaintext_s0[68]}), .O ({new_AGEMA_signal_2190, \stateArray/S13reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q13 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[93], ciphertext_s0[93]}), .I3 ({new_AGEMA_signal_1908, \stateArray/S13reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11_917 }), .I4 ({plaintext_s1[69], plaintext_s0[69]}), .O ({new_AGEMA_signal_2192, \stateArray/S13reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q13 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[94], ciphertext_s0[94]}), .I3 ({new_AGEMA_signal_1909, \stateArray/S13reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11_919 }), .I4 ({plaintext_s1[70], plaintext_s0[70]}), .O ({new_AGEMA_signal_2194, \stateArray/S13reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q13 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[95], ciphertext_s0[95]}), .I3 ({new_AGEMA_signal_1910, \stateArray/S13reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11_921 }), .I4 ({plaintext_s1[71], plaintext_s0[71]}), .O ({new_AGEMA_signal_2196, \stateArray/S13reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q13 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[48], ciphertext_s0[48]}), .I3 ({new_AGEMA_signal_1911, \stateArray/S23reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11_923 }), .I4 ({plaintext_s1[32], plaintext_s0[32]}), .O ({new_AGEMA_signal_2198, \stateArray/S23reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q14 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[49], ciphertext_s0[49]}), .I3 ({new_AGEMA_signal_1922, \stateArray/S23reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q12 }), .I4 ({plaintext_s1[33], plaintext_s0[33]}), .O ({new_AGEMA_signal_2200, \stateArray/S23reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q13 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({new_AGEMA_signal_1912, \stateArray/S23reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11_926 }), .I4 ({plaintext_s1[34], plaintext_s0[34]}), .O ({new_AGEMA_signal_2202, \stateArray/S23reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q14 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[51], ciphertext_s0[51]}), .I3 ({new_AGEMA_signal_1923, \stateArray/S23reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q12 }), .I4 ({plaintext_s1[35], plaintext_s0[35]}), .O ({new_AGEMA_signal_2204, \stateArray/S23reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q14 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[52], ciphertext_s0[52]}), .I3 ({new_AGEMA_signal_1924, \stateArray/S23reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q12 }), .I4 ({plaintext_s1[36], plaintext_s0[36]}), .O ({new_AGEMA_signal_2206, \stateArray/S23reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q13 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[53], ciphertext_s0[53]}), .I3 ({new_AGEMA_signal_1913, \stateArray/S23reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11_930 }), .I4 ({plaintext_s1[37], plaintext_s0[37]}), .O ({new_AGEMA_signal_2208, \stateArray/S23reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q13 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[54], ciphertext_s0[54]}), .I3 ({new_AGEMA_signal_1914, \stateArray/S23reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11_932 }), .I4 ({plaintext_s1[38], plaintext_s0[38]}), .O ({new_AGEMA_signal_2210, \stateArray/S23reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q13 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[55], ciphertext_s0[55]}), .I3 ({new_AGEMA_signal_1915, \stateArray/S23reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11_934 }), .I4 ({plaintext_s1[39], plaintext_s0[39]}), .O ({new_AGEMA_signal_2212, \stateArray/S23reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT6 #( .INIT ( 64'h0000000000000002 ) ) \ctrl/selSR1 ( .I0 (nReset_407), .I1 (\ctrl/seq6/GEN[0].SFF/Q_841 ), .I2 (\ctrl/seq6/GEN[4].SFF/Q_842 ), .I3 (\ctrl/seq6/GEN[3].SFF/Q_840 ), .I4 (\ctrl/seq6/GEN[1].SFF/Q_838 ), .I5 (\ctrl/seq6/GEN[2].SFF/Q_839 ), .O (selSR) ) ;
    LUT5 #( .INIT ( 32'hFFFF8880 ) ) \ctrl/CSselMC_rstpot ( .I0 (nReset_407), .I1 (\ctrl/CSselMC_835 ), .I2 (\ctrl/seq4/GEN[0].SFF/Q_836 ), .I3 (\ctrl/seq4/GEN[1].SFF/Q_837 ), .I4 (\ctrl/finalStep1 ), .O (\ctrl/CSselMC_rstpot_1330 ) ) ;
    LUT6 #( .INIT ( 64'hFFFFFFFFFFFEFFFF ) ) enKS1 ( .I0 (\ctrl/seq6/GEN[2].SFF/Q_839 ), .I1 (\ctrl/seq6/GEN[4].SFF/Q_842 ), .I2 (\ctrl/seq6/GEN[3].SFF/Q_840 ), .I3 (\ctrl/seq6/GEN[1].SFF/Q_838 ), .I4 (nReset_407), .I5 (\ctrl/seq6/GEN[0].SFF/Q_841 ), .O (enKS) ) ;
    INV \ctrl/nReset_inv1_INV_0 ( .I (nReset_407), .O (\calcRCon/nReset_inv ) ) ;
    INV nReset_rstpot1_INV_0 ( .I (start), .O (nReset_rstpot) ) ;
    ClockGatingController #(3) ClockGatingInst ( .clk (clk), .rst (start), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'h52379DE7B844E3E1 ) ) \Inst_bSbox/b7_3 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r ({Fresh[63], Fresh[62], Fresh[61], Fresh[60], Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48], Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30], Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .O ({new_AGEMA_signal_1861, \Inst_bSbox/b7 [3]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'h4CB3770196CA0329 ) ) \Inst_bSbox/b7_2 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r ({Fresh[127], Fresh[126], Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120], Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114], Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108], Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96], Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90], Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84], Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72], Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65], Fresh[64]}), .O ({new_AGEMA_signal_1862, \Inst_bSbox/b7 [2]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'hE7BAC28F866AAC82 ) ) \Inst_bSbox/b7_1 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186], Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180], Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174], Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168], Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162], Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156], Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150], Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144], Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138], Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132], Fresh[131], Fresh[130], Fresh[129], Fresh[128]}), .O ({new_AGEMA_signal_1863, \Inst_bSbox/b7 [1]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'h5CAA2EC7BF977090 ) ) \Inst_bSbox/b7_0 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r ({Fresh[255], Fresh[254], Fresh[253], Fresh[252], Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246], Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240], Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234], Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228], Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222], Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216], Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210], Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204], Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198], Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192]}), .O ({new_AGEMA_signal_1864, \Inst_bSbox/b7 [0]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'h21E0B83325591782 ) ) \Inst_bSbox/b6_3 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r ({Fresh[319], Fresh[318], Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312], Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306], Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300], Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294], Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288], Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282], Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276], Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270], Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264], Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258], Fresh[257], Fresh[256]}), .O ({new_AGEMA_signal_1865, \Inst_bSbox/b6 [3]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'h3F6BCB91B30DB559 ) ) \Inst_bSbox/b6_2 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378], Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372], Fresh[371], Fresh[370], Fresh[369], Fresh[368], Fresh[367], Fresh[366], Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360], Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354], Fresh[353], Fresh[352], Fresh[351], Fresh[350], Fresh[349], Fresh[348], Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342], Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336], Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330], Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324], Fresh[323], Fresh[322], Fresh[321], Fresh[320]}), .O ({new_AGEMA_signal_1866, \Inst_bSbox/b6 [2]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'hE4851B3BF3AB2560 ) ) \Inst_bSbox/b6_1 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r ({Fresh[447], Fresh[446], Fresh[445], Fresh[444], Fresh[443], Fresh[442], Fresh[441], Fresh[440], Fresh[439], Fresh[438], Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432], Fresh[431], Fresh[430], Fresh[429], Fresh[428], Fresh[427], Fresh[426], Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420], Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414], Fresh[413], Fresh[412], Fresh[411], Fresh[410], Fresh[409], Fresh[408], Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402], Fresh[401], Fresh[400], Fresh[399], Fresh[398], Fresh[397], Fresh[396], Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390], Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384]}), .O ({new_AGEMA_signal_1867, \Inst_bSbox/b6 [1]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'h980A3CC2C2FDB4FF ) ) \Inst_bSbox/b6_0 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r ({Fresh[511], Fresh[510], Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504], Fresh[503], Fresh[502], Fresh[501], Fresh[500], Fresh[499], Fresh[498], Fresh[497], Fresh[496], Fresh[495], Fresh[494], Fresh[493], Fresh[492], Fresh[491], Fresh[490], Fresh[489], Fresh[488], Fresh[487], Fresh[486], Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480], Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474], Fresh[473], Fresh[472], Fresh[471], Fresh[470], Fresh[469], Fresh[468], Fresh[467], Fresh[466], Fresh[465], Fresh[464], Fresh[463], Fresh[462], Fresh[461], Fresh[460], Fresh[459], Fresh[458], Fresh[457], Fresh[456], Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450], Fresh[449], Fresh[448]}), .O ({new_AGEMA_signal_1868, \Inst_bSbox/b6 [0]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'h54B248130B4F256F ) ) \Inst_bSbox/b5_3 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r ({Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570], Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564], Fresh[563], Fresh[562], Fresh[561], Fresh[560], Fresh[559], Fresh[558], Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552], Fresh[551], Fresh[550], Fresh[549], Fresh[548], Fresh[547], Fresh[546], Fresh[545], Fresh[544], Fresh[543], Fresh[542], Fresh[541], Fresh[540], Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534], Fresh[533], Fresh[532], Fresh[531], Fresh[530], Fresh[529], Fresh[528], Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522], Fresh[521], Fresh[520], Fresh[519], Fresh[518], Fresh[517], Fresh[516], Fresh[515], Fresh[514], Fresh[513], Fresh[512]}), .O ({new_AGEMA_signal_1869, \Inst_bSbox/b5 [3]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'h7D8DCC4706319E08 ) ) \Inst_bSbox/b5_2 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r ({Fresh[639], Fresh[638], Fresh[637], Fresh[636], Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630], Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624], Fresh[623], Fresh[622], Fresh[621], Fresh[620], Fresh[619], Fresh[618], Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612], Fresh[611], Fresh[610], Fresh[609], Fresh[608], Fresh[607], Fresh[606], Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600], Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594], Fresh[593], Fresh[592], Fresh[591], Fresh[590], Fresh[589], Fresh[588], Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582], Fresh[581], Fresh[580], Fresh[579], Fresh[578], Fresh[577], Fresh[576]}), .O ({new_AGEMA_signal_1870, \Inst_bSbox/b5 [2]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6BC2AA4E0D787AA4 ) ) \Inst_bSbox/b5_1 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r ({Fresh[703], Fresh[702], Fresh[701], Fresh[700], Fresh[699], Fresh[698], Fresh[697], Fresh[696], Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690], Fresh[689], Fresh[688], Fresh[687], Fresh[686], Fresh[685], Fresh[684], Fresh[683], Fresh[682], Fresh[681], Fresh[680], Fresh[679], Fresh[678], Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672], Fresh[671], Fresh[670], Fresh[669], Fresh[668], Fresh[667], Fresh[666], Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660], Fresh[659], Fresh[658], Fresh[657], Fresh[656], Fresh[655], Fresh[654], Fresh[653], Fresh[652], Fresh[651], Fresh[650], Fresh[649], Fresh[648], Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642], Fresh[641], Fresh[640]}), .O ({new_AGEMA_signal_1871, \Inst_bSbox/b5 [1]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'hF8045F7B6D98DD7F ) ) \Inst_bSbox/b5_0 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r ({Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762], Fresh[761], Fresh[760], Fresh[759], Fresh[758], Fresh[757], Fresh[756], Fresh[755], Fresh[754], Fresh[753], Fresh[752], Fresh[751], Fresh[750], Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744], Fresh[743], Fresh[742], Fresh[741], Fresh[740], Fresh[739], Fresh[738], Fresh[737], Fresh[736], Fresh[735], Fresh[734], Fresh[733], Fresh[732], Fresh[731], Fresh[730], Fresh[729], Fresh[728], Fresh[727], Fresh[726], Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720], Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714], Fresh[713], Fresh[712], Fresh[711], Fresh[710], Fresh[709], Fresh[708], Fresh[707], Fresh[706], Fresh[705], Fresh[704]}), .O ({new_AGEMA_signal_1872, \Inst_bSbox/b5 [0]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'hF210A3AECE472E53 ) ) \Inst_bSbox/b4_3 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r ({Fresh[831], Fresh[830], Fresh[829], Fresh[828], Fresh[827], Fresh[826], Fresh[825], Fresh[824], Fresh[823], Fresh[822], Fresh[821], Fresh[820], Fresh[819], Fresh[818], Fresh[817], Fresh[816], Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810], Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804], Fresh[803], Fresh[802], Fresh[801], Fresh[800], Fresh[799], Fresh[798], Fresh[797], Fresh[796], Fresh[795], Fresh[794], Fresh[793], Fresh[792], Fresh[791], Fresh[790], Fresh[789], Fresh[788], Fresh[787], Fresh[786], Fresh[785], Fresh[784], Fresh[783], Fresh[782], Fresh[781], Fresh[780], Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774], Fresh[773], Fresh[772], Fresh[771], Fresh[770], Fresh[769], Fresh[768]}), .O ({new_AGEMA_signal_1873, \Inst_bSbox/b4 [3]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'h2624B286BC48ECB4 ) ) \Inst_bSbox/b4_2 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r ({Fresh[895], Fresh[894], Fresh[893], Fresh[892], Fresh[891], Fresh[890], Fresh[889], Fresh[888], Fresh[887], Fresh[886], Fresh[885], Fresh[884], Fresh[883], Fresh[882], Fresh[881], Fresh[880], Fresh[879], Fresh[878], Fresh[877], Fresh[876], Fresh[875], Fresh[874], Fresh[873], Fresh[872], Fresh[871], Fresh[870], Fresh[869], Fresh[868], Fresh[867], Fresh[866], Fresh[865], Fresh[864], Fresh[863], Fresh[862], Fresh[861], Fresh[860], Fresh[859], Fresh[858], Fresh[857], Fresh[856], Fresh[855], Fresh[854], Fresh[853], Fresh[852], Fresh[851], Fresh[850], Fresh[849], Fresh[848], Fresh[847], Fresh[846], Fresh[845], Fresh[844], Fresh[843], Fresh[842], Fresh[841], Fresh[840], Fresh[839], Fresh[838], Fresh[837], Fresh[836], Fresh[835], Fresh[834], Fresh[833], Fresh[832]}), .O ({new_AGEMA_signal_1874, \Inst_bSbox/b4 [2]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'hF7F17A494CE30F58 ) ) \Inst_bSbox/b4_1 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r ({Fresh[959], Fresh[958], Fresh[957], Fresh[956], Fresh[955], Fresh[954], Fresh[953], Fresh[952], Fresh[951], Fresh[950], Fresh[949], Fresh[948], Fresh[947], Fresh[946], Fresh[945], Fresh[944], Fresh[943], Fresh[942], Fresh[941], Fresh[940], Fresh[939], Fresh[938], Fresh[937], Fresh[936], Fresh[935], Fresh[934], Fresh[933], Fresh[932], Fresh[931], Fresh[930], Fresh[929], Fresh[928], Fresh[927], Fresh[926], Fresh[925], Fresh[924], Fresh[923], Fresh[922], Fresh[921], Fresh[920], Fresh[919], Fresh[918], Fresh[917], Fresh[916], Fresh[915], Fresh[914], Fresh[913], Fresh[912], Fresh[911], Fresh[910], Fresh[909], Fresh[908], Fresh[907], Fresh[906], Fresh[905], Fresh[904], Fresh[903], Fresh[902], Fresh[901], Fresh[900], Fresh[899], Fresh[898], Fresh[897], Fresh[896]}), .O ({new_AGEMA_signal_1875, \Inst_bSbox/b4 [1]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'hC2B0F97752B8B11E ) ) \Inst_bSbox/b4_0 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r ({Fresh[1023], Fresh[1022], Fresh[1021], Fresh[1020], Fresh[1019], Fresh[1018], Fresh[1017], Fresh[1016], Fresh[1015], Fresh[1014], Fresh[1013], Fresh[1012], Fresh[1011], Fresh[1010], Fresh[1009], Fresh[1008], Fresh[1007], Fresh[1006], Fresh[1005], Fresh[1004], Fresh[1003], Fresh[1002], Fresh[1001], Fresh[1000], Fresh[999], Fresh[998], Fresh[997], Fresh[996], Fresh[995], Fresh[994], Fresh[993], Fresh[992], Fresh[991], Fresh[990], Fresh[989], Fresh[988], Fresh[987], Fresh[986], Fresh[985], Fresh[984], Fresh[983], Fresh[982], Fresh[981], Fresh[980], Fresh[979], Fresh[978], Fresh[977], Fresh[976], Fresh[975], Fresh[974], Fresh[973], Fresh[972], Fresh[971], Fresh[970], Fresh[969], Fresh[968], Fresh[967], Fresh[966], Fresh[965], Fresh[964], Fresh[963], Fresh[962], Fresh[961], Fresh[960]}), .O ({new_AGEMA_signal_1876, \Inst_bSbox/b4 [0]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'h4E9DDB76C892FB1B ) ) \Inst_bSbox/b3_3 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r ({Fresh[1087], Fresh[1086], Fresh[1085], Fresh[1084], Fresh[1083], Fresh[1082], Fresh[1081], Fresh[1080], Fresh[1079], Fresh[1078], Fresh[1077], Fresh[1076], Fresh[1075], Fresh[1074], Fresh[1073], Fresh[1072], Fresh[1071], Fresh[1070], Fresh[1069], Fresh[1068], Fresh[1067], Fresh[1066], Fresh[1065], Fresh[1064], Fresh[1063], Fresh[1062], Fresh[1061], Fresh[1060], Fresh[1059], Fresh[1058], Fresh[1057], Fresh[1056], Fresh[1055], Fresh[1054], Fresh[1053], Fresh[1052], Fresh[1051], Fresh[1050], Fresh[1049], Fresh[1048], Fresh[1047], Fresh[1046], Fresh[1045], Fresh[1044], Fresh[1043], Fresh[1042], Fresh[1041], Fresh[1040], Fresh[1039], Fresh[1038], Fresh[1037], Fresh[1036], Fresh[1035], Fresh[1034], Fresh[1033], Fresh[1032], Fresh[1031], Fresh[1030], Fresh[1029], Fresh[1028], Fresh[1027], Fresh[1026], Fresh[1025], Fresh[1024]}), .O ({new_AGEMA_signal_1877, \Inst_bSbox/b3 [3]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'hE9DA849CF6AC6C1B ) ) \Inst_bSbox/b3_2 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r ({Fresh[1151], Fresh[1150], Fresh[1149], Fresh[1148], Fresh[1147], Fresh[1146], Fresh[1145], Fresh[1144], Fresh[1143], Fresh[1142], Fresh[1141], Fresh[1140], Fresh[1139], Fresh[1138], Fresh[1137], Fresh[1136], Fresh[1135], Fresh[1134], Fresh[1133], Fresh[1132], Fresh[1131], Fresh[1130], Fresh[1129], Fresh[1128], Fresh[1127], Fresh[1126], Fresh[1125], Fresh[1124], Fresh[1123], Fresh[1122], Fresh[1121], Fresh[1120], Fresh[1119], Fresh[1118], Fresh[1117], Fresh[1116], Fresh[1115], Fresh[1114], Fresh[1113], Fresh[1112], Fresh[1111], Fresh[1110], Fresh[1109], Fresh[1108], Fresh[1107], Fresh[1106], Fresh[1105], Fresh[1104], Fresh[1103], Fresh[1102], Fresh[1101], Fresh[1100], Fresh[1099], Fresh[1098], Fresh[1097], Fresh[1096], Fresh[1095], Fresh[1094], Fresh[1093], Fresh[1092], Fresh[1091], Fresh[1090], Fresh[1089], Fresh[1088]}), .O ({new_AGEMA_signal_1878, \Inst_bSbox/b3 [2]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'h2568EA2EFFA8527D ) ) \Inst_bSbox/b3_1 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r ({Fresh[1215], Fresh[1214], Fresh[1213], Fresh[1212], Fresh[1211], Fresh[1210], Fresh[1209], Fresh[1208], Fresh[1207], Fresh[1206], Fresh[1205], Fresh[1204], Fresh[1203], Fresh[1202], Fresh[1201], Fresh[1200], Fresh[1199], Fresh[1198], Fresh[1197], Fresh[1196], Fresh[1195], Fresh[1194], Fresh[1193], Fresh[1192], Fresh[1191], Fresh[1190], Fresh[1189], Fresh[1188], Fresh[1187], Fresh[1186], Fresh[1185], Fresh[1184], Fresh[1183], Fresh[1182], Fresh[1181], Fresh[1180], Fresh[1179], Fresh[1178], Fresh[1177], Fresh[1176], Fresh[1175], Fresh[1174], Fresh[1173], Fresh[1172], Fresh[1171], Fresh[1170], Fresh[1169], Fresh[1168], Fresh[1167], Fresh[1166], Fresh[1165], Fresh[1164], Fresh[1163], Fresh[1162], Fresh[1161], Fresh[1160], Fresh[1159], Fresh[1158], Fresh[1157], Fresh[1156], Fresh[1155], Fresh[1154], Fresh[1153], Fresh[1152]}), .O ({new_AGEMA_signal_1879, \Inst_bSbox/b3 [1]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'h109020A2193D586A ) ) \Inst_bSbox/b3_0 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r ({Fresh[1279], Fresh[1278], Fresh[1277], Fresh[1276], Fresh[1275], Fresh[1274], Fresh[1273], Fresh[1272], Fresh[1271], Fresh[1270], Fresh[1269], Fresh[1268], Fresh[1267], Fresh[1266], Fresh[1265], Fresh[1264], Fresh[1263], Fresh[1262], Fresh[1261], Fresh[1260], Fresh[1259], Fresh[1258], Fresh[1257], Fresh[1256], Fresh[1255], Fresh[1254], Fresh[1253], Fresh[1252], Fresh[1251], Fresh[1250], Fresh[1249], Fresh[1248], Fresh[1247], Fresh[1246], Fresh[1245], Fresh[1244], Fresh[1243], Fresh[1242], Fresh[1241], Fresh[1240], Fresh[1239], Fresh[1238], Fresh[1237], Fresh[1236], Fresh[1235], Fresh[1234], Fresh[1233], Fresh[1232], Fresh[1231], Fresh[1230], Fresh[1229], Fresh[1228], Fresh[1227], Fresh[1226], Fresh[1225], Fresh[1224], Fresh[1223], Fresh[1222], Fresh[1221], Fresh[1220], Fresh[1219], Fresh[1218], Fresh[1217], Fresh[1216]}), .O ({new_AGEMA_signal_1880, \Inst_bSbox/b3 [0]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'hAC39B6C0D6CE2EFC ) ) \Inst_bSbox/b2_3 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r ({Fresh[1343], Fresh[1342], Fresh[1341], Fresh[1340], Fresh[1339], Fresh[1338], Fresh[1337], Fresh[1336], Fresh[1335], Fresh[1334], Fresh[1333], Fresh[1332], Fresh[1331], Fresh[1330], Fresh[1329], Fresh[1328], Fresh[1327], Fresh[1326], Fresh[1325], Fresh[1324], Fresh[1323], Fresh[1322], Fresh[1321], Fresh[1320], Fresh[1319], Fresh[1318], Fresh[1317], Fresh[1316], Fresh[1315], Fresh[1314], Fresh[1313], Fresh[1312], Fresh[1311], Fresh[1310], Fresh[1309], Fresh[1308], Fresh[1307], Fresh[1306], Fresh[1305], Fresh[1304], Fresh[1303], Fresh[1302], Fresh[1301], Fresh[1300], Fresh[1299], Fresh[1298], Fresh[1297], Fresh[1296], Fresh[1295], Fresh[1294], Fresh[1293], Fresh[1292], Fresh[1291], Fresh[1290], Fresh[1289], Fresh[1288], Fresh[1287], Fresh[1286], Fresh[1285], Fresh[1284], Fresh[1283], Fresh[1282], Fresh[1281], Fresh[1280]}), .O ({new_AGEMA_signal_1881, \Inst_bSbox/b2 [3]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'h577D64E03B0C3FFB ) ) \Inst_bSbox/b2_2 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r ({Fresh[1407], Fresh[1406], Fresh[1405], Fresh[1404], Fresh[1403], Fresh[1402], Fresh[1401], Fresh[1400], Fresh[1399], Fresh[1398], Fresh[1397], Fresh[1396], Fresh[1395], Fresh[1394], Fresh[1393], Fresh[1392], Fresh[1391], Fresh[1390], Fresh[1389], Fresh[1388], Fresh[1387], Fresh[1386], Fresh[1385], Fresh[1384], Fresh[1383], Fresh[1382], Fresh[1381], Fresh[1380], Fresh[1379], Fresh[1378], Fresh[1377], Fresh[1376], Fresh[1375], Fresh[1374], Fresh[1373], Fresh[1372], Fresh[1371], Fresh[1370], Fresh[1369], Fresh[1368], Fresh[1367], Fresh[1366], Fresh[1365], Fresh[1364], Fresh[1363], Fresh[1362], Fresh[1361], Fresh[1360], Fresh[1359], Fresh[1358], Fresh[1357], Fresh[1356], Fresh[1355], Fresh[1354], Fresh[1353], Fresh[1352], Fresh[1351], Fresh[1350], Fresh[1349], Fresh[1348], Fresh[1347], Fresh[1346], Fresh[1345], Fresh[1344]}), .O ({new_AGEMA_signal_1882, \Inst_bSbox/b2 [2]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'h23A869A2A428C424 ) ) \Inst_bSbox/b2_1 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r ({Fresh[1471], Fresh[1470], Fresh[1469], Fresh[1468], Fresh[1467], Fresh[1466], Fresh[1465], Fresh[1464], Fresh[1463], Fresh[1462], Fresh[1461], Fresh[1460], Fresh[1459], Fresh[1458], Fresh[1457], Fresh[1456], Fresh[1455], Fresh[1454], Fresh[1453], Fresh[1452], Fresh[1451], Fresh[1450], Fresh[1449], Fresh[1448], Fresh[1447], Fresh[1446], Fresh[1445], Fresh[1444], Fresh[1443], Fresh[1442], Fresh[1441], Fresh[1440], Fresh[1439], Fresh[1438], Fresh[1437], Fresh[1436], Fresh[1435], Fresh[1434], Fresh[1433], Fresh[1432], Fresh[1431], Fresh[1430], Fresh[1429], Fresh[1428], Fresh[1427], Fresh[1426], Fresh[1425], Fresh[1424], Fresh[1423], Fresh[1422], Fresh[1421], Fresh[1420], Fresh[1419], Fresh[1418], Fresh[1417], Fresh[1416], Fresh[1415], Fresh[1414], Fresh[1413], Fresh[1412], Fresh[1411], Fresh[1410], Fresh[1409], Fresh[1408]}), .O ({new_AGEMA_signal_1883, \Inst_bSbox/b2 [1]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'hA16387FB3B48B4C6 ) ) \Inst_bSbox/b2_0 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r ({Fresh[1535], Fresh[1534], Fresh[1533], Fresh[1532], Fresh[1531], Fresh[1530], Fresh[1529], Fresh[1528], Fresh[1527], Fresh[1526], Fresh[1525], Fresh[1524], Fresh[1523], Fresh[1522], Fresh[1521], Fresh[1520], Fresh[1519], Fresh[1518], Fresh[1517], Fresh[1516], Fresh[1515], Fresh[1514], Fresh[1513], Fresh[1512], Fresh[1511], Fresh[1510], Fresh[1509], Fresh[1508], Fresh[1507], Fresh[1506], Fresh[1505], Fresh[1504], Fresh[1503], Fresh[1502], Fresh[1501], Fresh[1500], Fresh[1499], Fresh[1498], Fresh[1497], Fresh[1496], Fresh[1495], Fresh[1494], Fresh[1493], Fresh[1492], Fresh[1491], Fresh[1490], Fresh[1489], Fresh[1488], Fresh[1487], Fresh[1486], Fresh[1485], Fresh[1484], Fresh[1483], Fresh[1482], Fresh[1481], Fresh[1480], Fresh[1479], Fresh[1478], Fresh[1477], Fresh[1476], Fresh[1475], Fresh[1474], Fresh[1473], Fresh[1472]}), .O ({new_AGEMA_signal_1884, \Inst_bSbox/b2 [0]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'hC870974094EAD8A9 ) ) \Inst_bSbox/b1_3 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r ({Fresh[1599], Fresh[1598], Fresh[1597], Fresh[1596], Fresh[1595], Fresh[1594], Fresh[1593], Fresh[1592], Fresh[1591], Fresh[1590], Fresh[1589], Fresh[1588], Fresh[1587], Fresh[1586], Fresh[1585], Fresh[1584], Fresh[1583], Fresh[1582], Fresh[1581], Fresh[1580], Fresh[1579], Fresh[1578], Fresh[1577], Fresh[1576], Fresh[1575], Fresh[1574], Fresh[1573], Fresh[1572], Fresh[1571], Fresh[1570], Fresh[1569], Fresh[1568], Fresh[1567], Fresh[1566], Fresh[1565], Fresh[1564], Fresh[1563], Fresh[1562], Fresh[1561], Fresh[1560], Fresh[1559], Fresh[1558], Fresh[1557], Fresh[1556], Fresh[1555], Fresh[1554], Fresh[1553], Fresh[1552], Fresh[1551], Fresh[1550], Fresh[1549], Fresh[1548], Fresh[1547], Fresh[1546], Fresh[1545], Fresh[1544], Fresh[1543], Fresh[1542], Fresh[1541], Fresh[1540], Fresh[1539], Fresh[1538], Fresh[1537], Fresh[1536]}), .O ({new_AGEMA_signal_1885, \Inst_bSbox/b1 [3]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6A450B2EF33486B4 ) ) \Inst_bSbox/b1_2 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r ({Fresh[1663], Fresh[1662], Fresh[1661], Fresh[1660], Fresh[1659], Fresh[1658], Fresh[1657], Fresh[1656], Fresh[1655], Fresh[1654], Fresh[1653], Fresh[1652], Fresh[1651], Fresh[1650], Fresh[1649], Fresh[1648], Fresh[1647], Fresh[1646], Fresh[1645], Fresh[1644], Fresh[1643], Fresh[1642], Fresh[1641], Fresh[1640], Fresh[1639], Fresh[1638], Fresh[1637], Fresh[1636], Fresh[1635], Fresh[1634], Fresh[1633], Fresh[1632], Fresh[1631], Fresh[1630], Fresh[1629], Fresh[1628], Fresh[1627], Fresh[1626], Fresh[1625], Fresh[1624], Fresh[1623], Fresh[1622], Fresh[1621], Fresh[1620], Fresh[1619], Fresh[1618], Fresh[1617], Fresh[1616], Fresh[1615], Fresh[1614], Fresh[1613], Fresh[1612], Fresh[1611], Fresh[1610], Fresh[1609], Fresh[1608], Fresh[1607], Fresh[1606], Fresh[1605], Fresh[1604], Fresh[1603], Fresh[1602], Fresh[1601], Fresh[1600]}), .O ({new_AGEMA_signal_1886, \Inst_bSbox/b1 [2]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'hE61A4C5E97816F7A ) ) \Inst_bSbox/b1_1 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r ({Fresh[1727], Fresh[1726], Fresh[1725], Fresh[1724], Fresh[1723], Fresh[1722], Fresh[1721], Fresh[1720], Fresh[1719], Fresh[1718], Fresh[1717], Fresh[1716], Fresh[1715], Fresh[1714], Fresh[1713], Fresh[1712], Fresh[1711], Fresh[1710], Fresh[1709], Fresh[1708], Fresh[1707], Fresh[1706], Fresh[1705], Fresh[1704], Fresh[1703], Fresh[1702], Fresh[1701], Fresh[1700], Fresh[1699], Fresh[1698], Fresh[1697], Fresh[1696], Fresh[1695], Fresh[1694], Fresh[1693], Fresh[1692], Fresh[1691], Fresh[1690], Fresh[1689], Fresh[1688], Fresh[1687], Fresh[1686], Fresh[1685], Fresh[1684], Fresh[1683], Fresh[1682], Fresh[1681], Fresh[1680], Fresh[1679], Fresh[1678], Fresh[1677], Fresh[1676], Fresh[1675], Fresh[1674], Fresh[1673], Fresh[1672], Fresh[1671], Fresh[1670], Fresh[1669], Fresh[1668], Fresh[1667], Fresh[1666], Fresh[1665], Fresh[1664]}), .O ({new_AGEMA_signal_1887, \Inst_bSbox/b1 [1]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'h7BAE007D4C53FC7D ) ) \Inst_bSbox/b1_0 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r ({Fresh[1791], Fresh[1790], Fresh[1789], Fresh[1788], Fresh[1787], Fresh[1786], Fresh[1785], Fresh[1784], Fresh[1783], Fresh[1782], Fresh[1781], Fresh[1780], Fresh[1779], Fresh[1778], Fresh[1777], Fresh[1776], Fresh[1775], Fresh[1774], Fresh[1773], Fresh[1772], Fresh[1771], Fresh[1770], Fresh[1769], Fresh[1768], Fresh[1767], Fresh[1766], Fresh[1765], Fresh[1764], Fresh[1763], Fresh[1762], Fresh[1761], Fresh[1760], Fresh[1759], Fresh[1758], Fresh[1757], Fresh[1756], Fresh[1755], Fresh[1754], Fresh[1753], Fresh[1752], Fresh[1751], Fresh[1750], Fresh[1749], Fresh[1748], Fresh[1747], Fresh[1746], Fresh[1745], Fresh[1744], Fresh[1743], Fresh[1742], Fresh[1741], Fresh[1740], Fresh[1739], Fresh[1738], Fresh[1737], Fresh[1736], Fresh[1735], Fresh[1734], Fresh[1733], Fresh[1732], Fresh[1731], Fresh[1730], Fresh[1729], Fresh[1728]}), .O ({new_AGEMA_signal_1888, \Inst_bSbox/b1 [0]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'h4F1EAD396F247A04 ) ) \Inst_bSbox/b0_3 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r ({Fresh[1855], Fresh[1854], Fresh[1853], Fresh[1852], Fresh[1851], Fresh[1850], Fresh[1849], Fresh[1848], Fresh[1847], Fresh[1846], Fresh[1845], Fresh[1844], Fresh[1843], Fresh[1842], Fresh[1841], Fresh[1840], Fresh[1839], Fresh[1838], Fresh[1837], Fresh[1836], Fresh[1835], Fresh[1834], Fresh[1833], Fresh[1832], Fresh[1831], Fresh[1830], Fresh[1829], Fresh[1828], Fresh[1827], Fresh[1826], Fresh[1825], Fresh[1824], Fresh[1823], Fresh[1822], Fresh[1821], Fresh[1820], Fresh[1819], Fresh[1818], Fresh[1817], Fresh[1816], Fresh[1815], Fresh[1814], Fresh[1813], Fresh[1812], Fresh[1811], Fresh[1810], Fresh[1809], Fresh[1808], Fresh[1807], Fresh[1806], Fresh[1805], Fresh[1804], Fresh[1803], Fresh[1802], Fresh[1801], Fresh[1800], Fresh[1799], Fresh[1798], Fresh[1797], Fresh[1796], Fresh[1795], Fresh[1794], Fresh[1793], Fresh[1792]}), .O ({new_AGEMA_signal_1889, \Inst_bSbox/b0 [3]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'h10BDB210C006EAB5 ) ) \Inst_bSbox/b0_2 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r ({Fresh[1919], Fresh[1918], Fresh[1917], Fresh[1916], Fresh[1915], Fresh[1914], Fresh[1913], Fresh[1912], Fresh[1911], Fresh[1910], Fresh[1909], Fresh[1908], Fresh[1907], Fresh[1906], Fresh[1905], Fresh[1904], Fresh[1903], Fresh[1902], Fresh[1901], Fresh[1900], Fresh[1899], Fresh[1898], Fresh[1897], Fresh[1896], Fresh[1895], Fresh[1894], Fresh[1893], Fresh[1892], Fresh[1891], Fresh[1890], Fresh[1889], Fresh[1888], Fresh[1887], Fresh[1886], Fresh[1885], Fresh[1884], Fresh[1883], Fresh[1882], Fresh[1881], Fresh[1880], Fresh[1879], Fresh[1878], Fresh[1877], Fresh[1876], Fresh[1875], Fresh[1874], Fresh[1873], Fresh[1872], Fresh[1871], Fresh[1870], Fresh[1869], Fresh[1868], Fresh[1867], Fresh[1866], Fresh[1865], Fresh[1864], Fresh[1863], Fresh[1862], Fresh[1861], Fresh[1860], Fresh[1859], Fresh[1858], Fresh[1857], Fresh[1856]}), .O ({new_AGEMA_signal_1890, \Inst_bSbox/b0 [2]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'h68AB4BFA8ACB7A13 ) ) \Inst_bSbox/b0_1 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r ({Fresh[1983], Fresh[1982], Fresh[1981], Fresh[1980], Fresh[1979], Fresh[1978], Fresh[1977], Fresh[1976], Fresh[1975], Fresh[1974], Fresh[1973], Fresh[1972], Fresh[1971], Fresh[1970], Fresh[1969], Fresh[1968], Fresh[1967], Fresh[1966], Fresh[1965], Fresh[1964], Fresh[1963], Fresh[1962], Fresh[1961], Fresh[1960], Fresh[1959], Fresh[1958], Fresh[1957], Fresh[1956], Fresh[1955], Fresh[1954], Fresh[1953], Fresh[1952], Fresh[1951], Fresh[1950], Fresh[1949], Fresh[1948], Fresh[1947], Fresh[1946], Fresh[1945], Fresh[1944], Fresh[1943], Fresh[1942], Fresh[1941], Fresh[1940], Fresh[1939], Fresh[1938], Fresh[1937], Fresh[1936], Fresh[1935], Fresh[1934], Fresh[1933], Fresh[1932], Fresh[1931], Fresh[1930], Fresh[1929], Fresh[1928], Fresh[1927], Fresh[1926], Fresh[1925], Fresh[1924], Fresh[1923], Fresh[1922], Fresh[1921], Fresh[1920]}), .O ({new_AGEMA_signal_1891, \Inst_bSbox/b0 [1]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'hB14EDE67096C6EED ) ) \Inst_bSbox/b0_0 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r ({Fresh[2047], Fresh[2046], Fresh[2045], Fresh[2044], Fresh[2043], Fresh[2042], Fresh[2041], Fresh[2040], Fresh[2039], Fresh[2038], Fresh[2037], Fresh[2036], Fresh[2035], Fresh[2034], Fresh[2033], Fresh[2032], Fresh[2031], Fresh[2030], Fresh[2029], Fresh[2028], Fresh[2027], Fresh[2026], Fresh[2025], Fresh[2024], Fresh[2023], Fresh[2022], Fresh[2021], Fresh[2020], Fresh[2019], Fresh[2018], Fresh[2017], Fresh[2016], Fresh[2015], Fresh[2014], Fresh[2013], Fresh[2012], Fresh[2011], Fresh[2010], Fresh[2009], Fresh[2008], Fresh[2007], Fresh[2006], Fresh[2005], Fresh[2004], Fresh[2003], Fresh[2002], Fresh[2001], Fresh[2000], Fresh[1999], Fresh[1998], Fresh[1997], Fresh[1996], Fresh[1995], Fresh[1994], Fresh[1993], Fresh[1992], Fresh[1991], Fresh[1990], Fresh[1989], Fresh[1988], Fresh[1987], Fresh[1986], Fresh[1985], Fresh[1984]}), .O ({new_AGEMA_signal_1892, \Inst_bSbox/b0 [0]}) ) ;

    /* cells in depth 2 */
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hAAAAF0CC ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hAAAAF0CC ) ) \stateArray/gen33ser[7].Inst1 ( .I0 ({new_AGEMA_signal_1900, StateInMC[7]}), .I1 ({new_AGEMA_signal_2157, SboxOut[7]}), .I2 ({new_AGEMA_signal_1351, StateOutXORroundKey[7]}), .I3 ({1'b0, intFinal}), .I4 ({1'b0, selMC}), .O ({new_AGEMA_signal_2213, \stateArray/input_MC [7]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hAAAAF0CC ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hAAAAF0CC ) ) \stateArray/gen33ser[6].Inst1 ( .I0 ({new_AGEMA_signal_1899, StateInMC[6]}), .I1 ({new_AGEMA_signal_2158, SboxOut[6]}), .I2 ({new_AGEMA_signal_1354, StateOutXORroundKey[6]}), .I3 ({1'b0, intFinal}), .I4 ({1'b0, selMC}), .O ({new_AGEMA_signal_2214, \stateArray/input_MC [6]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hAAAAF0CC ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hAAAAF0CC ) ) \stateArray/gen33ser[5].Inst1 ( .I0 ({new_AGEMA_signal_1898, StateInMC[5]}), .I1 ({new_AGEMA_signal_2159, SboxOut[5]}), .I2 ({new_AGEMA_signal_1357, StateOutXORroundKey[5]}), .I3 ({1'b0, intFinal}), .I4 ({1'b0, selMC}), .O ({new_AGEMA_signal_2215, \stateArray/input_MC [5]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hAAAAF0CC ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hAAAAF0CC ) ) \stateArray/gen33ser[4].Inst1 ( .I0 ({new_AGEMA_signal_1897, StateInMC[4]}), .I1 ({new_AGEMA_signal_2160, SboxOut[4]}), .I2 ({new_AGEMA_signal_1360, StateOutXORroundKey[4]}), .I3 ({1'b0, intFinal}), .I4 ({1'b0, selMC}), .O ({new_AGEMA_signal_2216, \stateArray/input_MC [4]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hAAAAF0CC ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hAAAAF0CC ) ) \stateArray/gen33ser[3].Inst1 ( .I0 ({new_AGEMA_signal_1896, StateInMC[3]}), .I1 ({new_AGEMA_signal_2161, SboxOut[3]}), .I2 ({new_AGEMA_signal_1363, StateOutXORroundKey[3]}), .I3 ({1'b0, intFinal}), .I4 ({1'b0, selMC}), .O ({new_AGEMA_signal_2217, \stateArray/input_MC [3]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hAAAAF0CC ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hAAAAF0CC ) ) \stateArray/gen33ser[2].Inst1 ( .I0 ({new_AGEMA_signal_1895, StateInMC[2]}), .I1 ({new_AGEMA_signal_2162, SboxOut[2]}), .I2 ({new_AGEMA_signal_1366, StateOutXORroundKey[2]}), .I3 ({1'b0, intFinal}), .I4 ({1'b0, selMC}), .O ({new_AGEMA_signal_2218, \stateArray/input_MC [2]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hAAAAF0CC ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hAAAAF0CC ) ) \stateArray/gen33ser[1].Inst1 ( .I0 ({new_AGEMA_signal_1894, StateInMC[1]}), .I1 ({new_AGEMA_signal_2163, SboxOut[1]}), .I2 ({new_AGEMA_signal_1369, StateOutXORroundKey[1]}), .I3 ({1'b0, intFinal}), .I4 ({1'b0, selMC}), .O ({new_AGEMA_signal_2219, \stateArray/input_MC [1]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hAAAAF0CC ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hAAAAF0CC ) ) \stateArray/gen33ser[0].Inst1 ( .I0 ({new_AGEMA_signal_1893, StateInMC[0]}), .I1 ({new_AGEMA_signal_2164, SboxOut[0]}), .I2 ({new_AGEMA_signal_1372, StateOutXORroundKey[0]}), .I3 ({1'b0, intFinal}), .I4 ({1'b0, selMC}), .O ({new_AGEMA_signal_2220, \stateArray/input_MC [0]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \Inst_bSbox/b7_4 ( .I0 ({new_AGEMA_signal_1864, \Inst_bSbox/b7 [0]}), .I1 ({new_AGEMA_signal_1863, \Inst_bSbox/b7 [1]}), .I2 ({new_AGEMA_signal_1862, \Inst_bSbox/b7 [2]}), .I3 ({new_AGEMA_signal_1861, \Inst_bSbox/b7 [3]}), .I4 ({new_AGEMA_signal_1438, SboxIn[6]}), .I5 ({new_AGEMA_signal_1436, SboxIn[7]}), .clk (clk), .r ({Fresh[2111], Fresh[2110], Fresh[2109], Fresh[2108], Fresh[2107], Fresh[2106], Fresh[2105], Fresh[2104], Fresh[2103], Fresh[2102], Fresh[2101], Fresh[2100], Fresh[2099], Fresh[2098], Fresh[2097], Fresh[2096], Fresh[2095], Fresh[2094], Fresh[2093], Fresh[2092], Fresh[2091], Fresh[2090], Fresh[2089], Fresh[2088], Fresh[2087], Fresh[2086], Fresh[2085], Fresh[2084], Fresh[2083], Fresh[2082], Fresh[2081], Fresh[2080], Fresh[2079], Fresh[2078], Fresh[2077], Fresh[2076], Fresh[2075], Fresh[2074], Fresh[2073], Fresh[2072], Fresh[2071], Fresh[2070], Fresh[2069], Fresh[2068], Fresh[2067], Fresh[2066], Fresh[2065], Fresh[2064], Fresh[2063], Fresh[2062], Fresh[2061], Fresh[2060], Fresh[2059], Fresh[2058], Fresh[2057], Fresh[2056], Fresh[2055], Fresh[2054], Fresh[2053], Fresh[2052], Fresh[2051], Fresh[2050], Fresh[2049], Fresh[2048]}), .O ({new_AGEMA_signal_2157, SboxOut[7]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \Inst_bSbox/b6_4 ( .I0 ({new_AGEMA_signal_1868, \Inst_bSbox/b6 [0]}), .I1 ({new_AGEMA_signal_1867, \Inst_bSbox/b6 [1]}), .I2 ({new_AGEMA_signal_1866, \Inst_bSbox/b6 [2]}), .I3 ({new_AGEMA_signal_1865, \Inst_bSbox/b6 [3]}), .I4 ({new_AGEMA_signal_1438, SboxIn[6]}), .I5 ({new_AGEMA_signal_1436, SboxIn[7]}), .clk (clk), .r ({Fresh[2175], Fresh[2174], Fresh[2173], Fresh[2172], Fresh[2171], Fresh[2170], Fresh[2169], Fresh[2168], Fresh[2167], Fresh[2166], Fresh[2165], Fresh[2164], Fresh[2163], Fresh[2162], Fresh[2161], Fresh[2160], Fresh[2159], Fresh[2158], Fresh[2157], Fresh[2156], Fresh[2155], Fresh[2154], Fresh[2153], Fresh[2152], Fresh[2151], Fresh[2150], Fresh[2149], Fresh[2148], Fresh[2147], Fresh[2146], Fresh[2145], Fresh[2144], Fresh[2143], Fresh[2142], Fresh[2141], Fresh[2140], Fresh[2139], Fresh[2138], Fresh[2137], Fresh[2136], Fresh[2135], Fresh[2134], Fresh[2133], Fresh[2132], Fresh[2131], Fresh[2130], Fresh[2129], Fresh[2128], Fresh[2127], Fresh[2126], Fresh[2125], Fresh[2124], Fresh[2123], Fresh[2122], Fresh[2121], Fresh[2120], Fresh[2119], Fresh[2118], Fresh[2117], Fresh[2116], Fresh[2115], Fresh[2114], Fresh[2113], Fresh[2112]}), .O ({new_AGEMA_signal_2158, SboxOut[6]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \Inst_bSbox/b5_4 ( .I0 ({new_AGEMA_signal_1872, \Inst_bSbox/b5 [0]}), .I1 ({new_AGEMA_signal_1871, \Inst_bSbox/b5 [1]}), .I2 ({new_AGEMA_signal_1870, \Inst_bSbox/b5 [2]}), .I3 ({new_AGEMA_signal_1869, \Inst_bSbox/b5 [3]}), .I4 ({new_AGEMA_signal_1438, SboxIn[6]}), .I5 ({new_AGEMA_signal_1436, SboxIn[7]}), .clk (clk), .r ({Fresh[2239], Fresh[2238], Fresh[2237], Fresh[2236], Fresh[2235], Fresh[2234], Fresh[2233], Fresh[2232], Fresh[2231], Fresh[2230], Fresh[2229], Fresh[2228], Fresh[2227], Fresh[2226], Fresh[2225], Fresh[2224], Fresh[2223], Fresh[2222], Fresh[2221], Fresh[2220], Fresh[2219], Fresh[2218], Fresh[2217], Fresh[2216], Fresh[2215], Fresh[2214], Fresh[2213], Fresh[2212], Fresh[2211], Fresh[2210], Fresh[2209], Fresh[2208], Fresh[2207], Fresh[2206], Fresh[2205], Fresh[2204], Fresh[2203], Fresh[2202], Fresh[2201], Fresh[2200], Fresh[2199], Fresh[2198], Fresh[2197], Fresh[2196], Fresh[2195], Fresh[2194], Fresh[2193], Fresh[2192], Fresh[2191], Fresh[2190], Fresh[2189], Fresh[2188], Fresh[2187], Fresh[2186], Fresh[2185], Fresh[2184], Fresh[2183], Fresh[2182], Fresh[2181], Fresh[2180], Fresh[2179], Fresh[2178], Fresh[2177], Fresh[2176]}), .O ({new_AGEMA_signal_2159, SboxOut[5]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \Inst_bSbox/b4_4 ( .I0 ({new_AGEMA_signal_1876, \Inst_bSbox/b4 [0]}), .I1 ({new_AGEMA_signal_1875, \Inst_bSbox/b4 [1]}), .I2 ({new_AGEMA_signal_1874, \Inst_bSbox/b4 [2]}), .I3 ({new_AGEMA_signal_1873, \Inst_bSbox/b4 [3]}), .I4 ({new_AGEMA_signal_1438, SboxIn[6]}), .I5 ({new_AGEMA_signal_1436, SboxIn[7]}), .clk (clk), .r ({Fresh[2303], Fresh[2302], Fresh[2301], Fresh[2300], Fresh[2299], Fresh[2298], Fresh[2297], Fresh[2296], Fresh[2295], Fresh[2294], Fresh[2293], Fresh[2292], Fresh[2291], Fresh[2290], Fresh[2289], Fresh[2288], Fresh[2287], Fresh[2286], Fresh[2285], Fresh[2284], Fresh[2283], Fresh[2282], Fresh[2281], Fresh[2280], Fresh[2279], Fresh[2278], Fresh[2277], Fresh[2276], Fresh[2275], Fresh[2274], Fresh[2273], Fresh[2272], Fresh[2271], Fresh[2270], Fresh[2269], Fresh[2268], Fresh[2267], Fresh[2266], Fresh[2265], Fresh[2264], Fresh[2263], Fresh[2262], Fresh[2261], Fresh[2260], Fresh[2259], Fresh[2258], Fresh[2257], Fresh[2256], Fresh[2255], Fresh[2254], Fresh[2253], Fresh[2252], Fresh[2251], Fresh[2250], Fresh[2249], Fresh[2248], Fresh[2247], Fresh[2246], Fresh[2245], Fresh[2244], Fresh[2243], Fresh[2242], Fresh[2241], Fresh[2240]}), .O ({new_AGEMA_signal_2160, SboxOut[4]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \Inst_bSbox/b3_4 ( .I0 ({new_AGEMA_signal_1880, \Inst_bSbox/b3 [0]}), .I1 ({new_AGEMA_signal_1879, \Inst_bSbox/b3 [1]}), .I2 ({new_AGEMA_signal_1878, \Inst_bSbox/b3 [2]}), .I3 ({new_AGEMA_signal_1877, \Inst_bSbox/b3 [3]}), .I4 ({new_AGEMA_signal_1438, SboxIn[6]}), .I5 ({new_AGEMA_signal_1436, SboxIn[7]}), .clk (clk), .r ({Fresh[2367], Fresh[2366], Fresh[2365], Fresh[2364], Fresh[2363], Fresh[2362], Fresh[2361], Fresh[2360], Fresh[2359], Fresh[2358], Fresh[2357], Fresh[2356], Fresh[2355], Fresh[2354], Fresh[2353], Fresh[2352], Fresh[2351], Fresh[2350], Fresh[2349], Fresh[2348], Fresh[2347], Fresh[2346], Fresh[2345], Fresh[2344], Fresh[2343], Fresh[2342], Fresh[2341], Fresh[2340], Fresh[2339], Fresh[2338], Fresh[2337], Fresh[2336], Fresh[2335], Fresh[2334], Fresh[2333], Fresh[2332], Fresh[2331], Fresh[2330], Fresh[2329], Fresh[2328], Fresh[2327], Fresh[2326], Fresh[2325], Fresh[2324], Fresh[2323], Fresh[2322], Fresh[2321], Fresh[2320], Fresh[2319], Fresh[2318], Fresh[2317], Fresh[2316], Fresh[2315], Fresh[2314], Fresh[2313], Fresh[2312], Fresh[2311], Fresh[2310], Fresh[2309], Fresh[2308], Fresh[2307], Fresh[2306], Fresh[2305], Fresh[2304]}), .O ({new_AGEMA_signal_2161, SboxOut[3]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \Inst_bSbox/b2_4 ( .I0 ({new_AGEMA_signal_1884, \Inst_bSbox/b2 [0]}), .I1 ({new_AGEMA_signal_1883, \Inst_bSbox/b2 [1]}), .I2 ({new_AGEMA_signal_1882, \Inst_bSbox/b2 [2]}), .I3 ({new_AGEMA_signal_1881, \Inst_bSbox/b2 [3]}), .I4 ({new_AGEMA_signal_1438, SboxIn[6]}), .I5 ({new_AGEMA_signal_1436, SboxIn[7]}), .clk (clk), .r ({Fresh[2431], Fresh[2430], Fresh[2429], Fresh[2428], Fresh[2427], Fresh[2426], Fresh[2425], Fresh[2424], Fresh[2423], Fresh[2422], Fresh[2421], Fresh[2420], Fresh[2419], Fresh[2418], Fresh[2417], Fresh[2416], Fresh[2415], Fresh[2414], Fresh[2413], Fresh[2412], Fresh[2411], Fresh[2410], Fresh[2409], Fresh[2408], Fresh[2407], Fresh[2406], Fresh[2405], Fresh[2404], Fresh[2403], Fresh[2402], Fresh[2401], Fresh[2400], Fresh[2399], Fresh[2398], Fresh[2397], Fresh[2396], Fresh[2395], Fresh[2394], Fresh[2393], Fresh[2392], Fresh[2391], Fresh[2390], Fresh[2389], Fresh[2388], Fresh[2387], Fresh[2386], Fresh[2385], Fresh[2384], Fresh[2383], Fresh[2382], Fresh[2381], Fresh[2380], Fresh[2379], Fresh[2378], Fresh[2377], Fresh[2376], Fresh[2375], Fresh[2374], Fresh[2373], Fresh[2372], Fresh[2371], Fresh[2370], Fresh[2369], Fresh[2368]}), .O ({new_AGEMA_signal_2162, SboxOut[2]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \Inst_bSbox/b1_4 ( .I0 ({new_AGEMA_signal_1888, \Inst_bSbox/b1 [0]}), .I1 ({new_AGEMA_signal_1887, \Inst_bSbox/b1 [1]}), .I2 ({new_AGEMA_signal_1886, \Inst_bSbox/b1 [2]}), .I3 ({new_AGEMA_signal_1885, \Inst_bSbox/b1 [3]}), .I4 ({new_AGEMA_signal_1438, SboxIn[6]}), .I5 ({new_AGEMA_signal_1436, SboxIn[7]}), .clk (clk), .r ({Fresh[2495], Fresh[2494], Fresh[2493], Fresh[2492], Fresh[2491], Fresh[2490], Fresh[2489], Fresh[2488], Fresh[2487], Fresh[2486], Fresh[2485], Fresh[2484], Fresh[2483], Fresh[2482], Fresh[2481], Fresh[2480], Fresh[2479], Fresh[2478], Fresh[2477], Fresh[2476], Fresh[2475], Fresh[2474], Fresh[2473], Fresh[2472], Fresh[2471], Fresh[2470], Fresh[2469], Fresh[2468], Fresh[2467], Fresh[2466], Fresh[2465], Fresh[2464], Fresh[2463], Fresh[2462], Fresh[2461], Fresh[2460], Fresh[2459], Fresh[2458], Fresh[2457], Fresh[2456], Fresh[2455], Fresh[2454], Fresh[2453], Fresh[2452], Fresh[2451], Fresh[2450], Fresh[2449], Fresh[2448], Fresh[2447], Fresh[2446], Fresh[2445], Fresh[2444], Fresh[2443], Fresh[2442], Fresh[2441], Fresh[2440], Fresh[2439], Fresh[2438], Fresh[2437], Fresh[2436], Fresh[2435], Fresh[2434], Fresh[2433], Fresh[2432]}), .O ({new_AGEMA_signal_2163, SboxOut[1]}) ) ;
    LUT6_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \Inst_bSbox/b0_4 ( .I0 ({new_AGEMA_signal_1892, \Inst_bSbox/b0 [0]}), .I1 ({new_AGEMA_signal_1891, \Inst_bSbox/b0 [1]}), .I2 ({new_AGEMA_signal_1890, \Inst_bSbox/b0 [2]}), .I3 ({new_AGEMA_signal_1889, \Inst_bSbox/b0 [3]}), .I4 ({new_AGEMA_signal_1438, SboxIn[6]}), .I5 ({new_AGEMA_signal_1436, SboxIn[7]}), .clk (clk), .r ({Fresh[2559], Fresh[2558], Fresh[2557], Fresh[2556], Fresh[2555], Fresh[2554], Fresh[2553], Fresh[2552], Fresh[2551], Fresh[2550], Fresh[2549], Fresh[2548], Fresh[2547], Fresh[2546], Fresh[2545], Fresh[2544], Fresh[2543], Fresh[2542], Fresh[2541], Fresh[2540], Fresh[2539], Fresh[2538], Fresh[2537], Fresh[2536], Fresh[2535], Fresh[2534], Fresh[2533], Fresh[2532], Fresh[2531], Fresh[2530], Fresh[2529], Fresh[2528], Fresh[2527], Fresh[2526], Fresh[2525], Fresh[2524], Fresh[2523], Fresh[2522], Fresh[2521], Fresh[2520], Fresh[2519], Fresh[2518], Fresh[2517], Fresh[2516], Fresh[2515], Fresh[2514], Fresh[2513], Fresh[2512], Fresh[2511], Fresh[2510], Fresh[2509], Fresh[2508], Fresh[2507], Fresh[2506], Fresh[2505], Fresh[2504], Fresh[2503], Fresh[2502], Fresh[2501], Fresh[2500], Fresh[2499], Fresh[2498], Fresh[2497], Fresh[2496]}), .O ({new_AGEMA_signal_2164, SboxOut[0]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hCAFACA0A ) , .MASK ( 5'b01100 ), .INIT2 ( 32'hCAFACA0A ) ) \stateArray/S33reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({plaintext_s1[0], plaintext_s0[0]}), .I1 ({ciphertext_s1[8], ciphertext_s0[8]}), .I2 ({1'b0, nReset_407}), .I3 ({1'b0, \ctrl/finalStep1 }), .I4 ({new_AGEMA_signal_2220, \stateArray/input_MC [0]}), .O ({new_AGEMA_signal_2246, \stateArray/S33reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hCAFACA0A ) , .MASK ( 5'b01100 ), .INIT2 ( 32'hCAFACA0A ) ) \stateArray/S33reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({plaintext_s1[1], plaintext_s0[1]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({1'b0, nReset_407}), .I3 ({1'b0, \ctrl/finalStep1 }), .I4 ({new_AGEMA_signal_2219, \stateArray/input_MC [1]}), .O ({new_AGEMA_signal_2248, \stateArray/S33reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hCAFACA0A ) , .MASK ( 5'b01100 ), .INIT2 ( 32'hCAFACA0A ) ) \stateArray/S33reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({plaintext_s1[2], plaintext_s0[2]}), .I1 ({ciphertext_s1[10], ciphertext_s0[10]}), .I2 ({1'b0, nReset_407}), .I3 ({1'b0, \ctrl/finalStep1 }), .I4 ({new_AGEMA_signal_2218, \stateArray/input_MC [2]}), .O ({new_AGEMA_signal_2250, \stateArray/S33reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hCAFACA0A ) , .MASK ( 5'b01100 ), .INIT2 ( 32'hCAFACA0A ) ) \stateArray/S33reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({plaintext_s1[3], plaintext_s0[3]}), .I1 ({ciphertext_s1[11], ciphertext_s0[11]}), .I2 ({1'b0, nReset_407}), .I3 ({1'b0, \ctrl/finalStep1 }), .I4 ({new_AGEMA_signal_2217, \stateArray/input_MC [3]}), .O ({new_AGEMA_signal_2252, \stateArray/S33reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hCAFACA0A ) , .MASK ( 5'b01100 ), .INIT2 ( 32'hCAFACA0A ) ) \stateArray/S33reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({plaintext_s1[4], plaintext_s0[4]}), .I1 ({ciphertext_s1[12], ciphertext_s0[12]}), .I2 ({1'b0, nReset_407}), .I3 ({1'b0, \ctrl/finalStep1 }), .I4 ({new_AGEMA_signal_2216, \stateArray/input_MC [4]}), .O ({new_AGEMA_signal_2254, \stateArray/S33reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hCAFACA0A ) , .MASK ( 5'b01100 ), .INIT2 ( 32'hCAFACA0A ) ) \stateArray/S33reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({plaintext_s1[5], plaintext_s0[5]}), .I1 ({ciphertext_s1[13], ciphertext_s0[13]}), .I2 ({1'b0, nReset_407}), .I3 ({1'b0, \ctrl/finalStep1 }), .I4 ({new_AGEMA_signal_2215, \stateArray/input_MC [5]}), .O ({new_AGEMA_signal_2256, \stateArray/S33reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hCAFACA0A ) , .MASK ( 5'b01100 ), .INIT2 ( 32'hCAFACA0A ) ) \stateArray/S33reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({plaintext_s1[6], plaintext_s0[6]}), .I1 ({ciphertext_s1[14], ciphertext_s0[14]}), .I2 ({1'b0, nReset_407}), .I3 ({1'b0, \ctrl/finalStep1 }), .I4 ({new_AGEMA_signal_2214, \stateArray/input_MC [6]}), .O ({new_AGEMA_signal_2258, \stateArray/S33reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hCAFACA0A ) , .MASK ( 5'b01100 ), .INIT2 ( 32'hCAFACA0A ) ) \stateArray/S33reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({plaintext_s1[7], plaintext_s0[7]}), .I1 ({ciphertext_s1[15], ciphertext_s0[15]}), .I2 ({1'b0, nReset_407}), .I3 ({1'b0, \ctrl/finalStep1 }), .I4 ({new_AGEMA_signal_2213, \stateArray/input_MC [7]}), .O ({new_AGEMA_signal_2260, \stateArray/S33reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hFCAA0CAA0CAAFCAA ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h0CAAFCAAFCAA0CAA ) ) \KeyArray/S30reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q1 ( .I0 ({key_s1[24], key_s0[24]}), .I1 ({new_AGEMA_signal_1733, \KeyArray/S31reg/gen_ff[1].gff/GEN[0].SFF/Q_603 }), .I2 ({1'b0, \ctrl/CSselMC_835 }), .I3 ({1'b0, nReset_407}), .I4 ({new_AGEMA_signal_1415, N18}), .I5 ({new_AGEMA_signal_2164, SboxOut[0]}), .O ({new_AGEMA_signal_2222, \KeyArray/S30reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hFCAA0CAA0CAAFCAA ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h0CAAFCAAFCAA0CAA ) ) \KeyArray/S30reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q1 ( .I0 ({key_s1[25], key_s0[25]}), .I1 ({new_AGEMA_signal_1736, \KeyArray/S31reg/gen_ff[1].gff/GEN[1].SFF/Q_604 }), .I2 ({1'b0, \ctrl/CSselMC_835 }), .I3 ({1'b0, nReset_407}), .I4 ({new_AGEMA_signal_1416, N20}), .I5 ({new_AGEMA_signal_2163, SboxOut[1]}), .O ({new_AGEMA_signal_2224, \KeyArray/S30reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hFCAA0CAA0CAAFCAA ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h0CAAFCAAFCAA0CAA ) ) \KeyArray/S30reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q1 ( .I0 ({key_s1[26], key_s0[26]}), .I1 ({new_AGEMA_signal_1739, \KeyArray/S31reg/gen_ff[1].gff/GEN[2].SFF/Q_605 }), .I2 ({1'b0, \ctrl/CSselMC_835 }), .I3 ({1'b0, nReset_407}), .I4 ({new_AGEMA_signal_1417, N22}), .I5 ({new_AGEMA_signal_2162, SboxOut[2]}), .O ({new_AGEMA_signal_2226, \KeyArray/S30reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hFCAA0CAA0CAAFCAA ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h0CAAFCAAFCAA0CAA ) ) \KeyArray/S30reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q1 ( .I0 ({key_s1[27], key_s0[27]}), .I1 ({new_AGEMA_signal_1742, \KeyArray/S31reg/gen_ff[1].gff/GEN[3].SFF/Q_606 }), .I2 ({1'b0, \ctrl/CSselMC_835 }), .I3 ({1'b0, nReset_407}), .I4 ({new_AGEMA_signal_1418, N24}), .I5 ({new_AGEMA_signal_2161, SboxOut[3]}), .O ({new_AGEMA_signal_2228, \KeyArray/S30reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hFCAA0CAA0CAAFCAA ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h0CAAFCAAFCAA0CAA ) ) \KeyArray/S30reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q1 ( .I0 ({key_s1[28], key_s0[28]}), .I1 ({new_AGEMA_signal_1745, \KeyArray/S31reg/gen_ff[1].gff/GEN[4].SFF/Q_607 }), .I2 ({1'b0, \ctrl/CSselMC_835 }), .I3 ({1'b0, nReset_407}), .I4 ({new_AGEMA_signal_1419, N26}), .I5 ({new_AGEMA_signal_2160, SboxOut[4]}), .O ({new_AGEMA_signal_2230, \KeyArray/S30reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hFCAA0CAA0CAAFCAA ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h0CAAFCAAFCAA0CAA ) ) \KeyArray/S30reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q1 ( .I0 ({key_s1[29], key_s0[29]}), .I1 ({new_AGEMA_signal_1748, \KeyArray/S31reg/gen_ff[1].gff/GEN[5].SFF/Q_608 }), .I2 ({1'b0, \ctrl/CSselMC_835 }), .I3 ({1'b0, nReset_407}), .I4 ({new_AGEMA_signal_1420, N28}), .I5 ({new_AGEMA_signal_2159, SboxOut[5]}), .O ({new_AGEMA_signal_2232, \KeyArray/S30reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hFCAA0CAA0CAAFCAA ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h0CAAFCAAFCAA0CAA ) ) \KeyArray/S30reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q1 ( .I0 ({key_s1[30], key_s0[30]}), .I1 ({new_AGEMA_signal_1751, \KeyArray/S31reg/gen_ff[1].gff/GEN[6].SFF/Q_609 }), .I2 ({1'b0, \ctrl/CSselMC_835 }), .I3 ({1'b0, nReset_407}), .I4 ({new_AGEMA_signal_1421, N30}), .I5 ({new_AGEMA_signal_2158, SboxOut[6]}), .O ({new_AGEMA_signal_2234, \KeyArray/S30reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hFCAA0CAA0CAAFCAA ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h0CAAFCAAFCAA0CAA ) ) \KeyArray/S30reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q1 ( .I0 ({key_s1[31], key_s0[31]}), .I1 ({new_AGEMA_signal_1754, \KeyArray/S31reg/gen_ff[1].gff/GEN[7].SFF/Q_610 }), .I2 ({1'b0, \ctrl/CSselMC_835 }), .I3 ({1'b0, nReset_407}), .I4 ({new_AGEMA_signal_1422, N32}), .I5 ({new_AGEMA_signal_2157, SboxOut[7]}), .O ({new_AGEMA_signal_2236, \KeyArray/S30reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;

    /* register cells */
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S00reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1927, \stateArray/S00reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[120], ciphertext_s0[120]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S00reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1930, \stateArray/S00reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[121], ciphertext_s0[121]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S00reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1933, \stateArray/S00reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[122], ciphertext_s0[122]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S00reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1936, \stateArray/S00reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[123], ciphertext_s0[123]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S00reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1939, \stateArray/S00reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[124], ciphertext_s0[124]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S00reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1942, \stateArray/S00reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[125], ciphertext_s0[125]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S00reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1945, \stateArray/S00reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[126], ciphertext_s0[126]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S00reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1948, \stateArray/S00reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[127], ciphertext_s0[127]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S01reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1951, \stateArray/S01reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[112], ciphertext_s0[112]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S01reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1954, \stateArray/S01reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[113], ciphertext_s0[113]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S01reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1957, \stateArray/S01reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[114], ciphertext_s0[114]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S01reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1960, \stateArray/S01reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[115], ciphertext_s0[115]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S01reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1963, \stateArray/S01reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[116], ciphertext_s0[116]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S01reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1966, \stateArray/S01reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[117], ciphertext_s0[117]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S01reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1969, \stateArray/S01reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[118], ciphertext_s0[118]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S01reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1972, \stateArray/S01reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[119], ciphertext_s0[119]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S02reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1975, \stateArray/S02reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[104], ciphertext_s0[104]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S02reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1978, \stateArray/S02reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[105], ciphertext_s0[105]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S02reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1981, \stateArray/S02reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[106], ciphertext_s0[106]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S02reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1984, \stateArray/S02reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[107], ciphertext_s0[107]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S02reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1987, \stateArray/S02reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[108], ciphertext_s0[108]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S02reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1990, \stateArray/S02reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[109], ciphertext_s0[109]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S02reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1993, \stateArray/S02reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[110], ciphertext_s0[110]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S02reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1996, \stateArray/S02reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[111], ciphertext_s0[111]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S03reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_2166, \stateArray/S03reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[96], ciphertext_s0[96]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S03reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_2168, \stateArray/S03reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[97], ciphertext_s0[97]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S03reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_2170, \stateArray/S03reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[98], ciphertext_s0[98]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S03reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_2172, \stateArray/S03reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[99], ciphertext_s0[99]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S03reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_2174, \stateArray/S03reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[100], ciphertext_s0[100]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S03reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_2176, \stateArray/S03reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[101], ciphertext_s0[101]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S03reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_2178, \stateArray/S03reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[102], ciphertext_s0[102]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S03reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_2180, \stateArray/S03reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[103], ciphertext_s0[103]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S10reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1455, \stateArray/S10reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[88], ciphertext_s0[88]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S10reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1458, \stateArray/S10reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[89], ciphertext_s0[89]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S10reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1461, \stateArray/S10reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[90], ciphertext_s0[90]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S10reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1464, \stateArray/S10reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[91], ciphertext_s0[91]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S10reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1467, \stateArray/S10reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[92], ciphertext_s0[92]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S10reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1470, \stateArray/S10reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[93], ciphertext_s0[93]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S10reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1473, \stateArray/S10reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[94], ciphertext_s0[94]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S10reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1476, \stateArray/S10reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[95], ciphertext_s0[95]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S11reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1479, \stateArray/S11reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[80], ciphertext_s0[80]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S11reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1482, \stateArray/S11reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[81], ciphertext_s0[81]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S11reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1485, \stateArray/S11reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[82], ciphertext_s0[82]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S11reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1488, \stateArray/S11reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[83], ciphertext_s0[83]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S11reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1491, \stateArray/S11reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[84], ciphertext_s0[84]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S11reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1494, \stateArray/S11reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[85], ciphertext_s0[85]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S11reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1497, \stateArray/S11reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[86], ciphertext_s0[86]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S11reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1500, \stateArray/S11reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[87], ciphertext_s0[87]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S12reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1503, \stateArray/S12reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[72], ciphertext_s0[72]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S12reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1506, \stateArray/S12reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[73], ciphertext_s0[73]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S12reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1509, \stateArray/S12reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[74], ciphertext_s0[74]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S12reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1512, \stateArray/S12reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[75], ciphertext_s0[75]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S12reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1515, \stateArray/S12reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[76], ciphertext_s0[76]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S12reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1518, \stateArray/S12reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[77], ciphertext_s0[77]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S12reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1521, \stateArray/S12reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[78], ciphertext_s0[78]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S12reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1524, \stateArray/S12reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[79], ciphertext_s0[79]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S13reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_2182, \stateArray/S13reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[64], ciphertext_s0[64]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S13reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_2184, \stateArray/S13reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[65], ciphertext_s0[65]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S13reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_2186, \stateArray/S13reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[66], ciphertext_s0[66]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S13reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_2188, \stateArray/S13reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[67], ciphertext_s0[67]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S13reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_2190, \stateArray/S13reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[68], ciphertext_s0[68]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S13reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_2192, \stateArray/S13reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[69], ciphertext_s0[69]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S13reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_2194, \stateArray/S13reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[70], ciphertext_s0[70]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S13reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_2196, \stateArray/S13reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[71], ciphertext_s0[71]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S20reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_2000, \stateArray/S20reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S20reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_2004, \stateArray/S20reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S20reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_2008, \stateArray/S20reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S20reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_2012, \stateArray/S20reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S20reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_2016, \stateArray/S20reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S20reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_2020, \stateArray/S20reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S20reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_2024, \stateArray/S20reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S20reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_2028, \stateArray/S20reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S21reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_2031, \stateArray/S21reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S21reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_2034, \stateArray/S21reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S21reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_2037, \stateArray/S21reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S21reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_2040, \stateArray/S21reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S21reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_2043, \stateArray/S21reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S21reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_2046, \stateArray/S21reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S21reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_2049, \stateArray/S21reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S21reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_2052, \stateArray/S21reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S22reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_2054, \stateArray/S22reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S22reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_2056, \stateArray/S22reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S22reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_2058, \stateArray/S22reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S22reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_2060, \stateArray/S22reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S22reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_2062, \stateArray/S22reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S22reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_2064, \stateArray/S22reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S22reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_2066, \stateArray/S22reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S22reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_2068, \stateArray/S22reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S23reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_2198, \stateArray/S23reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S23reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_2200, \stateArray/S23reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S23reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_2202, \stateArray/S23reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S23reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_2204, \stateArray/S23reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S23reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_2206, \stateArray/S23reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S23reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_2208, \stateArray/S23reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S23reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_2210, \stateArray/S23reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S23reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_2212, \stateArray/S23reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S30reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_2072, \stateArray/S30reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S30reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_2076, \stateArray/S30reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S30reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_2080, \stateArray/S30reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S30reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_2084, \stateArray/S30reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S30reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_2088, \stateArray/S30reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S30reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_2092, \stateArray/S30reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S30reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_2096, \stateArray/S30reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S30reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_2100, \stateArray/S30reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S31reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_2103, \stateArray/S31reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S31reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_2106, \stateArray/S31reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S31reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_2109, \stateArray/S31reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S31reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_2112, \stateArray/S31reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S31reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_2115, \stateArray/S31reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S31reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_2118, \stateArray/S31reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S31reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_2121, \stateArray/S31reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S31reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_2124, \stateArray/S31reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S32reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_2126, \stateArray/S32reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S32reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_2128, \stateArray/S32reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S32reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_2130, \stateArray/S32reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S32reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_2132, \stateArray/S32reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S32reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_2134, \stateArray/S32reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S32reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_2136, \stateArray/S32reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S32reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_2138, \stateArray/S32reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S32reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_2140, \stateArray/S32reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S33reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_2246, \stateArray/S33reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S33reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_2248, \stateArray/S33reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S33reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_2250, \stateArray/S33reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S33reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_2252, \stateArray/S33reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S33reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_2254, \stateArray/S33reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S33reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_2256, \stateArray/S33reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S33reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_2258, \stateArray/S33reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \stateArray/S33reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_2260, \stateArray/S33reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S00reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_2237, \KeyArray/S00reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1371, \KeyArray/S00reg/gen_ff[1].gff/GEN[0].SFF/Q_401 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S00reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_2238, \KeyArray/S00reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1368, \KeyArray/S00reg/gen_ff[1].gff/GEN[1].SFF/Q_400 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S00reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_2239, \KeyArray/S00reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1365, \KeyArray/S00reg/gen_ff[1].gff/GEN[2].SFF/Q_399 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S00reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_2240, \KeyArray/S00reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1362, \KeyArray/S00reg/gen_ff[1].gff/GEN[3].SFF/Q_398 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S00reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_2241, \KeyArray/S00reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1359, \KeyArray/S00reg/gen_ff[1].gff/GEN[4].SFF/Q_397 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S00reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_2242, \KeyArray/S00reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1356, \KeyArray/S00reg/gen_ff[1].gff/GEN[5].SFF/Q_396 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S00reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_2243, \KeyArray/S00reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1353, \KeyArray/S00reg/gen_ff[1].gff/GEN[6].SFF/Q_395 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S00reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_2244, \KeyArray/S00reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1350, \KeyArray/S00reg/gen_ff[1].gff/GEN[7].SFF/Q_394 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S01reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1528, \KeyArray/S01reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1805, \KeyArray/S01reg/gen_ff[1].gff/GEN[0].SFF/Q_691 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S01reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1532, \KeyArray/S01reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1808, \KeyArray/S01reg/gen_ff[1].gff/GEN[1].SFF/Q_692 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S01reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1536, \KeyArray/S01reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1811, \KeyArray/S01reg/gen_ff[1].gff/GEN[2].SFF/Q_693 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S01reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1540, \KeyArray/S01reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1814, \KeyArray/S01reg/gen_ff[1].gff/GEN[3].SFF/Q_694 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S01reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1544, \KeyArray/S01reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1817, \KeyArray/S01reg/gen_ff[1].gff/GEN[4].SFF/Q_695 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S01reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1548, \KeyArray/S01reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1820, \KeyArray/S01reg/gen_ff[1].gff/GEN[5].SFF/Q_696 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S01reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1552, \KeyArray/S01reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1823, \KeyArray/S01reg/gen_ff[1].gff/GEN[6].SFF/Q_697 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S01reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1556, \KeyArray/S01reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1826, \KeyArray/S01reg/gen_ff[1].gff/GEN[7].SFF/Q_698 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S02reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1560, \KeyArray/S02reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1526, \KeyArray/S02reg/gen_ff[1].gff/GEN[0].SFF/Q_683 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S02reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1564, \KeyArray/S02reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1530, \KeyArray/S02reg/gen_ff[1].gff/GEN[1].SFF/Q_684 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S02reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1568, \KeyArray/S02reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1534, \KeyArray/S02reg/gen_ff[1].gff/GEN[2].SFF/Q_685 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S02reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1572, \KeyArray/S02reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1538, \KeyArray/S02reg/gen_ff[1].gff/GEN[3].SFF/Q_686 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S02reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1576, \KeyArray/S02reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1542, \KeyArray/S02reg/gen_ff[1].gff/GEN[4].SFF/Q_687 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S02reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1580, \KeyArray/S02reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1546, \KeyArray/S02reg/gen_ff[1].gff/GEN[5].SFF/Q_688 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S02reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1584, \KeyArray/S02reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1550, \KeyArray/S02reg/gen_ff[1].gff/GEN[6].SFF/Q_689 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S02reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1588, \KeyArray/S02reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1554, \KeyArray/S02reg/gen_ff[1].gff/GEN[7].SFF/Q_690 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S03reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1591, \KeyArray/S03reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1558, \KeyArray/S03reg/gen_ff[1].gff/GEN[0].SFF/Q_675 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S03reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1594, \KeyArray/S03reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1562, \KeyArray/S03reg/gen_ff[1].gff/GEN[1].SFF/Q_676 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S03reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1597, \KeyArray/S03reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1566, \KeyArray/S03reg/gen_ff[1].gff/GEN[2].SFF/Q_677 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S03reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1600, \KeyArray/S03reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1570, \KeyArray/S03reg/gen_ff[1].gff/GEN[3].SFF/Q_678 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S03reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1603, \KeyArray/S03reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1574, \KeyArray/S03reg/gen_ff[1].gff/GEN[4].SFF/Q_679 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S03reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1606, \KeyArray/S03reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1578, \KeyArray/S03reg/gen_ff[1].gff/GEN[5].SFF/Q_680 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S03reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1609, \KeyArray/S03reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1582, \KeyArray/S03reg/gen_ff[1].gff/GEN[6].SFF/Q_681 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S03reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1612, \KeyArray/S03reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1586, \KeyArray/S03reg/gen_ff[1].gff/GEN[7].SFF/Q_682 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S10reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1615, \KeyArray/S10reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1589, \KeyArray/S10reg/gen_ff[1].gff/GEN[0].SFF/Q_667 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S10reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1618, \KeyArray/S10reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1592, \KeyArray/S10reg/gen_ff[1].gff/GEN[1].SFF/Q_668 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S10reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1621, \KeyArray/S10reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1595, \KeyArray/S10reg/gen_ff[1].gff/GEN[2].SFF/Q_669 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S10reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1624, \KeyArray/S10reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1598, \KeyArray/S10reg/gen_ff[1].gff/GEN[3].SFF/Q_670 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S10reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1627, \KeyArray/S10reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1601, \KeyArray/S10reg/gen_ff[1].gff/GEN[4].SFF/Q_671 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S10reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1630, \KeyArray/S10reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1604, \KeyArray/S10reg/gen_ff[1].gff/GEN[5].SFF/Q_672 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S10reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1633, \KeyArray/S10reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1607, \KeyArray/S10reg/gen_ff[1].gff/GEN[6].SFF/Q_673 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S10reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1636, \KeyArray/S10reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1610, \KeyArray/S10reg/gen_ff[1].gff/GEN[7].SFF/Q_674 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S11reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1639, \KeyArray/S11reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1525, \KeyArray/S11reg/gen_ff[1].gff/GEN[0].SFF/Q_659 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S11reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1642, \KeyArray/S11reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1529, \KeyArray/S11reg/gen_ff[1].gff/GEN[1].SFF/Q_660 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S11reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1645, \KeyArray/S11reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1533, \KeyArray/S11reg/gen_ff[1].gff/GEN[2].SFF/Q_661 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S11reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1648, \KeyArray/S11reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1537, \KeyArray/S11reg/gen_ff[1].gff/GEN[3].SFF/Q_662 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S11reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1651, \KeyArray/S11reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1541, \KeyArray/S11reg/gen_ff[1].gff/GEN[4].SFF/Q_663 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S11reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1654, \KeyArray/S11reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1545, \KeyArray/S11reg/gen_ff[1].gff/GEN[5].SFF/Q_664 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S11reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1657, \KeyArray/S11reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1549, \KeyArray/S11reg/gen_ff[1].gff/GEN[6].SFF/Q_665 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S11reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1660, \KeyArray/S11reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1553, \KeyArray/S11reg/gen_ff[1].gff/GEN[7].SFF/Q_666 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S12reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1663, \KeyArray/S12reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1557, \KeyArray/S12reg/gen_ff[1].gff/GEN[0].SFF/Q_651 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S12reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1666, \KeyArray/S12reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1561, \KeyArray/S12reg/gen_ff[1].gff/GEN[1].SFF/Q_652 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S12reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1669, \KeyArray/S12reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1565, \KeyArray/S12reg/gen_ff[1].gff/GEN[2].SFF/Q_653 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S12reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1672, \KeyArray/S12reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1569, \KeyArray/S12reg/gen_ff[1].gff/GEN[3].SFF/Q_654 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S12reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1675, \KeyArray/S12reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1573, \KeyArray/S12reg/gen_ff[1].gff/GEN[4].SFF/Q_655 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S12reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1678, \KeyArray/S12reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1577, \KeyArray/S12reg/gen_ff[1].gff/GEN[5].SFF/Q_656 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S12reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1681, \KeyArray/S12reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1581, \KeyArray/S12reg/gen_ff[1].gff/GEN[6].SFF/Q_657 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S12reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1684, \KeyArray/S12reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1585, \KeyArray/S12reg/gen_ff[1].gff/GEN[7].SFF/Q_658 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S13reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1687, \KeyArray/S13reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1433, \KeyArray/S13reg/gen_ff[1].gff/GEN[0].SFF/Q_393 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S13reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1690, \KeyArray/S13reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1431, \KeyArray/S13reg/gen_ff[1].gff/GEN[1].SFF/Q_392 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S13reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1693, \KeyArray/S13reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1429, \KeyArray/S13reg/gen_ff[1].gff/GEN[2].SFF/Q_391 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S13reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1696, \KeyArray/S13reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1427, \KeyArray/S13reg/gen_ff[1].gff/GEN[3].SFF/Q_390 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S13reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1699, \KeyArray/S13reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1425, \KeyArray/S13reg/gen_ff[1].gff/GEN[4].SFF/Q_389 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S13reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1702, \KeyArray/S13reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1423, \KeyArray/S13reg/gen_ff[1].gff/GEN[5].SFF/Q_388 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S13reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1705, \KeyArray/S13reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1437, \KeyArray/S13reg/gen_ff[1].gff/GEN[6].SFF/Q_387 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S13reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1708, \KeyArray/S13reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1435, \KeyArray/S13reg/gen_ff[1].gff/GEN[7].SFF/Q_386 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S20reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1711, \KeyArray/S20reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1613, \KeyArray/S20reg/gen_ff[1].gff/GEN[0].SFF/Q_643 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S20reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1714, \KeyArray/S20reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1616, \KeyArray/S20reg/gen_ff[1].gff/GEN[1].SFF/Q_644 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S20reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1717, \KeyArray/S20reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1619, \KeyArray/S20reg/gen_ff[1].gff/GEN[2].SFF/Q_645 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S20reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1720, \KeyArray/S20reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1622, \KeyArray/S20reg/gen_ff[1].gff/GEN[3].SFF/Q_646 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S20reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1723, \KeyArray/S20reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1625, \KeyArray/S20reg/gen_ff[1].gff/GEN[4].SFF/Q_647 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S20reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1726, \KeyArray/S20reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1628, \KeyArray/S20reg/gen_ff[1].gff/GEN[5].SFF/Q_648 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S20reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1729, \KeyArray/S20reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1631, \KeyArray/S20reg/gen_ff[1].gff/GEN[6].SFF/Q_649 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S20reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1732, \KeyArray/S20reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1634, \KeyArray/S20reg/gen_ff[1].gff/GEN[7].SFF/Q_650 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S21reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1735, \KeyArray/S21reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1637, \KeyArray/S21reg/gen_ff[1].gff/GEN[0].SFF/Q_635 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S21reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1738, \KeyArray/S21reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1640, \KeyArray/S21reg/gen_ff[1].gff/GEN[1].SFF/Q_636 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S21reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1741, \KeyArray/S21reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1643, \KeyArray/S21reg/gen_ff[1].gff/GEN[2].SFF/Q_637 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S21reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1744, \KeyArray/S21reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1646, \KeyArray/S21reg/gen_ff[1].gff/GEN[3].SFF/Q_638 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S21reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1747, \KeyArray/S21reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1649, \KeyArray/S21reg/gen_ff[1].gff/GEN[4].SFF/Q_639 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S21reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1750, \KeyArray/S21reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1652, \KeyArray/S21reg/gen_ff[1].gff/GEN[5].SFF/Q_640 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S21reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1753, \KeyArray/S21reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1655, \KeyArray/S21reg/gen_ff[1].gff/GEN[6].SFF/Q_641 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S21reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1756, \KeyArray/S21reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1658, \KeyArray/S21reg/gen_ff[1].gff/GEN[7].SFF/Q_642 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S22reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1759, \KeyArray/S22reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1661, \KeyArray/S22reg/gen_ff[1].gff/GEN[0].SFF/Q_627 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S22reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1762, \KeyArray/S22reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1664, \KeyArray/S22reg/gen_ff[1].gff/GEN[1].SFF/Q_628 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S22reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1765, \KeyArray/S22reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1667, \KeyArray/S22reg/gen_ff[1].gff/GEN[2].SFF/Q_629 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S22reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1768, \KeyArray/S22reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1670, \KeyArray/S22reg/gen_ff[1].gff/GEN[3].SFF/Q_630 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S22reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1771, \KeyArray/S22reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1673, \KeyArray/S22reg/gen_ff[1].gff/GEN[4].SFF/Q_631 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S22reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1774, \KeyArray/S22reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1676, \KeyArray/S22reg/gen_ff[1].gff/GEN[5].SFF/Q_632 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S22reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1777, \KeyArray/S22reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1679, \KeyArray/S22reg/gen_ff[1].gff/GEN[6].SFF/Q_633 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S22reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1780, \KeyArray/S22reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1682, \KeyArray/S22reg/gen_ff[1].gff/GEN[7].SFF/Q_634 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S23reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1783, \KeyArray/S23reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1685, \KeyArray/S23reg/gen_ff[1].gff/GEN[0].SFF/Q_619 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S23reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1786, \KeyArray/S23reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1688, \KeyArray/S23reg/gen_ff[1].gff/GEN[1].SFF/Q_620 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S23reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1789, \KeyArray/S23reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1691, \KeyArray/S23reg/gen_ff[1].gff/GEN[2].SFF/Q_621 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S23reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1792, \KeyArray/S23reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1694, \KeyArray/S23reg/gen_ff[1].gff/GEN[3].SFF/Q_622 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S23reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1795, \KeyArray/S23reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1697, \KeyArray/S23reg/gen_ff[1].gff/GEN[4].SFF/Q_623 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S23reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1798, \KeyArray/S23reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1700, \KeyArray/S23reg/gen_ff[1].gff/GEN[5].SFF/Q_624 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S23reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1801, \KeyArray/S23reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1703, \KeyArray/S23reg/gen_ff[1].gff/GEN[6].SFF/Q_625 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S23reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1804, \KeyArray/S23reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1706, \KeyArray/S23reg/gen_ff[1].gff/GEN[7].SFF/Q_626 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S30reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_2222, \KeyArray/S30reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1709, \KeyArray/S30reg/gen_ff[1].gff/GEN[0].SFF/Q_611 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S30reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_2224, \KeyArray/S30reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1712, \KeyArray/S30reg/gen_ff[1].gff/GEN[1].SFF/Q_612 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S30reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_2226, \KeyArray/S30reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1715, \KeyArray/S30reg/gen_ff[1].gff/GEN[2].SFF/Q_613 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S30reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_2228, \KeyArray/S30reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1718, \KeyArray/S30reg/gen_ff[1].gff/GEN[3].SFF/Q_614 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S30reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_2230, \KeyArray/S30reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1721, \KeyArray/S30reg/gen_ff[1].gff/GEN[4].SFF/Q_615 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S30reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_2232, \KeyArray/S30reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1724, \KeyArray/S30reg/gen_ff[1].gff/GEN[5].SFF/Q_616 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S30reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_2234, \KeyArray/S30reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1727, \KeyArray/S30reg/gen_ff[1].gff/GEN[6].SFF/Q_617 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S30reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_2236, \KeyArray/S30reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1730, \KeyArray/S30reg/gen_ff[1].gff/GEN[7].SFF/Q_618 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S31reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1807, \KeyArray/S31reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1733, \KeyArray/S31reg/gen_ff[1].gff/GEN[0].SFF/Q_603 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S31reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1810, \KeyArray/S31reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1736, \KeyArray/S31reg/gen_ff[1].gff/GEN[1].SFF/Q_604 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S31reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1813, \KeyArray/S31reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1739, \KeyArray/S31reg/gen_ff[1].gff/GEN[2].SFF/Q_605 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S31reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1816, \KeyArray/S31reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1742, \KeyArray/S31reg/gen_ff[1].gff/GEN[3].SFF/Q_606 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S31reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1819, \KeyArray/S31reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1745, \KeyArray/S31reg/gen_ff[1].gff/GEN[4].SFF/Q_607 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S31reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1822, \KeyArray/S31reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1748, \KeyArray/S31reg/gen_ff[1].gff/GEN[5].SFF/Q_608 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S31reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1825, \KeyArray/S31reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1751, \KeyArray/S31reg/gen_ff[1].gff/GEN[6].SFF/Q_609 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S31reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1828, \KeyArray/S31reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1754, \KeyArray/S31reg/gen_ff[1].gff/GEN[7].SFF/Q_610 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S32reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1830, \KeyArray/S32reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1757, \KeyArray/S32reg/gen_ff[1].gff/GEN[0].SFF/Q_595 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S32reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1832, \KeyArray/S32reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1760, \KeyArray/S32reg/gen_ff[1].gff/GEN[1].SFF/Q_596 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S32reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1834, \KeyArray/S32reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1763, \KeyArray/S32reg/gen_ff[1].gff/GEN[2].SFF/Q_597 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S32reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1836, \KeyArray/S32reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1766, \KeyArray/S32reg/gen_ff[1].gff/GEN[3].SFF/Q_598 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S32reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1838, \KeyArray/S32reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1769, \KeyArray/S32reg/gen_ff[1].gff/GEN[4].SFF/Q_599 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S32reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1840, \KeyArray/S32reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1772, \KeyArray/S32reg/gen_ff[1].gff/GEN[5].SFF/Q_600 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S32reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1842, \KeyArray/S32reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1775, \KeyArray/S32reg/gen_ff[1].gff/GEN[6].SFF/Q_601 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S32reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1844, \KeyArray/S32reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1778, \KeyArray/S32reg/gen_ff[1].gff/GEN[7].SFF/Q_602 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S33reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1846, \KeyArray/S33reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1781, \KeyArray/S33reg/gen_ff[1].gff/GEN[0].SFF/Q_587 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S33reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1848, \KeyArray/S33reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1784, \KeyArray/S33reg/gen_ff[1].gff/GEN[1].SFF/Q_588 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S33reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1850, \KeyArray/S33reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1787, \KeyArray/S33reg/gen_ff[1].gff/GEN[2].SFF/Q_589 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S33reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1852, \KeyArray/S33reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1790, \KeyArray/S33reg/gen_ff[1].gff/GEN[3].SFF/Q_590 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S33reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1854, \KeyArray/S33reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1793, \KeyArray/S33reg/gen_ff[1].gff/GEN[4].SFF/Q_591 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S33reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1856, \KeyArray/S33reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1796, \KeyArray/S33reg/gen_ff[1].gff/GEN[5].SFF/Q_592 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S33reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1858, \KeyArray/S33reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1799, \KeyArray/S33reg/gen_ff[1].gff/GEN[6].SFF/Q_593 }) ) ;
    FDE_masked #(.low_latency(1), .pipeline(0)) \KeyArray/S33reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1860, \KeyArray/S33reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1802, \KeyArray/S33reg/gen_ff[1].gff/GEN[7].SFF/Q_594 }) ) ;
    FD \ctrl/seq4/GEN[1].SFF/Q ( .D (\ctrl/seq4/GEN[1].SFF/QD ), .C (clk_gated), .Q (\ctrl/seq4/GEN[1].SFF/Q_837 ) ) ;
    FD \ctrl/seq4/GEN[0].SFF/Q ( .D (\ctrl/seq4/GEN[0].SFF/QD ), .C (clk_gated), .Q (\ctrl/seq4/GEN[0].SFF/Q_836 ) ) ;
    FD \ctrl/seq6/GEN[4].SFF/Q ( .D (\ctrl/seq6/GEN[4].SFF/QD ), .C (clk_gated), .Q (\ctrl/seq6/GEN[4].SFF/Q_842 ) ) ;
    FD \ctrl/seq6/GEN[3].SFF/Q ( .D (\ctrl/seq6/GEN[3].SFF/QD ), .C (clk_gated), .Q (\ctrl/seq6/GEN[3].SFF/Q_840 ) ) ;
    FD \ctrl/seq6/GEN[2].SFF/Q ( .D (\ctrl/seq6/GEN[2].SFF/QD ), .C (clk_gated), .Q (\ctrl/seq6/GEN[2].SFF/Q_839 ) ) ;
    FD \ctrl/seq6/GEN[1].SFF/Q ( .D (\ctrl/seq6/GEN[1].SFF/QD ), .C (clk_gated), .Q (\ctrl/seq6/GEN[1].SFF/Q_838 ) ) ;
    FD \ctrl/seq6/GEN[0].SFF/Q ( .D (\ctrl/seq6/GEN[0].SFF/QD ), .C (clk_gated), .Q (\ctrl/seq6/GEN[0].SFF/Q_841 ) ) ;
    FDR \ctrl/CSenRC ( .D (\ctrl/finalStep1 ), .C (clk_gated), .R (\calcRCon/nReset_inv ), .Q (\ctrl/CSenRC_405 ) ) ;
    FDSE \calcRCon/s_current_state_7 ( .D (\calcRCon/s_current_state [6]), .C (clk_gated), .CE (selSR), .S (\calcRCon/nReset_inv ), .Q (\calcRCon/s_current_state [7]) ) ;
    FDRE \calcRCon/s_current_state_6 ( .D (\calcRCon/s_current_state [5]), .C (clk_gated), .CE (selSR), .R (\calcRCon/nReset_inv ), .Q (\calcRCon/s_current_state [6]) ) ;
    FDRE \calcRCon/s_current_state_5 ( .D (\calcRCon/s_current_state [4]), .C (clk_gated), .CE (selSR), .R (\calcRCon/nReset_inv ), .Q (\calcRCon/s_current_state [5]) ) ;
    FDRE \calcRCon/s_current_state_4 ( .D (\calcRCon/MSB_s_current_state[3]_XOR_19_o ), .C (clk_gated), .CE (selSR), .R (\calcRCon/nReset_inv ), .Q (\calcRCon/s_current_state [4]) ) ;
    FDSE \calcRCon/s_current_state_3 ( .D (\calcRCon/MSB_s_current_state[2]_XOR_20_o ), .C (clk_gated), .CE (selSR), .S (\calcRCon/nReset_inv ), .Q (\calcRCon/s_current_state [3]) ) ;
    FDSE \calcRCon/s_current_state_2 ( .D (\calcRCon/s_current_state [1]), .C (clk_gated), .CE (selSR), .S (\calcRCon/nReset_inv ), .Q (\calcRCon/s_current_state [2]) ) ;
    FDRE \calcRCon/s_current_state_1 ( .D (\calcRCon/MSB_s_current_state[0]_XOR_21_o ), .C (clk_gated), .CE (selSR), .R (\calcRCon/nReset_inv ), .Q (\calcRCon/s_current_state [1]) ) ;
    FDSE \calcRCon/s_current_state_0 ( .D (\calcRCon/s_current_state [7]), .C (clk_gated), .CE (selSR), .S (\calcRCon/nReset_inv ), .Q (\calcRCon/s_current_state [0]) ) ;
    FDR \ctrl/CSselMC ( .D (\ctrl/CSselMC_rstpot_1330 ), .C (clk_gated), .R (\calcRCon/nReset_inv ), .Q (\ctrl/CSselMC_835 ) ) ;
    FD nReset ( .D (nReset_rstpot), .C (clk_gated), .Q (nReset_407) ) ;
    FD nReset_1 ( .D (nReset_rstpot), .C (clk_gated), .Q (nReset_1_1341) ) ;
    FDR \ctrl/CSselMC_1 ( .D (\ctrl/CSselMC_rstpot_1330 ), .C (clk_gated), .R (\calcRCon/nReset_inv ), .Q (\ctrl/CSselMC_1_1342 ) ) ;
endmodule
